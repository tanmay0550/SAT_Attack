module b14_c (key_124, pi055, pi233, pi152, key_123, pi025, key_0, key_103, key_53, key_95, pi277, pi238, pi030, pi003, key_55, pi209, pi122, key_82, pi172, pi225, key_85, pi056, pi004, pi053, pi222, pi181, pi080, key_92, pi073, pi162, pi249, pi102, pi151, pi226, pi244, pi200, pi067, key_113, pi119, pi107, pi248, pi063, key_58, pi160, pi228, pi011, pi000, pi240, pi024, pi016, pi079, pi274, pi118, pi116, pi157, pi177, key_44, pi001, pi220, pi180, pi094, pi147, pi048, pi066, key_90, key_52, pi114, pi188, pi123, pi149, pi256, pi031, key_98, pi137, key_97, pi236, pi133, key_62, pi027, pi266, pi065, pi198, key_29, key_78, pi093, pi171, pi271, pi202, key_73, pi251, pi213, pi129, key_6, pi154, key_23, pi159, pi212, key_111, pi207, pi097, pi108, pi121, pi099, pi245, pi084, pi237, key_42, pi275, key_49, key_81, key_127, pi128, key_79, pi218, key_76, pi221, pi106, pi044, pi223, pi098, pi216, pi096, pi179, key_48, pi126, pi047, pi113, pi205, pi243, key_57, key_84, pi270, pi092, pi006, pi101, pi214, pi005, pi242, key_71, pi258, key_118, pi026, key_100, pi259, key_46, key_56, pi206, pi075, pi131, pi071, pi196, pi002, key_102, pi230, key_20, pi183, pi022, pi211, pi234, pi132, pi034, pi199, key_14, key_25, pi130, pi197, pi095, key_9, pi058, key_22, pi190, pi032, pi057, pi260, pi148, key_26, key_106, pi265, pi269, pi232, pi253, pi061, key_86, key_34, pi029, pi201, pi224, pi117, pi146, pi276, pi164, key_3, key_1, pi009, pi125, pi104, key_51, pi010, key_96, pi115, pi062, key_54, pi247, pi150, pi081, key_66, key_91, key_31, key_40, pi017, pi127, key_60, pi219, key_101, pi167, key_122, pi241, pi135, pi134, pi111, pi054, key_74, pi268, key_18, pi174, pi007, key_12, key_87, pi227, pi090, pi077, pi020, pi109, pi076, key_109, key_108, key_115, pi087, key_37, pi273, pi239, key_105, pi086, pi215, pi195, pi050, pi136, key_99, pi124, pi175, pi141, key_120, key_7, pi250, pi046, pi252, pi043, key_35, key_64, pi153, pi110, pi204, pi038, key_93, pi083, key_125, pi161, key_104, key_59, pi182, pi089, key_65, pi235, key_89, key_32, pi142, pi156, pi035, pi138, pi008, pi120, pi184, key_63, key_21, key_43, pi264, pi143, pi015, pi033, pi165, key_83, key_41, pi021, pi208, pi045, pi082, pi052, pi014, key_114, pi186, pi049, key_13, pi069, key_77, pi068, pi255, key_126, key_5, pi178, pi192, pi064, key_107, pi041, key_112, pi019, pi170, key_110, key_75, pi072, pi173, pi012, pi189, key_94, pi217, pi091, pi039, pi185, pi229, key_70, pi085, key_38, key_116, pi078, key_33, key_15, pi193, pi144, key_17, key_4, pi105, pi145, pi018, key_72, pi261, pi267, pi028, key_80, pi257, key_119, key_121, pi168, pi187, key_50, key_117, key_36, pi042, key_61, key_16, pi139, key_45, pi074, pi051, pi194, pi191, pi059, pi023, pi203, pi176, key_10, pi103, pi013, key_67, pi037, pi169, pi210, key_69, pi060, pi100, pi112, key_88, pi272, pi254, key_30, pi040, key_24, key_39, pi036, key_27, pi070, pi088, key_19, pi262, key_2, key_8, pi263, pi231, pi155, key_68, pi166, pi163, key_47, pi158, key_11, key_28, pi140, pi246, po131, po242, po255, po153, po121, po298, po286, po209, po007, po175, po295, po280, po269, po243, po181, po192, po139, po003, po200, po253, po056, po290, po249, po024, po041, po066, po138, po045, po282, po005, po241, po135, po002, po073, po164, po189, po070, po188, po165, po010, po094, po231, po142, po207, po236, po186, po177, po220, po157, po074, po271, po085, po163, po229, po173, po266, po247, po054, po162, po180, po127, po133, po225, po219, po090, po159, po093, po086, po075, po014, po050, po223, po061, po289, po263, po016, po122, po167, po096, po136, po176, po254, po020, po106, po117, po018, po203, po276, po288, po196, po152, po281, po216, po055, po035, po051, po033, po124, po046, po060, po026, po279, po047, po083, po224, po065, po259, po022, po036, po063, po168, po184, po091, po030, po037, po006, po208, po058, po049, po234, po155, po277, po150, po227, po143, po119, po272, po008, po178, po068, po004, po252, po078, po023, po161, po108, po154, po206, po204, po213, po250, po267, po011, po017, po183, po042, po071, po239, po048, po098, po021, po062, po221, po262, po202, po028, po171, po187, po287, po103, po115, po230, po232, po240, po278, po097, po087, po053, po233, po248, po214, po100, po256, po116, po251, po092, po081, po118, po015, po000, po009, po012, po112, po275, po120, po258, po025, po274, po195, po193, po273, po113, po257, po027, po179, po137, po140, po218, po141, po109, po151, po210, po105, po235, po264, po268, po043, po114, po190, po072, po031, po201, po284, po082, po194, po246, po032, po019, po169, po158, po059, po244, po270, po039, po101, po222, po228, po129, po148, po089, po077, po001, po174, po095, po110, po293, po198, po052, po013, po185, po261, po069, po226, po283, po166, po170, po146, po147, po029, po217, po199, po044, po126, po237, po102, po292, po156, po057, po297, po260, po172, po145, po079, po238, po191, po182, po034, po125, po291, po067, po088, po197, po205, po132, po107, po076, po064, po111, po215, po134, po160, po080, po149, po104, po296, po130, po212, po128, po294, po123, po040, po038, po144, po285, po084, po265, po099, po211, po245);
  input key_124;
  input pi055;
  input pi233;
  input pi152;
  input key_123;
  input pi025;
  input key_0;
  input key_103;
  input key_53;
  input key_95;
  input pi277;
  input pi238;
  input pi030;
  input pi003;
  input key_55;
  input pi209;
  input pi122;
  input key_82;
  input pi172;
  input pi225;
  input key_85;
  input pi056;
  input pi004;
  input pi053;
  input pi222;
  input pi181;
  input pi080;
  input key_92;
  input pi073;
  input pi162;
  input pi249;
  input pi102;
  input pi151;
  input pi226;
  input pi244;
  input pi200;
  input pi067;
  input key_113;
  input pi119;
  input pi107;
  input pi248;
  input pi063;
  input key_58;
  input pi160;
  input pi228;
  input pi011;
  input pi000;
  input pi240;
  input pi024;
  input pi016;
  input pi079;
  input pi274;
  input pi118;
  input pi116;
  input pi157;
  input pi177;
  input key_44;
  input pi001;
  input pi220;
  input pi180;
  input pi094;
  input pi147;
  input pi048;
  input pi066;
  input key_90;
  input key_52;
  input pi114;
  input pi188;
  input pi123;
  input pi149;
  input pi256;
  input pi031;
  input key_98;
  input pi137;
  input key_97;
  input pi236;
  input pi133;
  input key_62;
  input pi027;
  input pi266;
  input pi065;
  input pi198;
  input key_29;
  input key_78;
  input pi093;
  input pi171;
  input pi271;
  input pi202;
  input key_73;
  input pi251;
  input pi213;
  input pi129;
  input key_6;
  input pi154;
  input key_23;
  input pi159;
  input pi212;
  input key_111;
  input pi207;
  input pi097;
  input pi108;
  input pi121;
  input pi099;
  input pi245;
  input pi084;
  input pi237;
  input key_42;
  input pi275;
  input key_49;
  input key_81;
  input key_127;
  input pi128;
  input key_79;
  input pi218;
  input key_76;
  input pi221;
  input pi106;
  input pi044;
  input pi223;
  input pi098;
  input pi216;
  input pi096;
  input pi179;
  input key_48;
  input pi126;
  input pi047;
  input pi113;
  input pi205;
  input pi243;
  input key_57;
  input key_84;
  input pi270;
  input pi092;
  input pi006;
  input pi101;
  input pi214;
  input pi005;
  input pi242;
  input key_71;
  input pi258;
  input key_118;
  input pi026;
  input key_100;
  input pi259;
  input key_46;
  input key_56;
  input pi206;
  input pi075;
  input pi131;
  input pi071;
  input pi196;
  input pi002;
  input key_102;
  input pi230;
  input key_20;
  input pi183;
  input pi022;
  input pi211;
  input pi234;
  input pi132;
  input pi034;
  input pi199;
  input key_14;
  input key_25;
  input pi130;
  input pi197;
  input pi095;
  input key_9;
  input pi058;
  input key_22;
  input pi190;
  input pi032;
  input pi057;
  input pi260;
  input pi148;
  input key_26;
  input key_106;
  input pi265;
  input pi269;
  input pi232;
  input pi253;
  input pi061;
  input key_86;
  input key_34;
  input pi029;
  input pi201;
  input pi224;
  input pi117;
  input pi146;
  input pi276;
  input pi164;
  input key_3;
  input key_1;
  input pi009;
  input pi125;
  input pi104;
  input key_51;
  input pi010;
  input key_96;
  input pi115;
  input pi062;
  input key_54;
  input pi247;
  input pi150;
  input pi081;
  input key_66;
  input key_91;
  input key_31;
  input key_40;
  input pi017;
  input pi127;
  input key_60;
  input pi219;
  input key_101;
  input pi167;
  input key_122;
  input pi241;
  input pi135;
  input pi134;
  input pi111;
  input pi054;
  input key_74;
  input pi268;
  input key_18;
  input pi174;
  input pi007;
  input key_12;
  input key_87;
  input pi227;
  input pi090;
  input pi077;
  input pi020;
  input pi109;
  input pi076;
  input key_109;
  input key_108;
  input key_115;
  input pi087;
  input key_37;
  input pi273;
  input pi239;
  input key_105;
  input pi086;
  input pi215;
  input pi195;
  input pi050;
  input pi136;
  input key_99;
  input pi124;
  input pi175;
  input pi141;
  input key_120;
  input key_7;
  input pi250;
  input pi046;
  input pi252;
  input pi043;
  input key_35;
  input key_64;
  input pi153;
  input pi110;
  input pi204;
  input pi038;
  input key_93;
  input pi083;
  input key_125;
  input pi161;
  input key_104;
  input key_59;
  input pi182;
  input pi089;
  input key_65;
  input pi235;
  input key_89;
  input key_32;
  input pi142;
  input pi156;
  input pi035;
  input pi138;
  input pi008;
  input pi120;
  input pi184;
  input key_63;
  input key_21;
  input key_43;
  input pi264;
  input pi143;
  input pi015;
  input pi033;
  input pi165;
  input key_83;
  input key_41;
  input pi021;
  input pi208;
  input pi045;
  input pi082;
  input pi052;
  input pi014;
  input key_114;
  input pi186;
  input pi049;
  input key_13;
  input pi069;
  input key_77;
  input pi068;
  input pi255;
  input key_126;
  input key_5;
  input pi178;
  input pi192;
  input pi064;
  input key_107;
  input pi041;
  input key_112;
  input pi019;
  input pi170;
  input key_110;
  input key_75;
  input pi072;
  input pi173;
  input pi012;
  input pi189;
  input key_94;
  input pi217;
  input pi091;
  input pi039;
  input pi185;
  input pi229;
  input key_70;
  input pi085;
  input key_38;
  input key_116;
  input pi078;
  input key_33;
  input key_15;
  input pi193;
  input pi144;
  input key_17;
  input key_4;
  input pi105;
  input pi145;
  input pi018;
  input key_72;
  input pi261;
  input pi267;
  input pi028;
  input key_80;
  input pi257;
  input key_119;
  input key_121;
  input pi168;
  input pi187;
  input key_50;
  input key_117;
  input key_36;
  input pi042;
  input key_61;
  input key_16;
  input pi139;
  input key_45;
  input pi074;
  input pi051;
  input pi194;
  input pi191;
  input pi059;
  input pi023;
  input pi203;
  input pi176;
  input key_10;
  input pi103;
  input pi013;
  input key_67;
  input pi037;
  input pi169;
  input pi210;
  input key_69;
  input pi060;
  input pi100;
  input pi112;
  input key_88;
  input pi272;
  input pi254;
  input key_30;
  input pi040;
  input key_24;
  input key_39;
  input pi036;
  input key_27;
  input pi070;
  input pi088;
  input key_19;
  input pi262;
  input key_2;
  input key_8;
  input pi263;
  input pi231;
  input pi155;
  input key_68;
  input pi166;
  input pi163;
  input key_47;
  input pi158;
  input key_11;
  input key_28;
  input pi140;
  input pi246;

  output po131;
  output po242;
  output po255;
  output po153;
  output po121;
  output po298;
  output po286;
  output po209;
  output po007;
  output po175;
  output po295;
  output po280;
  output po269;
  output po243;
  output po181;
  output po192;
  output po139;
  output po003;
  output po200;
  output po253;
  output po056;
  output po290;
  output po249;
  output po024;
  output po041;
  output po066;
  output po138;
  output po045;
  output po282;
  output po005;
  output po241;
  output po135;
  output po002;
  output po073;
  output po164;
  output po189;
  output po070;
  output po188;
  output po165;
  output po010;
  output po094;
  output po231;
  output po142;
  output po207;
  output po236;
  output po186;
  output po177;
  output po220;
  output po157;
  output po074;
  output po271;
  output po085;
  output po163;
  output po229;
  output po173;
  output po266;
  output po247;
  output po054;
  output po162;
  output po180;
  output po127;
  output po133;
  output po225;
  output po219;
  output po090;
  output po159;
  output po093;
  output po086;
  output po075;
  output po014;
  output po050;
  output po223;
  output po061;
  output po289;
  output po263;
  output po016;
  output po122;
  output po167;
  output po096;
  output po136;
  output po176;
  output po254;
  output po020;
  output po106;
  output po117;
  output po018;
  output po203;
  output po276;
  output po288;
  output po196;
  output po152;
  output po281;
  output po216;
  output po055;
  output po035;
  output po051;
  output po033;
  output po124;
  output po046;
  output po060;
  output po026;
  output po279;
  output po047;
  output po083;
  output po224;
  output po065;
  output po259;
  output po022;
  output po036;
  output po063;
  output po168;
  output po184;
  output po091;
  output po030;
  output po037;
  output po006;
  output po208;
  output po058;
  output po049;
  output po234;
  output po155;
  output po277;
  output po150;
  output po227;
  output po143;
  output po119;
  output po272;
  output po008;
  output po178;
  output po068;
  output po004;
  output po252;
  output po078;
  output po023;
  output po161;
  output po108;
  output po154;
  output po206;
  output po204;
  output po213;
  output po250;
  output po267;
  output po011;
  output po017;
  output po183;
  output po042;
  output po071;
  output po239;
  output po048;
  output po098;
  output po021;
  output po062;
  output po221;
  output po262;
  output po202;
  output po028;
  output po171;
  output po187;
  output po287;
  output po103;
  output po115;
  output po230;
  output po232;
  output po240;
  output po278;
  output po097;
  output po087;
  output po053;
  output po233;
  output po248;
  output po214;
  output po100;
  output po256;
  output po116;
  output po251;
  output po092;
  output po081;
  output po118;
  output po015;
  output po000;
  output po009;
  output po012;
  output po112;
  output po275;
  output po120;
  output po258;
  output po025;
  output po274;
  output po195;
  output po193;
  output po273;
  output po113;
  output po257;
  output po027;
  output po179;
  output po137;
  output po140;
  output po218;
  output po141;
  output po109;
  output po151;
  output po210;
  output po105;
  output po235;
  output po264;
  output po268;
  output po043;
  output po114;
  output po190;
  output po072;
  output po031;
  output po201;
  output po284;
  output po082;
  output po194;
  output po246;
  output po032;
  output po019;
  output po169;
  output po158;
  output po059;
  output po244;
  output po270;
  output po039;
  output po101;
  output po222;
  output po228;
  output po129;
  output po148;
  output po089;
  output po077;
  output po001;
  output po174;
  output po095;
  output po110;
  output po293;
  output po198;
  output po052;
  output po013;
  output po185;
  output po261;
  output po069;
  output po226;
  output po283;
  output po166;
  output po170;
  output po146;
  output po147;
  output po029;
  output po217;
  output po199;
  output po044;
  output po126;
  output po237;
  output po102;
  output po292;
  output po156;
  output po057;
  output po297;
  output po260;
  output po172;
  output po145;
  output po079;
  output po238;
  output po191;
  output po182;
  output po034;
  output po125;
  output po291;
  output po067;
  output po088;
  output po197;
  output po205;
  output po132;
  output po107;
  output po076;
  output po064;
  output po111;
  output po215;
  output po134;
  output po160;
  output po080;
  output po149;
  output po104;
  output po296;
  output po130;
  output po212;
  output po128;
  output po294;
  output po123;
  output po040;
  output po038;
  output po144;
  output po285;
  output po084;
  output po265;
  output po099;
  output po211;
  output po245;

  wire not_new_n606__10;
  wire not_new_n5274_;
  wire or_not_new_n8595__not_new_n8593_;
  wire new_n1462_;
  wire not_new_n1604__8235430;
  wire not_new_n7527_;
  wire not_new_n7662__1;
  wire not_new_n1536__6;
  wire new_n6543_;
  wire new_n9836_;
  wire not_new_n1053__6782230728490;
  wire not_new_n626__1176490;
  wire not_new_n597__10;
  wire not_new_n1057__3;
  wire not_new_n3375__3;
  wire new_n9101_;
  wire not_new_n587__168070;
  wire not_new_n7988_;
  wire new_n5783_;
  wire not_new_n4169_;
  wire new_n4782_;
  wire not_new_n4764__0;
  wire not_new_n4420__0;
  wire not_new_n6810_;
  wire not_new_n606_;
  wire not_new_n647__8235430;
  wire new_n7680_;
  wire not_new_n7687_;
  wire new_n6471_;
  wire new_n8437_;
  wire not_new_n4817_;
  wire not_new_n965_;
  wire not_new_n962_;
  wire new_n2638_;
  wire not_new_n1597__168070;
  wire new_n1838_;
  wire new_n5737_;
  wire not_new_n8197_;
  wire not_new_n1596__113988951853731430;
  wire not_new_n6722_;
  wire new_n5308_;
  wire new_n5030_;
  wire new_n1355_;
  wire not_new_n5806__0;
  wire new_n3171_;
  wire not_new_n8720_;
  wire new_n1504_;
  wire new_n6559_;
  wire not_new_n7012_;
  wire not_new_n4907_;
  wire not_new_n9608_;
  wire not_new_n1067__70;
  wire not_new_n9565_;
  wire new_n10067_;
  wire not_new_n3099_;
  wire not_new_n7038_;
  wire and_new_n6362__new_n6430_;
  wire not_new_n1018__4;
  wire new_n10300_;
  wire not_new_n597__47475615099430;
  wire not_new_n594__24010;
  wire new_n1996_;
  wire not_new_n8837_;
  wire new_n8300_;
  wire new_n6168_;
  wire not_new_n4012_;
  wire new_n773_;
  wire not_new_n1233_;
  wire not_new_n4929__0;
  wire new_n9412_;
  wire not_new_n7395_;
  wire new_n3853_;
  wire new_n9050_;
  wire new_n7429_;
  wire new_n8566_;
  wire new_n4401_;
  wire not_new_n9205_;
  wire new_n8867_;
  wire not_new_n2852_;
  wire not_new_n1728__1176490;
  wire not_new_n4714_;
  wire not_po296_29286449308136415160327158440136953416342323212091034008010;
  wire not_new_n1269_;
  wire not_new_n593__3;
  wire not_new_n4559_;
  wire new_n7206_;
  wire new_n2722_;
  wire new_n8132_;
  wire new_n1158_;
  wire new_n7576_;
  wire and_new_n9879__new_n10247_;
  wire not_new_n6503_;
  wire not_new_n1602__332329305696010;
  wire not_new_n5085_;
  wire not_new_n6266_;
  wire not_new_n632__3;
  wire new_n5414_;
  wire not_new_n6484_;
  wire new_n6750_;
  wire not_new_n7215_;
  wire or_not_new_n6240__not_new_n6330_;
  wire new_n6326_;
  wire not_new_n9868__0;
  wire not_new_n5879_;
  wire and_and_new_n3804__new_n3807__new_n3813_;
  wire not_new_n638__968890104070;
  wire new_n5846_;
  wire po005;
  wire new_n693_;
  wire new_n2450_;
  wire not_new_n3008_;
  wire not_new_n5857_;
  wire not_new_n627__10;
  wire not_new_n8122_;
  wire new_n765_;
  wire not_new_n606__8235430;
  wire not_new_n9241_;
  wire not_new_n615__0;
  wire new_n6234_;
  wire not_new_n1017__5;
  wire not_new_n1422_;
  wire or_not_new_n2928__not_new_n2931_;
  wire not_new_n7641__0;
  wire not_new_n633__19773267430;
  wire not_new_n4930__0;
  wire new_n8926_;
  wire new_n3030_;
  wire new_n7634_;
  wire new_n1540_;
  wire new_n7082_;
  wire not_new_n7233_;
  wire new_n7282_;
  wire not_pi016_0;
  wire new_n5510_;
  wire not_new_n7651__1;
  wire new_n689_;
  wire new_n7034_;
  wire not_new_n5956_;
  wire not_new_n8244__0;
  wire not_pi192_0;
  wire new_n9197_;
  wire new_n9850_;
  wire new_n8349_;
  wire po078;
  wire new_n1790_;
  wire not_new_n9911_;
  wire not_new_n636__2;
  wire new_n5493_;
  wire new_n2712_;
  wire not_new_n6789_;
  wire not_new_n10144_;
  wire not_pi168_1;
  wire new_n9010_;
  wire new_n6414_;
  wire new_n4917_;
  wire not_new_n6635__5;
  wire not_new_n5046_;
  wire not_po298_0;
  wire not_new_n7086_;
  wire not_new_n3832_;
  wire new_n6933_;
  wire new_n6526_;
  wire new_n8480_;
  wire not_new_n6532__0;
  wire not_new_n4611_;
  wire and_new_n3729__new_n3726_;
  wire not_new_n637__47475615099430;
  wire not_new_n634__70;
  wire new_n3165_;
  wire new_n9933_;
  wire new_n4661_;
  wire not_new_n1061__10;
  wire new_n6635_;
  wire new_n4469_;
  wire new_n9056_;
  wire new_n10065_;
  wire not_pi128_0;
  wire not_new_n607__70;
  wire not_new_n630__47475615099430;
  wire new_n5300_;
  wire not_new_n10016__0;
  wire not_new_n9627_;
  wire new_n4424_;
  wire new_n6826_;
  wire not_new_n629__4;
  wire not_new_n3958_;
  wire not_new_n3184__968890104070;
  wire not_new_n1065__7;
  wire not_new_n8011_;
  wire not_new_n8104_;
  wire not_new_n7421__1;
  wire not_new_n1607_;
  wire not_new_n591__19773267430;
  wire new_n8947_;
  wire new_n9025_;
  wire not_new_n5515__0;
  wire not_new_n596__3;
  wire not_new_n6002__0;
  wire not_new_n6515_;
  wire new_n7139_;
  wire not_new_n5878__2;
  wire not_new_n9675_;
  wire po133;
  wire not_new_n9398__0;
  wire not_new_n5150_;
  wire new_n4838_;
  wire not_new_n1387_;
  wire not_new_n3228_;
  wire new_n7334_;
  wire new_n1646_;
  wire new_n6209_;
  wire new_n4084_;
  wire not_new_n8325_;
  wire not_new_n1601__1176490;
  wire new_n4799_;
  wire new_n5909_;
  wire not_new_n632__138412872010;
  wire not_new_n7697_;
  wire new_n9981_;
  wire not_new_n10213_;
  wire not_new_n1536__39098210485829880490;
  wire not_new_n994__8;
  wire not_new_n5597_;
  wire not_new_n7040_;
  wire new_n8503_;
  wire new_n5468_;
  wire not_new_n8022_;
  wire not_new_n1176_;
  wire new_n7412_;
  wire not_new_n633__5585458640832840070;
  wire new_n9709_;
  wire new_n8664_;
  wire not_new_n7265_;
  wire new_n5577_;
  wire not_new_n646__168070;
  wire not_new_n4127__0;
  wire new_n4234_;
  wire not_po296_302268019717750559482470516839540966128657419430;
  wire new_n9090_;
  wire not_new_n598__168070;
  wire not_new_n8951_;
  wire not_new_n9491__1;
  wire new_n5366_;
  wire new_n7657_;
  wire not_pi145_0;
  wire not_pi113_0;
  wire not_new_n6048_;
  wire new_n956_;
  wire not_new_n5266_;
  wire new_n7230_;
  wire or_not_new_n1806__not_new_n1807_;
  wire new_n1684_;
  wire not_new_n5446__0;
  wire not_new_n5898__1;
  wire new_n5832_;
  wire new_n8869_;
  wire new_n3632_;
  wire new_n7805_;
  wire not_new_n5563_;
  wire new_n959_;
  wire new_n1222_;
  wire or_or_not_new_n2964__not_new_n2967__not_new_n2966_;
  wire not_new_n9420_;
  wire not_new_n6944_;
  wire new_n2021_;
  wire not_new_n1017__7;
  wire not_new_n8501_;
  wire not_new_n1003__4;
  wire not_new_n5157_;
  wire new_n8602_;
  wire new_n9506_;
  wire new_n6333_;
  wire and_new_n2521__new_n2520_;
  wire new_n8734_;
  wire po066;
  wire not_new_n6242__2;
  wire not_new_n1591__3430;
  wire not_new_n3149_;
  wire not_new_n1003__1;
  wire new_n7833_;
  wire key_gate_22;
  wire not_new_n4725__0;
  wire not_new_n1028__70;
  wire not_new_n1071__490;
  wire po225;
  wire not_new_n9358__0;
  wire new_n9146_;
  wire not_new_n7379_;
  wire new_n4622_;
  wire new_n3385_;
  wire new_n1549_;
  wire not_new_n8118__2;
  wire not_new_n1612__3;
  wire not_po296_597682638941559493067901192655856192170251494124306816490;
  wire not_new_n775__8;
  wire new_n2838_;
  wire not_new_n6928_;
  wire not_new_n639__24010;
  wire or_not_pi269_1_not_pi260_1;
  wire not_new_n3996_;
  wire new_n8207_;
  wire not_new_n634__138412872010;
  wire not_new_n3454_;
  wire new_n8603_;
  wire new_n3998_;
  wire not_pi110_0;
  wire new_n10243_;
  wire not_new_n4549_;
  wire not_new_n589__1;
  wire not_new_n646__19773267430;
  wire new_n6924_;
  wire new_n9209_;
  wire not_new_n5991_;
  wire not_new_n9121_;
  wire not_new_n1583__1;
  wire not_new_n1537__113988951853731430;
  wire not_new_n10103__0;
  wire new_n8331_;
  wire not_new_n8162__0;
  wire new_n1740_;
  wire not_new_n2913_;
  wire not_new_n1235_;
  wire not_new_n587__10;
  wire new_n2506_;
  wire not_pi046_1;
  wire not_new_n2655_;
  wire new_n6249_;
  wire or_not_new_n3088__not_new_n3087_;
  wire new_n1731_;
  wire not_new_n6152_;
  wire not_new_n1037__403536070;
  wire not_pi028;
  wire not_new_n5890__1;
  wire or_not_pi064_5585458640832840070_not_new_n4019__0;
  wire new_n7201_;
  wire not_new_n1560_;
  wire or_or_not_new_n1255__not_new_n1253__not_new_n1907_;
  wire not_new_n10214_;
  wire new_n10018_;
  wire new_n2064_;
  wire new_n9151_;
  wire not_pi120_0;
  wire not_new_n6818_;
  wire not_new_n10321_;
  wire not_new_n5413_;
  wire not_new_n7219_;
  wire and_and_new_n3768__new_n3771__new_n3777_;
  wire new_n9210_;
  wire or_or_not_new_n1554__not_new_n2429__not_new_n1377_;
  wire new_n5693_;
  wire not_new_n6686_;
  wire new_n2801_;
  wire not_new_n5517__0;
  wire new_n7346_;
  wire not_pi115;
  wire new_n3886_;
  wire new_n6558_;
  wire new_n3225_;
  wire not_new_n6890_;
  wire not_new_n7903_;
  wire new_n6281_;
  wire not_new_n1045__39098210485829880490;
  wire not_new_n9512_;
  wire new_n2208_;
  wire not_new_n7258_;
  wire not_new_n7755__0;
  wire new_n8269_;
  wire new_n5009_;
  wire not_new_n6568_;
  wire not_new_n8886__0;
  wire not_new_n611__138412872010;
  wire new_n9185_;
  wire new_n7701_;
  wire not_new_n3435_;
  wire not_new_n605__0;
  wire not_new_n3227_;
  wire new_n3233_;
  wire not_new_n5878_;
  wire not_new_n1372_;
  wire not_new_n4014__3;
  wire new_n6429_;
  wire not_new_n9497_;
  wire not_new_n7924_;
  wire not_new_n1361_;
  wire not_new_n7921_;
  wire not_new_n581__17984650426474121466202803405696493492512490;
  wire not_new_n5812__0;
  wire or_not_new_n4831__not_new_n4789_;
  wire po073;
  wire not_new_n8812_;
  wire or_not_new_n2831__not_new_n1481_;
  wire not_new_n6443__8235430;
  wire new_n7561_;
  wire new_n7519_;
  wire new_n6888_;
  wire not_new_n617__1915812313805664144010;
  wire new_n3035_;
  wire new_n1533_;
  wire not_new_n5721_;
  wire new_n6844_;
  wire and_new_n3085__new_n998_;
  wire not_new_n6617__1;
  wire new_n4142_;
  wire not_po296_16284135979104490;
  wire not_new_n1601__2326305139872070;
  wire or_or_not_new_n1327__not_new_n1325__not_new_n2249_;
  wire new_n1028_;
  wire not_new_n1591__490;
  wire not_new_n1574_;
  wire new_n2392_;
  wire not_new_n4959_;
  wire new_n5700_;
  wire not_new_n1829_;
  wire not_new_n6233__2;
  wire new_n7834_;
  wire not_new_n9425__0;
  wire not_new_n4384_;
  wire not_new_n1607__403536070;
  wire new_n7395_;
  wire new_n2699_;
  wire not_new_n2345_;
  wire not_new_n1631__9;
  wire new_n611_;
  wire not_new_n10038_;
  wire not_new_n7562_;
  wire not_new_n5439__0;
  wire new_n5793_;
  wire not_pi093;
  wire not_pi151_0;
  wire new_n4827_;
  wire not_new_n6821_;
  wire not_new_n3782_;
  wire not_new_n7015_;
  wire not_new_n9427__1;
  wire not_new_n7605_;
  wire new_n7213_;
  wire not_new_n8582_;
  wire new_n9719_;
  wire new_n3085_;
  wire not_new_n593__1;
  wire not_new_n1051__5;
  wire not_new_n8772_;
  wire new_n8287_;
  wire not_new_n7643__0;
  wire not_new_n1728__7;
  wire not_new_n4752_;
  wire not_pi064_6782230728490;
  wire new_n8717_;
  wire new_n3693_;
  wire not_new_n5440__1;
  wire not_new_n4419_;
  wire not_new_n7811_;
  wire not_pi155;
  wire not_new_n4135__2;
  wire not_new_n1606__7;
  wire new_n606_;
  wire new_n6731_;
  wire new_n3829_;
  wire not_new_n6473__0;
  wire new_n6705_;
  wire not_new_n8272_;
  wire not_new_n8227_;
  wire or_not_new_n6343__not_new_n6344_;
  wire new_n4381_;
  wire new_n9830_;
  wire not_new_n4267_;
  wire not_new_n3164_;
  wire new_n8125_;
  wire not_new_n7812_;
  wire not_new_n6990__0;
  wire not_new_n9186_;
  wire new_n8367_;
  wire not_new_n2017_;
  wire new_n4613_;
  wire new_n1636_;
  wire not_new_n607__168070;
  wire new_n3076_;
  wire new_n5415_;
  wire not_new_n1534__70;
  wire new_n8299_;
  wire not_new_n1588__9;
  wire new_n5735_;
  wire not_po296_47475615099430;
  wire not_new_n4750_;
  wire not_new_n9998_;
  wire new_n7778_;
  wire not_new_n643__0;
  wire new_n3218_;
  wire new_n3125_;
  wire not_new_n1654_;
  wire new_n7443_;
  wire or_not_new_n6160__not_new_n6161_;
  wire new_n4110_;
  wire new_n7035_;
  wire new_n8974_;
  wire new_n1243_;
  wire not_new_n589__63668057609090279857414351392240010;
  wire new_n6643_;
  wire not_new_n4234_;
  wire or_not_new_n1287__not_new_n1285_;
  wire not_pi058_0;
  wire not_new_n6637_;
  wire not_new_n625__6;
  wire new_n6368_;
  wire new_n2380_;
  wire new_n7070_;
  wire not_new_n4954_;
  wire new_n4065_;
  wire new_n4676_;
  wire not_pi035_3;
  wire not_new_n7088_;
  wire new_n690_;
  wire not_pi171;
  wire not_new_n595__10;
  wire new_n6866_;
  wire new_n742_;
  wire not_new_n1371_;
  wire new_n6608_;
  wire new_n8674_;
  wire not_new_n1049__16284135979104490;
  wire not_new_n3219_;
  wire not_new_n1596__9;
  wire new_n7047_;
  wire new_n4853_;
  wire new_n8914_;
  wire new_n8004_;
  wire new_n3563_;
  wire new_n4373_;
  wire new_n5913_;
  wire not_new_n5457__0;
  wire new_n3850_;
  wire new_n8671_;
  wire new_n9586_;
  wire new_n6610_;
  wire not_new_n635__2824752490;
  wire not_new_n3322_;
  wire new_n3154_;
  wire not_new_n4956__0;
  wire or_or_or_not_new_n8528__not_new_n8429__not_new_n8457__not_new_n8458_;
  wire new_n5747_;
  wire not_new_n7859_;
  wire new_n7045_;
  wire not_new_n7603__0;
  wire new_n8930_;
  wire new_n4709_;
  wire or_not_new_n2865__not_new_n2868_;
  wire not_new_n6250_;
  wire not_new_n1576__2326305139872070;
  wire po244;
  wire not_new_n9750_;
  wire not_new_n5719_;
  wire not_new_n638__168070;
  wire new_n6270_;
  wire new_n1030_;
  wire not_new_n1729_;
  wire not_new_n989__490;
  wire not_new_n6345_;
  wire not_new_n4139_;
  wire not_new_n7643__2;
  wire key_gate_34;
  wire not_new_n9176_;
  wire key_gate_53;
  wire or_or_or_not_new_n2803__not_new_n2806__not_new_n2805__not_new_n2807_;
  wire not_new_n9915__0;
  wire new_n8765_;
  wire not_new_n4269_;
  wire new_n6561_;
  wire not_new_n604__968890104070;
  wire not_new_n8942_;
  wire not_new_n6036_;
  wire not_new_n587__5;
  wire not_new_n736__0;
  wire new_n3143_;
  wire not_new_n1571_;
  wire not_new_n4545_;
  wire not_new_n7134_;
  wire not_new_n3764_;
  wire not_new_n6782_;
  wire new_n2890_;
  wire not_new_n581__1299348114471230201171721456984490;
  wire new_n5614_;
  wire not_new_n2339_;
  wire not_new_n4798_;
  wire not_new_n7011__0;
  wire not_new_n2434_;
  wire not_new_n10178_;
  wire new_n10215_;
  wire po046;
  wire not_new_n1492_;
  wire new_n4505_;
  wire new_n9792_;
  wire not_new_n3257_;
  wire new_n5304_;
  wire or_not_new_n7664__0_not_new_n618__6782230728490;
  wire not_new_n757_;
  wire not_new_n3208_;
  wire new_n4260_;
  wire not_new_n8111__0;
  wire not_new_n5560_;
  wire new_n8965_;
  wire not_new_n5598_;
  wire new_n9525_;
  wire not_new_n8982__0;
  wire not_new_n5630__0;
  wire not_new_n1601__39098210485829880490;
  wire not_new_n6468_;
  wire new_n7693_;
  wire new_n4185_;
  wire new_n9127_;
  wire new_n2593_;
  wire not_new_n5528_;
  wire not_pi005_0;
  wire new_n1218_;
  wire not_new_n5900__0;
  wire new_n5148_;
  wire new_n8754_;
  wire not_pi274_1;
  wire new_n10280_;
  wire new_n2901_;
  wire new_n10275_;
  wire new_n4751_;
  wire new_n2668_;
  wire not_new_n617__5585458640832840070;
  wire or_not_new_n9469__not_new_n9339_;
  wire new_n5770_;
  wire and_and_new_n1953__new_n1956__new_n1954_;
  wire not_new_n8547_;
  wire not_new_n1041__168070;
  wire not_new_n7711_;
  wire not_new_n2533_;
  wire new_n4138_;
  wire not_new_n7451__0;
  wire new_n2385_;
  wire new_n4781_;
  wire not_new_n5768_;
  wire new_n2176_;
  wire new_n1644_;
  wire new_n8743_;
  wire new_n2670_;
  wire new_n3008_;
  wire new_n5206_;
  wire new_n9984_;
  wire new_n2698_;
  wire not_new_n9412__1;
  wire not_new_n10035_;
  wire new_n3627_;
  wire new_n9935_;
  wire new_n4785_;
  wire new_n9814_;
  wire new_n4366_;
  wire new_n1713_;
  wire not_pi142_3;
  wire new_n2375_;
  wire not_new_n6927_;
  wire not_new_n1631__138412872010;
  wire not_new_n3916_;
  wire not_new_n9291_;
  wire not_new_n10045__0;
  wire not_new_n624__19773267430;
  wire not_new_n3501_;
  wire new_n1474_;
  wire not_new_n8160_;
  wire not_new_n3277_;
  wire not_new_n2606_;
  wire new_n1380_;
  wire not_new_n2229_;
  wire not_new_n9541_;
  wire new_n2571_;
  wire not_new_n6991__0;
  wire not_new_n4313_;
  wire not_new_n9166_;
  wire not_new_n8527_;
  wire not_new_n7418_;
  wire new_n1874_;
  wire new_n4512_;
  wire not_new_n1035__10;
  wire not_new_n6546_;
  wire new_n4791_;
  wire not_new_n2819_;
  wire not_new_n601__8235430;
  wire not_new_n600__3;
  wire not_new_n9356_;
  wire new_n5769_;
  wire not_new_n2039_;
  wire not_new_n5700_;
  wire new_n7958_;
  wire new_n3741_;
  wire not_new_n9953__0;
  wire not_new_n1043__490;
  wire new_n3894_;
  wire not_new_n645__968890104070;
  wire or_not_new_n2946__not_new_n2949_;
  wire new_n7506_;
  wire new_n8443_;
  wire not_pi075;
  wire not_new_n1613__2824752490;
  wire not_new_n641__3430;
  wire new_n3695_;
  wire new_n4081_;
  wire not_new_n3961_;
  wire not_new_n1366_;
  wire not_pi064_113988951853731430;
  wire not_new_n2047_;
  wire not_new_n1603__8;
  wire new_n8325_;
  wire not_new_n1059__332329305696010;
  wire new_n10169_;
  wire not_new_n594__10;
  wire not_new_n634__168070;
  wire and_new_n1053__new_n6232_;
  wire new_n6235_;
  wire not_new_n625__273687473400809163430;
  wire new_n644_;
  wire new_n5809_;
  wire new_n2160_;
  wire new_n2811_;
  wire not_new_n6113_;
  wire new_n2501_;
  wire new_n7271_;
  wire not_new_n6490__0;
  wire new_n7423_;
  wire not_new_n4728__0;
  wire new_n6232_;
  wire not_new_n6941_;
  wire new_n6779_;
  wire new_n2979_;
  wire new_n6112_;
  wire not_new_n4993_;
  wire new_n1409_;
  wire not_new_n1049__2824752490;
  wire not_new_n678_;
  wire new_n2864_;
  wire not_new_n8267__0;
  wire not_new_n7927_;
  wire not_new_n9272_;
  wire po197;
  wire new_n4702_;
  wire not_new_n3363_;
  wire not_new_n8315_;
  wire not_new_n1598__332329305696010;
  wire not_new_n1589__1176490;
  wire not_new_n598__6782230728490;
  wire not_new_n7461_;
  wire new_n2074_;
  wire not_new_n3310__8;
  wire not_new_n5415_;
  wire new_n9875_;
  wire not_new_n7393_;
  wire new_n7315_;
  wire new_n9088_;
  wire new_n4317_;
  wire not_new_n8973_;
  wire new_n989_;
  wire new_n7375_;
  wire new_n5831_;
  wire not_new_n603__968890104070;
  wire not_new_n1061__1176490;
  wire not_new_n3550_;
  wire new_n3390_;
  wire not_new_n2132_;
  wire not_new_n9473_;
  wire new_n2086_;
  wire not_new_n4986_;
  wire not_new_n10160_;
  wire not_new_n7122_;
  wire not_new_n1728__490;
  wire not_new_n6234__0;
  wire not_new_n628__3;
  wire not_new_n4730_;
  wire not_new_n640__403536070;
  wire not_new_n1055__797922662976120010;
  wire not_new_n5292_;
  wire new_n7228_;
  wire new_n3209_;
  wire and_new_n7791__new_n7786_;
  wire not_new_n4387_;
  wire not_new_n8809_;
  wire not_new_n10153_;
  wire not_new_n648__6;
  wire or_not_new_n2944__not_new_n2943_;
  wire not_new_n5481_;
  wire not_new_n7014__2;
  wire not_new_n1602__7;
  wire not_new_n4248_;
  wire not_new_n8265_;
  wire not_new_n1051__6782230728490;
  wire new_n4966_;
  wire not_new_n8526_;
  wire and_and_new_n1896__new_n1899__new_n1897_;
  wire new_n7441_;
  wire new_n619_;
  wire new_n9260_;
  wire not_new_n1057__4;
  wire and_new_n1539__new_n2356_;
  wire and_new_n8837__new_n9203_;
  wire new_n6518_;
  wire not_new_n3811_;
  wire not_new_n1601__2824752490;
  wire po273;
  wire not_new_n5740_;
  wire not_new_n9376__0;
  wire not_pi275_1;
  wire not_new_n7477_;
  wire new_n6181_;
  wire not_new_n605__4;
  wire not_new_n6558_;
  wire new_n5454_;
  wire new_n5326_;
  wire new_n1051_;
  wire not_new_n3205_;
  wire not_new_n1596__24010;
  wire new_n4321_;
  wire not_new_n612_;
  wire new_n8924_;
  wire new_n8764_;
  wire new_n10334_;
  wire new_n1496_;
  wire not_new_n734_;
  wire new_n9254_;
  wire new_n2485_;
  wire new_n2797_;
  wire not_new_n639__5;
  wire new_n7556_;
  wire not_new_n4756__0;
  wire not_new_n10058_;
  wire not_new_n1018__1;
  wire not_new_n5082__0;
  wire new_n4713_;
  wire po067;
  wire not_new_n4304_;
  wire not_new_n4115__2;
  wire new_n10295_;
  wire not_new_n3311__3430;
  wire not_pi255_1;
  wire not_new_n9057_;
  wire not_new_n6023_;
  wire not_new_n1061__24010;
  wire new_n2695_;
  wire not_new_n937_;
  wire new_n8361_;
  wire not_new_n931_;
  wire new_n7225_;
  wire new_n7340_;
  wire not_new_n1603__3430;
  wire not_new_n7127_;
  wire new_n6793_;
  wire new_n3822_;
  wire new_n2568_;
  wire not_new_n5870_;
  wire not_new_n1014__5;
  wire new_n6735_;
  wire not_new_n1605__3;
  wire new_n9124_;
  wire not_new_n3221_;
  wire new_n8514_;
  wire new_n7099_;
  wire not_new_n1534__968890104070;
  wire key_gate_94;
  wire not_new_n6516_;
  wire new_n4188_;
  wire new_n1379_;
  wire new_n3122_;
  wire not_new_n2924_;
  wire not_new_n2834_;
  wire new_n7852_;
  wire not_new_n7109__0;
  wire or_or_not_new_n2973__not_new_n2976__not_new_n2975_;
  wire new_n1313_;
  wire new_n7814_;
  wire not_new_n7582_;
  wire not_new_n9921_;
  wire not_new_n9035_;
  wire not_new_n7731_;
  wire not_new_n3258_;
  wire new_n4759_;
  wire not_new_n7030_;
  wire new_n2823_;
  wire not_new_n2882_;
  wire not_new_n6136_;
  wire not_new_n9354_;
  wire not_new_n9879__0;
  wire not_new_n1005__3;
  wire and_new_n3016__new_n998_;
  wire not_new_n770_;
  wire not_new_n4737__0;
  wire not_new_n7501_;
  wire not_new_n1154__0;
  wire new_n8274_;
  wire not_new_n7155_;
  wire not_new_n1013_;
  wire new_n709_;
  wire new_n2907_;
  wire not_new_n4679_;
  wire new_n6057_;
  wire not_new_n1588__6;
  wire not_pi038_3;
  wire new_n2345_;
  wire not_new_n1184_;
  wire not_new_n7278_;
  wire not_new_n3447_;
  wire not_new_n6520__0;
  wire not_new_n1020__2;
  wire not_new_n5847_;
  wire po293;
  wire not_new_n3242_;
  wire new_n3697_;
  wire not_new_n1616__57648010;
  wire new_n1173_;
  wire new_n7019_;
  wire not_new_n3142_;
  wire not_new_n6281_;
  wire new_n761_;
  wire not_new_n3693_;
  wire not_new_n4422_;
  wire new_n7580_;
  wire new_n8676_;
  wire not_new_n3223_;
  wire not_new_n593__0;
  wire not_new_n5727_;
  wire new_n8204_;
  wire new_n8719_;
  wire not_new_n8539_;
  wire not_new_n9530__0;
  wire and_new_n1735__new_n1736_;
  wire not_new_n9208_;
  wire new_n2508_;
  wire not_new_n3330_;
  wire not_new_n775__16284135979104490;
  wire not_new_n8679_;
  wire new_n9427_;
  wire new_n9681_;
  wire not_new_n648__6782230728490;
  wire not_new_n9971_;
  wire new_n1426_;
  wire not_new_n584_;
  wire not_pi272;
  wire not_new_n632__47475615099430;
  wire not_new_n2884_;
  wire new_n3743_;
  wire or_not_new_n618__2326305139872070_not_new_n8496_;
  wire new_n7220_;
  wire new_n9692_;
  wire new_n2614_;
  wire new_n10259_;
  wire not_new_n3293_;
  wire not_new_n2302_;
  wire not_new_n5836_;
  wire not_new_n4508__0;
  wire not_new_n4187_;
  wire not_new_n4119__2;
  wire new_n3266_;
  wire new_n4156_;
  wire not_new_n1810_;
  wire not_new_n581__39098210485829880490;
  wire not_new_n2151_;
  wire new_n6349_;
  wire not_new_n7710_;
  wire not_new_n2350_;
  wire new_n2349_;
  wire not_new_n1588__10;
  wire not_new_n3372__6;
  wire new_n3664_;
  wire not_new_n3127_;
  wire new_n8079_;
  wire new_n5341_;
  wire not_new_n645__2326305139872070;
  wire new_n8827_;
  wire new_n942_;
  wire not_new_n1057__5;
  wire not_new_n589__5;
  wire not_new_n2720_;
  wire not_new_n8157__0;
  wire not_new_n1599_;
  wire not_new_n1594__1;
  wire not_new_n3355_;
  wire not_new_n4759_;
  wire not_new_n4140_;
  wire or_or_or_not_new_n2749__not_new_n2752__not_new_n2751__not_new_n2753_;
  wire not_new_n4746_;
  wire not_new_n5761__0;
  wire not_pi251_1;
  wire not_new_n3493_;
  wire not_new_n4763_;
  wire not_new_n4250_;
  wire and_new_n9402__new_n9804_;
  wire not_new_n611__2;
  wire not_new_n1588__24010;
  wire not_pi143_3;
  wire not_new_n7914_;
  wire not_new_n9961__0;
  wire key_gate_0;
  wire new_n3355_;
  wire new_n7525_;
  wire new_n8127_;
  wire not_new_n9317_;
  wire not_new_n3224_;
  wire not_pi168_3;
  wire not_new_n1981_;
  wire and_new_n1896__new_n1899_;
  wire new_n3031_;
  wire new_n5494_;
  wire new_n1204_;
  wire not_new_n1588__5585458640832840070;
  wire new_n3616_;
  wire new_n698_;
  wire new_n2461_;
  wire not_new_n6987_;
  wire not_pi023_0;
  wire new_n987_;
  wire or_or_not_new_n2246__not_new_n2243__not_new_n2244_;
  wire new_n6552_;
  wire not_new_n1027__1915812313805664144010;
  wire new_n6203_;
  wire not_new_n7491_;
  wire new_n2327_;
  wire not_new_n2266_;
  wire new_n9954_;
  wire not_new_n7012__0;
  wire not_new_n4458_;
  wire not_new_n8831_;
  wire not_new_n588__1;
  wire new_n7652_;
  wire not_new_n3707_;
  wire not_new_n630_;
  wire or_not_new_n1405__not_new_n616_;
  wire not_new_n1591__6;
  wire not_new_n984__7;
  wire not_new_n624__6;
  wire not_new_n4173_;
  wire new_n4833_;
  wire not_new_n3996__0;
  wire not_new_n1536__19773267430;
  wire not_new_n643__10;
  wire new_n6073_;
  wire new_n8340_;
  wire not_new_n5465_;
  wire not_pi111;
  wire not_new_n1611__968890104070;
  wire new_n2909_;
  wire po004;
  wire not_new_n5942__0;
  wire not_new_n2509__4;
  wire not_new_n6072_;
  wire new_n8893_;
  wire not_po296_403536070;
  wire not_new_n9340_;
  wire not_new_n3139_;
  wire not_new_n639__3;
  wire new_n4773_;
  wire new_n7104_;
  wire or_or_or_not_new_n2865__not_new_n2868__not_new_n2867__not_new_n2869_;
  wire not_new_n681_;
  wire not_new_n632__797922662976120010;
  wire not_new_n6207_;
  wire not_new_n3716_;
  wire not_new_n10097_;
  wire new_n8552_;
  wire not_new_n5759__0;
  wire new_n8233_;
  wire not_new_n9387_;
  wire new_n8841_;
  wire not_new_n8294__0;
  wire po072;
  wire new_n3382_;
  wire not_new_n4404_;
  wire not_new_n613__6;
  wire not_new_n1601__332329305696010;
  wire new_n3022_;
  wire not_new_n9389_;
  wire not_new_n3751_;
  wire new_n4665_;
  wire not_new_n8103_;
  wire new_n5014_;
  wire not_new_n5190_;
  wire not_pi222;
  wire not_new_n1169_;
  wire new_n9218_;
  wire new_n3587_;
  wire not_new_n6291_;
  wire new_n1878_;
  wire not_new_n7354__0;
  wire not_new_n3372__8;
  wire new_n7573_;
  wire not_new_n1065__5585458640832840070;
  wire not_pi177_1;
  wire not_new_n7520_;
  wire not_new_n1580__797922662976120010;
  wire not_new_n3233_;
  wire not_new_n9704_;
  wire new_n4712_;
  wire new_n5123_;
  wire new_n8116_;
  wire not_new_n4908_;
  wire new_n7731_;
  wire new_n7085_;
  wire not_new_n5938__0;
  wire not_po298_168070;
  wire new_n8182_;
  wire new_n2645_;
  wire new_n4748_;
  wire not_new_n7637_;
  wire not_new_n7739__0;
  wire not_new_n628__1;
  wire new_n6634_;
  wire not_new_n6539__0;
  wire new_n4663_;
  wire not_new_n7889_;
  wire not_new_n4712_;
  wire new_n6723_;
  wire new_n3123_;
  wire new_n4393_;
  wire not_new_n8683_;
  wire not_new_n9061_;
  wire not_new_n1523_;
  wire new_n10028_;
  wire not_new_n8120__0;
  wire not_new_n1027__0;
  wire new_n2730_;
  wire not_new_n8888_;
  wire not_new_n7341_;
  wire not_new_n5255_;
  wire not_new_n9364_;
  wire not_new_n5675_;
  wire not_pi033_2;
  wire not_new_n7891_;
  wire not_new_n10304_;
  wire not_new_n4731_;
  wire new_n3423_;
  wire not_pi212;
  wire key_gate_37;
  wire new_n4550_;
  wire new_n4624_;
  wire not_new_n9869_;
  wire not_pi045_0;
  wire new_n8314_;
  wire not_new_n8542_;
  wire not_new_n10238_;
  wire not_new_n1584__9;
  wire not_new_n7463_;
  wire not_new_n9522_;
  wire new_n6537_;
  wire new_n1314_;
  wire not_new_n4560_;
  wire not_new_n994__9;
  wire new_n8715_;
  wire not_new_n4266_;
  wire not_new_n4876_;
  wire not_new_n605__7;
  wire not_new_n9156_;
  wire not_new_n1613__47475615099430;
  wire new_n10177_;
  wire new_n4159_;
  wire not_new_n6656_;
  wire not_new_n4149_;
  wire or_not_new_n2785__not_new_n2788_;
  wire new_n5697_;
  wire not_new_n7054_;
  wire not_new_n5763__1;
  wire new_n9567_;
  wire not_new_n7848_;
  wire new_n6391_;
  wire new_n1624_;
  wire new_n4017_;
  wire new_n3164_;
  wire not_new_n7324_;
  wire new_n2478_;
  wire new_n7706_;
  wire not_new_n1845_;
  wire and_new_n2687__new_n2688_;
  wire not_new_n6889_;
  wire not_new_n4830_;
  wire new_n4038_;
  wire new_n8551_;
  wire not_new_n7791__0;
  wire new_n1712_;
  wire and_new_n8731__new_n8730_;
  wire not_new_n1292_;
  wire not_new_n596__138412872010;
  wire or_not_new_n1571__not_new_n2504_;
  wire not_new_n3885_;
  wire not_new_n591__4;
  wire not_new_n605__57648010;
  wire not_pi039_1;
  wire new_n1777_;
  wire not_new_n5867_;
  wire not_new_n627__3;
  wire not_new_n10236_;
  wire new_n1480_;
  wire not_new_n3673_;
  wire not_new_n7061_;
  wire or_or_not_new_n1844__not_new_n1845__not_new_n1847_;
  wire new_n9841_;
  wire new_n2025_;
  wire not_new_n6073_;
  wire not_po296_1176490;
  wire new_n6762_;
  wire new_n2757_;
  wire new_n7719_;
  wire new_n7151_;
  wire not_new_n3871_;
  wire not_new_n3987__0;
  wire not_new_n3719_;
  wire not_new_n590_;
  wire new_n10327_;
  wire not_new_n605__8235430;
  wire not_new_n1596__968890104070;
  wire new_n3352_;
  wire and_new_n9356__new_n9738_;
  wire not_new_n4903_;
  wire new_n5860_;
  wire new_n7700_;
  wire new_n7621_;
  wire not_new_n1035__2;
  wire not_new_n8844__0;
  wire not_new_n6974__2824752490;
  wire new_n6100_;
  wire not_new_n1164_;
  wire not_new_n8785_;
  wire not_new_n582__0;
  wire not_new_n1158__0;
  wire not_new_n645__3;
  wire new_n6068_;
  wire not_new_n7628_;
  wire new_n8675_;
  wire new_n9929_;
  wire new_n7140_;
  wire new_n8677_;
  wire not_new_n7431_;
  wire not_pi178;
  wire new_n9494_;
  wire new_n7036_;
  wire not_new_n1059__16284135979104490;
  wire not_new_n6373__8;
  wire new_n3450_;
  wire not_new_n7426_;
  wire not_new_n1602__2326305139872070;
  wire not_new_n5821_;
  wire not_new_n607__7;
  wire new_n6672_;
  wire not_new_n7985_;
  wire new_n5678_;
  wire new_n6217_;
  wire new_n2454_;
  wire not_new_n3184__0;
  wire new_n5800_;
  wire not_pi179_0;
  wire not_new_n1812_;
  wire not_pi162_2;
  wire new_n4333_;
  wire new_n9801_;
  wire not_new_n9372_;
  wire new_n3720_;
  wire not_new_n9426_;
  wire new_n6947_;
  wire new_n9539_;
  wire not_new_n610__1;
  wire not_new_n1555_;
  wire new_n10286_;
  wire not_new_n2444_;
  wire not_new_n1057__968890104070;
  wire not_new_n7579_;
  wire not_new_n8118__0;
  wire not_new_n7123_;
  wire not_new_n5170_;
  wire not_new_n1061__8;
  wire new_n732_;
  wire not_new_n748_;
  wire new_n1172_;
  wire not_new_n596__797922662976120010;
  wire not_new_n7389_;
  wire not_new_n1604__2326305139872070;
  wire not_new_n9992_;
  wire not_new_n6227_;
  wire not_new_n637__16284135979104490;
  wire or_not_new_n1567__not_new_n2494_;
  wire not_new_n629__19773267430;
  wire new_n6392_;
  wire not_pi053_0;
  wire or_or_or_not_new_n1055__168070_not_new_n6325__not_new_n6373__1_not_new_n6317_;
  wire new_n7997_;
  wire new_n6727_;
  wire new_n4074_;
  wire new_n1369_;
  wire new_n1494_;
  wire not_new_n7279_;
  wire not_new_n9868_;
  wire new_n6534_;
  wire not_new_n6960_;
  wire not_new_n3122_;
  wire not_pi257_0;
  wire new_n7238_;
  wire new_n9752_;
  wire not_new_n625__8235430;
  wire not_new_n6461_;
  wire not_new_n8130__0;
  wire new_n9429_;
  wire not_pi167_0;
  wire new_n8466_;
  wire not_new_n1887_;
  wire not_new_n1616__2;
  wire not_new_n640__4;
  wire not_new_n5022_;
  wire not_new_n5360_;
  wire new_n10342_;
  wire not_new_n2321_;
  wire not_new_n7430__0;
  wire not_new_n589__113988951853731430;
  wire new_n4060_;
  wire not_new_n597__9;
  wire new_n5898_;
  wire new_n4360_;
  wire new_n2004_;
  wire not_new_n618__113988951853731430;
  wire not_new_n7714_;
  wire new_n5648_;
  wire not_new_n6232__1;
  wire key_gate_124;
  wire not_new_n1053__24010;
  wire new_n3611_;
  wire not_new_n1065__4;
  wire not_new_n730__1;
  wire new_n4275_;
  wire new_n1916_;
  wire new_n8358_;
  wire new_n3455_;
  wire not_new_n7984_;
  wire not_new_n5349_;
  wire not_new_n1604__2;
  wire not_new_n3341_;
  wire not_new_n9327_;
  wire new_n1228_;
  wire not_new_n2574_;
  wire not_new_n1014__2;
  wire not_new_n1028__8;
  wire not_new_n1061__490;
  wire not_new_n1589__6;
  wire not_new_n9881_;
  wire new_n5053_;
  wire po149;
  wire not_pi051_2;
  wire not_new_n634__2326305139872070;
  wire not_new_n1597__57648010;
  wire not_new_n1588__168070;
  wire po084;
  wire not_new_n8950_;
  wire not_new_n635__2326305139872070;
  wire not_new_n1049__8235430;
  wire new_n6885_;
  wire new_n9695_;
  wire not_new_n4567_;
  wire not_new_n5755__0;
  wire not_new_n629__3;
  wire not_new_n5758_;
  wire new_n7916_;
  wire not_new_n7846_;
  wire new_n1986_;
  wire not_new_n3088_;
  wire not_new_n644__9;
  wire new_n9839_;
  wire not_new_n8935_;
  wire not_new_n3522_;
  wire new_n2111_;
  wire new_n2863_;
  wire not_new_n5549_;
  wire not_new_n1728__2;
  wire new_n8243_;
  wire not_new_n8533_;
  wire not_new_n626__16284135979104490;
  wire not_new_n610__9;
  wire new_n8220_;
  wire new_n2893_;
  wire not_pi179_1;
  wire not_new_n8616_;
  wire not_new_n3773_;
  wire new_n6666_;
  wire not_new_n6823_;
  wire new_n4794_;
  wire not_new_n6998__0;
  wire not_new_n616__0;
  wire not_new_n6974_;
  wire new_n3550_;
  wire and_new_n2652__new_n2651_;
  wire new_n3734_;
  wire new_n9069_;
  wire new_n4667_;
  wire not_new_n3419_;
  wire not_new_n9922_;
  wire not_new_n621__168070;
  wire new_n7769_;
  wire not_new_n6334_;
  wire not_new_n3588_;
  wire new_n1235_;
  wire not_new_n5201_;
  wire not_new_n3156_;
  wire new_n3006_;
  wire not_new_n5476__0;
  wire not_new_n7070_;
  wire not_new_n4968_;
  wire not_new_n3015_;
  wire new_n2159_;
  wire not_new_n8359_;
  wire not_new_n9180_;
  wire not_new_n633__1;
  wire and_and_new_n1746__new_n1747__new_n1749_;
  wire not_new_n6443__3;
  wire not_new_n1039__797922662976120010;
  wire new_n6811_;
  wire or_or_not_new_n1565__not_new_n2484__not_new_n1399_;
  wire new_n3833_;
  wire not_new_n8968_;
  wire not_new_n8988_;
  wire not_new_n589__21838143759917965991093122527538323430;
  wire not_new_n10106_;
  wire new_n10217_;
  wire new_n8877_;
  wire not_new_n1180_;
  wire not_new_n6975__0;
  wire not_new_n3431_;
  wire new_n1502_;
  wire not_new_n591__24010;
  wire new_n6784_;
  wire not_new_n1594__3;
  wire not_new_n2033_;
  wire and_new_n1246__new_n1875_;
  wire not_new_n3343_;
  wire not_new_n586__2;
  wire not_new_n1041_;
  wire not_new_n9822_;
  wire not_new_n8244_;
  wire not_new_n8741_;
  wire not_new_n3513_;
  wire not_new_n8956_;
  wire not_new_n4421_;
  wire new_n8830_;
  wire new_n8842_;
  wire not_new_n5158_;
  wire new_n2612_;
  wire new_n7795_;
  wire not_new_n9330_;
  wire not_new_n5187_;
  wire not_new_n1015__6;
  wire not_new_n3714_;
  wire not_new_n604__57648010;
  wire not_new_n7753__2;
  wire not_new_n1489_;
  wire not_new_n683_;
  wire not_new_n4833__1;
  wire not_pi041_3;
  wire not_new_n4765_;
  wire not_new_n3842_;
  wire not_new_n6624_;
  wire not_new_n8849__0;
  wire not_new_n985_;
  wire not_pi033_3;
  wire not_new_n1609__0;
  wire not_new_n1047__0;
  wire not_new_n9376_;
  wire new_n9537_;
  wire new_n8713_;
  wire new_n1846_;
  wire not_new_n6138__0;
  wire not_new_n8358_;
  wire new_n2549_;
  wire not_new_n7084_;
  wire and_new_n9365__new_n9731_;
  wire new_n2726_;
  wire not_new_n713_;
  wire not_new_n4958_;
  wire not_new_n1152__0;
  wire not_new_n1039__4;
  wire not_new_n645__16284135979104490;
  wire new_n6482_;
  wire new_n6023_;
  wire not_new_n3372__1176490;
  wire new_n9825_;
  wire not_new_n6373__5;
  wire not_new_n1027__8;
  wire not_new_n9891_;
  wire new_n3045_;
  wire new_n1195_;
  wire not_new_n3185__57648010;
  wire not_new_n6985__1;
  wire not_new_n1175__1;
  wire not_pi163_1;
  wire not_new_n3315__168070;
  wire not_new_n1660_;
  wire new_n9443_;
  wire new_n3577_;
  wire not_new_n5421_;
  wire new_n6037_;
  wire new_n7783_;
  wire not_pi260;
  wire and_and_new_n6326__new_n6241__new_n6227_;
  wire not_pi246_1;
  wire not_new_n1598__0;
  wire not_new_n10256_;
  wire new_n3176_;
  wire not_new_n7260__0;
  wire new_n9641_;
  wire new_n1322_;
  wire new_n7756_;
  wire not_new_n5923_;
  wire not_new_n630__0;
  wire not_new_n1071__403536070;
  wire new_n5241_;
  wire not_new_n4539_;
  wire not_new_n8155__0;
  wire new_n8750_;
  wire new_n5583_;
  wire new_n9504_;
  wire not_new_n9288_;
  wire not_pi042_1;
  wire not_new_n9409_;
  wire not_new_n1449_;
  wire not_new_n9762_;
  wire not_new_n1601__4;
  wire not_new_n601__57648010;
  wire new_n8601_;
  wire new_n2268_;
  wire new_n6169_;
  wire new_n2639_;
  wire not_new_n5429_;
  wire not_new_n1337_;
  wire not_new_n3524_;
  wire not_new_n1611__403536070;
  wire new_n8453_;
  wire not_new_n647__968890104070;
  wire not_new_n7245_;
  wire not_new_n627__2326305139872070;
  wire not_new_n7087_;
  wire new_n7226_;
  wire not_new_n633__138412872010;
  wire not_new_n5488__0;
  wire not_new_n1613__797922662976120010;
  wire new_n3633_;
  wire new_n3907_;
  wire not_new_n7045__1;
  wire new_n2336_;
  wire not_new_n646__113988951853731430;
  wire new_n1650_;
  wire not_new_n1613__2;
  wire not_new_n1188_;
  wire not_pi130_0;
  wire not_new_n7309_;
  wire not_new_n8103__0;
  wire not_new_n7017__0;
  wire new_n6873_;
  wire new_n8872_;
  wire new_n5247_;
  wire not_po296_70;
  wire new_n2774_;
  wire not_new_n1059__2326305139872070;
  wire not_new_n3769_;
  wire not_new_n1588__968890104070;
  wire not_new_n994__2824752490;
  wire not_new_n10335_;
  wire not_new_n1067__403536070;
  wire new_n8268_;
  wire not_po298_6782230728490;
  wire not_new_n1602__6782230728490;
  wire not_new_n981_;
  wire not_new_n9705_;
  wire new_n4098_;
  wire new_n5408_;
  wire not_new_n8137_;
  wire not_new_n1607__490;
  wire not_new_n1576__6782230728490;
  wire new_n3565_;
  wire po026;
  wire new_n9475_;
  wire not_new_n595__8235430;
  wire not_new_n9444_;
  wire new_n8123_;
  wire new_n8246_;
  wire new_n2420_;
  wire not_new_n7357__1;
  wire new_n5829_;
  wire not_new_n9728_;
  wire po119;
  wire not_new_n5992_;
  wire not_new_n9466_;
  wire not_new_n642__6782230728490;
  wire not_pi181_0;
  wire new_n2885_;
  wire or_or_not_new_n9361__not_new_n9358__0_not_new_n9750_;
  wire not_new_n6773_;
  wire new_n4262_;
  wire not_new_n2267_;
  wire new_n5766_;
  wire new_n4090_;
  wire not_new_n7599__2;
  wire not_new_n6992__2;
  wire not_new_n1053__7;
  wire not_pi178_2;
  wire not_new_n1358_;
  wire new_n4024_;
  wire not_new_n1611__797922662976120010;
  wire new_n1225_;
  wire not_new_n1241_;
  wire not_new_n3933__0;
  wire new_n9913_;
  wire not_new_n4801__0;
  wire new_n4407_;
  wire new_n2530_;
  wire new_n6756_;
  wire not_new_n7608_;
  wire new_n3141_;
  wire not_new_n4109_;
  wire new_n7558_;
  wire not_new_n9615_;
  wire not_new_n4114_;
  wire not_new_n1588__57648010;
  wire not_new_n611__8235430;
  wire not_new_n9654_;
  wire not_new_n1237_;
  wire not_new_n4289_;
  wire not_new_n1601__6;
  wire new_n8046_;
  wire new_n9077_;
  wire not_new_n6557_;
  wire not_new_n1007__0;
  wire not_new_n3451_;
  wire new_n6993_;
  wire new_n1224_;
  wire new_n9893_;
  wire not_new_n6604_;
  wire new_n7052_;
  wire new_n3722_;
  wire new_n3790_;
  wire not_new_n1997_;
  wire new_n9283_;
  wire not_new_n630__4;
  wire new_n3472_;
  wire new_n7526_;
  wire not_new_n961_;
  wire not_new_n5264_;
  wire not_new_n7008__0;
  wire not_new_n5766__0;
  wire new_n6157_;
  wire new_n4228_;
  wire not_new_n8958_;
  wire po186;
  wire new_n9833_;
  wire po177;
  wire not_new_n4918_;
  wire new_n8879_;
  wire new_n6387_;
  wire not_new_n9933_;
  wire not_pi176_2;
  wire not_new_n4784__0;
  wire not_new_n600__8;
  wire new_n8459_;
  wire not_new_n3877_;
  wire new_n3638_;
  wire not_new_n9618_;
  wire new_n3480_;
  wire new_n5828_;
  wire not_new_n1599__8235430;
  wire new_n8335_;
  wire not_new_n5764__1;
  wire not_new_n1600__6782230728490;
  wire new_n3025_;
  wire not_new_n4319_;
  wire new_n8154_;
  wire not_new_n8899__2;
  wire not_new_n599__6;
  wire new_n9671_;
  wire new_n2154_;
  wire not_new_n1728_;
  wire new_n5528_;
  wire new_n1333_;
  wire not_new_n8674_;
  wire not_new_n623__5;
  wire not_new_n2869_;
  wire new_n4511_;
  wire not_new_n632__1;
  wire new_n5146_;
  wire new_n10073_;
  wire new_n7529_;
  wire new_n3147_;
  wire not_new_n626__70;
  wire new_n9071_;
  wire not_new_n8158__1;
  wire new_n8850_;
  wire new_n8992_;
  wire not_pi144;
  wire new_n750_;
  wire not_new_n1631__1176490;
  wire new_n7885_;
  wire not_new_n9902_;
  wire new_n3964_;
  wire new_n2494_;
  wire not_new_n4742_;
  wire not_new_n1027__168070;
  wire not_new_n9837_;
  wire not_pi216;
  wire not_new_n10244_;
  wire not_new_n742__0;
  wire new_n8419_;
  wire not_new_n1399_;
  wire not_new_n9184_;
  wire not_new_n3310__0;
  wire not_new_n638__2;
  wire not_new_n7011_;
  wire not_new_n9490_;
  wire not_pi003_0;
  wire not_new_n1536__8235430;
  wire new_n5812_;
  wire not_new_n1601_;
  wire new_n3859_;
  wire new_n8415_;
  wire not_new_n9958_;
  wire not_new_n2509__7;
  wire new_n6401_;
  wire not_new_n6778_;
  wire and_new_n4580__new_n4649_;
  wire not_new_n8909_;
  wire not_new_n6567_;
  wire not_new_n7741__0;
  wire new_n1012_;
  wire not_new_n637__5;
  wire not_new_n8240_;
  wire new_n2045_;
  wire not_new_n6472__0;
  wire not_new_n7742__0;
  wire new_n7224_;
  wire not_new_n1333_;
  wire not_new_n1053__57648010;
  wire not_new_n5359_;
  wire not_new_n1581__0;
  wire new_n9672_;
  wire new_n7760_;
  wire not_new_n2683_;
  wire not_new_n7092_;
  wire not_new_n6324_;
  wire po167;
  wire not_new_n720_;
  wire not_new_n736__2;
  wire not_new_n4308_;
  wire not_new_n4488_;
  wire not_new_n6974__6;
  wire new_n930_;
  wire not_new_n639__332329305696010;
  wire new_n1768_;
  wire new_n594_;
  wire new_n9463_;
  wire new_n8799_;
  wire not_new_n599__57648010;
  wire not_new_n5459__0;
  wire new_n5968_;
  wire not_new_n1581__968890104070;
  wire new_n7988_;
  wire not_new_n625__70;
  wire not_new_n2573_;
  wire not_new_n9204_;
  wire new_n2114_;
  wire new_n2290_;
  wire new_n1820_;
  wire not_new_n7490_;
  wire new_n9473_;
  wire not_new_n604__3430;
  wire not_new_n585__70;
  wire new_n2230_;
  wire not_new_n7535_;
  wire new_n10322_;
  wire not_new_n4297_;
  wire new_n2458_;
  wire new_n7004_;
  wire new_n6604_;
  wire new_n9682_;
  wire new_n7991_;
  wire not_new_n8033_;
  wire not_new_n2318_;
  wire new_n10216_;
  wire not_new_n594__57648010;
  wire new_n1290_;
  wire not_new_n590__2;
  wire not_new_n2499_;
  wire new_n1510_;
  wire not_new_n2077_;
  wire new_n7553_;
  wire new_n8397_;
  wire not_new_n10229_;
  wire not_new_n605__1;
  wire and_new_n4348__new_n4301_;
  wire new_n9252_;
  wire not_new_n4354_;
  wire not_new_n625__6782230728490;
  wire not_new_n7753__1;
  wire new_n3019_;
  wire not_new_n8645__0;
  wire new_n6143_;
  wire and_and_new_n3732__new_n3735__new_n3741_;
  wire not_new_n2816_;
  wire new_n10099_;
  wire not_new_n2804_;
  wire new_n3780_;
  wire not_new_n625__10;
  wire not_new_n2604_;
  wire new_n3105_;
  wire new_n9388_;
  wire new_n6119_;
  wire new_n9733_;
  wire not_new_n8250__0;
  wire not_pi141_3;
  wire new_n4828_;
  wire new_n9790_;
  wire not_pi105_0;
  wire not_new_n2019_;
  wire not_new_n4912_;
  wire new_n998_;
  wire new_n8446_;
  wire not_new_n9170_;
  wire not_new_n585__24010;
  wire not_new_n8132__0;
  wire new_n8737_;
  wire not_new_n1283_;
  wire not_new_n587_;
  wire not_new_n1051_;
  wire new_n7828_;
  wire not_new_n1059__5;
  wire not_new_n6796_;
  wire not_new_n9262_;
  wire not_new_n8148__0;
  wire not_pi118_0;
  wire not_new_n1589__0;
  wire new_n5358_;
  wire new_n7825_;
  wire new_n9212_;
  wire new_n4881_;
  wire new_n4953_;
  wire not_new_n8798__1;
  wire new_n4752_;
  wire new_n7156_;
  wire new_n2397_;
  wire not_new_n994__47475615099430;
  wire not_new_n6005_;
  wire not_new_n2897_;
  wire not_new_n5334_;
  wire not_new_n3311__5;
  wire not_new_n7036_;
  wire not_new_n3336_;
  wire not_new_n1547_;
  wire new_n2724_;
  wire new_n4052_;
  wire new_n5442_;
  wire not_new_n6310_;
  wire new_n1014_;
  wire new_n4253_;
  wire new_n1257_;
  wire not_pi268_1;
  wire not_pi041_2;
  wire not_new_n4452__0;
  wire not_pi112;
  wire not_new_n6632_;
  wire not_new_n1051__8;
  wire not_new_n8403_;
  wire and_new_n4984__new_n5390_;
  wire new_n9728_;
  wire not_new_n928__490;
  wire new_n6657_;
  wire new_n5848_;
  wire new_n2583_;
  wire not_new_n6156_;
  wire new_n6527_;
  wire not_new_n756_;
  wire not_new_n1536__113988951853731430;
  wire not_new_n6355_;
  wire new_n3562_;
  wire not_new_n5094_;
  wire not_pi070;
  wire not_pi220;
  wire not_new_n6599_;
  wire not_new_n581__3430;
  wire not_new_n1245_;
  wire new_n9053_;
  wire not_new_n1587_;
  wire new_n9136_;
  wire not_new_n3324_;
  wire not_new_n9194_;
  wire new_n6188_;
  wire not_new_n4826_;
  wire not_new_n3761_;
  wire not_new_n5994_;
  wire new_n6967_;
  wire new_n3566_;
  wire not_new_n10100__0;
  wire new_n5003_;
  wire or_or_not_new_n2847__not_new_n2850__not_new_n2849_;
  wire not_new_n601__6;
  wire not_new_n6537__0;
  wire not_new_n5020_;
  wire not_new_n1011__1;
  wire not_new_n3389_;
  wire not_new_n1051__4;
  wire not_new_n7736_;
  wire not_new_n7495_;
  wire new_n598_;
  wire not_new_n1003__2;
  wire not_new_n1580__1176490;
  wire or_not_new_n8528__not_new_n8429_;
  wire new_n6487_;
  wire new_n10247_;
  wire not_new_n2802_;
  wire not_new_n5520_;
  wire not_new_n9018_;
  wire new_n1511_;
  wire not_new_n1596__4;
  wire not_new_n626__1915812313805664144010;
  wire new_n5167_;
  wire po111;
  wire not_new_n3323_;
  wire or_not_new_n2838__not_new_n2841_;
  wire or_or_not_new_n2527__not_new_n2531__not_new_n1421_;
  wire not_new_n640__47475615099430;
  wire not_new_n632__70;
  wire or_not_new_n3113__not_new_n3112_;
  wire or_not_new_n1299__not_new_n1297_;
  wire not_new_n1229_;
  wire not_new_n5890__0;
  wire new_n9514_;
  wire not_new_n8979_;
  wire new_n4741_;
  wire new_n2323_;
  wire not_new_n5890__3;
  wire new_n9272_;
  wire new_n4347_;
  wire not_new_n5102_;
  wire new_n4778_;
  wire new_n7305_;
  wire new_n2653_;
  wire not_new_n3278_;
  wire not_new_n2773_;
  wire not_new_n7014__1;
  wire not_new_n8117_;
  wire not_new_n6283_;
  wire not_new_n589__32199057558131797268376070;
  wire not_new_n658_;
  wire not_new_n10149_;
  wire po016;
  wire not_new_n6340_;
  wire not_new_n994__490;
  wire not_new_n8221_;
  wire not_new_n5770__0;
  wire new_n2565_;
  wire new_n7632_;
  wire not_new_n1049__10;
  wire and_new_n3750__new_n3753_;
  wire new_n1027_;
  wire new_n9156_;
  wire new_n4973_;
  wire new_n1779_;
  wire not_new_n593__10;
  wire new_n6616_;
  wire not_new_n4079_;
  wire new_n3617_;
  wire not_new_n9434_;
  wire not_new_n9071_;
  wire new_n8648_;
  wire not_new_n4481__0;
  wire not_new_n622__16284135979104490;
  wire new_n7503_;
  wire not_pi102_0;
  wire not_new_n7401_;
  wire not_new_n1067__10;
  wire new_n2251_;
  wire not_new_n6995__0;
  wire not_new_n604__8235430;
  wire or_not_new_n2883__not_new_n2886_;
  wire not_new_n644__273687473400809163430;
  wire new_n4956_;
  wire not_new_n1616__168070;
  wire new_n9343_;
  wire key_gate_67;
  wire new_n9723_;
  wire not_new_n5440_;
  wire not_new_n656_;
  wire not_new_n6610_;
  wire and_new_n1274__new_n2008_;
  wire not_new_n8306_;
  wire new_n8317_;
  wire new_n6745_;
  wire not_new_n1516_;
  wire new_n8021_;
  wire new_n7089_;
  wire or_or_not_new_n1482__not_new_n2858__not_new_n2857_;
  wire not_new_n1524_;
  wire and_new_n3073__new_n998_;
  wire new_n4654_;
  wire not_new_n1012_;
  wire new_n9996_;
  wire not_new_n3418_;
  wire new_n7294_;
  wire not_new_n718_;
  wire not_new_n728__0;
  wire not_new_n1423_;
  wire new_n8362_;
  wire not_new_n7034_;
  wire new_n7158_;
  wire not_new_n610__8;
  wire not_new_n7113__0;
  wire not_new_n6210_;
  wire not_pi173_0;
  wire new_n8642_;
  wire not_new_n6598_;
  wire not_new_n2111_;
  wire not_new_n769_;
  wire and_new_n6403__new_n6402_;
  wire not_new_n7620_;
  wire new_n3080_;
  wire new_n10142_;
  wire or_not_new_n2935__not_new_n2934_;
  wire not_new_n4078_;
  wire not_new_n3372__0;
  wire not_new_n650_;
  wire new_n9663_;
  wire not_new_n5793_;
  wire not_new_n5852_;
  wire new_n6071_;
  wire not_new_n600__4;
  wire new_n9174_;
  wire new_n4073_;
  wire not_new_n5790__0;
  wire not_new_n7826_;
  wire or_or_not_new_n1287__not_new_n1285__not_new_n2059_;
  wire not_new_n2766_;
  wire new_n1452_;
  wire not_new_n5024_;
  wire not_new_n5878__3;
  wire new_n6828_;
  wire not_new_n4793_;
  wire new_n4340_;
  wire not_new_n3796_;
  wire new_n6720_;
  wire not_new_n1004_;
  wire or_not_new_n8609__not_new_n8595__0;
  wire not_new_n6995__2;
  wire not_new_n3914__1;
  wire not_new_n4944__0;
  wire not_new_n7266_;
  wire not_new_n5672_;
  wire not_new_n7375_;
  wire not_new_n5907_;
  wire not_new_n631__70;
  wire not_new_n6148_;
  wire not_new_n1583__3430;
  wire new_n5322_;
  wire not_new_n1321_;
  wire not_new_n2813_;
  wire new_n9577_;
  wire not_new_n4690_;
  wire not_new_n5920_;
  wire not_new_n9588_;
  wire not_new_n1998_;
  wire not_new_n1010__5;
  wire not_new_n2744_;
  wire new_n4183_;
  wire not_new_n7032__0;
  wire not_new_n5941_;
  wire key_gate_81;
  wire not_new_n3485_;
  wire not_new_n6226__0;
  wire not_new_n7771__0;
  wire not_new_n1305_;
  wire new_n7499_;
  wire not_new_n3809_;
  wire new_n7688_;
  wire not_new_n4416_;
  wire new_n9482_;
  wire new_n4160_;
  wire not_new_n7445__0;
  wire not_pi145_3;
  wire not_pi131_0;
  wire not_new_n641__70;
  wire not_new_n2584_;
  wire not_new_n3029_;
  wire not_pi115_0;
  wire and_and_new_n3780__new_n3783__new_n3789_;
  wire not_new_n585__1;
  wire new_n9780_;
  wire not_new_n593__7;
  wire not_new_n4589_;
  wire po198;
  wire new_n5252_;
  wire not_new_n3907_;
  wire not_new_n1053_;
  wire not_new_n3184__138412872010;
  wire new_n5743_;
  wire new_n6080_;
  wire new_n4070_;
  wire not_new_n2635_;
  wire not_new_n8828__0;
  wire not_new_n3106_;
  wire not_new_n589__657123623635342801395430;
  wire not_new_n597__6;
  wire not_new_n641__3;
  wire new_n633_;
  wire new_n9666_;
  wire new_n8168_;
  wire not_new_n10286_;
  wire not_new_n6466_;
  wire not_new_n2972_;
  wire new_n978_;
  wire not_new_n631__16284135979104490;
  wire not_new_n1597__3;
  wire not_new_n617__7;
  wire not_new_n2703_;
  wire not_new_n2943_;
  wire not_new_n3158_;
  wire not_new_n9869__0;
  wire new_n7210_;
  wire new_n4155_;
  wire new_n6311_;
  wire new_n2559_;
  wire not_new_n3201_;
  wire new_n6581_;
  wire not_new_n7673_;
  wire not_new_n9369_;
  wire new_n8184_;
  wire not_new_n4453_;
  wire new_n6854_;
  wire not_new_n599__24010;
  wire not_new_n651_;
  wire not_new_n1587__0;
  wire not_new_n1008__0;
  wire new_n5879_;
  wire not_new_n2228_;
  wire not_new_n588__3;
  wire or_or_not_new_n1259__not_new_n1257__not_new_n1926_;
  wire new_n9013_;
  wire not_new_n4336_;
  wire and_new_n2327__new_n2328_;
  wire not_po298_8235430;
  wire not_new_n626__93874803376477543056490;
  wire new_n1725_;
  wire new_n5271_;
  wire not_pi064_6;
  wire new_n8504_;
  wire not_pi050_3;
  wire new_n5368_;
  wire not_new_n3863_;
  wire not_new_n603__403536070;
  wire not_new_n5804__0;
  wire new_n4615_;
  wire new_n7274_;
  wire or_not_new_n4818__not_new_n4749_;
  wire new_n6145_;
  wire new_n9338_;
  wire not_pi269_5;
  wire new_n7446_;
  wire new_n6677_;
  wire or_not_new_n1844__not_new_n1845_;
  wire not_new_n3091_;
  wire not_new_n8270_;
  wire new_n2606_;
  wire new_n4459_;
  wire or_or_or_not_new_n2910__not_new_n2913__not_new_n2912__not_new_n2914_;
  wire not_new_n4787__1;
  wire not_new_n10029__1;
  wire not_new_n7152_;
  wire new_n7302_;
  wire not_pi082;
  wire not_new_n4126__2;
  wire not_new_n2685_;
  wire not_new_n7232_;
  wire new_n8793_;
  wire not_new_n984__8235430;
  wire new_n9529_;
  wire not_new_n5837_;
  wire not_new_n8807_;
  wire new_n4944_;
  wire new_n2361_;
  wire new_n9366_;
  wire new_n3925_;
  wire not_new_n5417_;
  wire not_new_n603__8235430;
  wire new_n2362_;
  wire not_new_n5768__0;
  wire not_new_n1010__6;
  wire not_new_n618__93874803376477543056490;
  wire not_new_n989__1;
  wire not_new_n645__0;
  wire new_n9093_;
  wire new_n4025_;
  wire new_n7714_;
  wire not_new_n593__138412872010;
  wire new_n6321_;
  wire not_pi243;
  wire not_new_n8266_;
  wire not_new_n7300_;
  wire new_n1439_;
  wire new_n7853_;
  wire or_not_new_n2962__not_new_n2961_;
  wire new_n6215_;
  wire not_new_n10103_;
  wire new_n3507_;
  wire not_new_n3746_;
  wire not_new_n8578_;
  wire new_n1920_;
  wire not_new_n638__70;
  wire new_n8951_;
  wire not_new_n4435_;
  wire not_new_n6779_;
  wire new_n3114_;
  wire not_new_n600__2326305139872070;
  wire or_not_new_n2792__not_new_n2791_;
  wire not_new_n4658_;
  wire not_new_n589__2326305139872070;
  wire not_new_n5504_;
  wire not_new_n6902_;
  wire not_pi185;
  wire new_n3098_;
  wire new_n5745_;
  wire not_new_n8637_;
  wire not_new_n8920_;
  wire new_n7350_;
  wire new_n3303_;
  wire not_new_n2135_;
  wire not_new_n1598__47475615099430;
  wire not_new_n3359_;
  wire not_new_n1435_;
  wire new_n6777_;
  wire not_new_n6926_;
  wire new_n632_;
  wire not_new_n7647_;
  wire not_new_n984__9;
  wire not_new_n8846__0;
  wire not_pi136;
  wire new_n4735_;
  wire not_new_n6481__1;
  wire new_n7003_;
  wire not_new_n730__0;
  wire new_n9547_;
  wire or_not_new_n1235__not_new_n1233_;
  wire new_n9166_;
  wire new_n3896_;
  wire new_n8520_;
  wire not_pi186;
  wire not_new_n679_;
  wire new_n8026_;
  wire new_n8385_;
  wire not_new_n3978_;
  wire new_n5932_;
  wire not_new_n3906_;
  wire po240;
  wire not_new_n8794_;
  wire new_n6250_;
  wire not_new_n1031__6;
  wire not_new_n2469_;
  wire not_new_n2738_;
  wire new_n1796_;
  wire not_new_n8900__0;
  wire not_new_n4558_;
  wire new_n9541_;
  wire not_new_n7032_;
  wire new_n10195_;
  wire not_new_n1597_;
  wire new_n4101_;
  wire not_new_n8250_;
  wire not_new_n984__5;
  wire not_new_n1005__2;
  wire new_n8431_;
  wire not_new_n8927_;
  wire new_n3251_;
  wire new_n5929_;
  wire not_new_n648__9;
  wire not_new_n989__797922662976120010;
  wire not_new_n6460_;
  wire and_new_n1270__new_n1989_;
  wire not_new_n2000_;
  wire not_new_n1589__8235430;
  wire new_n8991_;
  wire not_new_n636__2824752490;
  wire not_new_n9863_;
  wire new_n4555_;
  wire new_n5705_;
  wire not_new_n1596__332329305696010;
  wire not_new_n640__0;
  wire new_n4859_;
  wire not_new_n1588__1;
  wire not_new_n8543_;
  wire new_n9958_;
  wire not_new_n628__168070;
  wire new_n2008_;
  wire not_new_n645__24010;
  wire new_n7624_;
  wire new_n2922_;
  wire not_new_n7226_;
  wire not_new_n4651_;
  wire not_new_n589__4599865365447399609768010;
  wire not_pi228;
  wire not_new_n1041__47475615099430;
  wire not_pi163_0;
  wire new_n4548_;
  wire not_new_n8266__3;
  wire new_n6275_;
  wire new_n5567_;
  wire new_n9303_;
  wire or_or_not_new_n1562__not_new_n2469__not_new_n1393_;
  wire new_n6647_;
  wire not_new_n7016__0;
  wire not_new_n3116_;
  wire new_n4965_;
  wire po054;
  wire new_n6683_;
  wire new_n6818_;
  wire not_new_n1059__10;
  wire not_new_n648__273687473400809163430;
  wire new_n3974_;
  wire new_n7892_;
  wire new_n6576_;
  wire not_new_n5205_;
  wire and_and_and_new_n6422__new_n6426__new_n6360__new_n6359_;
  wire not_pi132_3;
  wire not_new_n2224_;
  wire not_pi050_2;
  wire new_n2671_;
  wire not_new_n1602__8235430;
  wire not_new_n5067_;
  wire new_n10038_;
  wire new_n8070_;
  wire not_new_n597__1176490;
  wire not_new_n738__1;
  wire not_new_n8053_;
  wire new_n2149_;
  wire new_n6813_;
  wire not_new_n1978_;
  wire new_n8000_;
  wire not_new_n7871_;
  wire not_new_n1675_;
  wire new_n9223_;
  wire not_new_n1027__273687473400809163430;
  wire new_n6373_;
  wire new_n1252_;
  wire not_new_n1591__168070;
  wire new_n2358_;
  wire not_new_n6285_;
  wire not_new_n3141_;
  wire not_new_n775__1176490;
  wire not_new_n1581__332329305696010;
  wire not_new_n3559_;
  wire not_pi140_3;
  wire not_new_n1536__968890104070;
  wire not_new_n611__3430;
  wire new_n9689_;
  wire not_pi057_3;
  wire new_n10187_;
  wire new_n2960_;
  wire new_n8245_;
  wire new_n1997_;
  wire new_n7531_;
  wire not_new_n1534_;
  wire not_new_n5808_;
  wire not_new_n7983_;
  wire not_new_n6243_;
  wire new_n4981_;
  wire new_n7542_;
  wire new_n7518_;
  wire not_new_n7327_;
  wire not_new_n5725_;
  wire not_new_n604__4;
  wire not_new_n6801_;
  wire not_new_n5546_;
  wire not_new_n7281_;
  wire new_n9310_;
  wire not_new_n631__797922662976120010;
  wire not_new_n4130__0;
  wire not_new_n8921_;
  wire new_n6653_;
  wire new_n4055_;
  wire new_n3462_;
  wire not_new_n1045__138412872010;
  wire not_new_n5025_;
  wire new_n4967_;
  wire not_new_n3392_;
  wire not_pi103_0;
  wire new_n2352_;
  wire new_n5628_;
  wire not_new_n8992__0;
  wire new_n6842_;
  wire new_n10041_;
  wire not_new_n4811_;
  wire not_new_n989__6782230728490;
  wire new_n6403_;
  wire not_new_n9925_;
  wire not_new_n585__8;
  wire not_new_n8429_;
  wire new_n10340_;
  wire not_new_n6480__0;
  wire new_n3595_;
  wire not_new_n3169_;
  wire new_n10005_;
  wire not_new_n3872_;
  wire not_new_n10290_;
  wire not_new_n2646_;
  wire new_n8587_;
  wire new_n9679_;
  wire not_new_n4252_;
  wire not_new_n2021_;
  wire not_pi170;
  wire not_pi063_1;
  wire new_n9451_;
  wire new_n10024_;
  wire new_n9976_;
  wire not_new_n8169__0;
  wire not_new_n3731_;
  wire not_new_n7764_;
  wire not_new_n3870_;
  wire new_n8490_;
  wire not_new_n5637_;
  wire not_new_n588__1176490;
  wire not_new_n5486_;
  wire not_new_n7354_;
  wire not_new_n7157_;
  wire new_n4408_;
  wire new_n4518_;
  wire new_n5998_;
  wire not_new_n3283_;
  wire new_n585_;
  wire not_new_n1601__403536070;
  wire not_new_n5257_;
  wire and_and_new_n2508__new_n2510__new_n2507_;
  wire not_new_n6201_;
  wire not_new_n1008__5;
  wire not_new_n1345_;
  wire key_gate_92;
  wire new_n6230_;
  wire not_new_n4571_;
  wire new_n5594_;
  wire new_n7388_;
  wire new_n7630_;
  wire not_new_n9158_;
  wire new_n3543_;
  wire not_new_n6222_;
  wire not_new_n9431_;
  wire not_new_n618__490;
  wire not_new_n4737_;
  wire not_new_n4749__1;
  wire not_new_n618__3430;
  wire not_pi205;
  wire not_new_n1598__24010;
  wire new_n9988_;
  wire not_new_n4017__2;
  wire not_new_n9213_;
  wire not_new_n629__16284135979104490;
  wire new_n9515_;
  wire not_new_n6278_;
  wire not_new_n618__3;
  wire new_n2503_;
  wire not_new_n597__19773267430;
  wire new_n2258_;
  wire not_new_n586_;
  wire not_pi147_4;
  wire new_n639_;
  wire not_pi100_0;
  wire not_new_n3297_;
  wire new_n9171_;
  wire not_new_n3185__70;
  wire new_n10220_;
  wire not_new_n6044_;
  wire not_new_n624__2326305139872070;
  wire not_new_n7695_;
  wire not_new_n705_;
  wire not_new_n4655_;
  wire not_new_n6578_;
  wire new_n2734_;
  wire new_n7450_;
  wire not_new_n2797_;
  wire key_gate_21;
  wire not_new_n10252_;
  wire new_n7768_;
  wire not_new_n6646_;
  wire not_new_n1601__47475615099430;
  wire not_new_n4121_;
  wire not_new_n597__1;
  wire not_new_n6807_;
  wire not_new_n3185__10;
  wire not_new_n3760_;
  wire not_new_n4429__0;
  wire not_new_n6571_;
  wire not_new_n638__8235430;
  wire new_n1472_;
  wire new_n8708_;
  wire not_new_n581__4599865365447399609768010;
  wire new_n6606_;
  wire new_n2534_;
  wire new_n9137_;
  wire not_new_n1522_;
  wire new_n2202_;
  wire new_n1347_;
  wire new_n3653_;
  wire or_not_new_n3124__not_new_n3125_;
  wire not_pi036_0;
  wire new_n2844_;
  wire po085;
  wire not_new_n8350_;
  wire or_not_new_n2892__not_new_n2895_;
  wire not_new_n5777__0;
  wire not_new_n10338_;
  wire new_n6922_;
  wire not_new_n635__10;
  wire not_new_n3089_;
  wire new_n9564_;
  wire or_or_not_new_n1560__not_new_n2459__not_new_n1389_;
  wire not_new_n4957_;
  wire not_new_n619__2;
  wire not_new_n5632_;
  wire not_new_n7730_;
  wire not_new_n633__1176490;
  wire not_new_n1536__6782230728490;
  wire new_n6718_;
  wire new_n10004_;
  wire not_new_n643__7;
  wire not_new_n5966_;
  wire new_n5535_;
  wire new_n1778_;
  wire new_n10193_;
  wire not_new_n1684_;
  wire new_n5635_;
  wire new_n1914_;
  wire not_new_n595__70;
  wire not_new_n4479__0;
  wire new_n6663_;
  wire new_n4994_;
  wire new_n6627_;
  wire not_new_n8134__2;
  wire not_new_n9823_;
  wire not_new_n7258__0;
  wire new_n769_;
  wire new_n1152_;
  wire not_new_n8478_;
  wire new_n4337_;
  wire new_n9807_;
  wire not_new_n3888_;
  wire new_n8145_;
  wire not_new_n1596__273687473400809163430;
  wire not_new_n7186_;
  wire not_new_n4163__0;
  wire not_new_n3461_;
  wire po275;
  wire not_new_n5561_;
  wire new_n1605_;
  wire new_n7656_;
  wire not_new_n5569_;
  wire not_new_n5032_;
  wire new_n999_;
  wire not_new_n6482__2;
  wire not_new_n4672_;
  wire not_new_n598_;
  wire new_n6691_;
  wire new_n5822_;
  wire new_n8144_;
  wire new_n1597_;
  wire new_n7311_;
  wire not_new_n9404_;
  wire new_n754_;
  wire not_new_n1027__8235430;
  wire new_n10097_;
  wire not_new_n586__7;
  wire not_new_n7218_;
  wire not_new_n1630_;
  wire not_new_n4450__0;
  wire new_n6381_;
  wire not_new_n3315__968890104070;
  wire not_pi048_2;
  wire not_new_n1838_;
  wire new_n3284_;
  wire not_new_n2828_;
  wire new_n8763_;
  wire not_new_n5776_;
  wire new_n3528_;
  wire not_new_n6708_;
  wire not_new_n628__332329305696010;
  wire not_new_n7939_;
  wire new_n2099_;
  wire not_new_n6062_;
  wire not_new_n986_;
  wire not_new_n2919_;
  wire not_new_n5811_;
  wire new_n5926_;
  wire new_n1461_;
  wire or_not_new_n2917__not_new_n2916_;
  wire not_new_n581__138412872010;
  wire new_n2486_;
  wire new_n4472_;
  wire not_new_n5892_;
  wire not_new_n1827_;
  wire new_n4869_;
  wire new_n6673_;
  wire not_new_n9457_;
  wire not_new_n984__403536070;
  wire new_n4968_;
  wire new_n5616_;
  wire po135;
  wire new_n5323_;
  wire new_n10205_;
  wire not_new_n6655__0;
  wire new_n1995_;
  wire not_new_n5813_;
  wire new_n4086_;
  wire not_new_n7967_;
  wire new_n948_;
  wire not_new_n6764_;
  wire new_n5646_;
  wire not_new_n653_;
  wire new_n9241_;
  wire new_n9478_;
  wire not_new_n6249_;
  wire not_new_n645__403536070;
  wire new_n2381_;
  wire not_new_n3315__1176490;
  wire po096;
  wire new_n3064_;
  wire new_n4170_;
  wire not_new_n4951_;
  wire or_not_new_n4814__not_new_n4734_;
  wire new_n8094_;
  wire not_new_n1613__6;
  wire not_new_n1618_;
  wire new_n8634_;
  wire not_new_n7806_;
  wire not_new_n3173_;
  wire not_new_n5877_;
  wire not_new_n604__7;
  wire not_new_n634__10;
  wire po184;
  wire new_n7722_;
  wire not_new_n1007__1;
  wire not_new_n7804_;
  wire new_n6360_;
  wire new_n10252_;
  wire not_new_n998_;
  wire not_new_n5019_;
  wire new_n3902_;
  wire new_n4191_;
  wire new_n3157_;
  wire new_n5689_;
  wire not_new_n10302_;
  wire new_n3482_;
  wire not_new_n5657_;
  wire not_new_n4777_;
  wire new_n8609_;
  wire not_new_n586__10;
  wire not_new_n3502_;
  wire not_new_n2038_;
  wire po258;
  wire new_n3103_;
  wire not_pi066_0;
  wire not_new_n1585__57648010;
  wire not_new_n3838_;
  wire new_n8899_;
  wire not_new_n1534__9;
  wire not_new_n589__93874803376477543056490;
  wire new_n1003_;
  wire not_new_n9487_;
  wire new_n7571_;
  wire new_n6216_;
  wire not_new_n588__57648010;
  wire new_n1269_;
  wire not_new_n633__490;
  wire not_new_n3775_;
  wire not_new_n8116_;
  wire not_new_n1562_;
  wire not_new_n7340_;
  wire not_new_n9867_;
  wire not_new_n1588__16284135979104490;
  wire not_new_n625__2326305139872070;
  wire not_new_n7837__0;
  wire not_new_n1450_;
  wire new_n10192_;
  wire not_new_n9573_;
  wire not_new_n9260_;
  wire not_new_n7980_;
  wire new_n9312_;
  wire not_new_n8457_;
  wire new_n3151_;
  wire new_n7162_;
  wire new_n10240_;
  wire not_new_n9400_;
  wire not_new_n4547_;
  wire new_n7057_;
  wire new_n10297_;
  wire new_n2005_;
  wire not_new_n7717_;
  wire new_n9424_;
  wire not_new_n2843_;
  wire not_new_n641__168070;
  wire new_n7329_;
  wire new_n6277_;
  wire not_new_n8418_;
  wire not_new_n8458_;
  wire new_n6318_;
  wire not_new_n5882__0;
  wire not_pi036_3;
  wire not_new_n7941_;
  wire not_new_n8187_;
  wire not_new_n1538__8;
  wire new_n6589_;
  wire not_new_n630__2;
  wire new_n5834_;
  wire not_new_n632__57648010;
  wire new_n5049_;
  wire not_new_n591__3430;
  wire new_n4163_;
  wire not_new_n6613__0;
  wire not_new_n8304_;
  wire new_n8802_;
  wire new_n5539_;
  wire not_new_n1568_;
  wire and_and_new_n6422__new_n6426__new_n6360_;
  wire not_new_n617__39098210485829880490;
  wire not_new_n631__6;
  wire new_n9454_;
  wire not_new_n6550_;
  wire not_new_n2474_;
  wire new_n7898_;
  wire not_new_n9459_;
  wire not_new_n5921_;
  wire po288;
  wire not_new_n1031__1176490;
  wire new_n5212_;
  wire not_new_n8143_;
  wire not_pi268_0;
  wire new_n2582_;
  wire not_new_n1028__5;
  wire not_new_n1047__1;
  wire new_n940_;
  wire not_new_n1155__0;
  wire and_and_not_pi040_1_not_pi039_1_not_pi042_1;
  wire not_new_n7363__0;
  wire not_new_n587__2326305139872070;
  wire new_n4716_;
  wire not_new_n617_;
  wire not_new_n5741__1;
  wire not_new_n5346_;
  wire not_new_n7035__1;
  wire not_pi217;
  wire not_new_n2921_;
  wire not_new_n5434_;
  wire not_new_n1316_;
  wire new_n2497_;
  wire not_new_n641__4;
  wire new_n3899_;
  wire new_n9859_;
  wire not_new_n6767_;
  wire not_new_n5911_;
  wire not_new_n5874_;
  wire not_new_n3185__8;
  wire or_not_new_n8799__0_not_new_n8996__0;
  wire new_n4750_;
  wire not_new_n1063__4;
  wire not_new_n7657_;
  wire not_pi144_1;
  wire not_new_n1598__3430;
  wire not_new_n1601__5585458640832840070;
  wire not_new_n1007__3;
  wire not_new_n606__6;
  wire not_new_n6969_;
  wire not_new_n595__168070;
  wire not_new_n1055__39098210485829880490;
  wire not_new_n1960_;
  wire new_n8098_;
  wire new_n2609_;
  wire not_new_n7059_;
  wire new_n5116_;
  wire not_new_n8560_;
  wire not_new_n7140_;
  wire not_new_n637__968890104070;
  wire new_n3940_;
  wire not_new_n8618__0;
  wire not_new_n1061__19773267430;
  wire and_and_new_n2181__new_n2184__new_n2182_;
  wire not_new_n5715_;
  wire new_n8774_;
  wire not_new_n1594__8;
  wire not_new_n1065__24010;
  wire new_n5150_;
  wire not_new_n1591__0;
  wire new_n1814_;
  wire not_new_n3743_;
  wire po102;
  wire not_new_n6371_;
  wire new_n5843_;
  wire new_n4106_;
  wire not_new_n5798__2;
  wire new_n4184_;
  wire new_n2171_;
  wire new_n9476_;
  wire new_n8971_;
  wire not_new_n4184_;
  wire new_n5224_;
  wire new_n8285_;
  wire or_or_not_new_n3914__not_new_n3969__not_new_n4014_;
  wire new_n6515_;
  wire key_gate_61;
  wire not_new_n3469_;
  wire new_n1987_;
  wire not_new_n9676_;
  wire new_n3941_;
  wire not_new_n9386__0;
  wire new_n5052_;
  wire not_new_n5256_;
  wire new_n3666_;
  wire not_new_n7105_;
  wire not_new_n1004__1;
  wire not_pi120;
  wire not_new_n8259_;
  wire not_new_n5842_;
  wire not_new_n2950_;
  wire not_new_n581__4;
  wire not_new_n3376_;
  wire not_new_n9634_;
  wire not_new_n994__2326305139872070;
  wire not_new_n7255_;
  wire new_n6938_;
  wire not_new_n10330_;
  wire new_n9612_;
  wire new_n7618_;
  wire new_n5869_;
  wire not_new_n7522_;
  wire new_n6649_;
  wire new_n4484_;
  wire not_new_n6147_;
  wire po075;
  wire new_n1886_;
  wire new_n1485_;
  wire not_new_n4073_;
  wire not_new_n4163_;
  wire not_new_n1600_;
  wire not_pi036_1;
  wire not_new_n8243_;
  wire new_n4922_;
  wire and_new_n3058__new_n998_;
  wire not_new_n627__2;
  wire not_new_n1581__70;
  wire new_n2228_;
  wire not_new_n5240__0;
  wire new_n7061_;
  wire new_n7129_;
  wire not_new_n6628_;
  wire not_new_n7611__0;
  wire new_n1365_;
  wire not_new_n629__138412872010;
  wire not_new_n2243_;
  wire new_n1797_;
  wire not_new_n1806_;
  wire new_n6474_;
  wire new_n4350_;
  wire not_new_n631__9;
  wire not_pi275_0;
  wire not_new_n8740_;
  wire not_new_n1594__6;
  wire not_new_n6713_;
  wire not_new_n4479_;
  wire not_new_n636__6;
  wire new_n8185_;
  wire not_new_n2674_;
  wire new_n4021_;
  wire not_new_n4550_;
  wire or_not_new_n1327__not_new_n1325_;
  wire new_n4194_;
  wire not_new_n5949_;
  wire new_n4858_;
  wire not_new_n1053__6;
  wire new_n6185_;
  wire po151;
  wire not_new_n6451_;
  wire and_new_n3732__new_n3735_;
  wire new_n5680_;
  wire new_n5242_;
  wire not_pi022;
  wire new_n3545_;
  wire new_n1699_;
  wire new_n4822_;
  wire not_new_n4157_;
  wire not_new_n3326_;
  wire new_n9708_;
  wire not_new_n1598__8235430;
  wire new_n5352_;
  wire new_n5872_;
  wire new_n4779_;
  wire new_n5140_;
  wire not_pi045;
  wire not_new_n1415_;
  wire not_pi174_0;
  wire not_new_n607__2;
  wire not_new_n5794__1;
  wire new_n3645_;
  wire new_n3747_;
  wire not_new_n647__113988951853731430;
  wire new_n2842_;
  wire not_new_n9755_;
  wire key_gate_104;
  wire not_new_n9446_;
  wire not_new_n8236_;
  wire or_or_not_new_n3397__not_new_n3398__not_new_n1761_;
  wire not_new_n6663__0;
  wire new_n10294_;
  wire new_n7199_;
  wire new_n7796_;
  wire not_new_n3017_;
  wire not_new_n2820_;
  wire new_n9511_;
  wire not_new_n7776_;
  wire not_new_n6412_;
  wire new_n6047_;
  wire not_new_n1067__1176490;
  wire new_n8849_;
  wire not_new_n641__10;
  wire not_new_n8266__2;
  wire new_n1301_;
  wire new_n10212_;
  wire not_new_n1031_;
  wire new_n3346_;
  wire new_n5633_;
  wire not_new_n2142_;
  wire not_new_n5042_;
  wire not_new_n10209_;
  wire not_new_n9149_;
  wire not_new_n620__3;
  wire new_n9902_;
  wire not_new_n9905_;
  wire new_n5345_;
  wire new_n3088_;
  wire not_new_n8983__0;
  wire not_new_n710_;
  wire not_new_n1895_;
  wire not_new_n6962_;
  wire new_n5858_;
  wire new_n660_;
  wire not_new_n619__19773267430;
  wire not_new_n9135_;
  wire new_n2761_;
  wire new_n5287_;
  wire not_new_n2727_;
  wire not_new_n1566_;
  wire new_n7841_;
  wire new_n6439_;
  wire not_pi052_3;
  wire not_new_n3204_;
  wire new_n3467_;
  wire not_new_n6860_;
  wire po011;
  wire not_new_n8131_;
  wire new_n4297_;
  wire new_n2424_;
  wire new_n7153_;
  wire not_new_n1594__168070;
  wire not_new_n4434__0;
  wire new_n4640_;
  wire not_new_n1538__332329305696010;
  wire new_n966_;
  wire new_n9332_;
  wire not_new_n3520_;
  wire po087;
  wire not_new_n1611__113988951853731430;
  wire new_n6193_;
  wire not_pi267_0;
  wire not_new_n625__332329305696010;
  wire not_new_n3184__47475615099430;
  wire not_pi170_2;
  wire new_n7200_;
  wire new_n3670_;
  wire new_n6156_;
  wire not_new_n8817_;
  wire new_n4976_;
  wire not_new_n1603__3;
  wire not_new_n4816_;
  wire new_n7290_;
  wire new_n9512_;
  wire new_n6127_;
  wire new_n751_;
  wire new_n1220_;
  wire not_new_n8194_;
  wire not_new_n1648_;
  wire not_new_n1538__797922662976120010;
  wire not_new_n9905__0;
  wire not_new_n5766_;
  wire not_new_n1608_;
  wire not_new_n8435_;
  wire and_new_n1222__new_n1223_;
  wire not_new_n1612__113988951853731430;
  wire not_new_n591__47475615099430;
  wire not_new_n5474_;
  wire new_n2082_;
  wire not_new_n4775__1;
  wire new_n2687_;
  wire new_n8056_;
  wire new_n8518_;
  wire not_new_n601__1176490;
  wire and_new_n9512__new_n9773_;
  wire not_pi137;
  wire not_new_n624__968890104070;
  wire not_new_n1613__968890104070;
  wire not_new_n6812__0;
  wire not_new_n6463_;
  wire not_new_n1447_;
  wire new_n5548_;
  wire new_n9347_;
  wire not_new_n5169_;
  wire not_pi264;
  wire not_pi132;
  wire not_new_n4840_;
  wire new_n2850_;
  wire new_n1900_;
  wire new_n6755_;
  wire new_n6416_;
  wire not_new_n5824_;
  wire not_pi045_2;
  wire not_new_n618__24010;
  wire or_not_new_n1545__not_new_n1360_;
  wire new_n1726_;
  wire not_new_n2956_;
  wire not_new_n8899_;
  wire not_new_n7073_;
  wire and_and_new_n2124__new_n2127__new_n2125_;
  wire new_n2619_;
  wire not_new_n4443_;
  wire not_new_n621__47475615099430;
  wire not_new_n1792_;
  wire not_new_n2793_;
  wire not_new_n2073_;
  wire not_new_n647__490;
  wire po168;
  wire not_new_n1063__3430;
  wire not_new_n3970_;
  wire not_po296_5080218607396233653221881976522165017724345248360010;
  wire not_new_n4032__0;
  wire new_n3876_;
  wire not_new_n7597__0;
  wire new_n4687_;
  wire new_n7125_;
  wire new_n2700_;
  wire new_n1783_;
  wire not_new_n3455_;
  wire not_new_n647__3430;
  wire not_new_n621__9;
  wire new_n2142_;
  wire new_n4745_;
  wire new_n3252_;
  wire po009;
  wire not_new_n1607__0;
  wire not_new_n1581_;
  wire not_new_n4114__2;
  wire not_new_n588__7;
  wire not_new_n7412__1;
  wire not_new_n8124__0;
  wire new_n5013_;
  wire new_n580_;
  wire new_n7607_;
  wire new_n3556_;
  wire not_new_n618__1;
  wire new_n6382_;
  wire not_new_n1585__24010;
  wire not_new_n621__8;
  wire not_new_n591__1;
  wire and_new_n8724__new_n8726_;
  wire not_new_n2926_;
  wire new_n1209_;
  wire not_new_n581__32199057558131797268376070;
  wire not_new_n3315__9;
  wire new_n6164_;
  wire po226;
  wire not_new_n5483__0;
  wire not_new_n1596__2326305139872070;
  wire not_new_n2731_;
  wire not_new_n3203_;
  wire not_new_n1160_;
  wire and_and_new_n2327__new_n2328__new_n2331_;
  wire or_not_new_n4829__not_new_n4794_;
  wire not_new_n4899_;
  wire not_new_n1055__113988951853731430;
  wire new_n6841_;
  wire not_new_n6635__3;
  wire not_new_n9955_;
  wire new_n8560_;
  wire new_n1901_;
  wire new_n4737_;
  wire not_new_n5219_;
  wire not_new_n727__1;
  wire new_n8252_;
  wire new_n2860_;
  wire not_new_n3981__1;
  wire not_new_n9886_;
  wire not_new_n7454__2;
  wire not_new_n5055_;
  wire not_new_n607__3430;
  wire not_new_n6753_;
  wire new_n3042_;
  wire or_not_new_n2565__not_new_n2564_;
  wire new_n3313_;
  wire new_n9520_;
  wire or_not_new_n1263__not_new_n1261_;
  wire not_new_n6830_;
  wire not_new_n624__3;
  wire not_new_n1443_;
  wire not_pi170_3;
  wire new_n6999_;
  wire not_new_n623_;
  wire new_n9489_;
  wire new_n9774_;
  wire not_new_n4788_;
  wire not_new_n5059__0;
  wire not_new_n1059__138412872010;
  wire new_n8167_;
  wire new_n3594_;
  wire not_new_n6221_;
  wire new_n8350_;
  wire new_n1489_;
  wire new_n2779_;
  wire new_n3763_;
  wire new_n6099_;
  wire new_n7165_;
  wire new_n9919_;
  wire new_n3839_;
  wire not_new_n613__2;
  wire not_new_n1006_;
  wire new_n1674_;
  wire not_new_n1045__8;
  wire and_new_n8692__new_n8691_;
  wire not_new_n8640_;
  wire new_n8034_;
  wire new_n6501_;
  wire not_new_n10250_;
  wire not_new_n9452_;
  wire po017;
  wire new_n691_;
  wire new_n3847_;
  wire not_new_n9905__1;
  wire not_new_n3109_;
  wire not_new_n1071__19773267430;
  wire po097;
  wire new_n3806_;
  wire not_new_n3546_;
  wire not_new_n5900__4;
  wire not_new_n4927_;
  wire new_n5040_;
  wire new_n9465_;
  wire not_new_n8113__0;
  wire new_n8645_;
  wire not_pi059;
  wire new_n1753_;
  wire not_new_n6846_;
  wire not_new_n3299_;
  wire new_n4599_;
  wire not_new_n631__8235430;
  wire new_n8955_;
  wire not_new_n5963_;
  wire not_new_n1728__24010;
  wire and_new_n10047__new_n10048_;
  wire new_n6109_;
  wire not_new_n10090_;
  wire not_new_n1201_;
  wire new_n5027_;
  wire not_new_n4631_;
  wire not_new_n639__1;
  wire not_new_n5829_;
  wire not_new_n598__8;
  wire not_pi138_0;
  wire new_n2325_;
  wire not_pi114_0;
  wire not_new_n640_;
  wire not_new_n5213_;
  wire not_new_n3048_;
  wire new_n7582_;
  wire not_new_n9631_;
  wire not_new_n6634__2;
  wire new_n2084_;
  wire not_new_n9888_;
  wire not_new_n642__1;
  wire not_new_n7439_;
  wire new_n7742_;
  wire or_not_new_n5184__not_new_n5183_;
  wire not_new_n4048_;
  wire not_new_n4717_;
  wire new_n4028_;
  wire new_n3717_;
  wire new_n8146_;
  wire not_new_n4762__0;
  wire not_new_n5777_;
  wire not_new_n5383_;
  wire new_n2126_;
  wire new_n9932_;
  wire not_new_n5878__0;
  wire not_new_n5271_;
  wire new_n8962_;
  wire new_n5249_;
  wire not_new_n8106__2;
  wire not_new_n3366_;
  wire new_n8058_;
  wire not_new_n3288_;
  wire not_new_n679__0;
  wire new_n9052_;
  wire not_new_n5789__0;
  wire not_new_n9805_;
  wire new_n10060_;
  wire new_n720_;
  wire not_new_n9352_;
  wire not_new_n5450__0;
  wire not_new_n6997_;
  wire not_new_n1601__7;
  wire not_new_n700_;
  wire new_n10228_;
  wire not_new_n5027_;
  wire not_new_n9119__0;
  wire not_new_n1545_;
  wire not_new_n5887_;
  wire new_n7482_;
  wire not_new_n603__3;
  wire not_new_n7041__1;
  wire not_new_n1849_;
  wire not_new_n5786__0;
  wire not_new_n638__13410686196639649008070;
  wire not_new_n6169_;
  wire not_new_n601__10;
  wire new_n2019_;
  wire new_n6484_;
  wire new_n7297_;
  wire not_new_n7418__1;
  wire not_new_n618__6782230728490;
  wire not_new_n8324_;
  wire not_new_n3917__0;
  wire not_po298_797922662976120010;
  wire new_n10214_;
  wire not_new_n3396_;
  wire new_n9693_;
  wire not_new_n5014_;
  wire not_new_n1900_;
  wire not_new_n629__168070;
  wire new_n8278_;
  wire not_po298_70;
  wire new_n9943_;
  wire not_new_n3315__24010;
  wire or_not_new_n4291__not_new_n4326_;
  wire new_n4410_;
  wire new_n6014_;
  wire not_new_n3140_;
  wire new_n5654_;
  wire new_n9110_;
  wire not_new_n3727_;
  wire new_n5576_;
  wire and_and_and_new_n1043__new_n6232__new_n6229__new_n6317_;
  wire not_new_n6974__1176490;
  wire new_n4740_;
  wire not_new_n7430__2;
  wire new_n6900_;
  wire new_n3377_;
  wire new_n1798_;
  wire new_n4181_;
  wire not_new_n9546_;
  wire not_new_n1028__7;
  wire not_new_n9978_;
  wire not_new_n1616__490;
  wire new_n2284_;
  wire not_new_n7007__1;
  wire new_n8771_;
  wire not_new_n1178_;
  wire not_new_n1581__10;
  wire new_n1951_;
  wire new_n6908_;
  wire not_new_n5895_;
  wire not_new_n6361_;
  wire not_new_n6871_;
  wire new_n9333_;
  wire and_and_new_n6244__new_n6372__new_n1596_;
  wire not_new_n624__24010;
  wire not_new_n3874_;
  wire not_new_n3213_;
  wire not_new_n641__19773267430;
  wire not_new_n10019_;
  wire not_pi125_0;
  wire not_new_n4091_;
  wire new_n7806_;
  wire new_n3021_;
  wire not_new_n8445_;
  wire new_n3932_;
  wire new_n10071_;
  wire not_new_n4155__1;
  wire not_new_n8852_;
  wire new_n2830_;
  wire new_n4371_;
  wire not_new_n1591__24010;
  wire new_n4650_;
  wire not_new_n7018_;
  wire key_gate_74;
  wire and_new_n3061__new_n998_;
  wire not_pi134_3;
  wire new_n7278_;
  wire new_n4249_;
  wire new_n6490_;
  wire not_new_n9510__0;
  wire not_new_n7813_;
  wire new_n4359_;
  wire new_n9219_;
  wire not_new_n1850_;
  wire not_new_n624_;
  wire new_n7265_;
  wire new_n7170_;
  wire new_n4257_;
  wire not_new_n8280_;
  wire new_n3307_;
  wire new_n3659_;
  wire not_new_n627__490;
  wire not_new_n7735__3;
  wire new_n8399_;
  wire new_n8390_;
  wire not_new_n5414_;
  wire new_n760_;
  wire not_new_n1163__0;
  wire new_n4063_;
  wire not_new_n631__968890104070;
  wire new_n7932_;
  wire not_new_n9743_;
  wire not_new_n10132_;
  wire not_new_n6538_;
  wire not_new_n6475__0;
  wire not_new_n9471_;
  wire not_new_n1315_;
  wire new_n5691_;
  wire not_new_n8166_;
  wire not_pi133;
  wire not_new_n10066_;
  wire new_n2574_;
  wire not_new_n3968_;
  wire new_n2377_;
  wire new_n5404_;
  wire or_or_not_new_n2208__not_new_n2205__not_new_n2206_;
  wire not_new_n3508_;
  wire not_new_n1049__490;
  wire not_new_n645__490;
  wire new_n1652_;
  wire not_new_n6271_;
  wire not_pi269;
  wire not_new_n1457_;
  wire not_new_n1008__2;
  wire new_n3422_;
  wire new_n7601_;
  wire not_new_n1063__10;
  wire not_pi270_1;
  wire not_new_n5749__1;
  wire not_new_n1047__968890104070;
  wire not_new_n6886_;
  wire not_new_n1768_;
  wire new_n8700_;
  wire not_new_n5297_;
  wire not_pi064;
  wire not_new_n3387__1;
  wire not_new_n3836_;
  wire not_pi257;
  wire not_new_n603__332329305696010;
  wire new_n7050_;
  wire new_n1764_;
  wire new_n9199_;
  wire not_pi109_0;
  wire not_new_n8179_;
  wire not_new_n2509__8235430;
  wire not_new_n3924__0;
  wire not_new_n6306_;
  wire not_new_n5096__0;
  wire new_n1730_;
  wire new_n6660_;
  wire new_n6428_;
  wire not_new_n7314_;
  wire not_new_n9763_;
  wire and_new_n2662__new_n2661_;
  wire new_n5029_;
  wire not_new_n589__5585458640832840070;
  wire not_new_n8286__1;
  wire new_n7022_;
  wire new_n7409_;
  wire not_new_n628__0;
  wire new_n3929_;
  wire not_new_n4825__1;
  wire new_n1545_;
  wire not_pi138_2;
  wire new_n4579_;
  wire new_n2213_;
  wire not_new_n4954__0;
  wire not_new_n1059__24010;
  wire new_n8800_;
  wire new_n4626_;
  wire not_new_n3578_;
  wire not_new_n7177_;
  wire new_n7176_;
  wire new_n4368_;
  wire not_new_n9177_;
  wire not_new_n5893_;
  wire not_new_n8996_;
  wire not_new_n3356_;
  wire not_new_n7058_;
  wire new_n3099_;
  wire not_new_n8118_;
  wire not_new_n10312_;
  wire not_new_n8866_;
  wire not_pi187_0;
  wire not_new_n989__2;
  wire not_new_n581__7;
  wire new_n1821_;
  wire not_new_n1010_;
  wire new_n9477_;
  wire not_new_n6584_;
  wire not_new_n9516_;
  wire not_new_n5109_;
  wire new_n1757_;
  wire not_new_n627__8235430;
  wire not_new_n6443__5;
  wire not_new_n8126_;
  wire new_n3079_;
  wire not_new_n1605__5;
  wire not_new_n595__332329305696010;
  wire new_n7071_;
  wire not_new_n2265_;
  wire not_new_n646__5;
  wire not_new_n1600__3430;
  wire not_new_n7082_;
  wire new_n8960_;
  wire not_new_n7487_;
  wire not_new_n8266__1;
  wire not_new_n8000_;
  wire not_new_n1045__2326305139872070;
  wire new_n4648_;
  wire new_n1574_;
  wire not_new_n9597_;
  wire not_new_n2857_;
  wire not_new_n5567_;
  wire not_new_n622__10;
  wire new_n3597_;
  wire new_n6669_;
  wire new_n2561_;
  wire not_new_n8857_;
  wire not_new_n989__113988951853731430;
  wire not_new_n8978__0;
  wire new_n3168_;
  wire not_new_n8140_;
  wire new_n9419_;
  wire and_and_new_n2276__new_n2279__new_n2277_;
  wire not_new_n8878__0;
  wire new_n1711_;
  wire new_n8892_;
  wire new_n8388_;
  wire not_new_n8451_;
  wire not_new_n9182_;
  wire and_new_n6374__new_n6372_;
  wire new_n1433_;
  wire not_new_n1071__5;
  wire new_n6852_;
  wire not_new_n1039__47475615099430;
  wire new_n8643_;
  wire and_new_n9915__new_n10334_;
  wire new_n7186_;
  wire not_new_n4415__0;
  wire new_n6039_;
  wire not_new_n1669_;
  wire not_new_n4967_;
  wire not_new_n933__0;
  wire new_n6521_;
  wire or_not_new_n4228__not_new_n4329_;
  wire not_new_n7664_;
  wire not_new_n1023__1;
  wire new_n9987_;
  wire not_new_n606__7;
  wire not_new_n10195_;
  wire new_n8105_;
  wire new_n7960_;
  wire new_n5788_;
  wire new_n9819_;
  wire not_new_n7836_;
  wire not_new_n6482_;
  wire not_new_n1049__6;
  wire new_n4166_;
  wire new_n4608_;
  wire not_new_n627__47475615099430;
  wire not_new_n1596__8;
  wire not_new_n8608_;
  wire key_gate_32;
  wire not_new_n3151_;
  wire not_new_n8035_;
  wire not_new_n1020__6;
  wire not_new_n581__52433383167563036344614587188619514555430;
  wire new_n5958_;
  wire not_new_n2981_;
  wire not_new_n9506__3;
  wire not_new_n6847_;
  wire not_new_n8139_;
  wire new_n986_;
  wire new_n7996_;
  wire new_n9944_;
  wire new_n7557_;
  wire new_n9628_;
  wire or_or_not_new_n8609__not_new_n8595__0_not_new_n1168__0;
  wire not_pi039_3;
  wire new_n4268_;
  wire not_new_n3660_;
  wire not_new_n1597__113988951853731430;
  wire not_new_n7571_;
  wire not_new_n8739_;
  wire new_n10135_;
  wire new_n4463_;
  wire not_new_n4032_;
  wire new_n2390_;
  wire not_new_n4013__0;
  wire new_n7023_;
  wire not_new_n618_;
  wire po220;
  wire or_not_new_n1565__not_new_n2484_;
  wire or_not_new_n4246__not_new_n4350_;
  wire new_n4753_;
  wire key_gate_64;
  wire new_n4015_;
  wire new_n6018_;
  wire not_new_n3310__9;
  wire new_n2746_;
  wire not_new_n6505__0;
  wire not_new_n1979_;
  wire not_new_n6443__19773267430;
  wire new_n5885_;
  wire not_new_n8392__0;
  wire new_n7537_;
  wire or_not_new_n2346__not_new_n2347_;
  wire new_n2692_;
  wire not_new_n4998__0;
  wire new_n7435_;
  wire not_new_n3184__2;
  wire not_new_n1043__3430;
  wire new_n4522_;
  wire or_not_new_n1882__not_new_n1883_;
  wire new_n2106_;
  wire new_n9073_;
  wire new_n1444_;
  wire new_n9346_;
  wire not_new_n10045_;
  wire new_n1984_;
  wire not_new_n7877_;
  wire new_n7014_;
  wire new_n9667_;
  wire not_new_n4172_;
  wire not_new_n1065__0;
  wire not_new_n9356__0;
  wire not_new_n7057_;
  wire not_new_n4704_;
  wire new_n5542_;
  wire not_new_n6791_;
  wire not_new_n6617_;
  wire new_n7109_;
  wire not_new_n581__168070;
  wire new_n9907_;
  wire not_new_n1596__5;
  wire new_n5134_;
  wire not_new_n4999__3;
  wire not_new_n6942_;
  wire not_new_n5124_;
  wire not_new_n5901__0;
  wire not_new_n4274_;
  wire new_n934_;
  wire not_pi064_3;
  wire new_n2709_;
  wire new_n1430_;
  wire new_n5655_;
  wire not_new_n1243_;
  wire not_new_n624__7;
  wire new_n8722_;
  wire not_new_n5573_;
  wire not_new_n4833_;
  wire new_n5373_;
  wire not_new_n633__8235430;
  wire new_n2107_;
  wire not_new_n8133_;
  wire new_n1660_;
  wire new_n4376_;
  wire not_new_n3495_;
  wire not_new_n5332_;
  wire or_not_new_n3134__not_new_n3133_;
  wire not_new_n1580__6782230728490;
  wire new_n6611_;
  wire new_n4284_;
  wire not_new_n5071_;
  wire not_new_n1604__6;
  wire not_po296_2115876138024253916377293617876786762900601936010;
  wire new_n9086_;
  wire not_new_n2962_;
  wire new_n2877_;
  wire new_n595_;
  wire new_n2802_;
  wire not_new_n626__5585458640832840070;
  wire not_new_n4923_;
  wire new_n5133_;
  wire not_new_n7276_;
  wire not_new_n9081_;
  wire not_new_n612__5;
  wire not_new_n934_;
  wire not_new_n637__403536070;
  wire not_new_n6876_;
  wire new_n8440_;
  wire not_new_n597__113988951853731430;
  wire not_new_n3185__2;
  wire new_n5658_;
  wire new_n2832_;
  wire not_new_n7633__0;
  wire not_new_n4439__0;
  wire not_new_n622__332329305696010;
  wire not_new_n5896_;
  wire new_n2665_;
  wire not_new_n625__13410686196639649008070;
  wire not_new_n999__0;
  wire new_n5711_;
  wire not_new_n7560_;
  wire new_n3878_;
  wire new_n9813_;
  wire new_n9035_;
  wire not_new_n1059__8235430;
  wire not_pi049_0;
  wire not_new_n599_;
  wire not_pi064_403536070;
  wire not_new_n9775_;
  wire not_new_n8168__0;
  wire not_new_n9953_;
  wire not_po296_2569235775210588780886114772242356213216070;
  wire not_new_n5455_;
  wire new_n9083_;
  wire not_new_n6614_;
  wire new_n8616_;
  wire new_n8956_;
  wire not_new_n928__2;
  wire not_pi214;
  wire new_n7698_;
  wire new_n6859_;
  wire not_new_n1280_;
  wire not_new_n9749_;
  wire not_new_n602__24010;
  wire not_new_n7316_;
  wire new_n8857_;
  wire not_new_n671_;
  wire new_n4263_;
  wire not_new_n9969_;
  wire not_new_n1594__24010;
  wire not_new_n2577_;
  wire not_new_n3790_;
  wire not_new_n1603__4;
  wire not_new_n4125__2;
  wire new_n8524_;
  wire new_n5256_;
  wire not_pi013;
  wire new_n7391_;
  wire not_new_n9392_;
  wire new_n2430_;
  wire new_n8158_;
  wire new_n3201_;
  wire new_n6577_;
  wire not_new_n581__9095436801298611408202050198891430;
  wire or_not_new_n2818__not_new_n2817_;
  wire not_new_n6242__5;
  wire not_new_n4017_;
  wire not_new_n3320_;
  wire new_n7103_;
  wire not_new_n6974__7;
  wire not_new_n6974__0;
  wire new_n5795_;
  wire new_n9645_;
  wire not_new_n8603_;
  wire not_new_n3372__2326305139872070;
  wire not_new_n4414_;
  wire not_new_n6022_;
  wire not_new_n640__332329305696010;
  wire new_n9060_;
  wire not_pi148_1;
  wire not_new_n1588__1176490;
  wire new_n2837_;
  wire not_pi256;
  wire not_new_n4789__0;
  wire not_new_n6894_;
  wire new_n7689_;
  wire not_new_n9578_;
  wire not_pi037_0;
  wire new_n9193_;
  wire new_n8206_;
  wire not_new_n605__9;
  wire new_n2013_;
  wire not_new_n1588__47475615099430;
  wire new_n5002_;
  wire and_new_n2295__new_n2298_;
  wire new_n2007_;
  wire not_new_n1024_;
  wire not_new_n602__2;
  wire new_n3851_;
  wire not_new_n7773__1;
  wire new_n3272_;
  wire not_new_n9090_;
  wire new_n5850_;
  wire not_new_n9911__0;
  wire not_new_n9836_;
  wire not_new_n8589_;
  wire or_not_new_n2595__not_new_n2594_;
  wire not_new_n4466_;
  wire new_n6379_;
  wire not_new_n5003_;
  wire not_pi146;
  wire not_new_n681__0;
  wire new_n4882_;
  wire not_new_n5899_;
  wire new_n4824_;
  wire po070;
  wire not_new_n1175__0;
  wire not_new_n6302_;
  wire new_n9055_;
  wire new_n8945_;
  wire not_new_n9689_;
  wire new_n3488_;
  wire not_new_n1469_;
  wire new_n5240_;
  wire not_new_n1598__2;
  wire not_pi140_2;
  wire not_new_n600__490;
  wire new_n2280_;
  wire new_n6861_;
  wire new_n10136_;
  wire or_new_n1031__new_n1037_;
  wire not_new_n5203__0;
  wire not_new_n9002_;
  wire not_new_n4290_;
  wire new_n5189_;
  wire new_n3959_;
  wire new_n2274_;
  wire new_n6111_;
  wire not_new_n6411_;
  wire not_pi245_0;
  wire not_new_n600__2824752490;
  wire not_new_n5883_;
  wire not_new_n9583_;
  wire new_n7550_;
  wire not_new_n8562_;
  wire not_new_n9790_;
  wire new_n7862_;
  wire key_gate_75;
  wire not_new_n600__16284135979104490;
  wire not_new_n4506__0;
  wire not_new_n8214_;
  wire not_new_n6032_;
  wire new_n1163_;
  wire new_n1799_;
  wire new_n8886_;
  wire new_n9926_;
  wire not_new_n4562_;
  wire not_new_n2736_;
  wire new_n8938_;
  wire not_new_n5740__1;
  wire not_new_n6192_;
  wire not_new_n3078_;
  wire new_n2787_;
  wire not_new_n5447_;
  wire not_new_n3184__1176490;
  wire new_n8781_;
  wire not_new_n6495_;
  wire new_n5873_;
  wire not_new_n637__9;
  wire not_new_n4448__0;
  wire not_new_n1053__8235430;
  wire new_n3985_;
  wire new_n6995_;
  wire not_new_n2818_;
  wire not_new_n6078_;
  wire and_new_n9888__new_n10254_;
  wire not_new_n5789_;
  wire new_n5949_;
  wire new_n8275_;
  wire new_n6702_;
  wire new_n1311_;
  wire not_new_n5224_;
  wire not_new_n1071__4;
  wire not_new_n602__3;
  wire not_new_n2429_;
  wire not_new_n617__490;
  wire new_n5367_;
  wire new_n3663_;
  wire not_new_n1041__490;
  wire po080;
  wire not_new_n9859_;
  wire not_new_n7509_;
  wire not_new_n7552_;
  wire not_new_n7229_;
  wire and_new_n1310__new_n2179_;
  wire key_gate_36;
  wire not_new_n633__70;
  wire not_pi051_1;
  wire new_n5153_;
  wire new_n5901_;
  wire new_n4265_;
  wire new_n2403_;
  wire not_new_n1581__2;
  wire new_n5108_;
  wire po010;
  wire new_n5679_;
  wire not_new_n10008__0;
  wire not_new_n636__6782230728490;
  wire new_n2102_;
  wire new_n10180_;
  wire new_n2679_;
  wire not_new_n1591__2;
  wire new_n6887_;
  wire not_new_n1047__16284135979104490;
  wire not_new_n2524_;
  wire not_new_n2665_;
  wire not_new_n597__7;
  wire not_new_n4743_;
  wire not_new_n10279_;
  wire not_new_n5964_;
  wire not_new_n633__3;
  wire new_n1942_;
  wire new_n5142_;
  wire new_n4496_;
  wire not_new_n1494_;
  wire not_new_n8203_;
  wire and_new_n9525__new_n9526_;
  wire or_not_new_n6226__not_new_n6323_;
  wire new_n747_;
  wire new_n9177_;
  wire key_gate_3;
  wire not_new_n3696_;
  wire not_new_n8127__0;
  wire not_new_n1028__0;
  wire new_n2231_;
  wire new_n6856_;
  wire not_pi059_0;
  wire not_new_n8904_;
  wire not_new_n975_;
  wire new_n5073_;
  wire not_new_n595__403536070;
  wire not_new_n4727_;
  wire and_new_n1463__new_n1465_;
  wire not_new_n3503_;
  wire not_new_n5348_;
  wire not_new_n581__273687473400809163430;
  wire new_n6889_;
  wire not_new_n1379_;
  wire not_new_n1589__16284135979104490;
  wire new_n6932_;
  wire not_new_n8449_;
  wire new_n9057_;
  wire not_new_n7045_;
  wire new_n3235_;
  wire not_new_n6293_;
  wire not_new_n9533_;
  wire new_n3655_;
  wire new_n3197_;
  wire not_new_n7810_;
  wire not_new_n4151_;
  wire not_new_n9929_;
  wire new_n2914_;
  wire new_n9605_;
  wire not_new_n608__168070;
  wire new_n4482_;
  wire new_n7169_;
  wire new_n7983_;
  wire new_n4349_;
  wire new_n3750_;
  wire new_n4456_;
  wire new_n8735_;
  wire new_n1000_;
  wire not_new_n2170_;
  wire not_new_n9212_;
  wire new_n6994_;
  wire new_n1873_;
  wire new_n3474_;
  wire not_new_n1612__9;
  wire not_new_n3849_;
  wire not_new_n4818__0;
  wire not_new_n2728_;
  wire po170;
  wire not_new_n609__57648010;
  wire not_new_n8776_;
  wire new_n5959_;
  wire not_new_n989__138412872010;
  wire not_new_n643__2824752490;
  wire not_new_n5072_;
  wire new_n3561_;
  wire not_new_n4644_;
  wire new_n4229_;
  wire new_n10299_;
  wire not_new_n4180_;
  wire new_n725_;
  wire not_new_n1598__57648010;
  wire or_not_new_n2955__not_new_n2958_;
  wire and_new_n3049__new_n998_;
  wire new_n8407_;
  wire new_n6005_;
  wire not_new_n10222_;
  wire not_new_n1433_;
  wire not_new_n8568_;
  wire new_n2898_;
  wire new_n4213_;
  wire not_new_n1031__2;
  wire new_n9997_;
  wire new_n7606_;
  wire new_n8644_;
  wire po209;
  wire po243;
  wire not_new_n8178__0;
  wire not_new_n952_;
  wire not_new_n6619_;
  wire new_n2022_;
  wire not_new_n5938_;
  wire new_n7562_;
  wire not_new_n602__70;
  wire new_n4707_;
  wire new_n1635_;
  wire not_pi129_1;
  wire new_n5316_;
  wire new_n4327_;
  wire not_new_n1534__168070;
  wire new_n5910_;
  wire new_n5174_;
  wire new_n671_;
  wire new_n6506_;
  wire not_new_n1596__7;
  wire not_new_n9514_;
  wire not_new_n585__0;
  wire new_n3503_;
  wire not_new_n1049__6782230728490;
  wire not_new_n644__138412872010;
  wire not_new_n6474__1;
  wire not_new_n1580__70;
  wire not_new_n4071__2;
  wire not_new_n6683_;
  wire new_n3046_;
  wire not_new_n9976_;
  wire new_n9963_;
  wire new_n8670_;
  wire not_new_n9363_;
  wire not_new_n3315__5585458640832840070;
  wire not_new_n1049__70;
  wire not_new_n7625__0;
  wire new_n4546_;
  wire not_new_n3844_;
  wire new_n5426_;
  wire not_new_n4123__2;
  wire not_new_n9614__0;
  wire not_new_n4975_;
  wire new_n6271_;
  wire key_gate_56;
  wire new_n6195_;
  wire new_n7068_;
  wire not_new_n5772_;
  wire not_new_n7351_;
  wire new_n9658_;
  wire not_new_n9320_;
  wire new_n6894_;
  wire new_n8913_;
  wire not_new_n6948_;
  wire new_n9371_;
  wire not_new_n5801__0;
  wire new_n7969_;
  wire new_n2085_;
  wire not_pi256_0;
  wire not_new_n1781__0;
  wire not_new_n3252_;
  wire not_pi211;
  wire new_n1626_;
  wire not_new_n6985_;
  wire not_new_n1277_;
  wire not_new_n7374_;
  wire new_n4048_;
  wire not_new_n9032_;
  wire new_n1557_;
  wire new_n2293_;
  wire not_new_n6809_;
  wire new_n1530_;
  wire new_n7907_;
  wire not_new_n7636_;
  wire not_new_n3259_;
  wire new_n3274_;
  wire not_new_n639__797922662976120010;
  wire or_or_not_new_n2300__not_new_n2301__not_new_n2303_;
  wire new_n1857_;
  wire new_n707_;
  wire new_n7605_;
  wire new_n6633_;
  wire new_n8792_;
  wire not_new_n2009_;
  wire new_n1219_;
  wire not_new_n8465_;
  wire new_n9062_;
  wire new_n5570_;
  wire new_n2026_;
  wire not_pi133_1;
  wire not_new_n1165__0;
  wire new_n4708_;
  wire new_n3904_;
  wire not_new_n9493_;
  wire new_n9832_;
  wire not_new_n1035__6;
  wire not_new_n611__1;
  wire not_new_n1003__3;
  wire new_n8280_;
  wire new_n9402_;
  wire new_n2536_;
  wire new_n2379_;
  wire new_n9455_;
  wire not_new_n4625_;
  wire new_n8996_;
  wire not_new_n3865_;
  wire new_n3609_;
  wire new_n10107_;
  wire not_new_n5466_;
  wire not_new_n7606__1;
  wire not_new_n8257_;
  wire new_n9411_;
  wire not_new_n1596__1;
  wire new_n6989_;
  wire new_n7285_;
  wire new_n4874_;
  wire not_new_n4207_;
  wire not_new_n2261__0;
  wire not_new_n1051__1176490;
  wire new_n8368_;
  wire not_new_n7654_;
  wire new_n9918_;
  wire not_new_n1521_;
  wire not_new_n8112_;
  wire not_new_n3954_;
  wire not_new_n611__70;
  wire not_new_n1584__332329305696010;
  wire and_and_new_n4295__new_n4334__new_n4338_;
  wire or_not_new_n2319__not_new_n2320_;
  wire not_new_n995_;
  wire not_new_n1538__1176490;
  wire new_n7193_;
  wire not_new_n775__0;
  wire not_new_n7349_;
  wire not_new_n3889_;
  wire not_new_n8878_;
  wire not_new_n4659_;
  wire new_n4227_;
  wire new_n7291_;
  wire not_new_n6693_;
  wire new_n1966_;
  wire new_n8424_;
  wire not_new_n1572_;
  wire not_new_n1583__24010;
  wire not_new_n6342_;
  wire new_n7073_;
  wire and_new_n6378__new_n6379_;
  wire not_new_n645__3430;
  wire not_new_n9760_;
  wire not_new_n1392_;
  wire new_n8303_;
  wire not_new_n3372__332329305696010;
  wire not_new_n2283_;
  wire new_n6488_;
  wire new_n3395_;
  wire new_n1715_;
  wire not_new_n7622__1;
  wire new_n7913_;
  wire new_n2257_;
  wire po077;
  wire not_new_n9426__1;
  wire not_new_n1071__1;
  wire not_new_n7625_;
  wire not_new_n1002__2;
  wire new_n4551_;
  wire not_new_n5794_;
  wire not_new_n3086_;
  wire not_new_n591__6782230728490;
  wire not_new_n928__1176490;
  wire new_n3379_;
  wire not_new_n8540_;
  wire not_new_n1607__8;
  wire not_new_n2617_;
  wire not_new_n6029_;
  wire new_n5259_;
  wire not_new_n5747__0;
  wire not_po296_881247870897231951843937366879128181133112010;
  wire not_new_n1627_;
  wire not_pi160;
  wire not_new_n7176_;
  wire not_new_n6485_;
  wire not_new_n9777_;
  wire new_n5563_;
  wire not_new_n5130_;
  wire or_not_new_n8781__not_new_n8701_;
  wire not_pi265_2;
  wire not_new_n1597__24010;
  wire not_new_n581__13410686196639649008070;
  wire not_new_n6098_;
  wire not_new_n10016__1;
  wire not_new_n624__3430;
  wire new_n1065_;
  wire not_new_n3848_;
  wire not_new_n2172_;
  wire new_n6954_;
  wire new_n8852_;
  wire new_n3246_;
  wire not_new_n3315__490;
  wire not_pi259_1;
  wire not_new_n4500_;
  wire not_new_n4836_;
  wire not_new_n1603__332329305696010;
  wire new_n4128_;
  wire not_new_n585__2824752490;
  wire and_and_new_n1934__new_n1937__new_n1935_;
  wire not_new_n4590_;
  wire not_new_n596__2824752490;
  wire new_n603_;
  wire not_new_n9373__2;
  wire new_n3359_;
  wire new_n5841_;
  wire not_new_n8195_;
  wire not_new_n5500__0;
  wire not_new_n7712_;
  wire new_n730_;
  wire new_n1911_;
  wire not_new_n626__7;
  wire not_new_n5921__0;
  wire new_n1965_;
  wire not_new_n1053__138412872010;
  wire new_n4573_;
  wire new_n4475_;
  wire not_new_n4467_;
  wire not_new_n1206_;
  wire not_new_n6473_;
  wire not_pi041_1;
  wire not_new_n3191_;
  wire new_n713_;
  wire not_new_n9405_;
  wire po098;
  wire not_new_n6172_;
  wire not_new_n633__2326305139872070;
  wire not_new_n9723_;
  wire not_new_n9637__0;
  wire new_n5967_;
  wire not_new_n7050_;
  wire not_new_n3311__8;
  wire not_new_n4944_;
  wire not_pi173_1;
  wire new_n7485_;
  wire new_n6918_;
  wire not_new_n971_;
  wire not_new_n6489__0;
  wire key_gate_42;
  wire not_new_n3433_;
  wire new_n10328_;
  wire or_or_not_new_n8833__not_new_n8830__0_not_new_n9222_;
  wire new_n4899_;
  wire not_pi122_0;
  wire not_new_n8661_;
  wire new_n9409_;
  wire new_n5552_;
  wire new_n1776_;
  wire not_new_n589__2824752490;
  wire new_n7072_;
  wire new_n6182_;
  wire not_new_n939_;
  wire new_n6726_;
  wire po052;
  wire or_not_new_n10126__not_new_n10125_;
  wire not_new_n4504_;
  wire not_new_n4947_;
  wire not_pi203;
  wire not_new_n640__3;
  wire not_new_n586__3;
  wire not_new_n1809_;
  wire new_n3365_;
  wire not_new_n1585__4;
  wire not_new_n9316_;
  wire not_new_n638__57648010;
  wire not_new_n7665_;
  wire not_new_n6138_;
  wire new_n8606_;
  wire not_new_n648__168070;
  wire not_new_n609__3;
  wire not_new_n1027__47475615099430;
  wire new_n6620_;
  wire not_pi147_0;
  wire not_new_n1607__9;
  wire new_n5205_;
  wire new_n10082_;
  wire not_new_n6974__57648010;
  wire new_n6890_;
  wire not_new_n1496_;
  wire new_n8389_;
  wire not_new_n1255_;
  wire not_new_n10028_;
  wire new_n5611_;
  wire not_new_n1584__138412872010;
  wire not_new_n5625_;
  wire new_n772_;
  wire new_n9885_;
  wire not_new_n4131__2;
  wire new_n1762_;
  wire not_new_n8802_;
  wire not_new_n7593_;
  wire new_n8773_;
  wire not_new_n7573_;
  wire not_new_n5751_;
  wire new_n9003_;
  wire new_n10125_;
  wire or_not_new_n2910__not_new_n2913_;
  wire new_n6815_;
  wire not_new_n994__403536070;
  wire not_new_n1193_;
  wire new_n10236_;
  wire or_not_new_n3176__not_new_n3175_;
  wire or_not_new_n2758__not_new_n2761_;
  wire new_n4488_;
  wire or_or_not_new_n1901__not_new_n1902__not_new_n1904_;
  wire new_n7495_;
  wire new_n3969_;
  wire not_new_n3424_;
  wire not_new_n2280__0;
  wire not_new_n4522_;
  wire new_n2138_;
  wire new_n7709_;
  wire new_n5870_;
  wire not_new_n7565_;
  wire new_n5019_;
  wire and_and_new_n6365__new_n6439__new_n6438_;
  wire not_pi271_1;
  wire new_n1071_;
  wire not_new_n4281_;
  wire not_new_n627__19773267430;
  wire new_n4796_;
  wire new_n7268_;
  wire not_new_n4999_;
  wire new_n2655_;
  wire new_n4114_;
  wire new_n1373_;
  wire new_n1657_;
  wire new_n8577_;
  wire po279;
  wire new_n10040_;
  wire new_n9699_;
  wire new_n1169_;
  wire new_n7469_;
  wire new_n4835_;
  wire not_new_n6625__0;
  wire not_new_n972_;
  wire not_new_n3159_;
  wire not_new_n1591__2326305139872070;
  wire or_or_not_new_n4228__not_new_n4329__not_new_n710_;
  wire not_new_n599__490;
  wire or_not_new_n3158__not_new_n3157_;
  wire not_new_n771_;
  wire not_new_n1047__5;
  wire not_new_n9164_;
  wire not_new_n6710_;
  wire not_new_n7742_;
  wire new_n1861_;
  wire not_new_n5468__0;
  wire new_n4886_;
  wire new_n7116_;
  wire not_new_n1602__797922662976120010;
  wire new_n3475_;
  wire not_new_n7048_;
  wire new_n5497_;
  wire not_new_n1728__19773267430;
  wire new_n8045_;
  wire new_n7905_;
  wire new_n3784_;
  wire po179;
  wire new_n9622_;
  wire new_n4072_;
  wire not_new_n10264_;
  wire not_new_n7652_;
  wire new_n8259_;
  wire not_new_n1728__70;
  wire and_and_not_pi037_2_not_pi036_2_not_pi039_3;
  wire not_new_n5480__0;
  wire not_new_n639__16284135979104490;
  wire new_n9097_;
  wire not_po296_26517308458596534717790233816010;
  wire new_n6953_;
  wire new_n5866_;
  wire new_n2180_;
  wire new_n8265_;
  wire not_new_n622__8;
  wire not_new_n7935_;
  wire not_new_n8285_;
  wire not_new_n1053__168070;
  wire new_n4582_;
  wire new_n5165_;
  wire new_n3596_;
  wire not_new_n7373_;
  wire not_new_n4720_;
  wire new_n1593_;
  wire new_n6038_;
  wire not_new_n3314_;
  wire not_new_n7037_;
  wire new_n3310_;
  wire not_new_n4123__1;
  wire not_new_n1785_;
  wire not_new_n5674__1;
  wire not_new_n9214_;
  wire not_new_n6884_;
  wire not_pi273_0;
  wire not_new_n7726_;
  wire new_n1164_;
  wire not_pi149;
  wire not_new_n5791_;
  wire not_new_n2716_;
  wire not_new_n9682_;
  wire not_new_n8537_;
  wire or_not_new_n2718__not_new_n2717_;
  wire not_new_n641__1176490;
  wire not_new_n9698_;
  wire not_new_n6922_;
  wire new_n2733_;
  wire not_new_n984__332329305696010;
  wire new_n6800_;
  wire new_n4122_;
  wire new_n9078_;
  wire new_n6760_;
  wire not_new_n994__6782230728490;
  wire not_new_n666_;
  wire not_new_n7016_;
  wire or_not_new_n2246__not_new_n2243_;
  wire new_n9483_;
  wire not_new_n8482_;
  wire not_new_n1289_;
  wire new_n5473_;
  wire new_n2030_;
  wire not_pi111_0;
  wire new_n1467_;
  wire new_n4989_;
  wire new_n9240_;
  wire new_n3782_;
  wire not_new_n1063__9;
  wire new_n9532_;
  wire not_new_n1395_;
  wire not_new_n7036__1;
  wire not_new_n1613__168070;
  wire new_n7418_;
  wire not_new_n625__5585458640832840070;
  wire not_pi261_0;
  wire new_n7091_;
  wire not_new_n9163_;
  wire not_new_n8684_;
  wire not_new_n2616_;
  wire not_new_n4017__1;
  wire new_n7330_;
  wire new_n3755_;
  wire new_n7425_;
  wire not_new_n3566_;
  wire not_new_n9441_;
  wire new_n4134_;
  wire not_new_n6737__0;
  wire new_n6981_;
  wire new_n2058_;
  wire or_not_new_n3116__not_new_n3115_;
  wire not_new_n1002__7;
  wire new_n1233_;
  wire not_new_n6443__57648010;
  wire new_n4567_;
  wire new_n1548_;
  wire new_n3256_;
  wire new_n2289_;
  wire new_n2603_;
  wire not_new_n634__3430;
  wire new_n9119_;
  wire not_new_n7221_;
  wire new_n8352_;
  wire not_new_n2587_;
  wire not_new_n10000_;
  wire not_pi017;
  wire not_new_n4974_;
  wire new_n8071_;
  wire new_n7591_;
  wire not_new_n5748__1;
  wire not_new_n7568_;
  wire not_new_n7137_;
  wire not_new_n5491_;
  wire not_new_n1051__24010;
  wire not_new_n7360__0;
  wire not_new_n6176_;
  wire not_new_n4095_;
  wire not_new_n8867_;
  wire not_new_n5036_;
  wire po013;
  wire not_new_n5670_;
  wire not_new_n7297_;
  wire new_n2759_;
  wire not_new_n3952_;
  wire not_new_n7291_;
  wire new_n7223_;
  wire not_new_n4302_;
  wire new_n1189_;
  wire new_n2994_;
  wire not_new_n588__3430;
  wire not_new_n3415_;
  wire not_new_n9651_;
  wire not_new_n8448_;
  wire new_n6246_;
  wire not_new_n4938__0;
  wire not_new_n5761_;
  wire not_new_n9453_;
  wire new_n7638_;
  wire not_new_n9496_;
  wire new_n3775_;
  wire new_n9072_;
  wire not_new_n9660_;
  wire not_new_n7158_;
  wire not_new_n6977_;
  wire not_new_n1197_;
  wire not_new_n626__8;
  wire new_n682_;
  wire not_new_n5512_;
  wire not_new_n1598__168070;
  wire not_new_n4834_;
  wire not_new_n9980_;
  wire not_new_n6076_;
  wire new_n6533_;
  wire not_new_n8170__1;
  wire not_new_n7880_;
  wire not_new_n9445_;
  wire not_new_n3717_;
  wire not_new_n3372__1;
  wire not_new_n622__6782230728490;
  wire not_new_n2839_;
  wire new_n3127_;
  wire and_new_n4337__new_n4336_;
  wire not_new_n3104_;
  wire new_n3280_;
  wire not_new_n593__5;
  wire not_new_n7136_;
  wire not_new_n9222_;
  wire not_new_n1023__2;
  wire not_new_n3372__2;
  wire not_new_n7295_;
  wire new_n1556_;
  wire new_n8315_;
  wire not_new_n10165__0;
  wire not_new_n591__1176490;
  wire new_n7097_;
  wire not_pi257_1;
  wire not_new_n3668_;
  wire new_n9791_;
  wire new_n7369_;
  wire not_new_n6552_;
  wire not_new_n1602__47475615099430;
  wire new_n1826_;
  wire not_new_n610_;
  wire not_new_n1902_;
  wire not_new_n3476_;
  wire new_n638_;
  wire po221;
  wire not_new_n3788_;
  wire not_new_n708_;
  wire new_n2288_;
  wire not_new_n608__8235430;
  wire new_n4860_;
  wire not_new_n6472_;
  wire not_new_n8673_;
  wire not_new_n1045__57648010;
  wire new_n7670_;
  wire not_new_n631__7;
  wire not_new_n7025_;
  wire not_new_n1607__1;
  wire not_new_n1043__1;
  wire not_new_n1588__5;
  wire not_new_n1576__2;
  wire new_n9065_;
  wire not_pi040_4;
  wire not_new_n9377_;
  wire new_n1495_;
  wire not_new_n5940_;
  wire not_new_n1597__39098210485829880490;
  wire not_new_n4127__2;
  wire new_n5432_;
  wire new_n1437_;
  wire not_new_n5444_;
  wire not_new_n1043__968890104070;
  wire not_new_n2918_;
  wire not_pi172;
  wire new_n7563_;
  wire new_n7980_;
  wire not_new_n1601__3430;
  wire not_new_n581__113988951853731430;
  wire not_new_n4684_;
  wire not_new_n5900_;
  wire not_new_n5971_;
  wire not_new_n9011__0;
  wire new_n4054_;
  wire not_new_n6650_;
  wire new_n6975_;
  wire new_n4016_;
  wire new_n2721_;
  wire new_n5623_;
  wire new_n9784_;
  wire not_new_n1346_;
  wire not_new_n648__138412872010;
  wire not_new_n593__57648010;
  wire new_n1831_;
  wire new_n2661_;
  wire or_not_new_n618__19773267430_not_new_n6865_;
  wire not_pi255_2;
  wire not_new_n6494_;
  wire new_n2547_;
  wire not_new_n2014__0;
  wire not_new_n630__5585458640832840070;
  wire not_new_n1728__6;
  wire new_n3427_;
  wire new_n1503_;
  wire new_n9781_;
  wire new_n2127_;
  wire not_new_n7855__0;
  wire new_n3943_;
  wire new_n7995_;
  wire po203;
  wire not_new_n7676_;
  wire not_new_n585__47475615099430;
  wire not_new_n8843_;
  wire not_new_n7168_;
  wire new_n10000_;
  wire not_new_n1616__1176490;
  wire new_n6176_;
  wire not_new_n2673_;
  wire not_new_n2706_;
  wire not_new_n7932_;
  wire new_n8338_;
  wire not_new_n6304_;
  wire new_n2060_;
  wire not_new_n1172_;
  wire new_n2666_;
  wire not_new_n1613__1176490;
  wire new_n2924_;
  wire not_new_n585_;
  wire new_n3696_;
  wire new_n3443_;
  wire new_n8024_;
  wire not_new_n4299_;
  wire not_new_n9154_;
  wire new_n7484_;
  wire new_n8262_;
  wire not_new_n994__968890104070;
  wire not_new_n5438_;
  wire not_new_n5518_;
  wire and_new_n2374__new_n2373_;
  wire not_new_n9427__2;
  wire not_po298_24010;
  wire not_pi049_2;
  wire new_n3961_;
  wire key_gate_127;
  wire not_new_n5418_;
  wire new_n3381_;
  wire new_n6276_;
  wire new_n4418_;
  wire new_n1349_;
  wire po190;
  wire new_n7247_;
  wire new_n4695_;
  wire new_n4894_;
  wire new_n2282_;
  wire not_new_n2489_;
  wire not_new_n936_;
  wire new_n5578_;
  wire not_new_n5745_;
  wire new_n9767_;
  wire not_new_n1544_;
  wire not_new_n1039__3430;
  wire new_n5452_;
  wire new_n7059_;
  wire not_new_n4131__1;
  wire not_new_n4182_;
  wire not_new_n8244__1;
  wire new_n1415_;
  wire not_new_n1053__9;
  wire po044;
  wire not_new_n643__5;
  wire new_n10242_;
  wire new_n6869_;
  wire not_new_n3692_;
  wire not_new_n10025_;
  wire new_n9771_;
  wire new_n9847_;
  wire not_new_n8082__0;
  wire not_pi189_0;
  wire new_n680_;
  wire not_new_n9435_;
  wire not_new_n5164_;
  wire new_n8170_;
  wire new_n5682_;
  wire not_new_n619__138412872010;
  wire new_n4298_;
  wire not_new_n6155_;
  wire new_n2767_;
  wire new_n4196_;
  wire new_n5109_;
  wire new_n9726_;
  wire new_n6148_;
  wire not_new_n1049__168070;
  wire or_or_not_new_n1552__not_new_n2419__not_new_n1373_;
  wire new_n597_;
  wire not_new_n1631__19773267430;
  wire not_new_n927__1;
  wire new_n4220_;
  wire not_new_n593__332329305696010;
  wire not_new_n8282__0;
  wire not_pi044_2;
  wire not_new_n2206_;
  wire not_new_n3921_;
  wire not_new_n593__4;
  wire new_n8082_;
  wire not_new_n613__7;
  wire not_new_n594__490;
  wire not_new_n594__332329305696010;
  wire new_n4915_;
  wire new_n10257_;
  wire new_n6432_;
  wire new_n8701_;
  wire or_not_new_n2982__not_new_n2985_;
  wire or_not_new_n2899__not_new_n2898_;
  wire new_n3687_;
  wire not_new_n930_;
  wire not_new_n5624_;
  wire new_n1547_;
  wire not_new_n602__2824752490;
  wire po083;
  wire not_new_n618__797922662976120010;
  wire not_new_n6105_;
  wire new_n6040_;
  wire not_new_n3318__1;
  wire new_n7055_;
  wire not_pi181;
  wire not_new_n4955__0;
  wire not_new_n1581__7;
  wire not_new_n6504_;
  wire not_new_n6079_;
  wire new_n6375_;
  wire not_new_n2844_;
  wire not_new_n1536__332329305696010;
  wire not_new_n7359_;
  wire not_new_n3315__2;
  wire new_n4850_;
  wire not_new_n1482_;
  wire new_n4701_;
  wire not_new_n645__8;
  wire not_new_n639__2326305139872070;
  wire new_n9265_;
  wire not_new_n9849_;
  wire not_new_n6493_;
  wire not_new_n1069__8235430;
  wire not_new_n7241_;
  wire new_n1181_;
  wire or_or_not_new_n1558__not_new_n2449__not_new_n1385_;
  wire new_n8258_;
  wire new_n3647_;
  wire new_n4059_;
  wire not_new_n9491__0;
  wire key_gate_112;
  wire new_n3661_;
  wire not_new_n7378_;
  wire not_new_n9864_;
  wire not_new_n601__2824752490;
  wire not_new_n1534__1;
  wire new_n4652_;
  wire new_n6846_;
  wire and_new_n10212__new_n10211_;
  wire new_n755_;
  wire or_or_not_new_n1319__not_new_n1317__not_new_n2211_;
  wire new_n3448_;
  wire and_new_n8667__new_n8666_;
  wire not_new_n1534__2824752490;
  wire not_new_n9524__0;
  wire not_new_n6516__0;
  wire not_new_n5462__0;
  wire new_n1165_;
  wire new_n1329_;
  wire new_n7167_;
  wire new_n1656_;
  wire not_pi103;
  wire not_new_n7610__0;
  wire new_n7399_;
  wire not_new_n5688_;
  wire not_new_n631__57648010;
  wire not_new_n7021__1;
  wire new_n2173_;
  wire not_new_n2872_;
  wire not_pi087;
  wire not_new_n1020__4;
  wire new_n8214_;
  wire not_new_n5040_;
  wire new_n8576_;
  wire not_new_n1055__3430;
  wire not_new_n644__0;
  wire not_new_n7614_;
  wire and_new_n2389__new_n2388_;
  wire not_new_n613__0;
  wire not_new_n8978__3;
  wire not_new_n6625__1;
  wire not_new_n5291_;
  wire not_new_n1018__5;
  wire new_n2553_;
  wire new_n1323_;
  wire new_n10096_;
  wire not_new_n969_;
  wire or_or_or_not_new_n2928__not_new_n2931__not_new_n2930__not_new_n2932_;
  wire not_new_n606__3;
  wire not_new_n9155_;
  wire not_new_n9476_;
  wire not_new_n7026__0;
  wire new_n3244_;
  wire not_new_n9625_;
  wire not_new_n8314_;
  wire new_n8898_;
  wire new_n9026_;
  wire new_n1836_;
  wire new_n1946_;
  wire not_new_n2509_;
  wire new_n6763_;
  wire not_new_n5993_;
  wire not_new_n1631__490;
  wire or_not_new_n2803__not_new_n2806_;
  wire not_new_n4766__0;
  wire not_new_n6151_;
  wire new_n8160_;
  wire new_n9205_;
  wire and_new_n1234__new_n1818_;
  wire not_new_n8162_;
  wire not_new_n2927_;
  wire not_new_n1065__2326305139872070;
  wire new_n6263_;
  wire new_n1824_;
  wire not_new_n588__8;
  wire or_not_new_n6538__1_not_new_n6877_;
  wire new_n8188_;
  wire not_new_n7727_;
  wire not_new_n5884_;
  wire new_n8753_;
  wire not_new_n7757_;
  wire not_new_n9939_;
  wire not_new_n1471_;
  wire not_new_n646__6782230728490;
  wire not_new_n927__0;
  wire new_n9373_;
  wire not_new_n1055__168070;
  wire not_new_n5361_;
  wire new_n6498_;
  wire new_n7477_;
  wire new_n5703_;
  wire new_n4449_;
  wire not_new_n8044_;
  wire not_pi107_0;
  wire new_n5458_;
  wire not_pi185_0;
  wire not_new_n2464_;
  wire not_new_n1061__5;
  wire not_new_n7043__1;
  wire not_new_n3892_;
  wire not_new_n7631__0;
  wire not_new_n7604_;
  wire not_new_n6626_;
  wire not_new_n9875__0;
  wire new_n2630_;
  wire not_new_n5540_;
  wire new_n4435_;
  wire not_new_n1596__5585458640832840070;
  wire not_new_n587__70;
  wire new_n4692_;
  wire new_n1992_;
  wire not_new_n1065__5;
  wire not_new_n7886_;
  wire not_new_n3207_;
  wire new_n8435_;
  wire new_n2417_;
  wire not_new_n9415__0;
  wire not_new_n605__5;
  wire new_n5530_;
  wire not_new_n608__5;
  wire not_new_n8832_;
  wire not_new_n9118_;
  wire new_n7906_;
  wire not_new_n8128__0;
  wire not_new_n6971_;
  wire new_n6291_;
  wire not_new_n10012_;
  wire new_n4238_;
  wire not_new_n1607__4;
  wire not_new_n7014_;
  wire not_new_n617__2824752490;
  wire new_n1229_;
  wire and_new_n1294__new_n2103_;
  wire not_new_n4418__0;
  wire not_new_n5467_;
  wire new_n9256_;
  wire not_new_n4167_;
  wire new_n6062_;
  wire not_new_n8698_;
  wire new_n4841_;
  wire or_not_new_n6373__9_not_new_n6237_;
  wire not_new_n4626_;
  wire new_n4784_;
  wire not_new_n586__168070;
  wire not_new_n6988__0;
  wire not_new_n8651_;
  wire new_n8020_;
  wire not_new_n7083_;
  wire not_new_n7887__0;
  wire new_n7707_;
  wire not_new_n984__113988951853731430;
  wire new_n8147_;
  wire not_new_n6122_;
  wire not_new_n8402_;
  wire key_gate_113;
  wire not_new_n1063__3;
  wire new_n2118_;
  wire new_n4921_;
  wire not_new_n636__0;
  wire new_n2150_;
  wire new_n9001_;
  wire not_new_n5810_;
  wire new_n4288_;
  wire new_n5556_;
  wire not_new_n617__2;
  wire new_n5350_;
  wire not_new_n2576_;
  wire new_n6697_;
  wire po183;
  wire not_new_n629__113988951853731430;
  wire not_new_n4557_;
  wire not_new_n927_;
  wire new_n7387_;
  wire not_new_n4794_;
  wire not_new_n628__10;
  wire new_n5008_;
  wire new_n2520_;
  wire not_new_n6560_;
  wire not_new_n10034_;
  wire not_new_n7954_;
  wire new_n3922_;
  wire new_n3183_;
  wire not_new_n7770__0;
  wire new_n7962_;
  wire not_new_n10052__0;
  wire not_new_n3981__0;
  wire new_n630_;
  wire new_n1622_;
  wire new_n8461_;
  wire po284;
  wire not_new_n601__19773267430;
  wire new_n2783_;
  wire new_n4998_;
  wire not_new_n589__3788186922656647816827176259430;
  wire not_new_n598__332329305696010;
  wire not_new_n7621_;
  wire new_n9727_;
  wire new_n2944_;
  wire new_n8228_;
  wire new_n3858_;
  wire new_n8658_;
  wire not_new_n5798_;
  wire not_new_n7239_;
  wire new_n1735_;
  wire not_new_n6343_;
  wire new_n6858_;
  wire not_new_n7750__0;
  wire not_new_n9714__0;
  wire not_new_n641__490;
  wire not_new_n3969_;
  wire new_n6262_;
  wire not_new_n5718_;
  wire not_new_n632__3430;
  wire not_new_n7586_;
  wire not_new_n7745_;
  wire not_new_n9686_;
  wire new_n920_;
  wire not_new_n8900_;
  wire new_n4504_;
  wire new_n9161_;
  wire new_n1998_;
  wire not_new_n9677_;
  wire not_new_n610__3;
  wire new_n5196_;
  wire not_pi262_1;
  wire new_n5166_;
  wire not_new_n9918__0;
  wire not_new_n9185_;
  wire new_n6529_;
  wire new_n6284_;
  wire not_new_n6064__0;
  wire not_new_n1049__9;
  wire not_new_n6817_;
  wire not_new_n5720_;
  wire not_new_n3192_;
  wire new_n7743_;
  wire not_new_n1589__10;
  wire or_not_new_n3944__not_new_n3914__1;
  wire not_new_n640__9;
  wire not_new_n3112_;
  wire new_n4673_;
  wire not_new_n9306_;
  wire new_n5688_;
  wire not_new_n3310__490;
  wire or_not_new_n10210__not_new_n10153_;
  wire not_new_n3408_;
  wire not_new_n984__2;
  wire not_new_n585__16284135979104490;
  wire new_n10027_;
  wire not_new_n631__273687473400809163430;
  wire new_n4656_;
  wire not_po298_332329305696010;
  wire not_new_n1577_;
  wire not_new_n5909_;
  wire new_n7788_;
  wire new_n3535_;
  wire new_n9018_;
  wire new_n2545_;
  wire not_new_n1580__968890104070;
  wire not_new_n8987__0;
  wire not_new_n1576__332329305696010;
  wire not_pi245;
  wire new_n9063_;
  wire not_new_n6863_;
  wire new_n8190_;
  wire new_n1425_;
  wire new_n7640_;
  wire not_new_n1474_;
  wire new_n3957_;
  wire new_n8035_;
  wire not_po296_248930711762415449007872216849586085868492917169640490;
  wire not_new_n1591__138412872010;
  wire new_n3689_;
  wire not_new_n8169__1;
  wire new_n2821_;
  wire new_n5218_;
  wire new_n7254_;
  wire not_new_n8806_;
  wire not_po296_725745515342319093317411710931737859674906464051430;
  wire not_new_n5754_;
  wire not_new_n5845_;
  wire not_new_n5173_;
  wire new_n9540_;
  wire new_n2488_;
  wire new_n981_;
  wire not_new_n7118_;
  wire not_new_n5366_;
  wire new_n3169_;
  wire not_new_n8380_;
  wire new_n7535_;
  wire not_new_n4898__2;
  wire new_n6906_;
  wire not_new_n7262_;
  wire new_n3043_;
  wire not_new_n8715_;
  wire not_new_n5805_;
  wire new_n7514_;
  wire new_n6475_;
  wire new_n3947_;
  wire not_new_n8253_;
  wire not_new_n635__16284135979104490;
  wire new_n4153_;
  wire not_new_n4766_;
  wire new_n1517_;
  wire new_n7848_;
  wire not_new_n989__968890104070;
  wire new_n2627_;
  wire not_new_n625__47475615099430;
  wire new_n10014_;
  wire new_n3016_;
  wire new_n4000_;
  wire new_n5918_;
  wire new_n2854_;
  wire new_n4884_;
  wire not_new_n4708_;
  wire new_n6674_;
  wire new_n7748_;
  wire not_new_n585__3430;
  wire not_new_n7156_;
  wire new_n5540_;
  wire new_n1400_;
  wire not_new_n6770_;
  wire new_n3593_;
  wire not_new_n1473_;
  wire new_n9406_;
  wire not_new_n624__8235430;
  wire and_and_new_n2067__new_n2070__new_n2068_;
  wire not_new_n692_;
  wire not_new_n8409_;
  wire not_pi272_1;
  wire new_n9079_;
  wire not_new_n7633_;
  wire not_new_n8034_;
  wire not_new_n5081_;
  wire new_n3319_;
  wire not_new_n7464_;
  wire new_n8811_;
  wire not_new_n4736_;
  wire not_new_n629__2824752490;
  wire new_n9413_;
  wire new_n9632_;
  wire new_n4684_;
  wire not_new_n589__1915812313805664144010;
  wire not_new_n5864_;
  wire new_n3324_;
  wire not_new_n609__70;
  wire not_new_n4390_;
  wire not_new_n1591__403536070;
  wire new_n5096_;
  wire not_new_n7260_;
  wire not_new_n2875_;
  wire not_new_n8821_;
  wire not_new_n646__70;
  wire new_n8051_;
  wire not_new_n9883_;
  wire not_new_n9872_;
  wire or_not_new_n1996__not_new_n1997_;
  wire new_n6623_;
  wire key_gate_33;
  wire new_n3271_;
  wire new_n4439_;
  wire new_n4338_;
  wire new_n4402_;
  wire not_new_n3375__4;
  wire not_new_n619__0;
  wire not_new_n1035__0;
  wire new_n3115_;
  wire new_n4413_;
  wire new_n7827_;
  wire new_n1737_;
  wire not_new_n4750__0;
  wire new_n4062_;
  wire new_n4949_;
  wire new_n2313_;
  wire new_n7517_;
  wire new_n10026_;
  wire not_new_n8955_;
  wire not_new_n8262__1;
  wire new_n8851_;
  wire not_new_n9111_;
  wire new_n2121_;
  wire not_pi037_2;
  wire and_new_n4298__new_n4341_;
  wire new_n1376_;
  wire and_new_n4327__new_n4331_;
  wire not_new_n639_;
  wire new_n7545_;
  wire new_n7611_;
  wire not_new_n5241_;
  wire not_new_n5853_;
  wire not_pi266_2;
  wire or_not_new_n999__1_not_new_n3377_;
  wire new_n7147_;
  wire not_new_n606__1176490;
  wire new_n1271_;
  wire new_n3242_;
  wire or_or_or_not_new_n2973__not_new_n2976__not_new_n2975__not_new_n2977_;
  wire not_new_n605__70;
  wire new_n9015_;
  wire not_new_n625__968890104070;
  wire not_new_n1591__4;
  wire new_n4786_;
  wire not_new_n5223_;
  wire not_new_n8595__2;
  wire new_n6142_;
  wire not_pi096;
  wire not_pi064_9;
  wire new_n4039_;
  wire new_n9927_;
  wire not_new_n581__63668057609090279857414351392240010;
  wire new_n5966_;
  wire not_new_n8833_;
  wire new_n10061_;
  wire new_n9499_;
  wire not_new_n7639__0;
  wire not_new_n6023__0;
  wire new_n9783_;
  wire not_new_n4329_;
  wire not_new_n7649_;
  wire not_new_n1606__3;
  wire not_new_n6606_;
  wire new_n2193_;
  wire or_or_not_new_n1235__not_new_n1233__not_new_n1812_;
  wire not_new_n5542_;
  wire not_new_n1612__19773267430;
  wire not_new_n1584__57648010;
  wire and_new_n2010__new_n2013_;
  wire not_new_n4249_;
  wire not_new_n637__113988951853731430;
  wire not_new_n1043__403536070;
  wire not_new_n617__10;
  wire not_new_n1602__968890104070;
  wire not_new_n4363_;
  wire not_new_n9519__0;
  wire not_new_n1004__4;
  wire new_n8652_;
  wire new_n6461_;
  wire not_new_n3311__1176490;
  wire not_new_n5574_;
  wire not_new_n4605_;
  wire not_new_n5080_;
  wire new_n8882_;
  wire not_new_n1067__8235430;
  wire not_pi049_3;
  wire not_new_n4483_;
  wire not_new_n6174_;
  wire not_new_n6949_;
  wire not_po296_490;
  wire not_new_n9702_;
  wire not_new_n5866_;
  wire new_n6335_;
  wire not_new_n8002_;
  wire not_new_n7959_;
  wire new_n2232_;
  wire not_new_n3914_;
  wire not_new_n6976__2;
  wire not_new_n3740_;
  wire not_new_n597__6782230728490;
  wire new_n6141_;
  wire key_gate_123;
  wire not_new_n5216_;
  wire new_n10123_;
  wire not_po298_113988951853731430;
  wire not_new_n6974__24010;
  wire not_pi265_4;
  wire not_new_n5489_;
  wire not_new_n4322_;
  wire not_new_n3911_;
  wire not_new_n7334_;
  wire not_new_n6553_;
  wire not_new_n4086_;
  wire not_new_n6897_;
  wire new_n1368_;
  wire new_n6133_;
  wire not_new_n7104_;
  wire not_new_n3373_;
  wire not_new_n5171_;
  wire not_new_n5178_;
  wire not_new_n1537__9;
  wire new_n3135_;
  wire not_pi163_2;
  wire not_new_n2595_;
  wire new_n4531_;
  wire not_new_n9463_;
  wire not_new_n744__1;
  wire not_pi064_490;
  wire not_new_n9234_;
  wire not_new_n3313_;
  wire new_n8984_;
  wire new_n5328_;
  wire new_n2070_;
  wire not_new_n1065__490;
  wire and_new_n5582__new_n5648_;
  wire not_new_n7961_;
  wire not_new_n8248__1;
  wire not_new_n9989_;
  wire not_new_n994__1176490;
  wire not_new_n635__9;
  wire new_n1904_;
  wire new_n2815_;
  wire not_pi092;
  wire not_new_n8995_;
  wire not_new_n591__138412872010;
  wire not_new_n4465__0;
  wire not_new_n630__8;
  wire new_n9503_;
  wire not_new_n2883_;
  wire not_new_n9140__0;
  wire new_n3836_;
  wire new_n7269_;
  wire not_new_n1576__113988951853731430;
  wire new_n3051_;
  wire not_new_n1065__9;
  wire not_new_n1059__9;
  wire new_n2355_;
  wire not_new_n4697_;
  wire not_new_n627__1176490;
  wire new_n7978_;
  wire not_new_n617__8;
  wire not_new_n9283_;
  wire not_new_n6619__0;
  wire not_new_n3346_;
  wire new_n8028_;
  wire and_new_n6385__new_n6386_;
  wire new_n9877_;
  wire not_new_n1585__403536070;
  wire new_n5484_;
  wire not_new_n2211_;
  wire not_new_n602__1;
  wire not_new_n3153_;
  wire not_new_n1602__57648010;
  wire not_new_n6877_;
  wire not_new_n5181_;
  wire not_new_n5030_;
  wire not_new_n1007__7;
  wire new_n8445_;
  wire or_or_not_new_n3965__not_new_n3966__not_new_n3968_;
  wire new_n7017_;
  wire new_n4541_;
  wire not_new_n10156__0;
  wire not_new_n2733_;
  wire not_new_n610__0;
  wire not_new_n7322_;
  wire not_new_n2746_;
  wire not_new_n3825_;
  wire not_new_n1631__57648010;
  wire new_n7272_;
  wire new_n7244_;
  wire not_new_n1430_;
  wire not_new_n4795_;
  wire not_new_n8447_;
  wire new_n7408_;
  wire new_n5757_;
  wire new_n7949_;
  wire not_new_n6242__0;
  wire or_or_not_new_n1315__not_new_n1313__not_new_n2192_;
  wire or_not_new_n6226__0_not_new_n6336_;
  wire new_n6013_;
  wire new_n9591_;
  wire new_n9530_;
  wire not_new_n7791_;
  wire not_new_n8593__0;
  wire new_n3194_;
  wire not_new_n5073_;
  wire not_new_n2509__6;
  wire new_n6847_;
  wire new_n1227_;
  wire new_n2157_;
  wire not_new_n5450_;
  wire not_new_n7631_;
  wire new_n3057_;
  wire not_new_n1045__168070;
  wire new_n5425_;
  wire new_n6086_;
  wire new_n1853_;
  wire new_n8740_;
  wire not_new_n1583_;
  wire not_pi129_3;
  wire new_n1387_;
  wire new_n1522_;
  wire not_new_n6711_;
  wire new_n9096_;
  wire not_new_n2301_;
  wire new_n4135_;
  wire not_new_n8343_;
  wire new_n4045_;
  wire not_pi054_2;
  wire not_new_n636__24010;
  wire not_new_n1203_;
  wire not_new_n622__113988951853731430;
  wire not_new_n10061__0;
  wire new_n736_;
  wire not_new_n585__10;
  wire new_n4096_;
  wire new_n7935_;
  wire not_new_n5002_;
  wire new_n5121_;
  wire not_new_n9871__0;
  wire not_new_n1186_;
  wire not_new_n9594_;
  wire not_new_n6068_;
  wire not_new_n7720_;
  wire not_new_n1037__332329305696010;
  wire key_gate_17;
  wire not_new_n3345_;
  wire or_or_or_not_new_n2964__not_new_n2967__not_new_n2966__not_new_n2968_;
  wire new_n5412_;
  wire new_n2793_;
  wire new_n4346_;
  wire not_new_n3184__490;
  wire not_new_n9048_;
  wire not_new_n5011_;
  wire new_n5500_;
  wire not_new_n1210_;
  wire new_n2683_;
  wire not_new_n3662_;
  wire po270;
  wire not_new_n5730_;
  wire not_new_n629__490;
  wire new_n4501_;
  wire new_n2464_;
  wire not_new_n595__47475615099430;
  wire not_new_n3730_;
  wire not_new_n1008__4;
  wire not_new_n7769__0;
  wire not_new_n1024__3;
  wire or_not_new_n2645__not_new_n2644_;
  wire or_or_not_new_n2151__not_new_n2148__not_new_n2149_;
  wire new_n2351_;
  wire not_new_n1584_;
  wire not_new_n591__5;
  wire not_new_n3441_;
  wire not_new_n7023__1;
  wire po130;
  wire not_new_n5526_;
  wire not_new_n6496_;
  wire or_not_new_n2343__not_new_n2344_;
  wire not_new_n5986_;
  wire new_n3383_;
  wire new_n710_;
  wire not_new_n10020_;
  wire not_new_n4121__2;
  wire new_n3494_;
  wire new_n5269_;
  wire new_n1752_;
  wire new_n10110_;
  wire new_n702_;
  wire not_new_n6737_;
  wire new_n7149_;
  wire new_n7570_;
  wire not_new_n7421__0;
  wire not_new_n3687_;
  wire new_n6332_;
  wire new_n3292_;
  wire not_new_n1256_;
  wire not_new_n1350_;
  wire new_n5930_;
  wire new_n2186_;
  wire not_pi269_4;
  wire new_n7381_;
  wire new_n10159_;
  wire not_pi267;
  wire not_new_n4347_;
  wire new_n5661_;
  wire not_new_n1588__273687473400809163430;
  wire new_n2875_;
  wire not_new_n7598_;
  wire new_n1564_;
  wire not_pi029;
  wire not_new_n5122_;
  wire not_new_n9428_;
  wire new_n9325_;
  wire not_new_n5329_;
  wire not_new_n5801_;
  wire not_new_n8038_;
  wire new_n9613_;
  wire not_new_n1453_;
  wire not_new_n9374__0;
  wire not_new_n626__138412872010;
  wire not_new_n9472_;
  wire po006;
  wire new_n8940_;
  wire new_n10291_;
  wire not_new_n984__4;
  wire new_n6380_;
  wire not_new_n6471_;
  wire new_n2199_;
  wire not_new_n1153_;
  wire new_n6019_;
  wire not_new_n6784_;
  wire not_pi225;
  wire not_new_n625__1915812313805664144010;
  wire not_new_n1367_;
  wire not_new_n6980_;
  wire new_n1981_;
  wire and_new_n2682__new_n2681_;
  wire new_n10010_;
  wire not_new_n2974_;
  wire not_new_n7411_;
  wire not_new_n1537__5;
  wire not_new_n3387__3;
  wire not_new_n1467_;
  wire not_new_n8829__0;
  wire not_new_n5483_;
  wire new_n3100_;
  wire not_po296_3119734822845423713013303218219760490;
  wire not_new_n1031__2824752490;
  wire new_n10106_;
  wire new_n2758_;
  wire not_new_n1728__138412872010;
  wire not_pi137_1;
  wire not_new_n626__403536070;
  wire not_pi057_2;
  wire new_n9965_;
  wire new_n4520_;
  wire not_new_n5218__0;
  wire not_pi264_1;
  wire not_new_n2930_;
  wire or_not_new_n1863__not_new_n1864_;
  wire not_new_n2780_;
  wire new_n2234_;
  wire not_new_n645__47475615099430;
  wire new_n7873_;
  wire not_new_n7060_;
  wire not_new_n587__2824752490;
  wire new_n8673_;
  wire not_new_n639__113988951853731430;
  wire not_new_n631__657123623635342801395430;
  wire not_new_n5462_;
  wire not_new_n8175__0;
  wire not_new_n5485__0;
  wire not_new_n1401_;
  wire new_n7740_;
  wire new_n7592_;
  wire not_new_n2760_;
  wire not_new_n609__4;
  wire not_new_n7213_;
  wire not_new_n7741_;
  wire new_n9763_;
  wire not_pi063;
  wire not_new_n9385_;
  wire new_n3152_;
  wire new_n5361_;
  wire not_new_n632__273687473400809163430;
  wire new_n4698_;
  wire new_n1747_;
  wire new_n3232_;
  wire new_n6083_;
  wire new_n8099_;
  wire new_n3217_;
  wire not_new_n9968_;
  wire not_pi141;
  wire not_new_n7457__0;
  wire new_n5320_;
  wire not_new_n3923__0;
  wire new_n9085_;
  wire not_new_n585__19773267430;
  wire new_n5629_;
  wire not_new_n6572_;
  wire not_new_n7920_;
  wire new_n5936_;
  wire and_new_n6251__new_n6371_;
  wire new_n4657_;
  wire new_n2940_;
  wire not_new_n1041__6782230728490;
  wire not_new_n1049__3430;
  wire not_new_n4136__2;
  wire new_n2953_;
  wire not_new_n629__2326305139872070;
  wire not_new_n10152_;
  wire new_n4294_;
  wire not_new_n6186_;
  wire new_n3398_;
  wire not_new_n8125_;
  wire not_new_n9511_;
  wire not_new_n4462_;
  wire new_n10183_;
  wire new_n4846_;
  wire not_new_n928__19773267430;
  wire new_n8133_;
  wire not_new_n6701_;
  wire new_n7845_;
  wire not_new_n9142_;
  wire new_n7851_;
  wire not_new_n5073__0;
  wire new_n9414_;
  wire not_new_n1059__19773267430;
  wire not_new_n597__0;
  wire not_new_n6700_;
  wire not_new_n6545_;
  wire new_n995_;
  wire not_new_n588__16284135979104490;
  wire not_new_n593__6782230728490;
  wire not_new_n10299_;
  wire new_n1459_;
  wire not_new_n6159__0;
  wire not_new_n8109__0;
  wire new_n7180_;
  wire not_new_n1596__1176490;
  wire new_n8527_;
  wire new_n977_;
  wire not_new_n8979__0;
  wire not_pi042_3;
  wire not_new_n4519_;
  wire not_new_n587__9;
  wire not_new_n10326_;
  wire not_new_n10184__0;
  wire new_n5351_;
  wire new_n7438_;
  wire not_new_n4350_;
  wire new_n9493_;
  wire not_new_n5362_;
  wire new_n2617_;
  wire new_n6648_;
  wire new_n10168_;
  wire new_n2181_;
  wire new_n2091_;
  wire not_new_n8513_;
  wire new_n10127_;
  wire or_or_not_new_n2883__not_new_n2886__not_new_n2885_;
  wire key_gate_24;
  wire new_n726_;
  wire not_new_n1611__5;
  wire not_new_n1065__16284135979104490;
  wire new_n8766_;
  wire new_n4497_;
  wire new_n8697_;
  wire not_new_n1626__1;
  wire not_new_n644__70;
  wire po129;
  wire not_po296_1299348114471230201171721456984490;
  wire new_n3161_;
  wire not_new_n6529__0;
  wire new_n10140_;
  wire not_new_n1405_;
  wire not_new_n3587_;
  wire not_new_n8634_;
  wire new_n2962_;
  wire new_n8982_;
  wire new_n8074_;
  wire or_not_new_n1331__not_new_n1329_;
  wire not_pi202;
  wire not_new_n10203_;
  wire not_new_n2509__10;
  wire new_n8348_;
  wire not_new_n7647__0;
  wire not_pi272_0;
  wire new_n9606_;
  wire not_new_n1591__8;
  wire new_n2444_;
  wire new_n1488_;
  wire new_n634_;
  wire new_n8816_;
  wire new_n1383_;
  wire new_n9099_;
  wire not_new_n9990_;
  wire or_not_new_n8221__not_new_n8220_;
  wire new_n8622_;
  wire new_n7600_;
  wire not_new_n1594__5;
  wire not_new_n643__6;
  wire not_new_n10291_;
  wire new_n1160_;
  wire not_new_n7794_;
  wire new_n9623_;
  wire new_n614_;
  wire not_new_n3337_;
  wire not_new_n1597__5585458640832840070;
  wire not_new_n7346_;
  wire not_new_n9857_;
  wire not_new_n600__47475615099430;
  wire not_new_n8940_;
  wire not_new_n6323_;
  wire not_new_n4428_;
  wire new_n8801_;
  wire not_new_n8124_;
  wire not_po296_657123623635342801395430;
  wire new_n1351_;
  wire new_n7993_;
  wire not_new_n1049__113988951853731430;
  wire not_new_n4775_;
  wire new_n2018_;
  wire new_n665_;
  wire not_new_n5754__0;
  wire new_n7105_;
  wire not_new_n9620__0;
  wire new_n1247_;
  wire new_n4932_;
  wire not_new_n7302_;
  wire not_new_n1027__10;
  wire not_new_n1585__10;
  wire new_n4088_;
  wire new_n6058_;
  wire not_new_n8461_;
  wire new_n3612_;
  wire new_n8110_;
  wire not_new_n4444_;
  wire not_new_n5920__1;
  wire new_n9365_;
  wire not_new_n5803_;
  wire not_new_n641__24010;
  wire new_n7215_;
  wire not_new_n7109_;
  wire not_new_n8332_;
  wire not_new_n7332_;
  wire not_new_n10206_;
  wire new_n9437_;
  wire not_new_n1308_;
  wire po039;
  wire new_n1537_;
  wire new_n9849_;
  wire not_new_n5347_;
  wire not_new_n5342_;
  wire new_n8902_;
  wire po283;
  wire not_po296_185621159210175743024531636712070;
  wire not_new_n630__490;
  wire not_new_n2881_;
  wire not_new_n4396_;
  wire new_n6155_;
  wire not_new_n1047__2824752490;
  wire not_new_n581__125892552985318850263419623839875454447587430;
  wire not_new_n617__657123623635342801395430;
  wire new_n9914_;
  wire not_new_n6909_;
  wire not_new_n673_;
  wire new_n1327_;
  wire new_n4107_;
  wire not_new_n1039__7;
  wire new_n10013_;
  wire not_new_n1576__1;
  wire not_new_n3335_;
  wire not_new_n3854_;
  wire not_new_n3544_;
  wire not_new_n588__6782230728490;
  wire or_or_not_new_n8781__not_new_n8701__not_new_n8780_;
  wire not_new_n5839_;
  wire new_n2789_;
  wire new_n10261_;
  wire new_n7785_;
  wire new_n5608_;
  wire new_n1706_;
  wire new_n5550_;
  wire not_new_n3460_;
  wire not_new_n9325_;
  wire not_new_n1604__4;
  wire not_new_n3835_;
  wire not_new_n6344_;
  wire new_n5088_;
  wire new_n9342_;
  wire new_n7720_;
  wire not_new_n1598__113988951853731430;
  wire and_new_n2399__new_n2398_;
  wire new_n4502_;
  wire not_new_n1043__10;
  wire new_n7801_;
  wire not_new_n5807__0;
  wire new_n5765_;
  wire new_n1913_;
  wire not_new_n1537__403536070;
  wire key_gate_51;
  wire new_n744_;
  wire not_new_n1900__0;
  wire not_new_n634__7;
  wire new_n2707_;
  wire new_n2363_;
  wire new_n8625_;
  wire new_n5955_;
  wire new_n9838_;
  wire not_new_n4243_;
  wire new_n5364_;
  wire not_new_n7581_;
  wire not_new_n8708_;
  wire new_n6049_;
  wire new_n1366_;
  wire not_new_n1613__138412872010;
  wire not_new_n3429_;
  wire new_n7718_;
  wire not_new_n2594_;
  wire new_n6383_;
  wire not_new_n9515_;
  wire not_new_n7249_;
  wire not_new_n630__113988951853731430;
  wire or_not_new_n8413__not_new_n8252_;
  wire not_new_n3555_;
  wire new_n8638_;
  wire new_n10308_;
  wire not_new_n8971_;
  wire not_new_n4802__1;
  wire not_new_n1061__57648010;
  wire not_pi274_0;
  wire not_new_n3506_;
  wire not_new_n6811_;
  wire po112;
  wire not_new_n1728__2824752490;
  wire not_new_n8866__0;
  wire not_new_n6745_;
  wire not_new_n1059__6;
  wire not_new_n1071__8235430;
  wire not_new_n1604__9;
  wire and_new_n3007__new_n998_;
  wire not_new_n598__1;
  wire new_n10128_;
  wire not_new_n1538__47475615099430;
  wire not_pi128;
  wire new_n7108_;
  wire new_n9339_;
  wire or_not_new_n4841__not_new_n4762_;
  wire not_new_n2341_;
  wire not_new_n632__4;
  wire not_new_n5748__0;
  wire not_new_n1047__168070;
  wire not_new_n6651__0;
  wire not_pi040_3;
  wire not_new_n7870_;
  wire not_new_n9059_;
  wire not_new_n1538__10;
  wire not_new_n4499_;
  wire new_n2575_;
  wire or_not_new_n5453__not_new_n5706__1;
  wire new_n1174_;
  wire not_new_n5499_;
  wire not_new_n2052__0;
  wire not_new_n7090_;
  wire new_n5396_;
  wire new_n1921_;
  wire not_new_n9326__0;
  wire new_n8986_;
  wire new_n5037_;
  wire new_n2083_;
  wire not_new_n1597__2;
  wire not_new_n8824_;
  wire not_new_n9535_;
  wire not_new_n8857__0;
  wire new_n7650_;
  wire not_pi051_3;
  wire not_new_n8131__0;
  wire new_n3600_;
  wire new_n5355_;
  wire not_new_n7590_;
  wire not_new_n9950_;
  wire new_n9683_;
  wire new_n6582_;
  wire new_n10219_;
  wire not_new_n6178_;
  wire new_n9765_;
  wire not_new_n8687_;
  wire not_new_n8155_;
  wire new_n3003_;
  wire new_n4797_;
  wire not_new_n3583_;
  wire not_new_n8209_;
  wire new_n2997_;
  wire not_new_n630__797922662976120010;
  wire not_new_n3375__0;
  wire not_new_n7597_;
  wire or_not_new_n1247__not_new_n1245_;
  wire new_n8493_;
  wire not_new_n595__1176490;
  wire not_new_n9611_;
  wire not_new_n5367_;
  wire new_n7142_;
  wire new_n5340_;
  wire not_new_n1190_;
  wire not_new_n648__47475615099430;
  wire not_new_n1600__403536070;
  wire not_new_n6771_;
  wire not_new_n6974__1;
  wire not_new_n7735__1;
  wire not_new_n641__57648010;
  wire not_new_n8125__0;
  wire not_new_n8027_;
  wire new_n6132_;
  wire new_n8721_;
  wire new_n8076_;
  wire not_new_n1363_;
  wire new_n2598_;
  wire new_n2905_;
  wire not_new_n6645_;
  wire not_new_n8601_;
  wire not_new_n1065__6782230728490;
  wire new_n9614_;
  wire new_n3657_;
  wire not_new_n7743_;
  wire new_n7867_;
  wire not_new_n1728__968890104070;
  wire not_new_n6842_;
  wire not_new_n5915__0;
  wire new_n4149_;
  wire not_pi172_3;
  wire not_new_n5459__1;
  wire not_new_n4333_;
  wire not_new_n1534__2326305139872070;
  wire not_new_n590__1;
  wire not_new_n1824__0;
  wire not_new_n5307_;
  wire new_n2326_;
  wire not_new_n3904_;
  wire new_n5726_;
  wire new_n3845_;
  wire new_n950_;
  wire not_new_n10069_;
  wire not_new_n7828_;
  wire not_new_n7107_;
  wire not_new_n8902_;
  wire not_new_n6543_;
  wire not_new_n9830_;
  wire not_new_n3966_;
  wire not_new_n8918_;
  wire not_new_n9467_;
  wire new_n9148_;
  wire not_pi246;
  wire not_new_n4446_;
  wire new_n3970_;
  wire and_not_pi048_2_not_pi047_2;
  wire not_new_n1045__6;
  wire new_n3236_;
  wire new_n3920_;
  wire not_new_n1591__10;
  wire new_n3136_;
  wire not_new_n3184__6;
  wire new_n10265_;
  wire not_new_n6370_;
  wire not_new_n1537__1;
  wire po146;
  wire new_n8321_;
  wire not_new_n6009_;
  wire not_new_n943_;
  wire new_n5060_;
  wire new_n1279_;
  wire new_n9669_;
  wire not_new_n8584_;
  wire not_new_n4640_;
  wire not_new_n3477_;
  wire not_new_n1003__6;
  wire not_new_n1601__8;
  wire not_new_n9957_;
  wire new_n9817_;
  wire not_new_n1576__968890104070;
  wire not_new_n7025__0;
  wire new_n2913_;
  wire new_n7183_;
  wire new_n8179_;
  wire new_n3952_;
  wire not_new_n8229_;
  wire not_new_n1057_;
  wire not_new_n7847_;
  wire not_new_n635__19773267430;
  wire not_new_n6760_;
  wire not_new_n9858_;
  wire not_new_n2523_;
  wire not_new_n3943_;
  wire not_new_n9558_;
  wire not_new_n4286__0;
  wire new_n6409_;
  wire new_n9198_;
  wire not_new_n8654_;
  wire not_new_n5875_;
  wire new_n10307_;
  wire new_n5455_;
  wire not_new_n9919__0;
  wire not_new_n977_;
  wire not_new_n9812_;
  wire not_new_n9378_;
  wire new_n2260_;
  wire not_pi028_0;
  wire new_n10206_;
  wire not_new_n7551_;
  wire new_n8037_;
  wire not_new_n1589__490;
  wire new_n4807_;
  wire not_new_n8066_;
  wire not_new_n623__3;
  wire new_n6074_;
  wire not_new_n1581__1;
  wire new_n1045_;
  wire and_new_n4351__new_n4350_;
  wire not_new_n1876_;
  wire or_or_not_new_n2170__not_new_n2167__not_new_n2168_;
  wire new_n7681_;
  wire not_new_n9481_;
  wire not_new_n9895_;
  wire key_gate_6;
  wire not_new_n4436__0;
  wire not_new_n9200_;
  wire new_n10278_;
  wire not_new_n1526_;
  wire new_n6819_;
  wire not_new_n2694_;
  wire new_n7567_;
  wire key_gate_57;
  wire new_n5199_;
  wire new_n10232_;
  wire not_new_n5115_;
  wire not_new_n8837__1;
  wire new_n8068_;
  wire not_new_n4598_;
  wire not_new_n637__2326305139872070;
  wire not_new_n1591__16284135979104490;
  wire not_new_n2282_;
  wire not_new_n3453_;
  wire not_new_n10116_;
  wire new_n8968_;
  wire new_n4689_;
  wire not_new_n2806_;
  wire not_new_n9949__0;
  wire new_n2275_;
  wire new_n3363_;
  wire not_new_n984__57648010;
  wire not_new_n4740_;
  wire new_n8301_;
  wire new_n1571_;
  wire not_new_n1014__4;
  wire not_new_n585__138412872010;
  wire not_new_n10217_;
  wire not_new_n1631__8;
  wire not_new_n6001_;
  wire new_n2459_;
  wire new_n1007_;
  wire new_n4269_;
  wire not_new_n6364_;
  wire not_new_n605__490;
  wire not_new_n3861_;
  wire not_new_n1596__47475615099430;
  wire not_new_n5665_;
  wire not_new_n7563_;
  wire not_new_n996_;
  wire not_new_n606__4;
  wire new_n2596_;
  wire not_new_n4570_;
  wire new_n6961_;
  wire new_n7522_;
  wire not_new_n636__113988951853731430;
  wire new_n10016_;
  wire not_new_n7355_;
  wire new_n6547_;
  wire not_new_n9847_;
  wire not_new_n994__3430;
  wire not_new_n7436__0;
  wire not_new_n1619__0;
  wire not_new_n8367_;
  wire not_new_n4442__0;
  wire not_new_n586__4;
  wire not_new_n7774_;
  wire new_n8232_;
  wire not_new_n1356_;
  wire new_n8575_;
  wire new_n3639_;
  wire new_n5989_;
  wire not_new_n8621_;
  wire not_new_n1628_;
  wire new_n4205_;
  wire new_n8140_;
  wire new_n8796_;
  wire not_new_n6983__0;
  wire new_n8884_;
  wire new_n9290_;
  wire new_n4845_;
  wire not_new_n9530_;
  wire new_n1463_;
  wire not_pi263_2;
  wire new_n6426_;
  wire or_not_new_n6327__not_new_n6373__2;
  wire new_n5566_;
  wire not_new_n775__8235430;
  wire not_new_n719__0;
  wire or_not_new_n2189__not_new_n2186_;
  wire not_new_n761_;
  wire new_n6191_;
  wire not_new_n9943__0;
  wire not_new_n1926_;
  wire new_n2937_;
  wire new_n3496_;
  wire not_new_n643__24010;
  wire new_n6462_;
  wire new_n7322_;
  wire not_new_n7611__1;
  wire not_new_n9196_;
  wire new_n2175_;
  wire new_n6378_;
  wire not_new_n6974__10;
  wire not_new_n4220_;
  wire new_n7426_;
  wire new_n8553_;
  wire new_n6541_;
  wire not_new_n8087_;
  wire not_new_n3539_;
  wire not_new_n6981__1;
  wire new_n4190_;
  wire not_new_n4130_;
  wire and_new_n5083__new_n5411_;
  wire not_new_n1611__9;
  wire not_new_n753_;
  wire not_new_n587__1;
  wire not_new_n5873_;
  wire or_not_new_n2015__not_new_n2016_;
  wire not_new_n10332_;
  wire not_new_n775__19773267430;
  wire not_new_n7041__0;
  wire new_n9546_;
  wire not_new_n3181_;
  wire new_n6495_;
  wire new_n5114_;
  wire not_new_n6477_;
  wire not_new_n6347_;
  wire not_new_n1067__3;
  wire not_new_n1589__19773267430;
  wire new_n8573_;
  wire not_new_n1393_;
  wire not_new_n7039_;
  wire new_n6350_;
  wire new_n6451_;
  wire new_n8578_;
  wire new_n3962_;
  wire not_new_n7708_;
  wire new_n3827_;
  wire not_new_n8304__0;
  wire new_n9892_;
  wire not_new_n3311__6;
  wire new_n1514_;
  wire not_new_n6539__2;
  wire new_n1293_;
  wire new_n2015_;
  wire not_new_n1012__7;
  wire new_n3891_;
  wire not_new_n595__9;
  wire new_n7899_;
  wire or_or_not_new_n2015__not_new_n2016__not_new_n2018_;
  wire not_new_n641__403536070;
  wire not_new_n941_;
  wire or_not_new_n1920__not_new_n1921_;
  wire new_n10304_;
  wire new_n7470_;
  wire and_new_n2692__new_n2691_;
  wire not_new_n994__332329305696010;
  wire not_po296_32199057558131797268376070;
  wire not_new_n5207_;
  wire or_or_not_new_n1303__not_new_n1301__not_new_n2135_;
  wire new_n1453_;
  wire new_n9956_;
  wire not_new_n7079_;
  wire new_n7836_;
  wire new_n2654_;
  wire not_new_n10298_;
  wire new_n1019_;
  wire new_n7789_;
  wire not_new_n8110__1;
  wire not_new_n6864_;
  wire new_n3748_;
  wire not_new_n9870__0;
  wire not_new_n4950_;
  wire not_new_n1589__4;
  wire po094;
  wire new_n10331_;
  wire new_n7304_;
  wire not_new_n1063__6782230728490;
  wire new_n5305_;
  wire not_new_n10082_;
  wire not_new_n4418_;
  wire not_new_n9786_;
  wire not_new_n9945__0;
  wire new_n9777_;
  wire new_n8510_;
  wire not_new_n595__3;
  wire not_new_n8282_;
  wire not_new_n4504__0;
  wire not_new_n8933_;
  wire not_new_n4917_;
  wire new_n4357_;
  wire not_new_n989__2824752490;
  wire new_n8141_;
  wire new_n3094_;
  wire new_n2387_;
  wire not_new_n9055_;
  wire not_new_n9592_;
  wire new_n10021_;
  wire not_new_n8863_;
  wire not_new_n4125__1;
  wire new_n1403_;
  wire not_new_n8925_;
  wire new_n9647_;
  wire not_new_n1349_;
  wire new_n3009_;
  wire new_n3821_;
  wire new_n7060_;
  wire not_new_n5861_;
  wire new_n3613_;
  wire new_n9941_;
  wire not_new_n4825__0;
  wire not_new_n3315__0;
  wire not_new_n4344__0;
  wire not_new_n640__3430;
  wire po230;
  wire new_n8589_;
  wire new_n5093_;
  wire not_new_n3766_;
  wire new_n10312_;
  wire new_n4144_;
  wire new_n5171_;
  wire not_new_n3315__332329305696010;
  wire new_n5467_;
  wire not_new_n3351_;
  wire or_or_not_new_n2928__not_new_n2931__not_new_n2930_;
  wire new_n8506_;
  wire not_new_n1005__6;
  wire not_new_n10133_;
  wire not_new_n618__57648010;
  wire not_new_n4796__0;
  wire not_new_n603__57648010;
  wire new_n7000_;
  wire new_n7497_;
  wire new_n2241_;
  wire not_new_n7408_;
  wire not_new_n10093_;
  wire new_n681_;
  wire new_n1216_;
  wire not_new_n594__70;
  wire not_new_n7854_;
  wire not_new_n4694_;
  wire new_n6624_;
  wire not_new_n7029_;
  wire not_new_n1027__113988951853731430;
  wire not_new_n4227__0;
  wire not_new_n8146_;
  wire not_new_n1629_;
  wire new_n9798_;
  wire not_new_n1045_;
  wire new_n9989_;
  wire not_new_n5948__0;
  wire new_n5777_;
  wire not_new_n1678_;
  wire not_new_n9089_;
  wire not_new_n3352_;
  wire not_new_n4457__0;
  wire not_new_n1612__16284135979104490;
  wire new_n1223_;
  wire new_n1434_;
  wire not_new_n731__0;
  wire new_n3672_;
  wire not_new_n1603__138412872010;
  wire not_new_n5439_;
  wire not_new_n6188_;
  wire new_n9200_;
  wire new_n1577_;
  wire new_n5754_;
  wire not_new_n5661_;
  wire not_new_n8331_;
  wire not_new_n591__332329305696010;
  wire new_n6734_;
  wire not_po296_4599865365447399609768010;
  wire new_n5826_;
  wire not_new_n7018__0;
  wire key_gate_12;
  wire not_po296_14811132966169777414641055325137507340304213552070;
  wire new_n4721_;
  wire new_n9611_;
  wire new_n9070_;
  wire not_new_n6947_;
  wire new_n2480_;
  wire not_new_n6515__0;
  wire not_new_n6139_;
  wire not_new_n3231_;
  wire not_new_n1616__3;
  wire not_new_n6974__19773267430;
  wire not_new_n6190_;
  wire new_n8998_;
  wire not_new_n603__24010;
  wire not_new_n2237_;
  wire not_new_n6523__0;
  wire new_n5560_;
  wire not_new_n3114_;
  wire not_new_n3171_;
  wire not_new_n8184_;
  wire new_n4805_;
  wire new_n9358_;
  wire new_n5990_;
  wire not_new_n5835_;
  wire not_new_n3395_;
  wire not_new_n4312_;
  wire new_n650_;
  wire new_n607_;
  wire not_new_n4603_;
  wire not_new_n619__168070;
  wire new_n3401_;
  wire not_new_n3982_;
  wire not_new_n4489_;
  wire not_new_n8466_;
  wire new_n3766_;
  wire new_n1033_;
  wire new_n7794_;
  wire not_new_n8718_;
  wire not_new_n1332_;
  wire not_new_n7311_;
  wire new_n3857_;
  wire new_n10162_;
  wire not_new_n1035_;
  wire not_new_n3276_;
  wire not_new_n7437_;
  wire not_po296_541169560379521116689596608490;
  wire not_new_n8025_;
  wire not_new_n2889_;
  wire new_n5272_;
  wire new_n8286_;
  wire new_n2769_;
  wire not_new_n8856__0;
  wire not_new_n8385_;
  wire new_n6345_;
  wire new_n2296_;
  wire new_n578_;
  wire new_n2982_;
  wire not_new_n5869_;
  wire not_new_n604__1176490;
  wire not_new_n1597__797922662976120010;
  wire new_n2166_;
  wire new_n2402_;
  wire not_new_n10262_;
  wire not_new_n7371_;
  wire new_n9287_;
  wire not_new_n9301_;
  wire new_n6264_;
  wire not_new_n589__9;
  wire not_new_n1607__168070;
  wire new_n2788_;
  wire not_new_n9356__1;
  wire not_new_n1616__403536070;
  wire not_new_n8339_;
  wire not_new_n1599__47475615099430;
  wire not_new_n1057__19773267430;
  wire and_new_n3792__new_n3795_;
  wire not_new_n5218_;
  wire not_new_n6974__403536070;
  wire new_n9869_;
  wire new_n8225_;
  wire not_new_n2978_;
  wire not_new_n3311__57648010;
  wire new_n8728_;
  wire not_new_n6655__1;
  wire new_n5919_;
  wire not_new_n2500_;
  wire not_new_n6443__70;
  wire new_n10329_;
  wire new_n699_;
  wire not_pi242;
  wire not_new_n618__1176490;
  wire new_n5154_;
  wire key_gate_2;
  wire new_n10258_;
  wire not_new_n4788__0;
  wire not_new_n643__2326305139872070;
  wire not_new_n982_;
  wire new_n4113_;
  wire not_new_n8186_;
  wire not_new_n7639_;
  wire new_n7163_;
  wire new_n3933_;
  wire and_new_n2335__new_n2336_;
  wire not_new_n1600__3;
  wire not_new_n634_;
  wire not_new_n2645_;
  wire not_new_n4904_;
  wire not_pi025;
  wire or_or_not_new_n2794__not_new_n2797__not_new_n2796_;
  wire new_n9232_;
  wire new_n7849_;
  wire new_n4729_;
  wire not_new_n7160_;
  wire or_not_new_n1550__not_new_n1370_;
  wire not_new_n4159__0;
  wire not_new_n9996_;
  wire new_n7660_;
  wire new_n4649_;
  wire not_new_n6874_;
  wire new_n2897_;
  wire not_new_n4477__0;
  wire not_pi067;
  wire new_n7699_;
  wire not_new_n591__10;
  wire new_n5214_;
  wire not_new_n635__57648010;
  wire new_n6253_;
  wire new_n6496_;
  wire not_new_n1625_;
  wire not_new_n606__24010;
  wire not_new_n639__9;
  wire not_new_n7141_;
  wire po155;
  wire not_new_n5634_;
  wire new_n5558_;
  wire not_new_n8888__0;
  wire not_new_n956_;
  wire not_new_n7651_;
  wire not_new_n1597__7;
  wire not_new_n5744__0;
  wire not_new_n623__2;
  wire not_po298_4;
  wire not_new_n6965_;
  wire not_pi137_3;
  wire new_n2776_;
  wire new_n5010_;
  wire new_n9754_;
  wire not_pi150_0;
  wire new_n10273_;
  wire new_n7930_;
  wire po141;
  wire not_new_n3944_;
  wire new_n1848_;
  wire not_pi141_1;
  wire not_new_n3372__6782230728490;
  wire and_new_n1290__new_n2084_;
  wire new_n4270_;
  wire new_n8860_;
  wire not_new_n7705_;
  wire not_new_n5233_;
  wire new_n6467_;
  wire not_new_n593__2824752490;
  wire not_new_n6721_;
  wire not_new_n1585__47475615099430;
  wire new_n3270_;
  wire not_new_n9945_;
  wire new_n3628_;
  wire not_new_n928__1;
  wire not_new_n3166_;
  wire not_new_n9774_;
  wire not_new_n7019__1;
  wire new_n593_;
  wire not_new_n8113__1;
  wire not_new_n6549_;
  wire not_new_n6556_;
  wire new_n2441_;
  wire not_po296_4183778472590916451475308348590993345191760458870147715430;
  wire not_new_n10124__0;
  wire new_n5058_;
  wire new_n1670_;
  wire new_n3071_;
  wire new_n1912_;
  wire not_new_n594__4;
  wire not_new_n9450_;
  wire not_new_n8326_;
  wire new_n7909_;
  wire po123;
  wire new_n9022_;
  wire not_pi040_0;
  wire not_new_n1181_;
  wire new_n3826_;
  wire new_n2374_;
  wire not_new_n2753_;
  wire not_new_n1069_;
  wire new_n2986_;
  wire not_new_n5792_;
  wire new_n6259_;
  wire new_n2334_;
  wire or_or_not_new_n6328__not_new_n6373__3_not_new_n6329_;
  wire not_new_n5053_;
  wire not_new_n933_;
  wire not_new_n989__16284135979104490;
  wire not_new_n5436_;
  wire new_n7250_;
  wire and_not_pi044_1_not_pi043_1;
  wire not_new_n639__138412872010;
  wire not_new_n5785__0;
  wire not_new_n620__5;
  wire new_n2646_;
  wire not_new_n5428_;
  wire not_new_n1585__1;
  wire new_n6337_;
  wire not_new_n8254_;
  wire not_new_n638__39098210485829880490;
  wire new_n4104_;
  wire not_new_n3119_;
  wire not_new_n3537_;
  wire new_n10237_;
  wire not_new_n10284_;
  wire new_n6632_;
  wire not_new_n619__6782230728490;
  wire not_new_n1276_;
  wire new_n6525_;
  wire not_new_n2763_;
  wire not_new_n6519__0;
  wire not_new_n2268_;
  wire not_new_n1045__403536070;
  wire or_or_not_new_n1231__not_new_n1229__not_new_n1793_;
  wire not_new_n9937_;
  wire not_new_n8308_;
  wire not_new_n6911_;
  wire not_new_n1611__8;
  wire not_new_n3270_;
  wire not_new_n8491_;
  wire new_n6121_;
  wire not_new_n1538__8235430;
  wire new_n8691_;
  wire not_new_n8486_;
  wire not_new_n1020__3;
  wire not_new_n1007__2;
  wire not_new_n626__5;
  wire not_new_n1537__2824752490;
  wire not_new_n636__3430;
  wire not_new_n2546_;
  wire new_n6915_;
  wire new_n6875_;
  wire not_new_n6795_;
  wire not_new_n1214_;
  wire not_new_n6540_;
  wire new_n9580_;
  wire not_new_n7498_;
  wire not_new_n2877_;
  wire not_new_n617__57648010;
  wire not_new_n685_;
  wire and_new_n9717__new_n9715_;
  wire new_n9712_;
  wire new_n7972_;
  wire not_new_n4523_;
  wire not_new_n6719__0;
  wire not_new_n3585_;
  wire new_n2046_;
  wire new_n9233_;
  wire not_new_n7222_;
  wire not_new_n9016_;
  wire not_new_n626__6782230728490;
  wire and_new_n6422__new_n6426_;
  wire new_n642_;
  wire not_new_n3674_;
  wire not_new_n1616__138412872010;
  wire new_n6299_;
  wire new_n7937_;
  wire not_new_n4171__0;
  wire not_new_n8939_;
  wire not_new_n9591_;
  wire not_new_n4004__0;
  wire new_n9453_;
  wire new_n7150_;
  wire or_not_new_n1275__not_new_n1273_;
  wire not_new_n9770_;
  wire not_new_n1576__490;
  wire new_n7430_;
  wire and_new_n4344__new_n4343_;
  wire not_new_n9485_;
  wire or_not_new_n1303__not_new_n1301_;
  wire new_n1435_;
  wire new_n5388_;
  wire not_new_n2735_;
  wire not_new_n6805_;
  wire new_n5779_;
  wire and_not_pi051_1_not_pi050_1;
  wire new_n8795_;
  wire not_new_n5066_;
  wire not_new_n1041__9;
  wire new_n10091_;
  wire not_new_n4116_;
  wire not_new_n2782_;
  wire new_n1061_;
  wire new_n1748_;
  wire not_new_n1055__6;
  wire new_n5502_;
  wire not_new_n7243_;
  wire new_n2532_;
  wire new_n6719_;
  wire not_new_n642__10;
  wire not_new_n5612_;
  wire not_new_n7425_;
  wire not_new_n4981_;
  wire not_new_n1051__6;
  wire new_n3129_;
  wire not_new_n5588_;
  wire not_new_n8266__5;
  wire not_pi176;
  wire not_new_n2752_;
  wire new_n9029_;
  wire new_n8669_;
  wire not_new_n622__3;
  wire not_new_n5420_;
  wire po051;
  wire new_n10003_;
  wire not_new_n594__403536070;
  wire new_n2442_;
  wire not_new_n5320_;
  wire new_n7349_;
  wire new_n4375_;
  wire not_pi050;
  wire not_new_n7779_;
  wire not_new_n2873_;
  wire not_new_n6102_;
  wire new_n8264_;
  wire new_n7797_;
  wire not_new_n9332_;
  wire not_new_n1723_;
  wire new_n9369_;
  wire new_n5042_;
  wire not_new_n7505_;
  wire new_n1182_;
  wire po062;
  wire new_n9160_;
  wire new_n7243_;
  wire not_new_n1598__16284135979104490;
  wire new_n7738_;
  wire not_new_n1805__0;
  wire not_new_n1576__138412872010;
  wire not_new_n7448__1;
  wire new_n7033_;
  wire not_new_n8830_;
  wire not_new_n631__24010;
  wire not_new_n928__0;
  wire not_new_n5394_;
  wire not_new_n2090_;
  wire not_new_n593__19773267430;
  wire new_n8464_;
  wire new_n10179_;
  wire not_new_n4980_;
  wire new_n668_;
  wire new_n9805_;
  wire new_n6686_;
  wire not_new_n621__138412872010;
  wire not_new_n7150_;
  wire new_n4627_;
  wire new_n8707_;
  wire new_n2874_;
  wire new_n3522_;
  wire not_new_n1179_;
  wire not_new_n7166_;
  wire new_n9566_;
  wire not_new_n7734_;
  wire not_pi199;
  wire not_new_n4718_;
  wire not_new_n1059__2824752490;
  wire not_new_n8555_;
  wire not_new_n4186_;
  wire not_new_n2014_;
  wire not_new_n1055__332329305696010;
  wire not_new_n601__24010;
  wire new_n5103_;
  wire or_or_not_new_n1920__not_new_n1921__not_new_n1923_;
  wire not_new_n1788_;
  wire new_n5983_;
  wire not_new_n7634_;
  wire not_new_n3381_;
  wire new_n6556_;
  wire not_new_n1045__113988951853731430;
  wire new_n6565_;
  wire not_pi156;
  wire not_new_n1065__2824752490;
  wire new_n9092_;
  wire not_new_n608__1176490;
  wire new_n5479_;
  wire new_n2040_;
  wire new_n8592_;
  wire new_n10054_;
  wire not_new_n6109_;
  wire not_new_n7317_;
  wire not_new_n4531_;
  wire not_new_n2305_;
  wire new_n4987_;
  wire new_n9769_;
  wire new_n3726_;
  wire not_new_n4925_;
  wire new_n5723_;
  wire not_new_n8029_;
  wire po247;
  wire not_new_n8519_;
  wire new_n5357_;
  wire not_new_n3310__168070;
  wire not_new_n4311_;
  wire new_n8521_;
  wire not_new_n5475_;
  wire new_n6990_;
  wire new_n10221_;
  wire not_new_n766_;
  wire not_new_n640__6782230728490;
  wire new_n3444_;
  wire new_n8923_;
  wire new_n5119_;
  wire and_and_new_n1735__new_n1736__new_n1738_;
  wire new_n2041_;
  wire not_new_n4831_;
  wire not_new_n743_;
  wire new_n5790_;
  wire not_new_n9916_;
  wire not_new_n2055_;
  wire new_n1170_;
  wire not_new_n8274_;
  wire not_new_n1047__57648010;
  wire not_new_n4211_;
  wire new_n6614_;
  wire new_n8344_;
  wire new_n5615_;
  wire not_new_n10045__1;
  wire not_new_n6443__138412872010;
  wire not_new_n8648_;
  wire or_not_new_n3128__not_new_n3127_;
  wire not_new_n9274_;
  wire new_n5482_;
  wire not_new_n621__0;
  wire new_n9527_;
  wire not_new_n8944_;
  wire not_new_n598__7;
  wire not_new_n7885_;
  wire not_new_n1325_;
  wire not_new_n617__968890104070;
  wire not_new_n8716_;
  wire not_new_n1035__490;
  wire not_new_n10014_;
  wire new_n5588_;
  wire new_n8941_;
  wire or_not_new_n2908__not_new_n2907_;
  wire not_new_n3118_;
  wire new_n9879_;
  wire new_n5506_;
  wire new_n6394_;
  wire not_new_n7029__1;
  wire not_new_n5756_;
  wire not_new_n733_;
  wire not_new_n601_;
  wire new_n8933_;
  wire not_new_n3987_;
  wire not_new_n9780_;
  wire new_n8030_;
  wire and_new_n8664__new_n8663_;
  wire new_n9024_;
  wire new_n3358_;
  wire not_new_n8415_;
  wire or_not_new_n3143__not_new_n3142_;
  wire not_new_n1065__8;
  wire not_new_n7875_;
  wire not_new_n7624_;
  wire new_n2209_;
  wire not_new_n6724_;
  wire not_new_n3370_;
  wire not_new_n935_;
  wire new_n5491_;
  wire new_n2856_;
  wire new_n7799_;
  wire not_new_n8838__0;
  wire new_n4635_;
  wire new_n8626_;
  wire not_new_n4115__0;
  wire new_n3320_;
  wire not_new_n9808_;
  wire not_new_n1067__9;
  wire new_n1500_;
  wire new_n9710_;
  wire not_new_n5849_;
  wire not_new_n4165__0;
  wire not_new_n3937_;
  wire not_new_n618__657123623635342801395430;
  wire new_n7353_;
  wire not_new_n984__24010;
  wire new_n2967_;
  wire not_new_n3926__0;
  wire new_n8215_;
  wire not_new_n7876__0;
  wire not_new_n5219__0;
  wire not_new_n599__9;
  wire not_new_n7686_;
  wire new_n5279_;
  wire not_new_n9843_;
  wire po128;
  wire new_n4217_;
  wire new_n5675_;
  wire new_n7939_;
  wire new_n5286_;
  wire new_n5902_;
  wire not_new_n7760_;
  wire new_n9278_;
  wire not_new_n5226_;
  wire not_new_n9504_;
  wire not_new_n1500_;
  wire not_new_n598__47475615099430;
  wire new_n5235_;
  wire new_n2594_;
  wire not_new_n9287_;
  wire not_po296_7490483309651862334944941026945644936490;
  wire new_n3772_;
  wire not_new_n637__1176490;
  wire new_n8216_;
  wire not_new_n4131__0;
  wire not_new_n7659_;
  wire not_new_n4454__0;
  wire new_n2315_;
  wire new_n5090_;
  wire not_new_n4517_;
  wire new_n10254_;
  wire not_new_n601__1;
  wire new_n9824_;
  wire not_pi034_3;
  wire not_pi044;
  wire not_new_n2020_;
  wire new_n1055_;
  wire not_new_n640__138412872010;
  wire new_n5781_;
  wire new_n5690_;
  wire not_new_n3184__4;
  wire not_new_n2256_;
  wire not_new_n986__0;
  wire not_new_n1360_;
  wire not_new_n4436_;
  wire new_n1910_;
  wire not_new_n627__4;
  wire new_n7713_;
  wire not_new_n6519__2;
  wire new_n4832_;
  wire not_new_n1389_;
  wire new_n2570_;
  wire not_new_n5174_;
  wire new_n1599_;
  wire new_n3421_;
  wire new_n975_;
  wire new_n9936_;
  wire new_n2807_;
  wire new_n4274_;
  wire not_new_n2092_;
  wire not_new_n9973_;
  wire not_new_n1049__4;
  wire new_n2360_;
  wire not_new_n8095_;
  wire po118;
  wire not_new_n5311_;
  wire new_n7629_;
  wire new_n5445_;
  wire not_new_n1307_;
  wire new_n5110_;
  wire new_n4867_;
  wire new_n9521_;
  wire new_n9704_;
  wire new_n7301_;
  wire not_new_n7160__0;
  wire new_n7231_;
  wire po148;
  wire new_n8810_;
  wire new_n2544_;
  wire not_new_n9993_;
  wire new_n712_;
  wire not_new_n10331_;
  wire not_new_n622__4;
  wire not_new_n8263_;
  wire new_n4643_;
  wire not_new_n9178_;
  wire not_new_n4000_;
  wire not_new_n7916_;
  wire new_n949_;
  wire not_new_n595__138412872010;
  wire new_n3060_;
  wire new_n5401_;
  wire not_new_n5676_;
  wire new_n1476_;
  wire not_new_n588__47475615099430;
  wire not_new_n1027__3;
  wire new_n3034_;
  wire not_new_n5492_;
  wire new_n7069_;
  wire not_new_n6749_;
  wire not_new_n9952_;
  wire not_new_n1027__24010;
  wire new_n7198_;
  wire and_new_n6227__new_n6232_;
  wire not_new_n1604__24010;
  wire new_n7941_;
  wire not_new_n6682_;
  wire not_new_n3315__3;
  wire not_new_n602__490;
  wire new_n3934_;
  wire new_n4290_;
  wire not_new_n4288_;
  wire not_new_n9564_;
  wire not_pi246_0;
  wire not_new_n1613__403536070;
  wire new_n6602_;
  wire not_pi143_0;
  wire not_new_n7754__1;
  wire not_new_n7478_;
  wire new_n6313_;
  wire not_new_n9030_;
  wire not_new_n1009__3;
  wire new_n7029_;
  wire not_new_n1612__1;
  wire not_new_n5900__3;
  wire new_n1868_;
  wire not_new_n6512_;
  wire new_n1559_;
  wire new_n6513_;
  wire not_new_n619__3430;
  wire not_new_n4792_;
  wire key_gate_95;
  wire not_new_n5878__1;
  wire new_n3802_;
  wire new_n5555_;
  wire new_n7587_;
  wire new_n2344_;
  wire new_n1587_;
  wire new_n5447_;
  wire not_new_n5904_;
  wire new_n4392_;
  wire not_new_n639__0;
  wire not_new_n646__332329305696010;
  wire new_n9740_;
  wire new_n1609_;
  wire new_n7807_;
  wire new_n3592_;
  wire not_new_n9840_;
  wire new_n2474_;
  wire not_new_n1063__403536070;
  wire not_new_n1657_;
  wire not_new_n1589__2824752490;
  wire not_new_n5545_;
  wire not_new_n9898_;
  wire not_new_n9936_;
  wire and_new_n7605__new_n7973_;
  wire or_not_new_n1548__not_new_n1366_;
  wire po019;
  wire new_n6208_;
  wire new_n9570_;
  wire new_n10045_;
  wire not_new_n635__8;
  wire not_pi152;
  wire new_n5164_;
  wire new_n3771_;
  wire new_n4813_;
  wire new_n5069_;
  wire new_n8126_;
  wire not_new_n602__47475615099430;
  wire not_new_n6069_;
  wire new_n9931_;
  wire new_n8804_;
  wire new_n5981_;
  wire not_new_n5860_;
  wire key_gate_87;
  wire new_n8568_;
  wire not_new_n3247_;
  wire not_new_n5565_;
  wire new_n7063_;
  wire not_new_n998__0;
  wire not_new_n1402_;
  wire not_new_n9727_;
  wire not_pi032_0;
  wire not_new_n5078__0;
  wire and_new_n1302__new_n2141_;
  wire new_n1396_;
  wire not_new_n1028__1;
  wire new_n2167_;
  wire not_new_n4074_;
  wire new_n4789_;
  wire not_new_n7040__0;
  wire not_new_n1059__113988951853731430;
  wire not_new_n3992_;
  wire not_new_n618__1915812313805664144010;
  wire new_n5787_;
  wire not_new_n10059_;
  wire new_n1267_;
  wire new_n9787_;
  wire not_new_n602__403536070;
  wire or_or_or_not_new_n6363__not_new_n6358__not_new_n6361__not_new_n6366_;
  wire not_new_n1002__0;
  wire not_new_n1049__8;
  wire not_new_n3222_;
  wire new_n1470_;
  wire and_new_n7159__new_n7547_;
  wire not_new_n3316_;
  wire not_new_n6443__797922662976120010;
  wire not_new_n1063__490;
  wire not_new_n8874__0;
  wire not_new_n2248_;
  wire not_new_n644__8;
  wire new_n1982_;
  wire not_new_n648__19773267430;
  wire not_new_n7220_;
  wire new_n2339_;
  wire po106;
  wire not_new_n1604__47475615099430;
  wire new_n7386_;
  wire not_new_n3483_;
  wire new_n2799_;
  wire not_new_n1011__6;
  wire new_n4162_;
  wire not_new_n1631__7;
  wire new_n6845_;
  wire new_n10270_;
  wire new_n2320_;
  wire not_new_n5927_;
  wire and_and_new_n1460__new_n1466__new_n1458_;
  wire new_n3951_;
  wire new_n674_;
  wire new_n3466_;
  wire not_new_n7439__0;
  wire not_new_n622__2;
  wire new_n3239_;
  wire new_n7946_;
  wire not_new_n9181_;
  wire not_new_n3449_;
  wire not_new_n7003__0;
  wire not_new_n10277_;
  wire not_new_n1041__57648010;
  wire new_n8310_;
  wire new_n5992_;
  wire new_n4493_;
  wire new_n7959_;
  wire new_n1509_;
  wire new_n6912_;
  wire new_n7218_;
  wire not_new_n4116__0;
  wire not_new_n8170__0;
  wire not_pi052_2;
  wire not_new_n9086__0;
  wire not_new_n721_;
  wire new_n7648_;
  wire not_new_n5075_;
  wire not_pi234;
  wire not_new_n3066_;
  wire not_new_n585__5;
  wire not_new_n1581__797922662976120010;
  wire not_pi165_3;
  wire not_new_n8966__0;
  wire new_n9251_;
  wire not_new_n7803_;
  wire new_n3895_;
  wire new_n1667_;
  wire and_new_n8082__new_n8430_;
  wire new_n2133_;
  wire not_new_n3704_;
  wire new_n10199_;
  wire new_n7382_;
  wire not_new_n609__8235430;
  wire new_n2515_;
  wire not_new_n7356_;
  wire new_n4018_;
  wire not_new_n2555_;
  wire new_n7461_;
  wire not_new_n6831_;
  wire not_new_n638__490;
  wire new_n6027_;
  wire not_new_n10272_;
  wire not_new_n5059_;
  wire not_new_n1195_;
  wire new_n2551_;
  wire new_n5802_;
  wire new_n6454_;
  wire not_new_n628__24010;
  wire po205;
  wire new_n990_;
  wire new_n2244_;
  wire not_pi080;
  wire new_n3912_;
  wire not_new_n8096_;
  wire new_n8162_;
  wire not_new_n4463_;
  wire new_n3268_;
  wire new_n3536_;
  wire new_n4809_;
  wire not_new_n8978__1;
  wire not_new_n7456_;
  wire new_n10245_;
  wire not_new_n3385_;
  wire not_new_n4998__1;
  wire new_n1791_;
  wire not_new_n5708_;
  wire or_not_new_n2794__not_new_n2797_;
  wire new_n3649_;
  wire not_new_n2933_;
  wire new_n7662_;
  wire not_new_n1765_;
  wire not_new_n5159_;
  wire new_n4905_;
  wire new_n2137_;
  wire new_n3540_;
  wire new_n2976_;
  wire not_new_n6905_;
  wire new_n7616_;
  wire new_n6032_;
  wire new_n3676_;
  wire not_new_n6373__9;
  wire new_n8369_;
  wire not_new_n6527__1;
  wire new_n1810_;
  wire new_n6507_;
  wire new_n6637_;
  wire not_new_n3758_;
  wire new_n7956_;
  wire not_new_n1049__5;
  wire not_new_n1043__6;
  wire not_new_n1588__490;
  wire not_new_n8319_;
  wire not_new_n4464__0;
  wire new_n2572_;
  wire not_new_n1043__168070;
  wire new_n10015_;
  wire not_new_n6330_;
  wire new_n9032_;
  wire new_n1572_;
  wire not_new_n5655_;
  wire not_new_n7139_;
  wire not_new_n5669_;
  wire not_new_n4372_;
  wire not_new_n628__93874803376477543056490;
  wire new_n7273_;
  wire not_new_n5919_;
  wire not_new_n6930_;
  wire not_new_n4411_;
  wire not_new_n6998__1;
  wire not_new_n5764_;
  wire not_new_n6813_;
  wire not_new_n6597_;
  wire not_new_n3514_;
  wire new_n1004_;
  wire new_n6798_;
  wire not_new_n646_;
  wire not_new_n629__24010;
  wire new_n5960_;
  wire not_pi254_1;
  wire not_new_n1585__6;
  wire not_new_n632__5;
  wire new_n7727_;
  wire new_n1389_;
  wire not_new_n1538__968890104070;
  wire new_n4680_;
  wire not_new_n7150__0;
  wire not_new_n1021_;
  wire not_new_n627__57648010;
  wire not_new_n8138__1;
  wire new_n8878_;
  wire or_not_new_n1556__not_new_n2439_;
  wire new_n4152_;
  wire not_new_n7357_;
  wire new_n9853_;
  wire not_new_n620__6;
  wire not_new_n6070_;
  wire not_new_n8550_;
  wire not_new_n6824_;
  wire not_new_n10179_;
  wire new_n8427_;
  wire not_new_n6338_;
  wire new_n3053_;
  wire not_new_n955_;
  wire not_new_n1696_;
  wire not_new_n6042_;
  wire not_new_n5244_;
  wire not_new_n1616__0;
  wire new_n8987_;
  wire new_n8939_;
  wire not_new_n3561_;
  wire not_new_n3387__4;
  wire new_n4647_;
  wire new_n9330_;
  wire new_n9133_;
  wire new_n8156_;
  wire not_new_n7119_;
  wire not_new_n1604__2824752490;
  wire not_new_n5105_;
  wire new_n2682_;
  wire not_new_n2745_;
  wire not_new_n2821_;
  wire new_n5772_;
  wire or_not_new_n2339__not_new_n2340_;
  wire new_n6460_;
  wire new_n7471_;
  wire not_new_n5779__0;
  wire not_new_n1039__168070;
  wire new_n8567_;
  wire new_n4938_;
  wire new_n4123_;
  wire new_n3569_;
  wire new_n3484_;
  wire new_n9125_;
  wire po127;
  wire not_new_n1065__403536070;
  wire not_new_n604__490;
  wire new_n6282_;
  wire new_n9392_;
  wire not_new_n9427__0;
  wire key_gate_121;
  wire new_n2847_;
  wire new_n10335_;
  wire not_new_n8117__1;
  wire new_n5067_;
  wire new_n1356_;
  wire not_new_n622__9;
  wire not_new_n8362_;
  wire not_new_n5703_;
  wire not_new_n5445__0;
  wire not_new_n9802_;
  wire not_new_n7217_;
  wire not_new_n5026_;
  wire not_new_n8744_;
  wire new_n3077_;
  wire not_new_n3507_;
  wire not_new_n732__0;
  wire not_new_n1059__3430;
  wire not_new_n8017_;
  wire not_new_n6786_;
  wire not_new_n643__4;
  wire not_pi249_0;
  wire not_new_n9617_;
  wire new_n9947_;
  wire new_n3924_;
  wire not_new_n622__2824752490;
  wire new_n8596_;
  wire new_n9385_;
  wire not_new_n1059__6782230728490;
  wire new_n4014_;
  wire new_n6020_;
  wire new_n7711_;
  wire not_new_n5530_;
  wire new_n8517_;
  wire not_new_n1354_;
  wire po169;
  wire not_pi008_0;
  wire not_new_n5056_;
  wire new_n6287_;
  wire not_new_n1602__10;
  wire new_n7420_;
  wire new_n1490_;
  wire new_n8855_;
  wire new_n9698_;
  wire not_new_n6565_;
  wire new_n1185_;
  wire not_new_n3315__403536070;
  wire not_new_n7247_;
  wire new_n5952_;
  wire not_new_n8121__0;
  wire new_n4941_;
  wire new_n1255_;
  wire not_new_n7306_;
  wire not_new_n1006__5;
  wire not_new_n2501_;
  wire new_n3810_;
  wire new_n3650_;
  wire new_n1631_;
  wire not_new_n7418__0;
  wire not_new_n6311_;
  wire new_n5430_;
  wire not_new_n1063__57648010;
  wire not_new_n4564_;
  wire not_new_n9073_;
  wire not_new_n8287_;
  wire not_new_n5771__0;
  wire or_not_new_n1283__not_new_n1281_;
  wire not_new_n5856_;
  wire new_n4115_;
  wire not_new_n5885__0;
  wire new_n3506_;
  wire not_new_n7161_;
  wire new_n5643_;
  wire new_n5728_;
  wire not_new_n6216_;
  wire new_n8776_;
  wire new_n6425_;
  wire new_n6066_;
  wire not_new_n1011__2;
  wire new_n8197_;
  wire not_new_n608__0;
  wire not_new_n8192_;
  wire not_new_n8286__0;
  wire new_n6658_;
  wire new_n3512_;
  wire new_n8957_;
  wire new_n2540_;
  wire not_new_n4018_;
  wire new_n8812_;
  wire not_new_n5763__0;
  wire not_new_n4835__0;
  wire not_new_n634__19773267430;
  wire new_n2183_;
  wire not_new_n9718_;
  wire not_new_n6125_;
  wire new_n7911_;
  wire new_n3418_;
  wire new_n5102_;
  wire new_n1343_;
  wire new_n2471_;
  wire new_n8550_;
  wire not_new_n7199_;
  wire new_n5519_;
  wire po204;
  wire not_new_n4747_;
  wire not_new_n661_;
  wire new_n4907_;
  wire new_n10063_;
  wire not_new_n3291_;
  wire new_n5784_;
  wire not_new_n5431_;
  wire not_new_n6376_;
  wire not_new_n3185__490;
  wire not_new_n9326__2;
  wire new_n5296_;
  wire new_n2586_;
  wire not_new_n9232_;
  wire new_n9595_;
  wire new_n4913_;
  wire not_new_n6759_;
  wire not_new_n4591_;
  wire new_n7372_;
  wire not_new_n585__8235430;
  wire not_new_n599__3430;
  wire not_new_n9734_;
  wire not_new_n3676_;
  wire new_n7854_;
  wire not_pi204;
  wire not_new_n5838_;
  wire not_new_n6518_;
  wire new_n7771_;
  wire new_n8814_;
  wire and_new_n4928__new_n5310_;
  wire not_new_n641__2;
  wire new_n6923_;
  wire new_n683_;
  wire not_new_n637__24010;
  wire new_n5536_;
  wire not_new_n7616_;
  wire not_new_n1581__47475615099430;
  wire new_n2635_;
  wire not_new_n2223_;
  wire new_n7723_;
  wire not_new_n10296_;
  wire new_n2618_;
  wire new_n6713_;
  wire and_and_new_n1731__new_n1732__new_n1734_;
  wire not_new_n695_;
  wire not_new_n3234_;
  wire not_new_n6931_;
  wire not_new_n1612__6;
  wire new_n3787_;
  wire new_n6788_;
  wire new_n9938_;
  wire new_n8714_;
  wire not_pi164_3;
  wire new_n4839_;
  wire not_new_n5462__1;
  wire new_n1903_;
  wire not_new_n1057__7;
  wire not_new_n7010__1;
  wire new_n4369_;
  wire not_new_n1020_;
  wire not_new_n6961_;
  wire not_new_n5197_;
  wire not_new_n2729_;
  wire new_n10105_;
  wire new_n5551_;
  wire not_new_n3310__3430;
  wire new_n1541_;
  wire not_new_n4495_;
  wire not_new_n7619__0;
  wire not_new_n4995_;
  wire not_new_n4513_;
  wire not_new_n5951_;
  wire new_n4678_;
  wire new_n5299_;
  wire not_new_n2798_;
  wire new_n9472_;
  wire not_new_n9629_;
  wire new_n8486_;
  wire and_new_n3004__new_n998_;
  wire not_pi166_3;
  wire not_new_n1065__10;
  wire not_new_n628__57648010;
  wire new_n9646_;
  wire not_new_n8341_;
  wire not_new_n775__70;
  wire not_new_n1252_;
  wire key_gate_5;
  wire not_new_n648__403536070;
  wire new_n7343_;
  wire not_new_n3271_;
  wire not_new_n586__5;
  wire new_n931_;
  wire new_n5044_;
  wire not_new_n1583__7;
  wire new_n7859_;
  wire not_new_n8404_;
  wire new_n9550_;
  wire not_new_n3372__19773267430;
  wire new_n6397_;
  wire not_new_n638__1577753820348458066150427430;
  wire not_new_n4787_;
  wire not_new_n2666_;
  wire not_new_n1601__70;
  wire not_new_n9420__0;
  wire new_n6934_;
  wire not_new_n6521__0;
  wire new_n6233_;
  wire not_new_n5797_;
  wire or_not_new_n9166__not_new_n9106_;
  wire new_n7664_;
  wire not_new_n10166__0;
  wire new_n8536_;
  wire new_n3679_;
  wire new_n4914_;
  wire new_n3305_;
  wire or_not_new_n4227__not_new_n1608_;
  wire not_new_n9913_;
  wire new_n1334_;
  wire not_new_n1011__7;
  wire not_new_n594__6782230728490;
  wire and_new_n2364__new_n2363_;
  wire not_new_n8614_;
  wire new_n1300_;
  wire not_new_n5095__1;
  wire new_n4035_;
  wire not_new_n925_;
  wire not_new_n8756_;
  wire not_new_n8170__2;
  wire new_n9785_;
  wire new_n1947_;
  wire or_or_or_not_new_n6239__not_new_n6350__not_new_n6232__3_not_new_n6317__0;
  wire not_new_n7754__4;
  wire not_new_n4432__0;
  wire or_not_new_n1028__8_not_new_n1622__1;
  wire new_n6586_;
  wire or_not_new_n1551__not_new_n1372_;
  wire not_new_n7664__1;
  wire new_n6717_;
  wire not_new_n6738_;
  wire not_new_n7838_;
  wire not_new_n2093_;
  wire not_new_n6501_;
  wire new_n9263_;
  wire not_new_n1536__7;
  wire not_new_n646__3430;
  wire not_new_n1589__168070;
  wire not_new_n4537_;
  wire not_new_n9375_;
  wire not_new_n6612_;
  wire new_n5143_;
  wire not_new_n587__6782230728490;
  wire not_new_n8961_;
  wire not_new_n1583__2;
  wire new_n5862_;
  wire not_new_n9247_;
  wire not_new_n581__5;
  wire not_new_n643__490;
  wire not_new_n994__7;
  wire new_n9100_;
  wire not_new_n4075_;
  wire not_pi031;
  wire not_new_n1017__6;
  wire new_n8597_;
  wire new_n4395_;
  wire new_n9281_;
  wire not_new_n1055__968890104070;
  wire and_and_new_n1915__new_n1918__new_n1916_;
  wire new_n648_;
  wire not_new_n4023_;
  wire new_n6008_;
  wire new_n1558_;
  wire new_n1016_;
  wire new_n6205_;
  wire new_n6832_;
  wire new_n2376_;
  wire not_new_n4832_;
  wire not_new_n7400_;
  wire not_new_n1065__332329305696010;
  wire new_n5627_;
  wire not_new_n7009__1;
  wire new_n1063_;
  wire not_new_n4357_;
  wire not_new_n631_;
  wire new_n3635_;
  wire not_new_n588__332329305696010;
  wire not_new_n1800_;
  wire not_new_n3567_;
  wire new_n1448_;
  wire not_new_n637__0;
  wire not_new_n2907_;
  wire not_new_n9753_;
  wire new_n7279_;
  wire new_n1471_;
  wire not_pi263_0;
  wire new_n1319_;
  wire new_n9513_;
  wire not_new_n4005_;
  wire not_new_n4093_;
  wire not_new_n3421_;
  wire new_n8944_;
  wire or_not_new_n2300__not_new_n2301_;
  wire not_new_n10033_;
  wire new_n2851_;
  wire new_n6609_;
  wire not_new_n613__1;
  wire not_new_n4814_;
  wire new_n9322_;
  wire not_new_n7733_;
  wire not_new_n10143_;
  wire new_n2029_;
  wire new_n7113_;
  wire not_new_n7407_;
  wire or_not_new_n3149__not_new_n3148_;
  wire new_n6524_;
  wire not_new_n5258_;
  wire new_n7858_;
  wire not_new_n1057__8;
  wire new_n6064_;
  wire not_new_n1027__19773267430;
  wire new_n1889_;
  wire new_n4803_;
  wire not_pi060;
  wire new_n5776_;
  wire not_new_n9355_;
  wire new_n4993_;
  wire not_new_n2509__3;
  wire not_new_n7666__0;
  wire not_new_n984__6782230728490;
  wire not_new_n3445_;
  wire new_n8426_;
  wire not_new_n9736_;
  wire not_new_n1067__968890104070;
  wire new_n2743_;
  wire not_new_n1454_;
  wire not_new_n1528_;
  wire not_new_n1037__2;
  wire not_new_n6451__0;
  wire not_po296_9;
  wire not_new_n1285_;
  wire not_new_n6508_;
  wire not_new_n4508_;
  wire not_new_n2218_;
  wire not_new_n1600__57648010;
  wire new_n7175_;
  wire new_n3248_;
  wire not_new_n7345_;
  wire or_not_new_n7311__not_new_n7203_;
  wire not_new_n5473_;
  wire new_n5349_;
  wire new_n7728_;
  wire not_new_n7063_;
  wire not_new_n7075_;
  wire not_new_n6522_;
  wire not_new_n7017_;
  wire new_n4926_;
  wire new_n8209_;
  wire not_pi062_2;
  wire new_n9697_;
  wire new_n4924_;
  wire not_new_n3249_;
  wire not_new_n4803_;
  wire new_n3869_;
  wire new_n2792_;
  wire not_new_n4978_;
  wire new_n10235_;
  wire new_n9334_;
  wire new_n7613_;
  wire not_new_n8631_;
  wire not_new_n3534_;
  wire new_n3106_;
  wire not_new_n2585_;
  wire not_new_n1616__19773267430;
  wire not_new_n4642_;
  wire new_n9778_;
  wire new_n2556_;
  wire not_new_n617__0;
  wire not_new_n6995_;
  wire new_n4307_;
  wire not_new_n581__77309937197074445241370944070;
  wire not_new_n2343_;
  wire new_n1934_;
  wire not_new_n1581__3;
  wire not_new_n4213_;
  wire new_n9479_;
  wire not_new_n4734_;
  wire not_new_n8840_;
  wire not_new_n9160_;
  wire new_n7812_;
  wire or_not_new_n2836__not_new_n2835_;
  wire not_new_n603__6782230728490;
  wire not_new_n4960_;
  wire new_n1283_;
  wire not_new_n641__8235430;
  wire not_new_n1599__9;
  wire not_new_n8398_;
  wire new_n7058_;
  wire not_new_n4478_;
  wire new_n2368_;
  wire or_or_or_not_new_n6240__not_new_n6330__not_new_n6331__not_new_n6242__1;
  wire not_pi068;
  wire not_new_n1047__1176490;
  wire not_new_n3971_;
  wire new_n4790_;
  wire not_new_n10013__0;
  wire not_new_n1015__5;
  wire new_n1766_;
  wire not_new_n1055__8235430;
  wire not_new_n646__47475615099430;
  wire not_new_n6237_;
  wire and_new_n4323__new_n4324_;
  wire not_new_n609_;
  wire not_new_n9021_;
  wire not_new_n8289_;
  wire new_n8236_;
  wire not_new_n5472_;
  wire not_new_n7566_;
  wire new_n9121_;
  wire new_n3636_;
  wire not_new_n626__6;
  wire not_new_n8305_;
  wire new_n7800_;
  wire po261;
  wire and_new_n8750__new_n8736_;
  wire not_new_n1173_;
  wire not_new_n1043__70;
  wire new_n6269_;
  wire new_n2253_;
  wire not_po296_8;
  wire not_new_n5616_;
  wire or_or_not_new_n1267__not_new_n1265__not_new_n1964_;
  wire new_n10253_;
  wire not_new_n4199_;
  wire new_n5045_;
  wire not_new_n1037__10;
  wire new_n7316_;
  wire new_n6477_;
  wire new_n2227_;
  wire not_new_n4014__1;
  wire not_new_n599__0;
  wire not_new_n622__403536070;
  wire new_n7088_;
  wire new_n7249_;
  wire not_new_n1598__2824752490;
  wire new_n6834_;
  wire new_n3651_;
  wire new_n10001_;
  wire not_new_n1028__6;
  wire new_n9037_;
  wire or_not_new_n8995__1_not_new_n8799__1;
  wire not_new_n619__5;
  wire not_new_n4244_;
  wire not_new_n4542_;
  wire new_n6458_;
  wire not_new_n599__8235430;
  wire new_n1813_;
  wire new_n9760_;
  wire not_new_n5639_;
  wire new_n3963_;
  wire new_n6816_;
  wire or_not_new_n2769__not_new_n1476_;
  wire new_n10072_;
  wire not_new_n1071__6;
  wire not_new_n10344_;
  wire not_new_n581__2;
  wire not_pi137_2;
  wire new_n3884_;
  wire new_n2999_;
  wire or_not_new_n4827__not_new_n4799_;
  wire not_new_n7631__1;
  wire new_n6754_;
  wire not_new_n10297_;
  wire and_new_n6440__new_n6441_;
  wire not_new_n1940_;
  wire new_n8244_;
  wire not_new_n1047__10;
  wire new_n3187_;
  wire not_new_n5232_;
  wire not_new_n994__797922662976120010;
  wire not_new_n7523_;
  wire not_new_n1534__19773267430;
  wire new_n3350_;
  wire not_new_n5517_;
  wire not_new_n6587_;
  wire not_new_n620__1;
  wire not_new_n629__3430;
  wire not_new_n4399_;
  wire not_new_n1596__3430;
  wire not_new_n4678_;
  wire not_new_n3310__8235430;
  wire not_new_n1613__3;
  wire not_new_n9294_;
  wire new_n6177_;
  wire new_n1804_;
  wire not_new_n9273_;
  wire new_n4386_;
  wire or_or_or_not_new_n2785__not_new_n2788__not_new_n2787__not_new_n2789_;
  wire not_new_n6605_;
  wire not_new_n3051_;
  wire not_new_n5899__2;
  wire and_and_new_n6388__new_n6313__new_n6224_;
  wire not_new_n2249_;
  wire new_n7233_;
  wire new_n2428_;
  wire not_new_n3922_;
  wire not_new_n8494_;
  wire new_n5731_;
  wire or_or_not_new_n2053__not_new_n2054__not_new_n2056_;
  wire not_new_n8167__0;
  wire new_n4164_;
  wire not_new_n639__6;
  wire not_new_n1031__3;
  wire new_n10200_;
  wire not_new_n6547__0;
  wire and_new_n2632__new_n2631_;
  wire not_new_n4255_;
  wire not_new_n6370__0;
  wire not_new_n2097_;
  wire not_new_n8006_;
  wire new_n3015_;
  wire new_n9407_;
  wire not_new_n629__6782230728490;
  wire not_new_n9427_;
  wire not_new_n8129__1;
  wire new_n1719_;
  wire new_n2566_;
  wire not_pi148_2;
  wire new_n6408_;
  wire new_n4382_;
  wire new_n7337_;
  wire not_new_n631__0;
  wire new_n8859_;
  wire new_n7910_;
  wire not_new_n6741_;
  wire not_new_n8060_;
  wire not_pi213;
  wire not_pi050_0;
  wire and_new_n1575__new_n938_;
  wire not_new_n4837_;
  wire not_new_n4497_;
  wire not_new_n9855_;
  wire not_new_n7795_;
  wire new_n5847_;
  wire not_new_n9449_;
  wire or_or_not_new_n4234__not_new_n4336__not_new_n675_;
  wire not_new_n4899__1;
  wire new_n1576_;
  wire new_n1817_;
  wire not_new_n9349_;
  wire new_n6369_;
  wire not_new_n8922_;
  wire not_new_n7246_;
  wire not_new_n7805_;
  wire not_new_n4428__0;
  wire new_n6077_;
  wire not_new_n1057__6782230728490;
  wire new_n6422_;
  wire not_new_n3262_;
  wire not_new_n3339_;
  wire not_new_n2879_;
  wire not_new_n589__8;
  wire new_n6110_;
  wire not_new_n8237_;
  wire new_n8379_;
  wire new_n3887_;
  wire not_new_n5942_;
  wire new_n7404_;
  wire new_n2095_;
  wire new_n6384_;
  wire new_n8591_;
  wire not_new_n4262_;
  wire new_n9230_;
  wire not_new_n4643_;
  wire not_new_n5166__0;
  wire and_not_pi034_1_not_pi033_3;
  wire new_n8598_;
  wire not_new_n8433_;
  wire new_n2310_;
  wire new_n7654_;
  wire not_new_n4505_;
  wire not_new_n9638_;
  wire not_new_n10223_;
  wire not_new_n1177_;
  wire not_new_n1616__8235430;
  wire new_n4547_;
  wire not_new_n7689_;
  wire new_n1745_;
  wire new_n7869_;
  wire not_new_n586__2326305139872070;
  wire not_new_n6640_;
  wire not_new_n3494_;
  wire or_or_not_new_n6318__not_new_n6373__0_not_new_n6319_;
  wire not_new_n1037__2824752490;
  wire not_new_n989__10;
  wire new_n9816_;
  wire not_new_n9394__0;
  wire not_pi252;
  wire new_n7633_;
  wire new_n3990_;
  wire not_new_n3357_;
  wire new_n1608_;
  wire not_new_n4639_;
  wire new_n3989_;
  wire not_new_n2915_;
  wire new_n9651_;
  wire not_new_n620_;
  wire new_n3317_;
  wire not_new_n3547_;
  wire not_new_n1006__3;
  wire not_new_n1613__10;
  wire new_n5276_;
  wire po101;
  wire or_not_new_n5426__not_new_n605_;
  wire not_new_n8444_;
  wire not_pi186_0;
  wire not_new_n3185__6;
  wire not_new_n7027_;
  wire not_new_n637__138412872010;
  wire new_n6772_;
  wire not_new_n7744__0;
  wire not_new_n3509_;
  wire new_n2410_;
  wire not_new_n662_;
  wire not_new_n9647_;
  wire not_po298_490;
  wire new_n5931_;
  wire not_new_n1059__1;
  wire not_new_n598__24010;
  wire new_n3481_;
  wire new_n5178_;
  wire new_n8267_;
  wire new_n8008_;
  wire new_n8973_;
  wire not_new_n4624_;
  wire new_n9795_;
  wire new_n9276_;
  wire not_new_n9639_;
  wire not_new_n589__10;
  wire new_n8414_;
  wire not_new_n586__6782230728490;
  wire not_new_n3124_;
  wire not_new_n1043__3;
  wire not_new_n7627_;
  wire new_n6937_;
  wire not_new_n8145__0;
  wire new_n8949_;
  wire not_new_n6487__1;
  wire not_new_n1534__113988951853731430;
  wire not_new_n7416_;
  wire new_n5694_;
  wire or_not_new_n1596__3430_not_new_n5729_;
  wire new_n618_;
  wire po231;
  wire and_new_n2029__new_n2032_;
  wire not_new_n4205_;
  wire new_n10154_;
  wire or_not_new_n2783__not_new_n2782_;
  wire new_n7421_;
  wire not_new_n1059__70;
  wire not_new_n1602__9;
  wire not_new_n3134_;
  wire new_n5620_;
  wire not_new_n1304_;
  wire new_n4409_;
  wire not_new_n600__6782230728490;
  wire not_new_n9064_;
  wire not_new_n7484_;
  wire not_new_n633__332329305696010;
  wire new_n5942_;
  wire not_new_n5508__0;
  wire new_n7775_;
  wire not_new_n1007__5;
  wire not_new_n3354_;
  wire new_n5817_;
  wire not_new_n9334_;
  wire not_new_n5021_;
  wire not_new_n3315__19773267430;
  wire new_n9562_;
  wire not_pi131;
  wire new_n10170_;
  wire not_new_n625_;
  wire not_new_n5029_;
  wire not_new_n3400_;
  wire key_gate_52;
  wire new_n3001_;
  wire new_n4219_;
  wire new_n5797_;
  wire not_new_n611__6;
  wire not_new_n7354__2;
  wire new_n2063_;
  wire not_new_n1606__1;
  wire new_n3739_;
  wire not_new_n5113_;
  wire not_new_n628__490;
  wire not_new_n9462_;
  wire not_new_n6494__0;
  wire not_new_n7121_;
  wire new_n1710_;
  wire not_new_n1603__113988951853731430;
  wire not_new_n1534__47475615099430;
  wire not_new_n4369_;
  wire new_n4793_;
  wire not_new_n6657_;
  wire not_new_n9281_;
  wire not_new_n4127_;
  wire not_new_n4496__0;
  wire not_new_n593__70;
  wire not_new_n9442_;
  wire not_new_n585__3;
  wire new_n2629_;
  wire not_new_n9856_;
  wire not_new_n4785_;
  wire not_new_n1537__24010;
  wire not_new_n4971_;
  wire not_new_n6613__2;
  wire not_new_n7430_;
  wire new_n1543_;
  wire not_new_n3328_;
  wire new_n5562_;
  wire new_n1226_;
  wire new_n9596_;
  wire new_n5537_;
  wire not_new_n9456_;
  wire new_n7928_;
  wire new_n2737_;
  wire not_new_n3375_;
  wire new_n7367_;
  wire not_new_n632__19773267430;
  wire not_new_n2192_;
  wire new_n3200_;
  wire not_new_n9175_;
  wire new_n3834_;
  wire new_n5031_;
  wire new_n9782_;
  wire or_not_new_n9191__not_new_n9190_;
  wire new_n6236_;
  wire not_new_n5464_;
  wire new_n9180_;
  wire new_n4870_;
  wire not_new_n7045__0;
  wire new_n6829_;
  wire not_new_n5872_;
  wire new_n5248_;
  wire new_n3159_;
  wire not_new_n1596_;
  wire not_new_n1884_;
  wire not_new_n9094_;
  wire new_n3637_;
  wire not_new_n628__1915812313805664144010;
  wire new_n8410_;
  wire not_new_n1027__6782230728490;
  wire new_n7131_;
  wire po249;
  wire new_n1983_;
  wire not_new_n4774__0;
  wire new_n2400_;
  wire new_n6029_;
  wire new_n4519_;
  wire new_n4266_;
  wire not_new_n1576__797922662976120010;
  wire not_new_n4133_;
  wire not_new_n8045_;
  wire not_new_n7120_;
  wire not_new_n9820_;
  wire not_new_n994__2;
  wire new_n5380_;
  wire not_new_n6235__1;
  wire new_n4085_;
  wire new_n1970_;
  wire not_new_n599__4;
  wire not_new_n3755_;
  wire not_new_n5783__0;
  wire new_n7971_;
  wire or_or_not_new_n1825__not_new_n1826__not_new_n1828_;
  wire new_n2283_;
  wire not_new_n4195_;
  wire not_new_n5774__1;
  wire new_n6742_;
  wire not_new_n7668_;
  wire new_n9558_;
  wire not_new_n3372__13410686196639649008070;
  wire new_n1478_;
  wire not_new_n643__47475615099430;
  wire new_n752_;
  wire not_new_n624__403536070;
  wire not_new_n1053__4;
  wire not_new_n4459__0;
  wire not_new_n611__168070;
  wire not_new_n1020__1;
  wire new_n6021_;
  wire not_new_n5757__0;
  wire new_n2179_;
  wire new_n4282_;
  wire not_new_n8390_;
  wire new_n2669_;
  wire not_new_n595__24010;
  wire not_new_n1170__0;
  wire new_n3469_;
  wire new_n2332_;
  wire not_pi148;
  wire new_n2056_;
  wire not_new_n9841_;
  wire new_n6500_;
  wire not_new_n629__6;
  wire not_new_n1055__16284135979104490;
  wire not_new_n9997_;
  wire not_new_n9295_;
  wire new_n9222_;
  wire not_new_n9074_;
  wire not_new_n3403_;
  wire not_new_n1055__3;
  wire new_n4095_;
  wire not_new_n8224_;
  wire new_n5933_;
  wire not_new_n646__9;
  wire new_n3185_;
  wire new_n3489_;
  wire new_n7067_;
  wire not_new_n9206_;
  wire not_new_n9407__0;
  wire new_n609_;
  wire not_new_n984__16284135979104490;
  wire new_n3769_;
  wire new_n6219_;
  wire new_n5291_;
  wire new_n5727_;
  wire not_new_n8220_;
  wire new_n2738_;
  wire not_new_n1335_;
  wire or_not_new_n4837__not_new_n4772_;
  wire not_pi060_0;
  wire not_new_n9627__0;
  wire not_new_n7068_;
  wire new_n2610_;
  wire not_new_n1015__1;
  wire not_new_n1866_;
  wire new_n8078_;
  wire new_n3081_;
  wire not_new_n625__0;
  wire not_new_n1596__3;
  wire not_new_n1600__8235430;
  wire and_new_n9511__new_n9839_;
  wire new_n3442_;
  wire not_new_n1612__24010;
  wire new_n9415_;
  wire not_new_n644__2326305139872070;
  wire not_new_n2223__0;
  wire not_new_n8172__0;
  wire not_new_n1067__3430;
  wire or_not_new_n2749__not_new_n2752_;
  wire not_new_n640__6;
  wire not_new_n4724_;
  wire not_new_n4812__0;
  wire not_new_n631__3;
  wire new_n8152_;
  wire not_new_n8517_;
  wire not_new_n5989_;
  wire new_n4318_;
  wire new_n7365_;
  wire new_n1431_;
  wire not_new_n2226_;
  wire new_n5406_;
  wire or_or_not_new_n1279__not_new_n1277__not_new_n2021_;
  wire new_n2062_;
  wire new_n7324_;
  wire not_new_n6892_;
  wire not_new_n2983_;
  wire not_new_n1263_;
  wire new_n9968_;
  wire new_n3832_;
  wire new_n2068_;
  wire new_n2299_;
  wire not_new_n2977_;
  wire not_new_n1011_;
  wire new_n1261_;
  wire not_new_n8127__1;
  wire new_n5771_;
  wire new_n2271_;
  wire not_new_n5671_;
  wire new_n2272_;
  wire not_new_n590__0;
  wire new_n9039_;
  wire not_new_n6622__0;
  wire not_pi081;
  wire new_n9548_;
  wire not_new_n7404_;
  wire not_new_n9002__0;
  wire not_new_n6542_;
  wire not_new_n3945_;
  wire not_new_n8643_;
  wire new_n5652_;
  wire new_n3330_;
  wire new_n9173_;
  wire not_new_n5504__0;
  wire not_new_n6540__0;
  wire new_n688_;
  wire not_new_n596__70;
  wire not_new_n9066_;
  wire not_new_n1502_;
  wire not_pi269_3;
  wire not_new_n3289_;
  wire not_new_n8079_;
  wire not_new_n608__57648010;
  wire po103;
  wire not_new_n2980_;
  wire not_new_n1039__16284135979104490;
  wire not_new_n1487_;
  wire new_n5475_;
  wire not_new_n5926_;
  wire new_n7895_;
  wire new_n4857_;
  wire not_new_n1525_;
  wire new_n6951_;
  wire new_n1570_;
  wire not_new_n1071__47475615099430;
  wire not_new_n618__225393402906922580878632490;
  wire not_new_n1051__968890104070;
  wire not_new_n7979_;
  wire not_new_n647__6;
  wire new_n2925_;
  wire new_n4770_;
  wire not_new_n4606_;
  wire not_new_n602__4;
  wire new_n8822_;
  wire new_n5923_;
  wire not_new_n7944_;
  wire not_new_n586__3430;
  wire not_new_n2947_;
  wire new_n9642_;
  wire new_n3800_;
  wire new_n3523_;
  wire and_new_n2359__new_n2358_;
  wire new_n2954_;
  wire not_new_n9641_;
  wire not_new_n3893_;
  wire not_new_n635__47475615099430;
  wire new_n2347_;
  wire new_n1671_;
  wire not_pi044_0;
  wire new_n8328_;
  wire not_new_n7222__0;
  wire new_n1395_;
  wire new_n9861_;
  wire not_new_n3575_;
  wire new_n9522_;
  wire new_n2648_;
  wire not_new_n1559_;
  wire not_pi124;
  wire not_new_n4483__0;
  wire not_new_n649__0;
  wire not_new_n6453_;
  wire not_new_n7023__0;
  wire not_new_n6292_;
  wire new_n3994_;
  wire new_n6539_;
  wire not_new_n1604__1176490;
  wire not_new_n3979__0;
  wire new_n4036_;
  wire new_n6805_;
  wire new_n6655_;
  wire new_n6730_;
  wire not_new_n4799_;
  wire new_n9604_;
  wire not_new_n624__138412872010;
  wire not_new_n8126__0;
  wire not_new_n1493_;
  wire new_n5063_;
  wire not_new_n7015__0;
  wire not_new_n4134__2;
  wire new_n3278_;
  wire new_n7234_;
  wire new_n1742_;
  wire not_new_n4445_;
  wire not_new_n989__3;
  wire new_n7967_;
  wire not_new_n585__403536070;
  wire not_new_n8171__0;
  wire new_n5453_;
  wire not_new_n5035_;
  wire not_new_n8551_;
  wire new_n4823_;
  wire po033;
  wire not_new_n2944_;
  wire not_new_n772_;
  wire not_new_n5673_;
  wire not_new_n4632_;
  wire not_new_n9631__0;
  wire new_n964_;
  wire not_new_n1631__1;
  wire not_new_n1728__797922662976120010;
  wire new_n583_;
  wire or_or_not_new_n1406__not_new_n1407__not_new_n1410_;
  wire not_new_n1027__6;
  wire not_new_n596__403536070;
  wire not_new_n4555_;
  wire po021;
  wire not_new_n8352_;
  wire new_n5378_;
  wire new_n8047_;
  wire new_n8565_;
  wire new_n7968_;
  wire not_new_n596__16284135979104490;
  wire not_new_n8440_;
  wire new_n9450_;
  wire new_n1693_;
  wire not_new_n1699_;
  wire new_n7479_;
  wire not_new_n604__5;
  wire not_new_n2837_;
  wire not_pi047;
  wire new_n9208_;
  wire not_new_n636__2326305139872070;
  wire new_n647_;
  wire not_new_n6794_;
  wire new_n8150_;
  wire new_n3863_;
  wire new_n2237_;
  wire new_n7431_;
  wire not_po296_39098210485829880490;
  wire new_n7345_;
  wire new_n8720_;
  wire and_new_n2672__new_n2671_;
  wire not_new_n5091_;
  wire new_n8650_;
  wire not_new_n8264__1;
  wire not_new_n3557_;
  wire not_new_n5628_;
  wire not_new_n4449_;
  wire not_new_n7366__2;
  wire and_and_new_n2295__new_n2298__new_n2296_;
  wire not_new_n1057__10;
  wire not_new_n608__6;
  wire new_n7414_;
  wire not_new_n4561_;
  wire new_n2489_;
  wire new_n5922_;
  wire not_new_n4166__0;
  wire not_new_n2705_;
  wire new_n9843_;
  wire new_n10089_;
  wire new_n4532_;
  wire new_n5888_;
  wire not_new_n5607_;
  wire not_new_n1031__57648010;
  wire not_new_n1005__1;
  wire not_new_n8142__0;
  wire and_and_new_n1750__new_n1751__new_n1753_;
  wire new_n4727_;
  wire not_new_n4492_;
  wire new_n2884_;
  wire new_n3844_;
  wire not_new_n9539_;
  wire new_n1516_;
  wire not_new_n4196_;
  wire not_new_n1616__6782230728490;
  wire not_new_n7365_;
  wire not_new_n1005__5;
  wire not_new_n9827_;
  wire not_new_n4980__0;
  wire new_n3968_;
  wire new_n4279_;
  wire not_new_n5830_;
  wire not_new_n8136__0;
  wire not_new_n4977_;
  wire key_gate_41;
  wire new_n8540_;
  wire po223;
  wire new_n3408_;
  wire or_or_not_new_n1291__not_new_n1289__not_new_n2078_;
  wire new_n3407_;
  wire new_n972_;
  wire and_new_n6373__new_n6401_;
  wire new_n6400_;
  wire new_n8289_;
  wire new_n7347_;
  wire not_new_n8623_;
  wire not_new_n10285_;
  wire not_new_n5955_;
  wire new_n2567_;
  wire new_n2869_;
  wire new_n2255_;
  wire new_n8689_;
  wire not_new_n621__5;
  wire new_n6549_;
  wire not_new_n1400_;
  wire not_new_n5962_;
  wire not_new_n984__797922662976120010;
  wire not_new_n6443__2;
  wire new_n3334_;
  wire not_pi233;
  wire not_new_n6508__1;
  wire not_new_n6236_;
  wire not_new_n6800_;
  wire not_new_n9006_;
  wire not_new_n7399_;
  wire new_n7784_;
  wire not_new_n6563_;
  wire not_new_n3113_;
  wire not_new_n597__3430;
  wire new_n5021_;
  wire not_pi038_2;
  wire new_n9887_;
  wire not_new_n619__70;
  wire not_new_n4273_;
  wire new_n8323_;
  wire not_new_n3815_;
  wire new_n4674_;
  wire not_new_n648__2326305139872070;
  wire po082;
  wire not_new_n7035_;
  wire not_new_n4429_;
  wire not_new_n5249_;
  wire new_n6741_;
  wire new_n3145_;
  wire not_new_n1538__57648010;
  wire new_n5780_;
  wire not_new_n2965_;
  wire not_new_n7909_;
  wire new_n2203_;
  wire not_new_n6514_;
  wire not_new_n9361_;
  wire new_n9245_;
  wire new_n1006_;
  wire or_or_not_new_n1564__not_new_n2479__not_new_n1397_;
  wire not_new_n8977_;
  wire new_n5034_;
  wire new_n9992_;
  wire not_new_n643__403536070;
  wire not_new_n5203_;
  wire new_n7401_;
  wire not_new_n5325_;
  wire not_new_n6487__0;
  wire not_new_n9916__0;
  wire not_new_n622__6;
  wire new_n5284_;
  wire not_new_n1603__16284135979104490;
  wire not_new_n8505_;
  wire not_new_n604__2824752490;
  wire not_new_n3375__2;
  wire new_n2184_;
  wire new_n3575_;
  wire not_new_n7769_;
  wire not_new_n1041__2;
  wire and_new_n1306__new_n2160_;
  wire not_new_n9252_;
  wire not_new_n8636_;
  wire and_new_n3067__new_n998_;
  wire new_n2956_;
  wire not_new_n581__185621159210175743024531636712070;
  wire or_not_new_n4322__0_not_new_n680__0;
  wire new_n5264_;
  wire new_n5448_;
  wire not_new_n7353_;
  wire not_new_n598__3;
  wire new_n8413_;
  wire not_new_n1185_;
  wire not_new_n8880_;
  wire new_n7890_;
  wire not_new_n5010_;
  wire not_new_n6574_;
  wire new_n1907_;
  wire not_new_n647__16284135979104490;
  wire or_not_new_n1482__not_new_n2858_;
  wire not_new_n5065_;
  wire new_n3910_;
  wire not_new_n632__0;
  wire new_n2784_;
  wire not_new_n1382_;
  wire new_n9808_;
  wire not_new_n3468_;
  wire new_n2409_;
  wire new_n6130_;
  wire not_new_n1594__57648010;
  wire new_n3104_;
  wire new_n4310_;
  wire new_n2882_;
  wire not_new_n5898_;
  wire not_new_n1537__138412872010;
  wire not_new_n608__3430;
  wire not_new_n3571_;
  wire new_n4812_;
  wire new_n9239_;
  wire new_n1877_;
  wire not_new_n3995_;
  wire new_n6179_;
  wire not_new_n10270_;
  wire not_new_n2914_;
  wire not_new_n3487_;
  wire key_gate_106;
  wire not_new_n8226_;
  wire new_n3828_;
  wire not_new_n5533_;
  wire not_new_n6213_;
  wire not_new_n636__332329305696010;
  wire not_new_n1039_;
  wire not_new_n2603_;
  wire not_new_n3478_;
  wire new_n2932_;
  wire new_n731_;
  wire or_or_not_new_n1556__not_new_n2439__not_new_n1381_;
  wire not_new_n10230_;
  wire new_n2531_;
  wire not_new_n5391_;
  wire not_new_n3533_;
  wire or_or_not_new_n2955__not_new_n2958__not_new_n2957_;
  wire new_n2342_;
  wire not_new_n1394_;
  wire new_n8679_;
  wire new_n2819_;
  wire new_n5610_;
  wire not_new_n1933_;
  wire not_new_n8171__1;
  wire new_n8293_;
  wire new_n3375_;
  wire new_n7659_;
  wire not_new_n2551_;
  wire new_n10030_;
  wire not_new_n4019__0;
  wire not_pi169_2;
  wire not_new_n3365_;
  wire new_n9621_;
  wire not_new_n3935_;
  wire not_new_n4938_;
  wire not_new_n9396_;
  wire new_n1178_;
  wire not_pi192;
  wire not_new_n2973_;
  wire key_gate_72;
  wire not_new_n2928_;
  wire not_pi146_1;
  wire not_new_n1612__5;
  wire new_n3809_;
  wire not_new_n587__0;
  wire not_new_n9483_;
  wire not_new_n594__2824752490;
  wire new_n5443_;
  wire new_n3120_;
  wire not_new_n667_;
  wire new_n6091_;
  wire new_n8488_;
  wire new_n1784_;
  wire not_new_n622__24010;
  wire not_new_n1597__332329305696010;
  wire new_n5173_;
  wire new_n5534_;
  wire new_n2744_;
  wire not_new_n5239_;
  wire new_n1422_;
  wire not_new_n8395_;
  wire new_n1563_;
  wire new_n10075_;
  wire new_n3193_;
  wire not_new_n1174_;
  wire not_new_n7202_;
  wire not_new_n6065_;
  wire new_n4856_;
  wire not_new_n9524_;
  wire not_new_n774_;
  wire not_new_n6695_;
  wire not_new_n6654__0;
  wire not_new_n7651__0;
  wire not_new_n3410_;
  wire not_new_n1155_;
  wire not_new_n7502_;
  wire not_new_n718__2;
  wire not_new_n1037__16284135979104490;
  wire new_n9668_;
  wire new_n4722_;
  wire po065;
  wire not_new_n5897_;
  wire not_new_n3589_;
  wire not_new_n1404_;
  wire not_new_n634__403536070;
  wire new_n9636_;
  wire not_new_n6907_;
  wire not_new_n9308_;
  wire not_new_n3523_;
  wire not_new_n1261_;
  wire new_n2516_;
  wire new_n7655_;
  wire not_new_n5160_;
  wire new_n5637_;
  wire new_n7021_;
  wire not_new_n10202_;
  wire new_n2650_;
  wire not_new_n600_;
  wire not_new_n3465_;
  wire not_new_n2016_;
  wire not_new_n4943_;
  wire new_n4864_;
  wire new_n5065_;
  wire new_n1250_;
  wire not_new_n8709_;
  wire not_new_n8164__0;
  wire not_new_n648__16284135979104490;
  wire new_n5644_;
  wire po012;
  wire not_new_n9722_;
  wire new_n6242_;
  wire new_n9320_;
  wire new_n6728_;
  wire not_new_n619__4;
  wire not_new_n7839_;
  wire not_new_n1537__0;
  wire new_n6331_;
  wire not_new_n7081_;
  wire not_new_n4586_;
  wire new_n5814_;
  wire new_n10037_;
  wire new_n3309_;
  wire new_n3428_;
  wire not_new_n608__1;
  wire not_new_n645__7;
  wire new_n6194_;
  wire not_new_n1537__6;
  wire new_n6085_;
  wire not_new_n8394_;
  wire not_new_n1498_;
  wire not_new_n9985_;
  wire new_n7732_;
  wire not_new_n6233__1;
  wire new_n677_;
  wire new_n9201_;
  wire not_new_n7864_;
  wire new_n7352_;
  wire new_n6196_;
  wire new_n9894_;
  wire not_new_n3185_;
  wire new_n4816_;
  wire not_new_n9779_;
  wire not_new_n3536_;
  wire not_new_n1005__7;
  wire not_new_n8069_;
  wire not_new_n634__16284135979104490;
  wire not_new_n4193_;
  wire new_n3770_;
  wire not_new_n1580__8;
  wire not_new_n6232__3;
  wire new_n10287_;
  wire not_pi008;
  wire new_n9351_;
  wire not_new_n6633_;
  wire not_new_n959_;
  wire not_new_n4279_;
  wire not_new_n5939_;
  wire not_po298_47475615099430;
  wire not_new_n4475__0;
  wire not_new_n1041__8;
  wire new_n1523_;
  wire or_or_not_new_n1567__not_new_n2494__not_new_n1403_;
  wire not_new_n4164_;
  wire not_new_n1602__8;
  wire new_n8907_;
  wire new_n6879_;
  wire new_n6568_;
  wire not_new_n600__332329305696010;
  wire new_n6336_;
  wire new_n8039_;
  wire new_n7536_;
  wire not_new_n1388_;
  wire new_n4908_;
  wire not_new_n9102_;
  wire not_new_n3372__3430;
  wire not_new_n5741__0;
  wire new_n10316_;
  wire key_gate_9;
  wire not_new_n605__3430;
  wire po176;
  wire not_new_n8861_;
  wire new_n10230_;
  wire new_n6982_;
  wire new_n8360_;
  wire new_n4355_;
  wire not_new_n8556_;
  wire not_new_n5770__1;
  wire key_gate_23;
  wire not_new_n599__2;
  wire new_n9184_;
  wire or_not_new_n4234__not_new_n4336_;
  wire not_new_n1059__8;
  wire not_new_n1051__3;
  wire not_new_n6997__0;
  wire new_n3335_;
  wire not_new_n10128_;
  wire not_pi219;
  wire not_pi041_0;
  wire not_po296_5;
  wire not_new_n1159__1;
  wire not_new_n1481_;
  wire not_pi171_0;
  wire not_new_n597__490;
  wire new_n5025_;
  wire not_new_n627__3430;
  wire not_new_n1005__0;
  wire new_n5234_;
  wire new_n9991_;
  wire new_n1961_;
  wire new_n6796_;
  wire new_n1180_;
  wire not_new_n7251_;
  wire not_new_n1622__0;
  wire not_new_n8391_;
  wire new_n6201_;
  wire new_n7889_;
  wire not_new_n4103_;
  wire not_new_n7047__0;
  wire not_new_n5760__0;
  wire not_new_n3957_;
  wire new_n1633_;
  wire or_not_new_n5460__not_new_n5686__1;
  wire not_new_n6887_;
  wire new_n5097_;
  wire new_n5485_;
  wire not_new_n8995__1;
  wire new_n4491_;
  wire new_n6128_;
  wire new_n6334_;
  wire not_new_n621__273687473400809163430;
  wire new_n3529_;
  wire new_n4372_;
  wire new_n9314_;
  wire new_n756_;
  wire not_new_n8969_;
  wire not_new_n10255_;
  wire new_n1568_;
  wire not_new_n8680_;
  wire new_n3332_;
  wire not_pi064_797922662976120010;
  wire not_new_n3310__24010;
  wire not_new_n7071_;
  wire new_n8583_;
  wire new_n7300_;
  wire not_new_n9408_;
  wire not_new_n9116_;
  wire not_new_n5754__1;
  wire not_new_n4978__0;
  wire new_n8544_;
  wire not_new_n645__138412872010;
  wire not_new_n4787__0;
  wire not_new_n6855_;
  wire new_n1200_;
  wire not_new_n2938_;
  wire not_new_n7601__0;
  wire not_new_n619__3;
  wire not_new_n5254_;
  wire not_new_n928_;
  wire not_new_n9060_;
  wire not_new_n4096_;
  wire not_pi167;
  wire not_new_n5912__0;
  wire key_gate_69;
  wire new_n7445_;
  wire new_n1734_;
  wire not_new_n7937_;
  wire not_new_n984__70;
  wire and_new_n2238__new_n2241_;
  wire new_n1047_;
  wire new_n2466_;
  wire new_n7364_;
  wire not_new_n6487_;
  wire new_n2923_;
  wire new_n1375_;
  wire not_new_n6373__1;
  wire not_pi088;
  wire new_n8958_;
  wire not_new_n9253_;
  wire new_n4690_;
  wire not_new_n1055__4;
  wire not_new_n5136_;
  wire not_new_n2601_;
  wire new_n6905_;
  wire not_new_n3700_;
  wire not_new_n4019__1;
  wire not_pi206;
  wire not_pi130_1;
  wire not_new_n638__403536070;
  wire new_n695_;
  wire not_new_n8707__0;
  wire new_n5986_;
  wire or_not_new_n2585__not_new_n2584_;
  wire new_n6075_;
  wire not_new_n5251_;
  wire new_n1001_;
  wire not_new_n1863_;
  wire not_new_n3444_;
  wire new_n9945_;
  wire not_pi047_1;
  wire not_new_n7338_;
  wire new_n6736_;
  wire not_pi133_2;
  wire new_n6548_;
  wire new_n10149_;
  wire not_new_n7767_;
  wire new_n2504_;
  wire not_new_n1047__24010;
  wire new_n4094_;
  wire new_n7524_;
  wire new_n4983_;
  wire not_new_n6239_;
  wire not_new_n2841_;
  wire new_n10155_;
  wire new_n1717_;
  wire not_new_n611__490;
  wire new_n3498_;
  wire not_new_n1606__0;
  wire new_n9524_;
  wire new_n5609_;
  wire not_new_n1603__168070;
  wire not_new_n4768_;
  wire not_new_n597__2;
  wire not_new_n5617_;
  wire new_n2845_;
  wire not_new_n2509__24010;
  wire new_n2415_;
  wire new_n2858_;
  wire not_new_n1057__1;
  wire new_n7384_;
  wire not_new_n1599__168070;
  wire not_new_n1601__1915812313805664144010;
  wire not_new_n4774_;
  wire new_n6795_;
  wire not_new_n10220_;
  wire not_new_n3552_;
  wire not_new_n611__2824752490;
  wire not_new_n630__3;
  wire new_n1207_;
  wire not_new_n7504_;
  wire not_new_n2188_;
  wire new_n9821_;
  wire new_n6853_;
  wire not_new_n596__4;
  wire not_new_n4315_;
  wire new_n7888_;
  wire new_n1420_;
  wire not_new_n595_;
  wire not_new_n5788__0;
  wire new_n1315_;
  wire new_n8751_;
  wire new_n5856_;
  wire new_n1905_;
  wire not_new_n1599__5;
  wire not_new_n8232_;
  wire new_n7020_;
  wire not_new_n4556_;
  wire new_n3298_;
  wire not_new_n644__2;
  wire not_pi260_1;
  wire new_n1612_;
  wire not_new_n8793_;
  wire not_new_n634__968890104070;
  wire not_new_n9672_;
  wire not_new_n10232_;
  wire new_n1493_;
  wire not_new_n5863_;
  wire not_new_n3866_;
  wire not_new_n1605__0;
  wire not_pi250_0;
  wire new_n6000_;
  wire new_n2633_;
  wire new_n9381_;
  wire new_n3919_;
  wire new_n9880_;
  wire not_new_n5511__0;
  wire not_new_n2169_;
  wire new_n6554_;
  wire not_new_n1613__5;
  wire not_new_n5916_;
  wire new_n8775_;
  wire not_new_n7663__0;
  wire not_new_n1049__47475615099430;
  wire not_new_n643_;
  wire new_n7745_;
  wire not_new_n1611__70;
  wire not_pi232;
  wire not_new_n7644_;
  wire new_n7378_;
  wire not_new_n4128__2;
  wire not_new_n5749_;
  wire not_new_n623__0;
  wire not_new_n3689_;
  wire not_new_n598__19773267430;
  wire not_new_n604__47475615099430;
  wire not_new_n8462_;
  wire not_new_n7293__0;
  wire new_n9229_;
  wire new_n6126_;
  wire new_n5547_;
  wire not_new_n4150_;
  wire not_new_n7003__1;
  wire new_n2652_;
  wire not_new_n9703_;
  wire not_new_n9747_;
  wire not_new_n5553_;
  wire not_new_n637__6782230728490;
  wire not_pi134_1;
  wire new_n4776_;
  wire new_n3524_;
  wire not_new_n7334__0;
  wire not_new_n6132_;
  wire not_new_n7855_;
  wire or_not_new_n5764__0_not_new_n618__8235430;
  wire not_new_n611__3;
  wire not_new_n625__24010;
  wire not_new_n1532_;
  wire not_new_n966_;
  wire new_n1151_;
  wire not_new_n1059__3;
  wire not_new_n5901_;
  wire new_n3944_;
  wire not_new_n1602__3;
  wire not_new_n7567_;
  wire not_new_n8106_;
  wire new_n10269_;
  wire new_n8097_;
  wire not_new_n1385_;
  wire not_new_n8575_;
  wire new_n3814_;
  wire new_n4849_;
  wire not_new_n1612__8235430;
  wire not_new_n7991_;
  wire new_n601_;
  wire and_new_n2647__new_n2648_;
  wire new_n9293_;
  wire new_n3013_;
  wire not_pi144_3;
  wire not_new_n3464_;
  wire not_new_n9610_;
  wire not_new_n2845_;
  wire new_n1812_;
  wire new_n9608_;
  wire po126;
  wire not_new_n2787_;
  wire new_n7062_;
  wire new_n2371_;
  wire not_new_n8984_;
  wire po238;
  wire not_new_n6854_;
  wire not_new_n3950_;
  wire not_new_n9427__3;
  wire not_new_n620__2;
  wire new_n8806_;
  wire new_n6078_;
  wire not_new_n2299_;
  wire not_new_n5159__0;
  wire not_pi142_1;
  wire not_new_n7517_;
  wire not_new_n7612__0;
  wire not_new_n8804_;
  wire not_new_n5388_;
  wire new_n3354_;
  wire new_n9599_;
  wire not_new_n1609__1;
  wire new_n4420_;
  wire new_n5733_;
  wire new_n5421_;
  wire new_n1427_;
  wire new_n7100_;
  wire not_new_n1589__6782230728490;
  wire not_new_n640__2824752490;
  wire not_new_n2848_;
  wire not_new_n624__2824752490;
  wire not_new_n3722_;
  wire not_new_n6982_;
  wire new_n8386_;
  wire new_n1241_;
  wire new_n2141_;
  wire not_new_n3372__9;
  wire not_new_n7646__0;
  wire not_new_n636__403536070;
  wire not_new_n5771_;
  wire not_new_n1594__1176490;
  wire not_new_n4167__0;
  wire new_n5984_;
  wire or_not_new_n2535__not_new_n2534_;
  wire not_new_n9888__1;
  wire new_n9326_;
  wire new_n3160_;
  wire not_pi166_2;
  wire new_n1538_;
  wire not_new_n4749__0;
  wire or_not_new_n8139__1_not_new_n8231_;
  wire not_new_n10102_;
  wire key_gate_111;
  wire new_n8193_;
  wire not_new_n5535_;
  wire not_new_n9783_;
  wire or_not_new_n1027__0_not_new_n3384_;
  wire not_new_n686_;
  wire not_new_n3664_;
  wire new_n5423_;
  wire not_new_n4628_;
  wire new_n6892_;
  wire not_new_n628__8235430;
  wire not_new_n597__16284135979104490;
  wire not_new_n8262_;
  wire new_n10011_;
  wire not_new_n8557_;
  wire new_n8221_;
  wire not_new_n621__6782230728490;
  wire not_new_n1037__490;
  wire not_new_n1157_;
  wire new_n5938_;
  wire new_n7289_;
  wire not_new_n6502_;
  wire not_new_n624__332329305696010;
  wire new_n3228_;
  wire not_new_n4294_;
  wire new_n9872_;
  wire not_new_n9341_;
  wire not_new_n7759__0;
  wire not_new_n587__4;
  wire not_new_n9045_;
  wire new_n4171_;
  wire not_new_n617__5;
  wire not_new_n5680__1;
  wire new_n5543_;
  wire not_new_n5129_;
  wire new_n8130_;
  wire new_n5882_;
  wire or_or_or_not_new_n2838__not_new_n2841__not_new_n2840__not_new_n2842_;
  wire not_new_n644__1176490;
  wire not_new_n626__9;
  wire new_n757_;
  wire not_new_n7183_;
  wire not_new_n1476_;
  wire not_new_n621__2;
  wire new_n6153_;
  wire not_new_n5753_;
  wire not_new_n10241_;
  wire new_n7146_;
  wire not_new_n1581__4;
  wire new_n1775_;
  wire new_n8073_;
  wire not_new_n4071__1;
  wire new_n4374_;
  wire new_n4099_;
  wire new_n7798_;
  wire not_new_n9890__0;
  wire not_new_n1057__0;
  wire not_new_n1776_;
  wire not_new_n10156_;
  wire not_new_n644__57648010;
  wire not_new_n6443__168070;
  wire not_new_n1043_;
  wire or_or_not_new_n2831__not_new_n1481__not_new_n2830_;
  wire new_n2212_;
  wire po215;
  wire not_new_n4198_;
  wire new_n6966_;
  wire new_n5857_;
  wire not_new_n7406__0;
  wire not_new_n6318_;
  wire new_n7024_;
  wire not_new_n5484__0;
  wire and_new_n2162__new_n2165_;
  wire not_new_n1585__19773267430;
  wire not_new_n603__3430;
  wire not_new_n617__6;
  wire not_new_n1152_;
  wire not_new_n2287_;
  wire new_n6555_;
  wire not_new_n4183_;
  wire po163;
  wire new_n9446_;
  wire not_new_n3311__490;
  wire new_n5193_;
  wire and_new_n6316__new_n6227_;
  wire new_n6998_;
  wire not_new_n5016_;
  wire new_n9794_;
  wire new_n4628_;
  wire not_new_n621__7;
  wire po254;
  wire or_not_new_n9855__0_not_new_n10046__0;
  wire not_new_n8003_;
  wire not_new_n1162_;
  wire new_n7560_;
  wire not_new_n1236_;
  wire not_new_n8091_;
  wire not_new_n6690_;
  wire not_new_n6084_;
  wire not_pi038_0;
  wire not_new_n589__24010;
  wire not_new_n599__2824752490;
  wire not_new_n9066__0;
  wire not_new_n6974__332329305696010;
  wire new_n1288_;
  wire not_new_n646__6;
  wire not_pi147_1;
  wire and_and_and_new_n6385__new_n6386__new_n6241__new_n6375_;
  wire not_new_n2909_;
  wire not_new_n9123_;
  wire not_new_n2900_;
  wire new_n5288_;
  wire not_pi039_0;
  wire new_n7881_;
  wire not_new_n6336_;
  wire not_new_n5051_;
  wire new_n9268_;
  wire not_new_n9649_;
  wire new_n3630_;
  wire new_n8178_;
  wire not_new_n643__138412872010;
  wire not_new_n3225_;
  wire not_new_n6590_;
  wire new_n4292_;
  wire not_new_n1198_;
  wire not_new_n1906_;
  wire po029;
  wire not_new_n4152_;
  wire not_new_n588__2;
  wire new_n9165_;
  wire not_new_n10292_;
  wire not_new_n718__1;
  wire not_new_n8210_;
  wire new_n3694_;
  wire new_n10053_;
  wire not_new_n630__168070;
  wire new_n1505_;
  wire not_new_n5209_;
  wire or_not_new_n4899__0_not_new_n5096__0;
  wire not_new_n4833__0;
  wire not_new_n4992_;
  wire not_new_n8401_;
  wire new_n9553_;
  wire not_new_n639__57648010;
  wire key_gate_88;
  wire not_new_n637__3430;
  wire new_n1447_;
  wire new_n6472_;
  wire not_new_n7684_;
  wire not_new_n1057__1176490;
  wire new_n2667_;
  wire not_new_n8850__0;
  wire new_n3665_;
  wire not_pi180_2;
  wire or_or_not_new_n2497__not_new_n1568__not_new_n2498_;
  wire new_n1539_;
  wire not_new_n5773__0;
  wire not_new_n5882__2;
  wire not_new_n581__8235430;
  wire not_new_n6655_;
  wire not_new_n4473_;
  wire not_new_n588__10;
  wire new_n1615_;
  wire new_n2222_;
  wire new_n8065_;
  wire not_new_n1065__3430;
  wire not_new_n1508_;
  wire not_new_n5770__2;
  wire not_new_n3358_;
  wire not_new_n1607__10;
  wire or_not_new_n2525__not_new_n2524_;
  wire new_n8006_;
  wire new_n1930_;
  wire not_new_n1369_;
  wire not_new_n1534__57648010;
  wire not_new_n1069__9;
  wire new_n2888_;
  wire not_new_n1581__8235430;
  wire not_new_n4941_;
  wire new_n8474_;
  wire not_new_n7451_;
  wire new_n5971_;
  wire not_new_n643__16284135979104490;
  wire not_new_n1037__1;
  wire new_n2446_;
  wire or_not_new_n6339__not_new_n6232__1;
  wire not_new_n9416_;
  wire not_new_n9174_;
  wire not_new_n7737_;
  wire not_new_n8040_;
  wire not_po298_16284135979104490;
  wire new_n6956_;
  wire not_new_n9778_;
  wire not_new_n3894_;
  wire not_new_n581__11044276742439206463052992010;
  wire new_n5483_;
  wire new_n9274_;
  wire not_new_n4491__0;
  wire not_new_n3701_;
  wire new_n5492_;
  wire not_new_n4437_;
  wire and_new_n2702__new_n2701_;
  wire not_new_n1063__2824752490;
  wire new_n1238_;
  wire not_new_n598__8235430;
  wire not_new_n5918__0;
  wire new_n6584_;
  wire not_new_n4536_;
  wire not_new_n7542_;
  wire not_new_n642__0;
  wire not_po296_24010;
  wire or_not_new_n2919__not_new_n2922_;
  wire not_new_n8953_;
  wire not_new_n2547_;
  wire not_new_n638__4;
  wire not_new_n6319_;
  wire new_n3885_;
  wire new_n8657_;
  wire new_n6685_;
  wire not_new_n7815_;
  wire new_n3880_;
  wire new_n2604_;
  wire new_n6724_;
  wire not_new_n636_;
  wire not_new_n4493_;
  wire not_pi049;
  wire not_pi227;
  wire not_new_n7898_;
  wire new_n7182_;
  wire new_n8581_;
  wire not_new_n3155_;
  wire new_n5906_;
  wire new_n10198_;
  wire new_n8927_;
  wire and_new_n2384__new_n2383_;
  wire not_new_n638__32199057558131797268376070;
  wire not_new_n589__7;
  wire not_new_n5902_;
  wire new_n8113_;
  wire new_n3714_;
  wire new_n7844_;
  wire not_new_n3184__2326305139872070;
  wire not_new_n646__8;
  wire not_new_n5584_;
  wire new_n5961_;
  wire or_not_new_n2740__not_new_n2743_;
  wire new_n4405_;
  wire not_new_n941__0;
  wire not_new_n8389_;
  wire new_n7126_;
  wire not_new_n4490__0;
  wire not_new_n5974_;
  wire not_new_n1604__70;
  wire not_new_n6496__0;
  wire new_n764_;
  wire not_new_n1601__8235430;
  wire not_new_n1342_;
  wire not_new_n581__657123623635342801395430;
  wire new_n8295_;
  wire not_pi105;
  wire not_new_n5783_;
  wire not_new_n7270_;
  wire not_new_n8278_;
  wire not_new_n1591__19773267430;
  wire not_new_n586__47475615099430;
  wire and_new_n934__new_n986_;
  wire not_new_n1843_;
  wire not_new_n1599__1;
  wire not_new_n8372_;
  wire new_n4525_;
  wire new_n9624_;
  wire not_new_n3380_;
  wire not_new_n1585__332329305696010;
  wire new_n6149_;
  wire or_not_new_n6335__not_new_n6373__4;
  wire not_new_n8712_;
  wire not_pi269_1;
  wire new_n655_;
  wire not_new_n4132__2;
  wire new_n10153_;
  wire not_new_n6085_;
  wire new_n626_;
  wire not_new_n6674_;
  wire new_n988_;
  wire not_new_n642__57648010;
  wire not_new_n4945__0;
  wire not_new_n5382_;
  wire not_new_n8622_;
  wire not_new_n7001__0;
  wire not_pi054_3;
  wire new_n8586_;
  wire new_n8554_;
  wire new_n4851_;
  wire not_new_n5155_;
  wire new_n4267_;
  wire new_n5624_;
  wire new_n9556_;
  wire not_pi161_3;
  wire new_n7331_;
  wire not_new_n994__6;
  wire new_n4875_;
  wire po063;
  wire new_n8033_;
  wire new_n4391_;
  wire new_n2109_;
  wire new_n2715_;
  wire not_new_n4014__0;
  wire new_n1159_;
  wire not_new_n8111_;
  wire new_n2043_;
  wire not_new_n9197_;
  wire not_new_n5766__1;
  wire new_n2513_;
  wire not_new_n2761_;
  wire not_new_n8814_;
  wire new_n1645_;
  wire new_n8917_;
  wire new_n6668_;
  wire not_new_n6647_;
  wire not_new_n9307_;
  wire or_not_new_n2227__not_new_n2224_;
  wire not_new_n643__1176490;
  wire not_new_n6707_;
  wire new_n1890_;
  wire new_n4659_;
  wire new_n2591_;
  wire not_new_n5922_;
  wire not_new_n8247_;
  wire not_new_n6489_;
  wire new_n9393_;
  wire new_n4804_;
  wire not_new_n7225_;
  wire or_not_new_n6349__not_new_n6373__7;
  wire not_new_n4634_;
  wire new_n5129_;
  wire new_n9620_;
  wire or_not_new_n8411__not_new_n8293_;
  wire not_new_n8155__1;
  wire not_new_n1027__797922662976120010;
  wire not_new_n1550_;
  wire not_new_n7595_;
  wire not_new_n6527__2;
  wire new_n6594_;
  wire new_n5398_;
  wire not_new_n4085_;
  wire not_new_n6327_;
  wire not_new_n7117_;
  wire not_new_n1728__1;
  wire new_n3938_;
  wire new_n7012_;
  wire not_pi248;
  wire not_pi010_0;
  wire new_n2169_;
  wire new_n6247_;
  wire not_new_n1517_;
  wire not_po296_152867006319425761937651857692768264010;
  wire not_po296_225393402906922580878632490;
  wire new_n4422_;
  wire new_n8210_;
  wire new_n5332_;
  wire not_new_n7618_;
  wire not_new_n10099_;
  wire not_new_n4945__2;
  wire not_new_n1538__490;
  wire not_new_n4108_;
  wire not_new_n4738_;
  wire new_n3229_;
  wire not_new_n635__1;
  wire not_new_n9706_;
  wire and_new_n5748__new_n6116_;
  wire not_new_n7902_;
  wire new_n1456_;
  wire new_n6094_;
  wire not_new_n4915_;
  wire not_new_n637__19773267430;
  wire new_n5973_;
  wire not_pi035_0;
  wire not_new_n6982__0;
  wire not_new_n2786_;
  wire new_n5024_;
  wire not_new_n1601__113988951853731430;
  wire po061;
  wire new_n1850_;
  wire not_new_n3859_;
  wire new_n1749_;
  wire not_new_n4212_;
  wire new_n10132_;
  wire not_new_n581__541169560379521116689596608490;
  wire new_n3531_;
  wire or_not_new_n2537__not_new_n2541_;
  wire not_new_n601__70;
  wire new_n7829_;
  wire not_new_n606__8;
  wire po117;
  wire not_new_n595__8;
  wire not_new_n5286_;
  wire new_n6566_;
  wire new_n676_;
  wire new_n9571_;
  wire not_new_n989__47475615099430;
  wire not_new_n3851_;
  wire not_new_n8165_;
  wire new_n9629_;
  wire new_n926_;
  wire not_new_n8031_;
  wire new_n5724_;
  wire not_new_n5784_;
  wire new_n2625_;
  wire not_new_n589__9095436801298611408202050198891430;
  wire not_new_n7001__1;
  wire new_n1611_;
  wire new_n5137_;
  wire new_n6767_;
  wire not_new_n2285_;
  wire not_new_n3063_;
  wire new_n4132_;
  wire not_new_n637__4;
  wire not_new_n6981_;
  wire not_new_n7021_;
  wire and_new_n7161__new_n7474_;
  wire key_gate_28;
  wire not_new_n4831__0;
  wire not_new_n6507__0;
  wire new_n3110_;
  wire not_new_n8948_;
  wire new_n1385_;
  wire new_n3267_;
  wire not_new_n9384_;
  wire not_new_n775__2326305139872070;
  wire not_new_n4423_;
  wire not_new_n7145_;
  wire new_n7639_;
  wire not_new_n3986_;
  wire not_new_n648__113988951853731430;
  wire new_n2599_;
  wire not_new_n8887_;
  wire new_n7327_;
  wire not_new_n9581_;
  wire new_n7920_;
  wire not_new_n3102_;
  wire not_new_n9309_;
  wire not_new_n3967_;
  wire new_n9105_;
  wire not_new_n1730_;
  wire not_new_n7323_;
  wire not_new_n626__3;
  wire new_n1263_;
  wire not_new_n4985_;
  wire not_new_n3812_;
  wire not_new_n3185__8235430;
  wire new_n7615_;
  wire not_new_n2066_;
  wire not_new_n1612__2824752490;
  wire not_pi139_0;
  wire not_new_n3185__0;
  wire new_n9806_;
  wire not_new_n8895_;
  wire new_n8339_;
  wire not_new_n994__24010;
  wire new_n7511_;
  wire new_n1221_;
  wire new_n6588_;
  wire not_new_n8228_;
  wire not_new_n1582_;
  wire not_new_n5437_;
  wire key_gate_101;
  wire not_new_n5077_;
  wire not_new_n7237_;
  wire new_n5677_;
  wire not_new_n6658__0;
  wire not_new_n5083_;
  wire and_and_new_n2105__new_n2108__new_n2106_;
  wire or_not_new_n9719__not_new_n9718_;
  wire not_new_n1014__0;
  wire not_new_n6536_;
  wire not_new_n4423__0;
  wire new_n7341_;
  wire not_new_n1865_;
  wire or_or_not_new_n934__not_new_n933__0_not_new_n941__0;
  wire not_new_n629__332329305696010;
  wire new_n6443_;
  wire not_new_n3372_;
  wire new_n4715_;
  wire new_n10084_;
  wire new_n1418_;
  wire new_n9379_;
  wire not_new_n8548_;
  wire new_n5411_;
  wire not_new_n9474_;
  wire new_n3341_;
  wire not_new_n4420_;
  wire not_new_n1631__2;
  wire new_n7544_;
  wire not_pi162_3;
  wire not_new_n5650_;
  wire not_new_n4360_;
  wire not_pi166;
  wire new_n4718_;
  wire not_new_n1583__4;
  wire new_n5460_;
  wire not_new_n4066_;
  wire not_new_n1035__1;
  wire not_po296_205005145156954906122290109080958673914396262484637238056070;
  wire not_new_n585__9;
  wire not_new_n1059__1176490;
  wire new_n8329_;
  wire not_new_n3154_;
  wire not_new_n1886_;
  wire not_new_n1602__1;
  wire not_new_n9854_;
  wire not_new_n8848_;
  wire new_n5618_;
  wire not_new_n1427_;
  wire not_new_n1603__1176490;
  wire not_new_n5937_;
  wire not_new_n6943_;
  wire not_new_n5217_;
  wire not_new_n3922__0;
  wire not_new_n7635_;
  wire not_pi029_0;
  wire new_n4539_;
  wire not_new_n7471_;
  wire not_new_n8102_;
  wire not_new_n7888_;
  wire new_n7449_;
  wire not_new_n5469_;
  wire new_n2918_;
  wire not_new_n8198_;
  wire not_new_n4924_;
  wire new_n7122_;
  wire not_new_n8157_;
  wire not_new_n8110__0;
  wire and_and_new_n6395__new_n6396__new_n6228_;
  wire not_new_n628__403536070;
  wire not_new_n2723_;
  wire not_new_n1536__24010;
  wire new_n9764_;
  wire new_n8903_;
  wire not_pi136_2;
  wire not_new_n630__9;
  wire new_n4660_;
  wire new_n1305_;
  wire new_n9497_;
  wire not_new_n9520__0;
  wire not_pi019_0;
  wire not_new_n6387_;
  wire not_new_n9370_;
  wire new_n9216_;
  wire new_n2418_;
  wire new_n1580_;
  wire not_new_n624__490;
  wire not_new_n4437__0;
  wire new_n7190_;
  wire not_new_n3793_;
  wire not_new_n9007_;
  wire new_n6076_;
  wire not_new_n1065__1;
  wire new_n8452_;
  wire new_n6180_;
  wire not_new_n8779__0;
  wire not_new_n3997__0;
  wire not_new_n743__0;
  wire not_new_n588__70;
  wire new_n5531_;
  wire new_n7603_;
  wire not_new_n3847_;
  wire not_new_n9413__0;
  wire not_new_n7159__0;
  wire not_pi175_1;
  wire or_not_new_n1470__not_new_n3824_;
  wire not_new_n8163__0;
  wire not_new_n4174_;
  wire new_n7460_;
  wire new_n9762_;
  wire new_n7872_;
  wire po159;
  wire not_new_n9776_;
  wire new_n10282_;
  wire not_new_n725__0;
  wire not_new_n4001__0;
  wire not_new_n8151__0;
  wire not_new_n1958_;
  wire not_new_n7537_;
  wire new_n5900_;
  wire not_new_n6635__0;
  wire new_n7332_;
  wire not_new_n595__6782230728490;
  wire new_n4192_;
  wire not_new_n2597_;
  wire not_new_n8559_;
  wire or_not_new_n3130__not_new_n3131_;
  wire not_new_n7755_;
  wire not_new_n7819_;
  wire new_n5517_;
  wire not_new_n6692_;
  wire new_n9095_;
  wire not_new_n1588__8;
  wire not_new_n1495_;
  wire not_new_n588__138412872010;
  wire new_n5195_;
  wire new_n7456_;
  wire not_new_n7047_;
  wire not_new_n3294_;
  wire not_new_n1588__797922662976120010;
  wire new_n7751_;
  wire not_new_n8408_;
  wire not_new_n4781_;
  wire not_new_n601__4;
  wire or_not_new_n1335__not_new_n1333_;
  wire not_new_n9709_;
  wire not_new_n636__490;
  wire not_new_n626__113988951853731430;
  wire new_n4001_;
  wire not_new_n2459_;
  wire new_n7516_;
  wire not_new_n1600__138412872010;
  wire new_n5663_;
  wire not_new_n7259_;
  wire new_n5876_;
  wire new_n10002_;
  wire new_n669_;
  wire new_n5125_;
  wire not_new_n7923_;
  wire not_new_n9113_;
  wire not_new_n978_;
  wire new_n8253_;
  wire po246;
  wire not_new_n6443__968890104070;
  wire and_new_n5740__new_n6096_;
  wire not_new_n628__19773267430;
  wire not_new_n8894__0;
  wire not_new_n984_;
  wire not_new_n4769__0;
  wire new_n2477_;
  wire new_n7255_;
  wire not_new_n8432_;
  wire new_n8298_;
  wire new_n7083_;
  wire po217;
  wire not_new_n3908_;
  wire new_n8114_;
  wire not_new_n4202_;
  wire not_new_n9887_;
  wire not_new_n9735_;
  wire not_new_n596__6782230728490;
  wire not_new_n6454_;
  wire not_new_n6551_;
  wire new_n6303_;
  wire new_n7999_;
  wire not_new_n1598__6;
  wire not_new_n7800_;
  wire new_n2348_;
  wire not_pi250_4;
  wire not_new_n3527_;
  wire new_n1316_;
  wire not_new_n8709__0;
  wire not_new_n9502_;
  wire not_new_n6524_;
  wire not_new_n1580__113988951853731430;
  wire new_n3903_;
  wire not_new_n10251_;
  wire new_n5266_;
  wire new_n3967_;
  wire po099;
  wire not_new_n5529_;
  wire new_n8654_;
  wire new_n4948_;
  wire not_new_n586__8;
  wire new_n6921_;
  wire new_n1940_;
  wire or_not_new_n4933__not_new_n4930__0;
  wire not_new_n5525_;
  wire not_new_n989__0;
  wire or_or_not_new_n2803__not_new_n2806__not_new_n2805_;
  wire new_n9500_;
  wire not_new_n10188_;
  wire not_new_n9131_;
  wire new_n5433_;
  wire not_new_n7469_;
  wire new_n4216_;
  wire not_new_n605__1176490;
  wire not_new_n1417_;
  wire not_new_n10310_;
  wire not_new_n3163_;
  wire not_new_n4482_;
  wire new_n5673_;
  wire not_pi064_8235430;
  wire new_n4603_;
  wire not_new_n8078_;
  wire key_gate_90;
  wire new_n4129_;
  wire not_pi150;
  wire new_n7106_;
  wire not_new_n4425_;
  wire new_n2140_;
  wire not_pi055_0;
  wire new_n3936_;
  wire not_new_n7062_;
  wire not_new_n1604__8;
  wire not_new_n8962_;
  wire not_new_n6255_;
  wire not_new_n6617__0;
  wire not_new_n630__3430;
  wire new_n10017_;
  wire new_n3686_;
  wire not_pi079;
  wire or_or_not_new_n2265__not_new_n2262__not_new_n2263_;
  wire new_n5086_;
  wire new_n6231_;
  wire new_n6285_;
  wire new_n8874_;
  wire not_new_n4415__1;
  wire not_new_n9972_;
  wire new_n1192_;
  wire not_new_n601__47475615099430;
  wire not_new_n638__657123623635342801395430;
  wire and_and_new_n6374__new_n6372__new_n6371_;
  wire not_new_n5765_;
  wire not_pi236;
  wire new_n3294_;
  wire not_new_n7093_;
  wire new_n1039_;
  wire or_not_new_n2820__not_new_n2823_;
  wire new_n6220_;
  wire new_n8745_;
  wire new_n2093_;
  wire not_new_n7827_;
  wire new_n2760_;
  wire not_new_n1596__490;
  wire not_new_n1901_;
  wire not_new_n2554_;
  wire not_new_n5063__0;
  wire not_new_n1035__3430;
  wire new_n2929_;
  wire not_new_n8042_;
  wire not_new_n622_;
  wire new_n5851_;
  wire not_pi074;
  wire or_not_new_n1977__not_new_n1978_;
  wire not_new_n1598__4;
  wire not_new_n4780__1;
  wire not_pi172_1;
  wire new_n8283_;
  wire po199;
  wire not_new_n596__2;
  wire new_n3316_;
  wire not_new_n8974_;
  wire new_n7486_;
  wire not_new_n5465__1;
  wire not_new_n5723_;
  wire new_n3643_;
  wire and_new_n1262__new_n1951_;
  wire new_n7826_;
  wire not_new_n9974_;
  wire new_n9262_;
  wire not_new_n9658_;
  wire new_n5575_;
  wire not_new_n9258_;
  wire not_new_n585__332329305696010;
  wire new_n2356_;
  wire new_n8821_;
  wire new_n6904_;
  wire not_new_n648__8;
  wire not_new_n5235_;
  wire not_new_n6989_;
  wire new_n8402_;
  wire new_n5156_;
  wire not_new_n8893__0;
  wire new_n4441_;
  wire not_new_n638__9;
  wire not_new_n1055__70;
  wire not_pi033_1;
  wire new_n6897_;
  wire not_new_n3526_;
  wire not_new_n2148_;
  wire not_new_n7337_;
  wire not_new_n9918_;
  wire po236;
  wire not_new_n1039__24010;
  wire new_n8013_;
  wire not_new_n994__3;
  wire new_n4800_;
  wire not_new_n984__8;
  wire not_new_n7095_;
  wire po162;
  wire new_n10035_;
  wire not_pi261;
  wire new_n7124_;
  wire not_new_n8932_;
  wire not_new_n727__0;
  wire new_n8611_;
  wire not_new_n8024_;
  wire not_new_n1596__70;
  wire new_n8791_;
  wire new_n2457_;
  wire new_n8637_;
  wire not_new_n1039__0;
  wire not_new_n5925_;
  wire new_n9549_;
  wire not_new_n1420_;
  wire new_n8972_;
  wire not_new_n4972_;
  wire new_n8468_;
  wire new_n3315_;
  wire not_new_n6851_;
  wire not_new_n9469_;
  wire new_n8416_;
  wire not_new_n1384_;
  wire new_n8382_;
  wire not_new_n5709_;
  wire not_new_n6570_;
  wire not_new_n8075_;
  wire not_new_n4770__1;
  wire not_new_n1728__8;
  wire new_n7790_;
  wire not_new_n1053__1176490;
  wire new_n2680_;
  wire not_pi274;
  wire not_new_n7946_;
  wire or_not_new_n2587__not_new_n2591_;
  wire not_new_n1055__2326305139872070;
  wire new_n4774_;
  wire new_n2961_;
  wire and_new_n9189__new_n9187_;
  wire not_new_n624__6782230728490;
  wire not_new_n4937__0;
  wire not_new_n9834_;
  wire new_n3520_;
  wire not_new_n8585_;
  wire new_n4560_;
  wire new_n8483_;
  wire new_n8291_;
  wire new_n4958_;
  wire not_new_n1020__0;
  wire and_new_n8789__new_n8784_;
  wire new_n2462_;
  wire new_n6225_;
  wire new_n1640_;
  wire not_new_n7037__0;
  wire not_new_n6523_;
  wire po185;
  wire not_new_n9412__0;
  wire not_new_n9865_;
  wire not_new_n648__2824752490;
  wire not_new_n1604__57648010;
  wire not_pi179_2;
  wire new_n7762_;
  wire new_n2003_;
  wire not_new_n5273_;
  wire not_new_n10108_;
  wire not_pi056;
  wire new_n9033_;
  wire new_n2964_;
  wire not_new_n3311__7;
  wire new_n3463_;
  wire new_n7694_;
  wire new_n6033_;
  wire not_new_n1591__70;
  wire not_new_n1534__8;
  wire new_n705_;
  wire new_n10167_;
  wire not_new_n8839_;
  wire new_n6835_;
  wire not_new_n586__332329305696010;
  wire new_n4744_;
  wire not_new_n9328_;
  wire not_new_n3977__0;
  wire new_n4589_;
  wire not_new_n1037__6;
  wire new_n8641_;
  wire new_n5501_;
  wire not_new_n595__490;
  wire new_n5676_;
  wire new_n1010_;
  wire new_n6442_;
  wire new_n9331_;
  wire new_n7839_;
  wire new_n4089_;
  wire new_n1830_;
  wire new_n4617_;
  wire not_new_n5965_;
  wire not_new_n7908_;
  wire not_new_n8129_;
  wire new_n6218_;
  wire new_n7236_;
  wire not_new_n4378_;
  wire not_new_n7165_;
  wire not_new_n2762_;
  wire not_new_n10033__0;
  wire new_n5431_;
  wire not_new_n994__113988951853731430;
  wire not_new_n596__9;
  wire not_new_n7548_;
  wire new_n3205_;
  wire not_new_n644__968890104070;
  wire not_new_n581__403536070;
  wire new_n9739_;
  wire not_new_n1065__797922662976120010;
  wire not_new_n3990_;
  wire not_new_n8898__0;
  wire not_new_n8960_;
  wire not_new_n6164_;
  wire not_new_n1584__490;
  wire not_new_n626__0;
  wire new_n5474_;
  wire not_new_n7366_;
  wire not_new_n603__2326305139872070;
  wire not_new_n1047__2;
  wire not_new_n8093_;
  wire not_new_n1599__24010;
  wire new_n8475_;
  wire not_new_n599__5;
  wire not_new_n5854_;
  wire new_n2694_;
  wire new_n2023_;
  wire not_new_n6675_;
  wire not_new_n1728__2326305139872070;
  wire new_n9962_;
  wire not_new_n588__113988951853731430;
  wire not_new_n8018_;
  wire not_new_n6746_;
  wire new_n7187_;
  wire not_new_n1151__0;
  wire not_new_n634__797922662976120010;
  wire not_new_n9047_;
  wire not_new_n8657_;
  wire not_new_n1589__7;
  wire not_new_n1019_;
  wire new_n3351_;
  wire new_n3288_;
  wire new_n2938_;
  wire not_new_n5378_;
  wire not_new_n5944_;
  wire not_new_n1537__8;
  wire new_n7287_;
  wire not_new_n9438_;
  wire not_new_n642__168070;
  wire not_new_n1995_;
  wire new_n9172_;
  wire not_pi047_0;
  wire not_new_n10074_;
  wire not_new_n581__3788186922656647816827176259430;
  wire not_po298_5;
  wire new_n3182_;
  wire new_n3553_;
  wire new_n1990_;
  wire not_new_n2625_;
  wire new_n3999_;
  wire not_new_n598__797922662976120010;
  wire new_n7994_;
  wire not_new_n6984_;
  wire not_new_n8310_;
  wire new_n9827_;
  wire not_new_n8152__0;
  wire new_n8374_;
  wire key_gate_66;
  wire not_new_n3117_;
  wire new_n4757_;
  wire not_new_n4949__0;
  wire and_new_n8112__new_n8484_;
  wire new_n5050_;
  wire not_new_n1035__3;
  wire not_new_n635__8235430;
  wire not_new_n2871_;
  wire new_n4766_;
  wire new_n5094_;
  wire new_n5157_;
  wire not_new_n631__1915812313805664144010;
  wire new_n8844_;
  wire new_n2205_;
  wire not_new_n6295_;
  wire not_new_n9342_;
  wire not_new_n4657_;
  wire not_new_n642__3430;
  wire and_not_pi036_1_not_pi037_1;
  wire not_new_n994__57648010;
  wire not_new_n7163_;
  wire new_n9559_;
  wire not_new_n3985__0;
  wire new_n5225_;
  wire not_new_n7099_;
  wire not_new_n7051_;
  wire new_n8547_;
  wire new_n4787_;
  wire not_pi140_0;
  wire not_pi054;
  wire not_new_n2823_;
  wire not_new_n5630__1;
  wire new_n7512_;
  wire new_n3728_;
  wire new_n739_;
  wire not_new_n8882_;
  wire not_new_n2984_;
  wire new_n5301_;
  wire not_new_n4120__0;
  wire not_new_n1169__0;
  wire not_new_n5461_;
  wire new_n6941_;
  wire or_not_new_n1231__not_new_n1229_;
  wire new_n2328_;
  wire not_new_n1053__2;
  wire new_n3139_;
  wire new_n2713_;
  wire new_n8880_;
  wire new_n4465_;
  wire new_n1928_;
  wire not_new_n1012__0;
  wire new_n971_;
  wire not_new_n3857_;
  wire new_n5504_;
  wire not_new_n2208_;
  wire new_n6948_;
  wire not_new_n9621_;
  wire new_n4058_;
  wire new_n7636_;
  wire not_new_n5722_;
  wire new_n6204_;
  wire not_new_n6974__9;
  wire new_n7389_;
  wire not_new_n3150_;
  wire new_n8839_;
  wire not_new_n5804_;
  wire not_new_n1612__6782230728490;
  wire new_n8148_;
  wire not_new_n4453__0;
  wire or_not_new_n1559__not_new_n2454_;
  wire new_n1718_;
  wire new_n7521_;
  wire new_n3101_;
  wire not_new_n7591__0;
  wire new_n7880_;
  wire new_n6516_;
  wire not_new_n8269_;
  wire not_new_n5507_;
  wire not_new_n597__403536070;
  wire new_n6862_;
  wire or_not_new_n1027__13410686196639649008070_not_new_n4227__0;
  wire not_new_n7190_;
  wire new_n2581_;
  wire not_new_n8105__2;
  wire new_n8530_;
  wire new_n5353_;
  wire not_new_n6481_;
  wire key_gate_68;
  wire not_new_n1596__138412872010;
  wire new_n4749_;
  wire not_pi253;
  wire not_new_n654_;
  wire new_n5791_;
  wire not_new_n3095_;
  wire new_n8556_;
  wire new_n6781_;
  wire new_n10064_;
  wire new_n7566_;
  wire not_new_n2509__1;
  wire not_new_n3384__5;
  wire new_n6419_;
  wire not_new_n1612__168070;
  wire not_new_n3353_;
  wire not_new_n2932_;
  wire not_new_n8100_;
  wire not_new_n624__47475615099430;
  wire new_n8313_;
  wire new_n4724_;
  wire new_n6011_;
  wire not_new_n2189_;
  wire new_n3669_;
  wire not_new_n6589_;
  wire not_new_n6974__16284135979104490;
  wire new_n8905_;
  wire new_n1697_;
  wire new_n9005_;
  wire not_new_n8302_;
  wire not_new_n10080_;
  wire not_new_n644__797922662976120010;
  wire not_new_n9413_;
  wire new_n8292_;
  wire not_new_n1053__70;
  wire new_n5702_;
  wire not_new_n596__6;
  wire new_n1856_;
  wire new_n5717_;
  wire not_new_n598__490;
  wire not_new_n2935_;
  wire not_new_n633__2;
  wire not_new_n6634__1;
  wire new_n5194_;
  wire not_new_n9103_;
  wire not_pi036;
  wire new_n3889_;
  wire new_n3544_;
  wire new_n4351_;
  wire not_new_n7765_;
  wire new_n8662_;
  wire new_n8997_;
  wire new_n4320_;
  wire new_n3286_;
  wire not_new_n10059__0;
  wire not_new_n1536__797922662976120010;
  wire not_new_n1613__9;
  wire new_n2092_;
  wire new_n9882_;
  wire not_new_n10271_;
  wire not_new_n5076_;
  wire not_new_n5498_;
  wire not_new_n7028_;
  wire new_n2440_;
  wire new_n4557_;
  wire not_new_n3372__403536070;
  wire new_n3960_;
  wire not_new_n7042_;
  wire or_not_new_n5484__not_new_n605__0;
  wire new_n928_;
  wire new_n8564_;
  wire not_new_n7413_;
  wire not_new_n8456_;
  wire not_new_n1538_;
  wire not_new_n1442_;
  wire new_n1727_;
  wire not_new_n1047__332329305696010;
  wire not_new_n1600__2824752490;
  wire not_new_n5585_;
  wire new_n3166_;
  wire not_new_n7878_;
  wire new_n1687_;
  wire not_new_n1057__138412872010;
  wire not_new_n7756_;
  wire not_new_n5685_;
  wire po286;
  wire not_new_n3965_;
  wire new_n2426_;
  wire not_new_n4610_;
  wire new_n4844_;
  wire not_new_n6991__1;
  wire not_pi172_0;
  wire not_new_n1031__8235430;
  wire not_new_n7508_;
  wire not_new_n6335_;
  wire not_new_n8171_;
  wire new_n3172_;
  wire new_n7716_;
  wire not_new_n637__57648010;
  wire or_not_new_n1001__not_new_n1000_;
  wire new_n9756_;
  wire new_n3024_;
  wire not_new_n989__7;
  wire not_new_n3868_;
  wire not_new_n5736_;
  wire not_new_n9623_;
  wire new_n7986_;
  wire new_n6607_;
  wire new_n7792_;
  wire not_new_n1791_;
  wire not_new_n2204__0;
  wire new_n8539_;
  wire not_new_n5340_;
  wire new_n1281_;
  wire not_new_n1031__1;
  wire new_n8835_;
  wire or_not_new_n5466__not_new_n5674__1;
  wire not_po298_2326305139872070;
  wire not_new_n9329_;
  wire new_n9543_;
  wire not_new_n1047__8;
  wire not_new_n5571_;
  wire not_new_n6730_;
  wire not_new_n636__968890104070;
  wire new_n3849_;
  wire new_n8953_;
  wire not_new_n9366__0;
  wire not_new_n8982_;
  wire new_n6874_;
  wire new_n4711_;
  wire new_n5507_;
  wire new_n9759_;
  wire not_new_n587__24010;
  wire not_new_n1047__4;
  wire not_new_n7674_;
  wire and_and_new_n2314__new_n2317__new_n2315_;
  wire not_new_n8914_;
  wire not_new_n5642_;
  wire new_n10039_;
  wire not_new_n1028__2;
  wire not_new_n9286_;
  wire not_new_n1600__968890104070;
  wire not_new_n4118__0;
  wire not_new_n1728__47475615099430;
  wire not_new_n7738_;
  wire new_n6497_;
  wire new_n3471_;
  wire not_new_n5034_;
  wire new_n2020_;
  wire not_new_n8890_;
  wire or_not_new_n2053__not_new_n2054_;
  wire new_n9192_;
  wire not_new_n4773_;
  wire not_new_n6031_;
  wire new_n5516_;
  wire new_n645_;
  wire not_new_n3953_;
  wire po134;
  wire not_new_n5355_;
  wire key_gate_7;
  wire not_pi251_0;
  wire new_n6082_;
  wire and_new_n1750__new_n1751_;
  wire not_new_n8885_;
  wire not_pi035;
  wire not_new_n644__168070;
  wire new_n2434_;
  wire new_n8509_;
  wire new_n7209_;
  wire new_n6162_;
  wire new_n7819_;
  wire and_not_pi060_1_not_pi059_1;
  wire not_new_n1580__16284135979104490;
  wire not_new_n1728__4;
  wire new_n6531_;
  wire and_new_n7160__new_n7500_;
  wire not_new_n1584__2326305139872070;
  wire new_n4075_;
  wire not_new_n5918_;
  wire new_n4587_;
  wire new_n4506_;
  wire not_new_n1611__4;
  wire key_gate_8;
  wire not_new_n6735_;
  wire not_pi168_2;
  wire or_not_new_n6328__not_new_n6373__3;
  wire new_n7197_;
  wire not_new_n3372__10;
  wire not_new_n1331_;
  wire not_new_n7033_;
  wire not_new_n7010__2;
  wire not_new_n2756_;
  wire new_n3073_;
  wire not_new_n775__113988951853731430;
  wire new_n5778_;
  wire not_new_n3518_;
  wire not_new_n8251__0;
  wire new_n2910_;
  wire new_n4923_;
  wire not_new_n1014__1;
  wire not_new_n762_;
  wire new_n1976_;
  wire not_new_n1633_;
  wire new_n6592_;
  wire new_n10272_;
  wire not_new_n6234_;
  wire not_new_n8605_;
  wire not_new_n7004_;
  wire new_n8585_;
  wire not_new_n1063__8;
  wire not_new_n5315_;
  wire or_not_new_n2734__not_new_n2733_;
  wire not_new_n625__8;
  wire not_new_n5711_;
  wire not_new_n9440_;
  wire new_n9114_;
  wire new_n9074_;
  wire not_new_n3348_;
  wire new_n1594_;
  wire not_new_n5745__0;
  wire not_new_n2191_;
  wire not_new_n2085_;
  wire not_new_n607__8;
  wire not_new_n3315__1;
  wire not_new_n5184_;
  wire not_new_n3411_;
  wire not_new_n1591__1176490;
  wire not_pi064_8;
  wire new_n592_;
  wire new_n8391_;
  wire new_n9742_;
  wire not_new_n7423_;
  wire new_n3606_;
  wire and_new_n1760__new_n1759_;
  wire not_new_n6968_;
  wire not_new_n8919_;
  wire new_n1527_;
  wire not_new_n2544_;
  wire new_n2681_;
  wire not_new_n5755_;
  wire not_new_n634__39098210485829880490;
  wire not_new_n2829_;
  wire not_new_n611__24010;
  wire not_new_n8160__0;
  wire new_n6519_;
  wire new_n1350_;
  wire not_new_n3152_;
  wire not_new_n5627_;
  wire new_n2210_;
  wire not_new_n4949_;
  wire new_n1499_;
  wire new_n5935_;
  wire not_new_n5746_;
  wire not_new_n2864_;
  wire and_new_n1282__new_n2046_;
  wire new_n5585_;
  wire not_new_n9999_;
  wire new_n9677_;
  wire new_n9306_;
  wire new_n6739_;
  wire new_n9068_;
  wire not_new_n4781__0;
  wire not_new_n6548_;
  wire new_n4764_;
  wire not_new_n10323_;
  wire new_n1166_;
  wire not_new_n4270_;
  wire not_new_n1584__8235430;
  wire not_pi175_0;
  wire new_n4161_;
  wire not_new_n7147_;
  wire not_new_n4485_;
  wire not_new_n5497_;
  wire not_new_n7267__0;
  wire not_new_n1067__8;
  wire not_new_n1600__5;
  wire new_n5001_;
  wire not_new_n8172__1;
  wire not_new_n6994_;
  wire not_new_n10311_;
  wire not_pi104;
  wire not_new_n6532_;
  wire new_n8912_;
  wire new_n5867_;
  wire not_po296_6168735096280623662907561568153897267931784070;
  wire and_and_not_pi051_1_not_pi050_1_not_pi049_1;
  wire and_new_n3079__new_n998_;
  wire new_n3353_;
  wire new_n7240_;
  wire not_new_n6246_;
  wire not_new_n7026__1;
  wire not_pi057;
  wire not_new_n6263_;
  wire not_new_n1045__6782230728490;
  wire new_n1231_;
  wire new_n1020_;
  wire new_n4076_;
  wire not_pi072;
  wire not_new_n1603__19773267430;
  wire not_new_n1581__2326305139872070;
  wire new_n2218_;
  wire not_new_n1039__39098210485829880490;
  wire or_not_new_n4825__not_new_n4804_;
  wire new_n5227_;
  wire not_new_n1045__19773267430;
  wire new_n2878_;
  wire new_n740_;
  wire new_n960_;
  wire or_not_new_n1782__not_new_n1783_;
  wire not_new_n9086_;
  wire key_gate_35;
  wire not_new_n1580__19773267430;
  wire new_n2468_;
  wire not_new_n9093_;
  wire not_new_n718__0;
  wire not_new_n5185_;
  wire new_n8222_;
  wire or_not_new_n5436__not_new_n5630__1;
  wire new_n5962_;
  wire new_n4783_;
  wire not_new_n1603__490;
  wire not_new_n610__168070;
  wire new_n4601_;
  wire new_n9659_;
  wire key_gate_71;
  wire new_n7452_;
  wire not_new_n1584__6782230728490;
  wire not_new_n7315__0;
  wire new_n7046_;
  wire new_n3314_;
  wire not_new_n5705_;
  wire new_n4868_;
  wire new_n3730_;
  wire new_n5945_;
  wire new_n8104_;
  wire not_new_n7438_;
  wire not_new_n2230_;
  wire not_new_n8178_;
  wire not_new_n7116_;
  wire not_new_n3939_;
  wire not_new_n617__47475615099430;
  wire not_new_n9510_;
  wire new_n9732_;
  wire not_new_n5957_;
  wire not_new_n2827_;
  wire not_new_n8978__2;
  wire new_n3953_;
  wire or_not_new_n2597__not_new_n2601_;
  wire new_n6569_;
  wire not_new_n3165_;
  wire not_new_n4138_;
  wire new_n3230_;
  wire and_and_new_n8753__new_n8754__new_n8761_;
  wire not_new_n7642_;
  wire not_new_n1613__24010;
  wire new_n10336_;
  wire not_pi064_332329305696010;
  wire new_n6504_;
  wire new_n4592_;
  wire not_new_n7442_;
  wire not_new_n10100_;
  wire new_n2552_;
  wire not_new_n9724_;
  wire not_new_n1017__1;
  wire not_new_n4099_;
  wire not_pi069;
  wire not_pi182;
  wire new_n5079_;
  wire not_new_n2130_;
  wire not_new_n2545_;
  wire not_new_n639__168070;
  wire not_new_n9748_;
  wire new_n6945_;
  wire not_new_n7966_;
  wire not_new_n707_;
  wire new_n10059_;
  wire new_n9426_;
  wire new_n2706_;
  wire and_and_new_n2238__new_n2241__new_n2239_;
  wire not_new_n4701_;
  wire not_new_n2509__0;
  wire not_new_n1622__1;
  wire not_new_n10265_;
  wire not_new_n10182_;
  wire not_new_n3256_;
  wire new_n5685_;
  wire not_new_n1578_;
  wire not_new_n7783_;
  wire not_pi001_0;
  wire new_n1560_;
  wire new_n6255_;
  wire not_new_n2987_;
  wire new_n5964_;
  wire not_new_n5487_;
  wire not_new_n3311__10;
  wire new_n7422_;
  wire new_n5400_;
  wire new_n7314_;
  wire not_pi163_3;
  wire not_new_n2153_;
  wire new_n2770_;
  wire not_new_n3311__9;
  wire not_new_n4441__0;
  wire or_or_not_new_n6353__not_new_n6232__5_not_new_n1069__3430;
  wire new_n5978_;
  wire new_n3731_;
  wire new_n5480_;
  wire not_new_n3218_;
  wire new_n4906_;
  wire not_new_n4803__0;
  wire new_n6732_;
  wire new_n6712_;
  wire not_new_n5247_;
  wire not_new_n8070_;
  wire not_new_n648__5585458640832840070;
  wire new_n3052_;
  wire new_n1551_;
  wire not_new_n596__57648010;
  wire not_new_n5358_;
  wire not_new_n1537__3430;
  wire not_new_n7636__0;
  wire not_new_n9745_;
  wire not_new_n648__1;
  wire new_n5183_;
  wire not_new_n625__93874803376477543056490;
  wire new_n6093_;
  wire not_new_n9924_;
  wire new_n6984_;
  wire not_new_n729_;
  wire not_new_n4948__0;
  wire not_new_n1057__403536070;
  wire or_not_new_n1939__not_new_n1940_;
  wire not_new_n642__2;
  wire not_new_n5123_;
  wire not_new_n4137__0;
  wire not_new_n4071_;
  wire not_new_n1439_;
  wire new_n4343_;
  wire not_new_n1585__113988951853731430;
  wire new_n3275_;
  wire not_new_n7111_;
  wire not_pi207;
  wire new_n6089_;
  wire new_n2613_;
  wire not_pi106;
  wire not_new_n588__4;
  wire not_new_n8825_;
  wire and_and_new_n6357__new_n6356__new_n6404_;
  wire new_n1035_;
  wire new_n6517_;
  wire not_new_n8470_;
  wire new_n4066_;
  wire not_new_n4438__0;
  wire not_new_n5714_;
  wire new_n5836_;
  wire new_n2729_;
  wire not_new_n5843_;
  wire not_new_n5522_;
  wire not_new_n7524_;
  wire and_new_n1934__new_n1937_;
  wire new_n2824_;
  wire new_n6757_;
  wire new_n9617_;
  wire not_new_n6333_;
  wire not_new_n639__490;
  wire not_new_n639__2824752490;
  wire not_new_n1598__1176490;
  wire not_new_n1971_;
  wire new_n5889_;
  wire new_n4734_;
  wire new_n7079_;
  wire not_new_n3864_;
  wire not_new_n1035__9;
  wire not_new_n6509_;
  wire not_new_n1011__0;
  wire new_n3191_;
  wire new_n8387_;
  wire not_new_n3846_;
  wire not_pi012_0;
  wire new_n4165_;
  wire not_new_n7206_;
  wire not_new_n8707_;
  wire not_new_n928__797922662976120010;
  wire new_n9993_;
  wire not_new_n4614_;
  wire not_new_n9521_;
  wire new_n4209_;
  wire new_n8091_;
  wire new_n2044_;
  wire not_new_n1599__138412872010;
  wire new_n2969_;
  wire not_new_n9388_;
  wire not_new_n595__1;
  wire not_pi270_2;
  wire new_n2509_;
  wire not_new_n2896_;
  wire not_new_n4916_;
  wire not_new_n4263_;
  wire not_pi247_1;
  wire not_new_n4101_;
  wire not_new_n9879_;
  wire new_n2958_;
  wire new_n8492_;
  wire new_n7671_;
  wire new_n8519_;
  wire not_new_n3991_;
  wire not_new_n5156__0;
  wire new_n3333_;
  wire new_n1943_;
  wire not_pi130;
  wire new_n2235_;
  wire not_new_n7858_;
  wire new_n8312_;
  wire not_pi042;
  wire new_n9436_;
  wire or_not_new_n2881__not_new_n2880_;
  wire new_n3982_;
  wire not_new_n9948_;
  wire new_n4842_;
  wire new_n3900_;
  wire not_new_n1584__1;
  wire new_n6580_;
  wire new_n9496_;
  wire and_new_n2181__new_n2184_;
  wire new_n9660_;
  wire not_new_n8318_;
  wire and_and_and_new_n1053__new_n6232__new_n6395__new_n6317_;
  wire new_n7976_;
  wire new_n6043_;
  wire new_n3500_;
  wire not_new_n10261_;
  wire new_n2014_;
  wire not_new_n7681_;
  wire not_new_n5489__0;
  wire not_new_n3023_;
  wire new_n2814_;
  wire not_new_n8112__0;
  wire new_n3690_;
  wire new_n2148_;
  wire not_new_n1626__0;
  wire new_n6358_;
  wire new_n6801_;
  wire not_new_n1061__968890104070;
  wire new_n5642_;
  wire new_n8688_;
  wire new_n1714_;
  wire new_n6267_;
  wire key_gate_59;
  wire not_new_n9860_;
  wire new_n4919_;
  wire not_new_n1037_;
  wire and_new_n8997__new_n8998_;
  wire new_n3588_;
  wire not_new_n8153__0;
  wire not_new_n6512__0;
  wire not_new_n9110_;
  wire new_n1049_;
  wire not_new_n589__11044276742439206463052992010;
  wire new_n5883_;
  wire not_new_n7773__0;
  wire not_new_n4236_;
  wire not_new_n6088_;
  wire new_n5456_;
  wire or_not_new_n3173__not_new_n3172_;
  wire new_n2624_;
  wire not_new_n2633_;
  wire new_n7427_;
  wire new_n9191_;
  wire not_pi197;
  wire new_n763_;
  wire new_n9583_;
  wire new_n8523_;
  wire new_n3301_;
  wire not_new_n9534_;
  wire new_n996_;
  wire new_n1722_;
  wire new_n8481_;
  wire new_n8712_;
  wire new_n8747_;
  wire new_n3926_;
  wire new_n8529_;
  wire not_new_n2654_;
  wire not_pi056_1;
  wire not_new_n3266_;
  wire not_new_n648__968890104070;
  wire not_new_n5515_;
  wire not_new_n642__490;
  wire not_pi134_2;
  wire po116;
  wire new_n9425_;
  wire not_pi040_1;
  wire not_new_n9012_;
  wire not_new_n2509__5;
  wire not_new_n8350__0;
  wire not_new_n9346_;
  wire new_n1682_;
  wire new_n9080_;
  wire new_n1450_;
  wire not_new_n585__6782230728490;
  wire not_new_n10155_;
  wire not_pi033;
  wire or_not_new_n1271__not_new_n1269_;
  wire not_new_n9268_;
  wire not_new_n672_;
  wire not_pi266_0;
  wire not_new_n5451_;
  wire new_n4480_;
  wire new_n5422_;
  wire not_new_n1828_;
  wire not_new_n8851__0;
  wire not_new_n9793_;
  wire new_n8608_;
  wire not_new_n1869_;
  wire new_n8380_;
  wire not_new_n8405_;
  wire not_pi043_1;
  wire not_new_n3251_;
  wire new_n4448_;
  wire not_new_n4909_;
  wire not_po296_797922662976120010;
  wire new_n9823_;
  wire new_n4621_;
  wire new_n10033_;
  wire new_n10103_;
  wire new_n8983_;
  wire not_new_n5384_;
  wire not_new_n5811__0;
  wire new_n4991_;
  wire new_n7018_;
  wire not_new_n596__113988951853731430;
  wire new_n2372_;
  wire and_new_n1230__new_n1799_;
  wire new_n4286_;
  wire not_new_n2898_;
  wire new_n1404_;
  wire not_new_n9659_;
  wire not_new_n10151_;
  wire not_new_n4178_;
  wire and_and_new_n2517__new_n2518__new_n2516_;
  wire not_new_n10210_;
  wire new_n3464_;
  wire not_new_n639__10;
  wire not_new_n5536_;
  wire not_new_n1612__138412872010;
  wire new_n5667_;
  wire not_new_n5079__0;
  wire not_new_n6933_;
  wire not_new_n1600__490;
  wire not_new_n1045__10;
  wire new_n7761_;
  wire new_n5662_;
  wire new_n1888_;
  wire not_new_n5038_;
  wire not_new_n7596__0;
  wire new_n1958_;
  wire new_n8706_;
  wire not_new_n1424_;
  wire new_n10156_;
  wire not_new_n3185__24010;
  wire new_n9701_;
  wire new_n1899_;
  wire not_new_n4782_;
  wire new_n6174_;
  wire new_n4215_;
  wire new_n1662_;
  wire not_new_n4487_;
  wire not_new_n6970_;
  wire new_n8101_;
  wire not_pi107;
  wire not_new_n1167_;
  wire new_n9738_;
  wire not_new_n622__3430;
  wire new_n2492_;
  wire not_new_n1478_;
  wire new_n6843_;
  wire new_n9523_;
  wire new_n1971_;
  wire not_new_n1576__403536070;
  wire not_new_n6582_;
  wire not_new_n7496_;
  wire not_new_n9796_;
  wire not_new_n5544_;
  wire not_new_n6547_;
  wire not_new_n1183_;
  wire not_new_n10013__1;
  wire and_new_n1820__new_n1823_;
  wire not_new_n5182__0;
  wire new_n2600_;
  wire new_n8055_;
  wire new_n3629_;
  wire not_new_n1063__70;
  wire not_new_n7016__1;
  wire not_new_n4251_;
  wire not_new_n7130_;
  wire not_new_n1313_;
  wire not_new_n637__168070;
  wire new_n6546_;
  wire new_n6864_;
  wire not_new_n2775_;
  wire new_n2069_;
  wire not_new_n7004__2;
  wire not_new_n1631__332329305696010;
  wire or_not_new_n6042__not_new_n5927_;
  wire new_n7754_;
  wire new_n7900_;
  wire not_new_n9910_;
  wire new_n9011_;
  wire not_new_n6803_;
  wire not_new_n1811_;
  wire new_n3916_;
  wire new_n7901_;
  wire new_n7138_;
  wire new_n7380_;
  wire not_new_n8399_;
  wire new_n6385_;
  wire not_new_n9963_;
  wire new_n5390_;
  wire new_n4226_;
  wire new_n5437_;
  wire po034;
  wire not_new_n8627_;
  wire new_n5632_;
  wire not_new_n1604__0;
  wire not_new_n5917_;
  wire not_new_n4685_;
  wire new_n3761_;
  wire new_n1377_;
  wire new_n2951_;
  wire not_new_n1003__0;
  wire not_new_n4124__1;
  wire not_new_n7386_;
  wire new_n4133_;
  wire not_new_n10343_;
  wire key_gate_43;
  wire new_n4214_;
  wire not_new_n1600__168070;
  wire not_new_n5007_;
  wire new_n6622_;
  wire not_new_n2313_;
  wire not_new_n595__7;
  wire new_n2024_;
  wire not_new_n3694_;
  wire or_not_new_n1560__not_new_n2459_;
  wire new_n4195_;
  wire not_pi131_3;
  wire new_n5006_;
  wire not_new_n1597__490;
  wire and_new_n9168__new_n9167_;
  wire not_new_n9520_;
  wire new_n6371_;
  wire new_n7623_;
  wire new_n8124_;
  wire new_n4222_;
  wire not_new_n2989_;
  wire not_new_n6869_;
  wire not_new_n609__2;
  wire not_new_n599__332329305696010;
  wire not_new_n8892__0;
  wire not_new_n629__10;
  wire not_new_n7658_;
  wire not_new_n628__797922662976120010;
  wire not_new_n1576__2824752490;
  wire new_n8610_;
  wire not_new_n9132_;
  wire new_n5612_;
  wire not_new_n9218_;
  wire not_pi209;
  wire new_n2214_;
  wire new_n1852_;
  wire not_new_n5503_;
  wire or_or_not_new_n2110__not_new_n2111__not_new_n2113_;
  wire not_new_n5095_;
  wire new_n9507_;
  wire new_n4232_;
  wire not_new_n6480_;
  wire not_new_n8115_;
  wire new_n4559_;
  wire new_n9405_;
  wire not_new_n8159__0;
  wire not_new_n2954_;
  wire not_new_n638__24010;
  wire not_new_n4044_;
  wire not_new_n593__2326305139872070;
  wire new_n6776_;
  wire not_new_n696_;
  wire not_new_n9907_;
  wire new_n9662_;
  wire not_new_n612__1;
  wire new_n2678_;
  wire not_new_n3319_;
  wire not_new_n3161_;
  wire new_n6059_;
  wire not_new_n1324_;
  wire not_new_n5082_;
  wire new_n5267_;
  wire not_new_n4576_;
  wire new_n4057_;
  wire new_n5198_;
  wire new_n5438_;
  wire not_new_n644__24010;
  wire or_not_new_n1259__not_new_n1257_;
  wire not_po296_6782230728490;
  wire not_new_n4120__2;
  wire not_new_n1051__8235430;
  wire new_n3445_;
  wire not_new_n1053__2824752490;
  wire not_new_n8938_;
  wire not_new_n7576_;
  wire not_new_n1041__3;
  wire not_new_n3957__0;
  wire new_n8582_;
  wire not_new_n2199_;
  wire not_new_n2695_;
  wire new_n4400_;
  wire new_n3874_;
  wire new_n9181_;
  wire not_new_n990_;
  wire not_new_n8106__1;
  wire not_new_n1164__0;
  wire new_n2254_;
  wire not_new_n1599__57648010;
  wire not_new_n646__2;
  wire new_n10339_;
  wire new_n8336_;
  wire new_n6920_;
  wire new_n10292_;
  wire not_new_n9365__1;
  wire not_new_n604__168070;
  wire not_new_n1588__0;
  wire not_pi053_1;
  wire not_new_n964_;
  wire not_new_n1063__7;
  wire not_new_n5747_;
  wire not_new_n4574_;
  wire new_n1584_;
  wire new_n5622_;
  wire not_new_n9321_;
  wire not_new_n2838_;
  wire new_n4861_;
  wire new_n10323_;
  wire not_new_n7809_;
  wire new_n1616_;
  wire not_new_n2150_;
  wire new_n1698_;
  wire not_new_n1061__2326305139872070;
  wire new_n2200_;
  wire new_n9687_;
  wire new_n7217_;
  wire new_n8788_;
  wire new_n9474_;
  wire not_pi007;
  wire new_n6481_;
  wire new_n6737_;
  wire not_new_n8696_;
  wire not_new_n4486_;
  wire not_new_n1008__6;
  wire new_n1416_;
  wire new_n1274_;
  wire new_n8346_;
  wire not_new_n5047_;
  wire not_new_n2129_;
  wire new_n4834_;
  wire new_n10249_;
  wire new_n9746_;
  wire not_new_n619__7;
  wire not_new_n5179_;
  wire not_new_n7942_;
  wire new_n8115_;
  wire new_n1760_;
  wire not_new_n6305_;
  wire new_n8627_;
  wire po060;
  wire not_new_n1536__57648010;
  wire not_new_n4758_;
  wire not_new_n5260_;
  wire new_n8989_;
  wire new_n8798_;
  wire new_n6248_;
  wire not_new_n581__1070069044235980333563563003849377848070;
  wire or_not_new_n2110__not_new_n2111_;
  wire new_n6036_;
  wire not_new_n1580__138412872010;
  wire new_n8334_;
  wire not_new_n3135_;
  wire not_new_n7630_;
  wire not_new_n5087_;
  wire new_n2836_;
  wire new_n10129_;
  wire new_n3872_;
  wire not_new_n3133_;
  wire not_new_n1071__24010;
  wire new_n4130_;
  wire not_new_n2961_;
  wire new_n2569_;
  wire not_new_n8454_;
  wire not_new_n3951_;
  wire not_new_n589__138412872010;
  wire not_new_n6816_;
  wire and_new_n2667__new_n2668_;
  wire not_pi190_0;
  wire not_new_n3311__1;
  wire or_or_not_new_n1307__not_new_n1305__not_new_n2154_;
  wire not_new_n10029__3;
  wire not_new_n599__10;
  wire not_new_n7587_;
  wire not_new_n589__1577753820348458066150427430;
  wire or_or_not_new_n1996__not_new_n1997__not_new_n1999_;
  wire not_new_n4105_;
  wire or_not_new_n2874__not_new_n2877_;
  wire or_or_not_new_n2567__not_new_n2571__not_new_n1429_;
  wire and_new_n2257__new_n2260_;
  wire new_n3033_;
  wire not_new_n5054_;
  wire not_new_n6648_;
  wire not_new_n697_;
  wire not_new_n5781__0;
  wire new_n957_;
  wire not_new_n7672_;
  wire or_or_not_new_n1339__not_new_n1337__not_new_n2306_;
  wire not_new_n7599__0;
  wire not_new_n3315__8235430;
  wire new_n2408_;
  wire not_new_n625__1176490;
  wire not_new_n1452_;
  wire not_new_n635__70;
  wire new_n9294_;
  wire or_not_new_n2939__not_new_n1485_;
  wire not_pi020;
  wire not_new_n7899_;
  wire new_n8948_;
  wire not_new_n5832_;
  wire not_new_n7205_;
  wire not_new_n1051__19773267430;
  wire new_n8175_;
  wire not_new_n581__225393402906922580878632490;
  wire not_new_n8368__0;
  wire not_new_n1002__4;
  wire new_n3867_;
  wire not_new_n4837__1;
  wire not_new_n1279_;
  wire key_gate_73;
  wire new_n9154_;
  wire or_or_not_new_n1563__not_new_n2474__not_new_n1395_;
  wire new_n3258_;
  wire not_new_n4321__0;
  wire not_new_n3554_;
  wire not_pi258_0;
  wire new_n8846_;
  wire or_or_not_new_n2892__not_new_n2895__not_new_n2894_;
  wire new_n6808_;
  wire or_not_new_n7939__not_new_n7913_;
  wire new_n3582_;
  wire po121;
  wire new_n1421_;
  wire not_new_n3440_;
  wire new_n2248_;
  wire new_n4895_;
  wire not_pi027_0;
  wire new_n2165_;
  wire new_n8351_;
  wire new_n8384_;
  wire po041;
  wire not_new_n9186__0;
  wire not_new_n3499_;
  wire new_n1751_;
  wire not_new_n5172_;
  wire not_new_n1039__273687473400809163430;
  wire not_new_n2712_;
  wire not_new_n1570_;
  wire not_new_n9828_;
  wire not_new_n1037__19773267430;
  wire new_n9120_;
  wire new_n2404_;
  wire new_n596_;
  wire new_n9743_;
  wire new_n8357_;
  wire not_new_n1035__8;
  wire not_new_n9422__0;
  wire not_new_n7275_;
  wire not_new_n1602__168070;
  wire new_n3706_;
  wire not_pi038;
  wire and_new_n2637__new_n2638_;
  wire not_new_n3310__1176490;
  wire not_new_n3699_;
  wire not_new_n4137_;
  wire new_n4363_;
  wire not_new_n3185__138412872010;
  wire not_new_n4206_;
  wire not_new_n1538__6782230728490;
  wire new_n6716_;
  wire new_n3452_;
  wire not_new_n1027__332329305696010;
  wire or_or_not_new_n1566__not_new_n2489__not_new_n1401_;
  wire new_n5509_;
  wire not_new_n2894_;
  wire not_new_n3420_;
  wire not_new_n8943_;
  wire new_n7951_;
  wire new_n6108_;
  wire not_new_n4543_;
  wire not_new_n5180_;
  wire not_pi002_0;
  wire not_new_n5106_;
  wire not_new_n1008_;
  wire and_new_n9696__new_n9695_;
  wire new_n5268_;
  wire new_n4143_;
  wire new_n10231_;
  wire new_n4929_;
  wire or_not_new_n3136__not_new_n3137_;
  wire new_n5950_;
  wire not_new_n5611_;
  wire new_n10086_;
  wire new_n3405_;
  wire new_n10148_;
  wire not_new_n2874_;
  wire not_new_n1538__3430;
  wire new_n5336_;
  wire not_new_n9909__0;
  wire new_n6212_;
  wire new_n7385_;
  wire not_new_n1364_;
  wire not_new_n1844_;
  wire not_new_n1600__9;
  wire not_new_n1014__3;
  wire not_new_n601__0;
  wire new_n3090_;
  wire new_n8782_;
  wire or_or_not_new_n6340__not_new_n6341__not_new_n6342_;
  wire new_n2239_;
  wire not_new_n1017__2;
  wire new_n9344_;
  wire not_new_n4127__1;
  wire not_new_n1583__138412872010;
  wire new_n8015_;
  wire new_n3702_;
  wire not_new_n7415__1;
  wire new_n3216_;
  wire po182;
  wire not_new_n5954_;
  wire not_new_n4258_;
  wire not_new_n605__8;
  wire new_n6004_;
  wire not_new_n2059_;
  wire not_new_n2509__57648010;
  wire not_new_n4520_;
  wire not_new_n4771__0;
  wire not_new_n5434__0;
  wire new_n8378_;
  wire new_n1929_;
  wire not_new_n660_;
  wire new_n8683_;
  wire not_new_n5509_;
  wire not_new_n8105__0;
  wire not_new_n9692_;
  wire not_new_n1039__57648010;
  wire new_n4890_;
  wire new_n8003_;
  wire not_new_n7472_;
  wire new_n5946_;
  wire not_new_n3184__10;
  wire new_n6356_;
  wire new_n3564_;
  wire new_n5905_;
  wire not_new_n1603__0;
  wire not_new_n643__39098210485829880490;
  wire not_new_n607__24010;
  wire not_new_n1027__1176490;
  wire new_n1232_;
  wire key_gate_46;
  wire not_pi004;
  wire not_new_n9995_;
  wire new_n7338_;
  wire new_n9706_;
  wire new_n1885_;
  wire not_new_n7970_;
  wire not_new_n5433_;
  wire not_new_n8234_;
  wire not_new_n6500__0;
  wire new_n1352_;
  wire new_n8919_;
  wire not_new_n4973_;
  wire not_new_n5281_;
  wire not_new_n5604_;
  wire new_n10283_;
  wire not_new_n9255_;
  wire new_n7154_;
  wire not_new_n5126_;
  wire new_n2990_;
  wire and_new_n6373__new_n6398_;
  wire new_n2000_;
  wire or_not_new_n9704__not_new_n9705_;
  wire not_new_n5831_;
  wire not_new_n1051__47475615099430;
  wire not_new_n1211_;
  wire po037;
  wire new_n7051_;
  wire not_new_n9165_;
  wire not_new_n8361_;
  wire not_new_n3721_;
  wire not_new_n600__8235430;
  wire not_new_n6677_;
  wire not_new_n3407_;
  wire not_pi198;
  wire not_new_n590__4;
  wire new_n2524_;
  wire not_new_n8152_;
  wire new_n7520_;
  wire not_new_n4984__0;
  wire new_n2436_;
  wire not_new_n4123__0;
  wire not_new_n1584__24010;
  wire new_n6598_;
  wire not_new_n2922_;
  wire not_new_n628__2;
  wire new_n6680_;
  wire not_new_n7613__0;
  wire not_new_n7817_;
  wire not_new_n727_;
  wire not_new_n1037__4;
  wire not_new_n1069__2;
  wire not_pi143;
  wire not_new_n6802_;
  wire not_new_n7503_;
  wire not_new_n8845__1;
  wire new_n9103_;
  wire not_new_n9941_;
  wire not_new_n9797_;
  wire not_new_n8879__0;
  wire new_n3654_;
  wire new_n2001_;
  wire not_new_n8218_;
  wire not_new_n607__1176490;
  wire new_n2564_;
  wire not_new_n634__5585458640832840070;
  wire not_new_n6834_;
  wire new_n9098_;
  wire not_pi248_2;
  wire not_new_n5259_;
  wire not_pi171_2;
  wire not_new_n1343_;
  wire or_or_not_new_n2129__not_new_n2130__not_new_n2132_;
  wire new_n5489_;
  wire or_not_new_n1479__not_new_n1480_;
  wire not_new_n612__6;
  wire not_new_n4808__0;
  wire new_n2498_;
  wire new_n3754_;
  wire new_n4452_;
  wire not_new_n9488_;
  wire new_n5418_;
  wire new_n6372_;
  wire not_new_n1049__24010;
  wire new_n3945_;
  wire not_new_n9009_;
  wire not_pi159;
  wire not_new_n645__113988951853731430;
  wire not_new_n639__968890104070;
  wire not_new_n601__2326305139872070;
  wire not_new_n4843_;
  wire not_new_n6758_;
  wire not_po296_17984650426474121466202803405696493492512490;
  wire not_new_n6974__138412872010;
  wire not_new_n10006__0;
  wire new_n2870_;
  wire not_new_n7351__0;
  wire not_new_n6503__2;
  wire key_gate_89;
  wire new_n1780_;
  wire new_n701_;
  wire new_n1566_;
  wire new_n8558_;
  wire and_new_n5084__new_n5345_;
  wire not_new_n3100_;
  wire not_new_n9826_;
  wire new_n6646_;
  wire not_new_n586__1176490;
  wire new_n2378_;
  wire not_new_n3984_;
  wire not_new_n7561_;
  wire new_n4471_;
  wire new_n6642_;
  wire not_new_n4004_;
  wire not_new_n1763_;
  wire new_n4995_;
  wire new_n5579_;
  wire new_n1803_;
  wire new_n5569_;
  wire not_new_n6815_;
  wire new_n3892_;
  wire new_n9132_;
  wire po216;
  wire not_new_n7853_;
  wire new_n7931_;
  wire new_n1390_;
  wire not_new_n7583_;
  wire new_n4911_;
  wire not_new_n1631__70;
  wire not_new_n9179_;
  wire not_new_n641__5;
  wire new_n3255_;
  wire not_new_n4829_;
  wire not_new_n7549_;
  wire not_new_n10049_;
  wire not_new_n7135_;
  wire not_new_n10011_;
  wire not_new_n3184__6782230728490;
  wire not_new_n6443__332329305696010;
  wire not_new_n637__490;
  wire new_n3871_;
  wire new_n7115_;
  wire not_new_n1071__1176490;
  wire new_n6931_;
  wire new_n2499_;
  wire not_new_n619_;
  wire not_new_n3697_;
  wire new_n7724_;
  wire new_n5603_;
  wire not_new_n5905__1;
  wire not_new_n6027_;
  wire not_new_n1612__0;
  wire new_n6979_;
  wire not_new_n745_;
  wire new_n10058_;
  wire not_pi123_0;
  wire not_new_n928__113988951853731430;
  wire not_new_n6913_;
  wire not_new_n3875_;
  wire not_new_n4128_;
  wire not_new_n6183_;
  wire not_pi271_0;
  wire not_new_n4733_;
  wire not_new_n640__57648010;
  wire new_n5158_;
  wire not_new_n9486_;
  wire not_new_n8342_;
  wire po125;
  wire new_n766_;
  wire not_new_n7619_;
  wire not_new_n638__16284135979104490;
  wire new_n4593_;
  wire not_new_n9938_;
  wire new_n5696_;
  wire or_not_new_n7463__not_new_n7312_;
  wire new_n7168_;
  wire new_n5750_;
  wire not_new_n2912_;
  wire new_n2904_;
  wire not_new_n6579_;
  wire not_new_n638__113988951853731430;
  wire new_n10202_;
  wire new_n2803_;
  wire not_new_n6992_;
  wire not_new_n1196_;
  wire new_n9008_;
  wire not_new_n8273_;
  wire not_new_n1069__19773267430;
  wire not_new_n1598__19773267430;
  wire new_n8064_;
  wire not_new_n1616__2824752490;
  wire not_new_n9119_;
  wire not_new_n627__138412872010;
  wire new_n5250_;
  wire new_n615_;
  wire new_n3838_;
  wire or_or_not_new_n1763__not_new_n1764__not_new_n1766_;
  wire not_new_n5506_;
  wire not_new_n6781_;
  wire not_new_n8641_;
  wire new_n9796_;
  wire not_new_n4770__0;
  wire not_new_n2173_;
  wire new_n5393_;
  wire not_new_n4790_;
  wire not_new_n8438_;
  wire not_new_n1534__6782230728490;
  wire new_n1417_;
  wire new_n767_;
  wire not_new_n5195_;
  wire or_not_new_n1027__not_new_n1028__0;
  wire new_n1583_;
  wire not_pi138_3;
  wire new_n7643_;
  wire new_n2674_;
  wire not_new_n628__2824752490;
  wire or_not_new_n3161__not_new_n3160_;
  wire not_new_n1019__3;
  wire not_new_n7292_;
  wire po143;
  wire new_n7734_;
  wire new_n4336_;
  wire new_n7886_;
  wire not_new_n4577__0;
  wire new_n9901_;
  wire new_n10093_;
  wire new_n6545_;
  wire new_n4124_;
  wire new_n1445_;
  wire not_new_n2001_;
  wire new_n9575_;
  wire new_n1948_;
  wire new_n2266_;
  wire not_new_n6511__0;
  wire new_n4455_;
  wire new_n1643_;
  wire not_new_n7510_;
  wire new_n3554_;
  wire not_new_n5194_;
  wire po027;
  wire or_not_new_n1825__not_new_n1826_;
  wire new_n3776_;
  wire not_new_n3311__2;
  wire not_new_n6974__2;
  wire new_n8234_;
  wire new_n3066_;
  wire not_new_n624__1176490;
  wire new_n953_;
  wire new_n8733_;
  wire not_new_n9973__0;
  wire not_new_n8697_;
  wire not_new_n9960_;
  wire new_n8200_;
  wire not_new_n10022_;
  wire not_new_n6978__0;
  wire not_new_n2960_;
  wire not_new_n9070_;
  wire new_n6789_;
  wire not_new_n3688_;
  wire not_new_n8967_;
  wire new_n9568_;
  wire new_n663_;
  wire new_n7293_;
  wire not_new_n634__6782230728490;
  wire or_not_new_n6354__not_new_n6373__8;
  wire not_po296_57648010;
  wire not_new_n6901_;
  wire new_n10244_;
  wire not_new_n6581_;
  wire not_new_n2908_;
  wire not_new_n9915_;
  wire new_n5457_;
  wire not_new_n1016__1;
  wire new_n8808_;
  wire not_new_n994__0;
  wire not_new_n7992_;
  wire new_n9142_;
  wire not_new_n633__10;
  wire new_n7975_;
  wire not_new_n4117__2;
  wire not_new_n3564_;
  wire new_n4300_;
  wire new_n6446_;
  wire not_new_n6259_;
  wire not_pi046;
  wire new_n1254_;
  wire not_new_n4133__0;
  wire not_new_n4120__1;
  wire not_pi098_0;
  wire new_n2716_;
  wire new_n9998_;
  wire not_new_n9568_;
  wire not_new_n3913_;
  wire new_n4079_;
  wire not_new_n599__19773267430;
  wire new_n1518_;
  wire new_n1187_;
  wire not_new_n6294_;
  wire new_n5819_;
  wire new_n7251_;
  wire not_new_n6317__0;
  wire not_new_n602__1176490;
  wire not_new_n643__5585458640832840070;
  wire new_n8993_;
  wire not_new_n1580__57648010;
  wire not_new_n7023_;
  wire not_new_n10163_;
  wire not_new_n9505_;
  wire new_n3993_;
  wire new_n7559_;
  wire not_new_n8384_;
  wire not_new_n1613__0;
  wire not_new_n646__403536070;
  wire new_n3263_;
  wire not_new_n8975_;
  wire not_new_n595__0;
  wire new_n5310_;
  wire new_n3581_;
  wire not_new_n8284_;
  wire not_new_n608_;
  wire not_new_n635__168070;
  wire new_n3361_;
  wire new_n6430_;
  wire new_n5130_;
  wire new_n3753_;
  wire not_new_n9951__1;
  wire not_new_n3831_;
  wire not_new_n4134__1;
  wire not_new_n621__39098210485829880490;
  wire new_n1521_;
  wire not_new_n6312_;
  wire new_n4146_;
  wire not_new_n638__3;
  wire not_new_n1067__47475615099430;
  wire new_n8090_;
  wire new_n9452_;
  wire not_new_n6443__8;
  wire new_n2487_;
  wire not_new_n9813_;
  wire not_new_n7772_;
  wire not_new_n1069__168070;
  wire new_n8016_;
  wire new_n5544_;
  wire po059;
  wire new_n9399_;
  wire not_new_n3182_;
  wire not_new_n1645_;
  wire new_n924_;
  wire not_new_n644__10;
  wire new_n7252_;
  wire new_n10330_;
  wire new_n9480_;
  wire not_new_n6888_;
  wire new_n10262_;
  wire new_n4299_;
  wire not_new_n2166_;
  wire not_new_n1043__332329305696010;
  wire not_new_n8049_;
  wire new_n5047_;
  wire new_n5763_;
  wire not_new_n940_;
  wire not_new_n7159_;
  wire not_new_n6498__1;
  wire not_new_n636__19773267430;
  wire new_n7489_;
  wire not_new_n589__968890104070;
  wire not_new_n6443__4;
  wire new_n1479_;
  wire not_new_n610__4;
  wire new_n9535_;
  wire not_new_n6647__0;
  wire not_new_n5779_;
  wire not_new_n10150_;
  wire new_n5715_;
  wire new_n3367_;
  wire not_new_n8275__0;
  wire new_n9750_;
  wire new_n8904_;
  wire new_n1399_;
  wire not_new_n1585__7;
  wire new_n9016_;
  wire not_new_n6917_;
  wire not_new_n1604__168070;
  wire new_n6882_;
  wire not_new_n598__57648010;
  wire new_n9194_;
  wire new_n8260_;
  wire not_new_n7022__1;
  wire not_new_n8021_;
  wire not_new_n3315_;
  wire not_new_n1601__10;
  wire not_new_n624__168070;
  wire not_new_n6609_;
  wire new_n620_;
  wire new_n2080_;
  wire not_pi158_0;
  wire new_n8672_;
  wire not_new_n3384__2;
  wire new_n1794_;
  wire not_new_n1039__70;
  wire new_n6983_;
  wire or_or_not_new_n1311__not_new_n1309__not_new_n2173_;
  wire new_n6327_;
  wire or_not_new_n2635__not_new_n2634_;
  wire new_n5565_;
  wire not_new_n641__6;
  wire not_new_n10207_;
  wire not_new_n3990__0;
  wire not_pi265;
  wire not_new_n2878_;
  wire not_pi153;
  wire po022;
  wire new_n5101_;
  wire not_new_n1047__2326305139872070;
  wire new_n1696_;
  wire new_n9634_;
  wire not_new_n1591__2824752490;
  wire not_new_n4791__0;
  wire not_new_n4969__0;
  wire new_n5261_;
  wire not_new_n1534__8235430;
  wire not_pi161_0;
  wire not_new_n6706_;
  wire new_n2333_;
  wire not_new_n6215_;
  wire not_new_n1055__138412872010;
  wire not_new_n2891_;
  wire not_new_n3586_;
  wire new_n3546_;
  wire not_new_n7344_;
  wire new_n5477_;
  wire po202;
  wire not_new_n3994_;
  wire new_n5077_;
  wire not_new_n5453_;
  wire new_n7950_;
  wire new_n753_;
  wire not_new_n7483_;
  wire not_new_n1045__2824752490;
  wire not_new_n634__113988951853731430;
  wire new_n3439_;
  wire not_new_n8443_;
  wire new_n9196_;
  wire not_new_n6585_;
  wire not_new_n621__10;
  wire not_new_n5726_;
  wire not_new_n9899__0;
  wire not_new_n928__57648010;
  wire not_new_n7144_;
  wire new_n3781_;
  wire new_n10131_;
  wire not_new_n4490_;
  wire po201;
  wire not_new_n593__168070;
  wire not_new_n589__6;
  wire new_n1801_;
  wire not_new_n3310_;
  wire new_n9867_;
  wire new_n5706_;
  wire new_n4167_;
  wire new_n2132_;
  wire new_n1833_;
  wire new_n8663_;
  wire not_new_n3188_;
  wire new_n5062_;
  wire and_new_n1953__new_n1956_;
  wire new_n9747_;
  wire not_new_n1588__2824752490;
  wire not_new_n3108_;
  wire not_new_n1035__70;
  wire not_new_n6348_;
  wire not_new_n5369_;
  wire new_n3295_;
  wire not_new_n8874_;
  wire not_new_n4170_;
  wire new_n1666_;
  wire not_new_n9951_;
  wire and_new_n8983__new_n9311_;
  wire new_n9213_;
  wire not_new_n9096_;
  wire new_n2883_;
  wire not_new_n4919_;
  wire not_new_n587__1176490;
  wire not_new_n7002__1;
  wire new_n5707_;
  wire not_new_n5930_;
  wire not_new_n1588__138412872010;
  wire not_new_n5713_;
  wire new_n8120_;
  wire new_n3113_;
  wire not_new_n8238_;
  wire new_n9167_;
  wire not_new_n1611__1176490;
  wire new_n1162_;
  wire not_new_n6673__0;
  wire not_new_n1599__0;
  wire new_n7177_;
  wire new_n6782_;
  wire new_n6707_;
  wire not_new_n1583__2326305139872070;
  wire not_new_n590__3;
  wire new_n5951_;
  wire not_new_n2057_;
  wire not_new_n3387__2;
  wire new_n2703_;
  wire not_new_n1061__2824752490;
  wire new_n3435_;
  wire not_new_n8323_;
  wire not_new_n2951_;
  wire not_new_n8388_;
  wire new_n9786_;
  wire not_new_n604__8;
  wire not_new_n8253__0;
  wire new_n8649_;
  wire new_n6860_;
  wire new_n2373_;
  wire not_new_n637__332329305696010;
  wire new_n5054_;
  wire not_new_n3174_;
  wire not_new_n5638_;
  wire new_n8085_;
  wire new_n1308_;
  wire not_new_n9556__0;
  wire not_new_n8010_;
  wire not_new_n7231_;
  wire new_n5768_;
  wire not_new_n581__152867006319425761937651857692768264010;
  wire new_n7111_;
  wire not_new_n7006__0;
  wire not_new_n645__2824752490;
  wire not_new_n925__0;
  wire new_n4145_;
  wire new_n6237_;
  wire not_new_n5440__0;
  wire not_new_n9889__0;
  wire not_new_n3997_;
  wire or_not_new_n7047__0_not_new_n3369__0;
  wire not_new_n5487__0;
  wire new_n4233_;
  wire new_n6123_;
  wire not_new_n6688_;
  wire not_new_n1923_;
  wire not_new_n1825_;
  wire not_new_n4132_;
  wire not_new_n598__2824752490;
  wire new_n7276_;
  wire not_new_n6026_;
  wire not_new_n5983_;
  wire new_n3321_;
  wire new_n1464_;
  wire new_n5591_;
  wire not_new_n5110_;
  wire not_pi042_2;
  wire new_n7227_;
  wire new_n8497_;
  wire new_n7260_;
  wire not_new_n8889_;
  wire or_not_new_n4319__0_not_new_n713_;
  wire not_pi044_3;
  wire new_n4990_;
  wire new_n685_;
  wire new_n1524_;
  wire not_new_n7310_;
  wire new_n2710_;
  wire not_new_n8156_;
  wire new_n3735_;
  wire not_new_n5086_;
  wire not_new_n8036_;
  wire new_n1675_;
  wire not_new_n6474__2;
  wire new_n605_;
  wire not_new_n4729_;
  wire not_pi099_0;
  wire not_new_n1589_;
  wire not_new_n9008_;
  wire new_n4020_;
  wire new_n6420_;
  wire not_new_n645__8235430;
  wire not_new_n1613__1;
  wire new_n1330_;
  wire not_new_n3347_;
  wire new_n7922_;
  wire not_pi191_0;
  wire new_n2421_;
  wire not_new_n1596__0;
  wire new_n2305_;
  wire new_n3667_;
  wire not_new_n1490_;
  wire new_n5464_;
  wire not_new_n985__0;
  wire and_new_n6473__new_n6833_;
  wire new_n4241_;
  wire not_pi271;
  wire not_new_n1609_;
  wire new_n7266_;
  wire new_n5382_;
  wire new_n7039_;
  wire not_new_n1339_;
  wire not_new_n1585__8235430;
  wire not_new_n5707_;
  wire new_n8478_;
  wire not_new_n9151_;
  wire not_new_n6988_;
  wire not_new_n6974__5;
  wire not_new_n1601__9;
  wire new_n1552_;
  wire not_new_n8099_;
  wire not_new_n9265_;
  wire new_n5631_;
  wire new_n4125_;
  wire new_n9466_;
  wire not_new_n5128__0;
  wire not_new_n643__57648010;
  wire not_new_n7622__0;
  wire not_new_n763_;
  wire new_n5232_;
  wire not_new_n6470_;
  wire new_n9684_;
  wire not_new_n10056_;
  wire new_n8257_;
  wire new_n1248_;
  wire or_or_not_new_n2982__not_new_n2985__not_new_n2984_;
  wire not_new_n6205_;
  wire new_n8741_;
  wire not_new_n5765__0;
  wire new_n4970_;
  wire not_new_n7762_;
  wire not_new_n8062_;
  wire not_new_n9971__0;
  wire new_n6352_;
  wire not_new_n1538__2326305139872070;
  wire not_new_n6974__490;
  wire not_new_n1603__57648010;
  wire not_new_n9458_;
  wire not_new_n599__2326305139872070;
  wire not_new_n2991_;
  wire not_pi235;
  wire not_new_n6623_;
  wire new_n1005_;
  wire new_n4495_;
  wire not_new_n1518_;
  wire not_new_n5062_;
  wire not_new_n4318_;
  wire not_new_n2071_;
  wire not_new_n6443__6782230728490;
  wire not_new_n1613__16284135979104490;
  wire new_n8943_;
  wire not_new_n8855__0;
  wire or_not_new_n2685__not_new_n2684_;
  wire not_new_n4797__0;
  wire not_new_n1027__5585458640832840070;
  wire new_n8950_;
  wire not_new_n609__8;
  wire new_n5752_;
  wire new_n2965_;
  wire po107;
  wire not_new_n6443__490;
  wire new_n7312_;
  wire not_new_n1611__1;
  wire new_n2451_;
  wire new_n2431_;
  wire not_new_n1616__10;
  wire new_n9292_;
  wire new_n2717_;
  wire not_new_n8675_;
  wire new_n4821_;
  wire new_n3551_;
  wire and_new_n1258__new_n1932_;
  wire new_n961_;
  wire not_new_n9324_;
  wire not_new_n3671_;
  wire not_new_n2724_;
  wire not_new_n6640__1;
  wire not_new_n4799__0;
  wire or_or_not_new_n2727__not_new_n2730__not_new_n2729_;
  wire not_new_n1055__1;
  wire not_new_n1593_;
  wire not_new_n9040_;
  wire not_new_n9903_;
  wire not_new_n5808__0;
  wire not_new_n6754_;
  wire not_new_n775__47475615099430;
  wire new_n768_;
  wire new_n9384_;
  wire not_new_n3315__6782230728490;
  wire not_new_n3490_;
  wire new_n5568_;
  wire not_new_n1410_;
  wire not_new_n2110_;
  wire not_new_n1957__0;
  wire not_new_n1059__168070;
  wire new_n7173_;
  wire not_new_n8554_;
  wire not_pi145_2;
  wire not_new_n1037__1176490;
  wire not_new_n7240__0;
  wire not_pi050_1;
  wire po196;
  wire new_n4664_;
  wire not_new_n633__6782230728490;
  wire not_new_n588__403536070;
  wire not_new_n1386_;
  wire not_new_n3184__3;
  wire not_new_n10052_;
  wire not_new_n3920_;
  wire po277;
  wire not_pi155_0;
  wire not_new_n4439_;
  wire not_new_n1194_;
  wire new_n3349_;
  wire not_new_n1611__138412872010;
  wire not_new_n645__332329305696010;
  wire new_n7143_;
  wire new_n5012_;
  wire not_new_n1616__7;
  wire not_new_n8138_;
  wire not_new_n595__19773267430;
  wire not_pi048;
  wire not_new_n1605__6;
  wire new_n7006_;
  wire not_new_n1846_;
  wire new_n9113_;
  wire not_new_n1604__3430;
  wire not_new_n9092_;
  wire new_n3855_;
  wire not_new_n5859_;
  wire not_new_n8158_;
  wire new_n9753_;
  wire not_new_n581__2326305139872070;
  wire not_new_n5767__0;
  wire new_n7733_;
  wire new_n1786_;
  wire not_new_n7178_;
  wire new_n4686_;
  wire not_new_n4727__0;
  wire not_new_n7926_;
  wire not_new_n4778_;
  wire not_pi030_0;
  wire new_n5920_;
  wire not_new_n9908_;
  wire not_new_n7465_;
  wire not_new_n5294_;
  wire new_n8659_;
  wire new_n2771_;
  wire not_new_n9897_;
  wire not_new_n1611__332329305696010;
  wire not_new_n6296_;
  wire not_new_n1705_;
  wire new_n6489_;
  wire not_new_n7617__0;
  wire new_n6279_;
  wire not_new_n1023__4;
  wire not_new_n1576__16284135979104490;
  wire new_n5755_;
  wire not_new_n4532_;
  wire not_new_n2509__490;
  wire not_new_n6973_;
  wire new_n9593_;
  wire not_new_n1069__490;
  wire new_n8319_;
  wire new_n3537_;
  wire not_new_n1980_;
  wire not_new_n636__57648010;
  wire not_new_n4419__0;
  wire not_new_n625__168070;
  wire new_n4498_;
  wire or_not_new_n4833__not_new_n4782_;
  wire not_new_n5386_;
  wire not_pi180_1;
  wire not_pi009;
  wire not_new_n10164_;
  wire new_n6786_;
  wire not_new_n6819_;
  wire not_new_n5435_;
  wire new_n5762_;
  wire new_n2337_;
  wire po200;
  wire new_n5122_;
  wire new_n4383_;
  wire new_n5859_;
  wire new_n1336_;
  wire new_n8316_;
  wire not_new_n643__273687473400809163430;
  wire not_new_n7096_;
  wire not_new_n2094_;
  wire new_n8687_;
  wire new_n2393_;
  wire or_not_new_n3164__not_new_n3163_;
  wire not_new_n8110_;
  wire not_new_n2565_;
  wire not_new_n1611__168070;
  wire not_new_n5778_;
  wire not_new_n3748_;
  wire po018;
  wire new_n10007_;
  wire not_new_n1191_;
  wire new_n8392_;
  wire not_new_n9117_;
  wire not_new_n589_;
  wire not_new_n5706__0;
  wire new_n8288_;
  wire not_new_n3094_;
  wire not_new_n7072_;
  wire new_n8044_;
  wire not_new_n9480_;
  wire not_new_n7013__0;
  wire new_n4563_;
  wire new_n8599_;
  wire not_new_n3794_;
  wire new_n4230_;
  wire po252;
  wire not_new_n2895_;
  wire not_new_n4161__0;
  wire new_n3634_;
  wire not_new_n604__9;
  wire new_n1466_;
  wire not_new_n603__168070;
  wire not_new_n6996_;
  wire new_n3671_;
  wire not_new_n9884_;
  wire not_new_n1010__2;
  wire po233;
  wire new_n7831_;
  wire new_n5798_;
  wire new_n10083_;
  wire new_n2185_;
  wire not_new_n958_;
  wire not_new_n4344_;
  wire not_new_n1027__57648010;
  wire not_new_n1606__6;
  wire new_n2826_;
  wire new_n10213_;
  wire not_new_n7406__1;
  wire new_n5152_;
  wire new_n5730_;
  wire new_n3774_;
  wire not_new_n2892_;
  wire new_n4918_;
  wire not_new_n8268_;
  wire not_new_n7019__0;
  wire not_new_n9395_;
  wire new_n8761_;
  wire or_not_new_n1787__not_new_n1788_;
  wire not_new_n4076_;
  wire new_n3552_;
  wire not_new_n945_;
  wire new_n2416_;
  wire new_n4943_;
  wire not_new_n6247_;
  wire new_n6056_;
  wire not_new_n6214_;
  wire new_n7397_;
  wire new_n4470_;
  wire new_n3203_;
  wire not_new_n1534__332329305696010;
  wire not_new_n6522__0;
  wire not_new_n6915_;
  wire new_n3370_;
  wire new_n9267_;
  wire not_new_n10068_;
  wire new_n9335_;
  wire new_n1870_;
  wire new_n1483_;
  wire not_new_n1831_;
  wire not_new_n5084_;
  wire new_n7141_;
  wire not_new_n594__168070;
  wire not_new_n1071__168070;
  wire not_new_n1057__57648010;
  wire not_new_n1611__10;
  wire new_n5389_;
  wire new_n3465_;
  wire not_new_n1061__332329305696010;
  wire or_not_new_n1572__0_not_new_n1028__6;
  wire new_n5496_;
  wire not_new_n8906_;
  wire new_n9555_;
  wire not_new_n9327__1;
  wire new_n6061_;
  wire new_n8451_;
  wire new_n7415_;
  wire or_not_new_n8172__0_not_new_n1596__138412872010;
  wire not_new_n9037_;
  wire new_n9270_;
  wire not_new_n9259_;
  wire not_new_n9063_;
  wire not_new_n4901_;
  wire not_new_n605_;
  wire not_new_n6979_;
  wire not_new_n2863_;
  wire new_n2153_;
  wire not_new_n7530_;
  wire not_new_n6729_;
  wire not_new_n1591__968890104070;
  wire not_new_n2071__0;
  wire not_new_n3993_;
  wire not_new_n1603__6782230728490;
  wire not_new_n1006__2;
  wire new_n7178_;
  wire not_new_n3379_;
  wire not_new_n1359_;
  wire not_new_n1603__8235430;
  wire new_n5835_;
  wire not_new_n1149_;
  wire not_new_n1536__168070;
  wire not_new_n4986__0;
  wire new_n4693_;
  wire new_n6831_;
  wire not_new_n1600__1176490;
  wire new_n9519_;
  wire not_new_n1606_;
  wire not_new_n1045__3430;
  wire new_n9815_;
  wire not_new_n7209_;
  wire not_new_n9501_;
  wire new_n1205_;
  wire not_new_n5064_;
  wire new_n2605_;
  wire not_new_n3521_;
  wire new_n2204_;
  wire new_n7306_;
  wire new_n5147_;
  wire new_n8093_;
  wire not_new_n601__968890104070;
  wire new_n10211_;
  wire po232;
  wire not_pi130_2;
  wire not_new_n2503_;
  wire not_pi066;
  wire not_new_n724__1;
  wire not_new_n3540_;
  wire not_new_n5091__0;
  wire not_new_n928__8;
  wire not_new_n7025__1;
  wire not_new_n4278_;
  wire not_new_n1002__5;
  wire new_n8405_;
  wire new_n9433_;
  wire not_new_n5882_;
  wire not_new_n6629_;
  wire not_new_n1045__490;
  wire new_n2423_;
  wire new_n6227_;
  wire not_new_n3896_;
  wire not_new_n735__1;
  wire not_new_n1611__2;
  wire not_new_n6812_;
  wire po228;
  wire not_new_n1601__19773267430;
  wire and_and_and_new_n2325__new_n2332__new_n2333__new_n2329_;
  wire not_new_n767_;
  wire new_n3397_;
  wire not_new_n7036__0;
  wire new_n4428_;
  wire not_new_n1580__7;
  wire new_n8848_;
  wire not_new_n6920_;
  wire po172;
  wire not_new_n1583__3;
  wire not_new_n3770_;
  wire not_new_n5617__1;
  wire new_n8096_;
  wire and_new_n3082__new_n998_;
  wire or_not_new_n7313__not_new_n7314_;
  wire or_or_or_not_new_n2883__not_new_n2886__not_new_n2885__not_new_n2887_;
  wire new_n4717_;
  wire not_new_n1041__10;
  wire or_not_new_n7908__not_new_n7743_;
  wire new_n6987_;
  wire not_new_n7419_;
  wire key_gate_58;
  wire not_new_n1581__138412872010;
  wire new_n3093_;
  wire not_new_n3486_;
  wire new_n4590_;
  wire not_new_n7448_;
  wire not_new_n3220_;
  wire not_new_n4160_;
  wire not_new_n7187_;
  wire not_new_n5488_;
  wire not_new_n8148_;
  wire not_new_n4592_;
  wire new_n5756_;
  wire new_n7121_;
  wire not_new_n632__968890104070;
  wire new_n1262_;
  wire not_new_n9944__0;
  wire and_and_new_n2219__new_n2222__new_n2220_;
  wire not_new_n1039__8;
  wire new_n8959_;
  wire new_n4203_;
  wire not_new_n3682_;
  wire new_n5621_;
  wire new_n1211_;
  wire new_n974_;
  wire new_n4315_;
  wire new_n1292_;
  wire not_new_n597__3;
  wire not_new_n8716__0;
  wire not_new_n8083_;
  wire not_new_n8117__0;
  wire new_n6002_;
  wire not_new_n6209_;
  wire not_new_n622__1176490;
  wire not_new_n3170_;
  wire new_n2656_;
  wire not_new_n6353_;
  wire not_new_n1537__6782230728490;
  wire not_new_n627__403536070;
  wire not_new_n7802_;
  wire not_new_n4307_;
  wire po023;
  wire new_n7860_;
  wire not_new_n3366__0;
  wire key_gate_120;
  wire new_n5387_;
  wire not_new_n581__5585458640832840070;
  wire not_new_n1538__2;
  wire new_n1032_;
  wire not_new_n4003__0;
  wire new_n5999_;
  wire new_n3259_;
  wire not_new_n1063__2;
  wire new_n7075_;
  wire not_new_n7873_;
  wire not_new_n2743_;
  wire not_new_n617__113988951853731430;
  wire or_not_new_n2845__not_new_n2844_;
  wire new_n7936_;
  wire new_n7897_;
  wire not_new_n618__5;
  wire new_n5664_;
  wire not_new_n607__9;
  wire new_n8183_;
  wire new_n4510_;
  wire not_new_n8987_;
  wire new_n5861_;
  wire new_n4136_;
  wire not_new_n6180_;
  wire not_new_n9416__0;
  wire new_n2311_;
  wire not_new_n4937_;
  wire new_n9565_;
  wire not_new_n1598__70;
  wire not_new_n10280_;
  wire not_new_n1536__0;
  wire not_new_n7085_;
  wire new_n8681_;
  wire not_new_n1016__6;
  wire new_n8862_;
  wire or_not_new_n2557__not_new_n2561_;
  wire not_new_n9713_;
  wire not_new_n588__2326305139872070;
  wire new_n1440_;
  wire new_n10095_;
  wire new_n1320_;
  wire not_pi189;
  wire not_new_n1027__2824752490;
  wire not_new_n4618_;
  wire or_not_new_n1552__not_new_n2419_;
  wire not_new_n640__10;
  wire not_new_n3344_;
  wire not_new_n1045__8235430;
  wire not_new_n8609_;
  wire not_new_n1069__3430;
  wire new_n3167_;
  wire new_n3245_;
  wire not_new_n1001__0;
  wire new_n5806_;
  wire new_n9153_;
  wire new_n7832_;
  wire not_new_n588__168070;
  wire not_new_n7584_;
  wire not_new_n7065_;
  wire not_pi027;
  wire not_new_n6497_;
  wire new_n1952_;
  wire not_new_n602__6782230728490;
  wire not_new_n2281_;
  wire new_n2243_;
  wire not_new_n636__168070;
  wire not_po298_7;
  wire not_new_n5153_;
  wire not_new_n4224_;
  wire not_new_n6591_;
  wire not_new_n4472_;
  wire new_n4538_;
  wire new_n1287_;
  wire not_new_n4246_;
  wire not_pi005;
  wire not_new_n639__403536070;
  wire not_pi030;
  wire not_new_n600__19773267430;
  wire new_n2806_;
  wire new_n6469_;
  wire new_n4631_;
  wire not_new_n1012__6;
  wire not_new_n7685_;
  wire not_new_n6924_;
  wire new_n8043_;
  wire new_n4986_;
  wire not_new_n1016__5;
  wire new_n3277_;
  wire not_new_n7793_;
  wire not_new_n1043__6782230728490;
  wire new_n8263_;
  wire not_new_n9439_;
  wire not_new_n1557_;
  wire not_new_n9710_;
  wire new_n4529_;
  wire new_n2435_;
  wire new_n3758_;
  wire not_new_n4952_;
  wire not_new_n594__3430;
  wire not_new_n7752__0;
  wire not_pi248_1;
  wire new_n1884_;
  wire not_new_n7690_;
  wire or_not_new_n1251__not_new_n1249_;
  wire not_pi064_2;
  wire new_n9940_;
  wire not_new_n5538_;
  wire new_n3403_;
  wire not_new_n5521_;
  wire new_n2550_;
  wire new_n9009_;
  wire not_new_n1039__3;
  wire not_new_n7415__2;
  wire not_new_n9484__0;
  wire new_n8537_;
  wire not_new_n3384_;
  wire not_new_n7277__0;
  wire new_n9036_;
  wire not_new_n5321_;
  wire not_new_n8649_;
  wire new_n7455_;
  wire new_n3877_;
  wire not_new_n7348_;
  wire not_pi084;
  wire not_new_n1061__2;
  wire not_new_n1583__968890104070;
  wire new_n3856_;
  wire new_n8279_;
  wire new_n4595_;
  wire new_n4507_;
  wire new_n10124_;
  wire not_new_n2058_;
  wire not_new_n1663_;
  wire not_new_n8138__0;
  wire not_new_n1576__19773267430;
  wire not_new_n622__19773267430;
  wire or_not_new_n1158__1_not_new_n8715__0;
  wire new_n5904_;
  wire not_new_n7557_;
  wire not_new_n1583__2824752490;
  wire new_n4978_;
  wire not_new_n581__57648010;
  wire new_n6696_;
  wire new_n9430_;
  wire not_new_n1071__968890104070;
  wire new_n9967_;
  wire not_new_n7751_;
  wire new_n4339_;
  wire not_new_n1612__1176490;
  wire not_new_n10322_;
  wire not_new_n1031__4;
  wire not_new_n8439_;
  wire not_new_n1051__9;
  wire new_n6884_;
  wire not_new_n1612__490;
  wire new_n3692_;
  wire not_new_n606__490;
  wire not_new_n1631__2824752490;
  wire not_new_n628__6782230728490;
  wire new_n7123_;
  wire new_n6540_;
  wire new_n6572_;
  wire not_new_n3311__70;
  wire not_new_n1179__0;
  wire not_new_n8090_;
  wire not_new_n5314_;
  wire or_not_new_n6541__0_not_new_n1596__1176490;
  wire new_n9884_;
  wire new_n4985_;
  wire not_new_n3881_;
  wire not_new_n5606_;
  wire new_n7957_;
  wire not_pi164_1;
  wire not_new_n5753__1;
  wire not_new_n581__1577753820348458066150427430;
  wire new_n6678_;
  wire not_new_n5973_;
  wire not_new_n587__47475615099430;
  wire new_n8494_;
  wire not_pi169_0;
  wire not_new_n4751_;
  wire new_n2948_;
  wire not_new_n6081_;
  wire or_not_new_n6352__not_new_n6242__5;
  wire new_n8894_;
  wire new_n3011_;
  wire not_new_n6662_;
  wire not_new_n579_;
  wire new_n10081_;
  wire new_n5977_;
  wire not_new_n8061_;
  wire not_new_n639__4;
  wire new_n5674_;
  wire not_new_n633__8;
  wire new_n1508_;
  wire not_new_n1336_;
  wire not_new_n9701_;
  wire new_n2514_;
  wire new_n7339_;
  wire not_new_n7442__0;
  wire new_n616_;
  wire new_n8620_;
  wire not_new_n8190_;
  wire not_new_n6635__1;
  wire new_n8083_;
  wire new_n5604_;
  wire not_new_n1244_;
  wire new_n7410_;
  wire new_n1614_;
  wire new_n8593_;
  wire new_n9118_;
  wire not_new_n9965_;
  wire not_new_n6506_;
  wire new_n10094_;
  wire new_n4329_;
  wire not_new_n6654_;
  wire not_new_n1631__403536070;
  wire new_n2917_;
  wire not_new_n7704_;
  wire not_new_n947_;
  wire new_n5645_;
  wire not_new_n7076_;
  wire new_n3777_;
  wire new_n9643_;
  wire new_n3950_;
  wire not_new_n5432_;
  wire not_new_n1166_;
  wire not_new_n7772__0;
  wire not_new_n775__9;
  wire not_new_n4671_;
  wire not_new_n629__57648010;
  wire new_n3440_;
  wire new_n9703_;
  wire not_new_n1598__490;
  wire not_new_n644__39098210485829880490;
  wire new_n9818_;
  wire and_new_n6433__new_n6432_;
  wire not_new_n3549_;
  wire not_new_n3843_;
  wire new_n9990_;
  wire new_n2414_;
  wire new_n1957_;
  wire not_new_n1603__70;
  wire not_new_n6223_;
  wire new_n1168_;
  wire not_new_n1885_;
  wire not_new_n4259_;
  wire new_n7685_;
  wire new_n5321_;
  wire not_new_n7424_;
  wire not_new_n1041__968890104070;
  wire or_not_new_n8169__1_not_new_n8508_;
  wire new_n4644_;
  wire not_new_n7141__0;
  wire not_new_n5524_;
  wire not_new_n9781_;
  wire new_n9112_;
  wire not_new_n1613__8235430;
  wire new_n1491_;
  wire new_n4289_;
  wire not_new_n7014__0;
  wire new_n3607_;
  wire not_new_n1583__6782230728490;
  wire not_new_n3898_;
  wire key_gate_117;
  wire new_n2880_;
  wire not_new_n6596_;
  wire not_new_n4134_;
  wire new_n4173_;
  wire and_new_n6373__new_n6386_;
  wire new_n5032_;
  wire new_n4792_;
  wire not_new_n3372__968890104070;
  wire new_n5386_;
  wire new_n3840_;
  wire not_new_n1311_;
  wire not_po296_10;
  wire not_new_n1045__1176490;
  wire not_new_n4100_;
  wire not_new_n5740__0;
  wire new_n1939_;
  wire new_n3725_;
  wire new_n1188_;
  wire not_new_n5069_;
  wire not_new_n634__2;
  wire not_new_n2868_;
  wire new_n8111_;
  wire new_n10241_;
  wire not_new_n9873__0;
  wire not_new_n4573_;
  wire new_n1332_;
  wire new_n3396_;
  wire not_new_n6153_;
  wire not_new_n8972_;
  wire new_n6438_;
  wire not_new_n1000_;
  wire not_new_n621__113988951853731430;
  wire new_n5466_;
  wire new_n8856_;
  wire not_new_n5763_;
  wire not_new_n9949_;
  wire not_new_n7816_;
  wire not_new_n10339_;
  wire new_n4312_;
  wire not_new_n581__26517308458596534717790233816010;
  wire new_n6114_;
  wire not_new_n1537__8235430;
  wire not_new_n7770_;
  wire new_n9341_;
  wire not_new_n6443__2326305139872070;
  wire not_new_n1976_;
  wire not_new_n7368_;
  wire new_n4736_;
  wire not_new_n1067__57648010;
  wire not_new_n3310__4;
  wire new_n5117_;
  wire not_new_n8524_;
  wire new_n10102_;
  wire new_n8172_;
  wire not_pi165;
  wire new_n8526_;
  wire not_new_n1597__5;
  wire not_new_n1027__490;
  wire new_n2168_;
  wire not_new_n8964_;
  wire not_new_n10023_;
  wire new_n5335_;
  wire not_new_n9109__0;
  wire not_new_n2280_;
  wire not_new_n8544_;
  wire new_n9900_;
  wire new_n6102_;
  wire new_n3177_;
  wire not_new_n9382_;
  wire not_new_n3492_;
  wire not_new_n3580_;
  wire new_n3044_;
  wire not_new_n1613__70;
  wire new_n1724_;
  wire not_new_n4430_;
  wire new_n5020_;
  wire not_new_n628__47475615099430;
  wire new_n721_;
  wire new_n8171_;
  wire new_n4301_;
  wire or_or_or_not_new_n2794__not_new_n2797__not_new_n2796__not_new_n2798_;
  wire not_new_n631__5;
  wire not_new_n636__1176490;
  wire new_n7850_;
  wire new_n5767_;
  wire new_n2677_;
  wire new_n6857_;
  wire not_new_n1039__403536070;
  wire new_n8809_;
  wire new_n4825_;
  wire not_new_n646__8235430;
  wire not_new_n621_;
  wire new_n1785_;
  wire or_not_new_n9176__not_new_n9177_;
  wire not_new_n4521_;
  wire not_new_n3728_;
  wire new_n3497_;
  wire not_new_n5468_;
  wire not_new_n618__403536070;
  wire not_new_n581__10;
  wire and_new_n3052__new_n998_;
  wire new_n951_;
  wire not_new_n4477_;
  wire not_new_n6058_;
  wire or_or_not_new_n6897__not_new_n6798__not_new_n6826_;
  wire not_pi002;
  wire new_n2983_;
  wire new_n8447_;
  wire not_new_n593__490;
  wire not_new_n642__138412872010;
  wire new_n3703_;
  wire new_n8725_;
  wire not_new_n4804_;
  wire not_new_n626__490;
  wire not_new_n2053_;
  wire new_n10268_;
  wire po161;
  wire not_pi061;
  wire not_new_n7623__0;
  wire new_n9578_;
  wire new_n7675_;
  wire not_new_n1010__4;
  wire not_new_n1533_;
  wire new_n4174_;
  wire new_n967_;
  wire and_new_n3070__new_n998_;
  wire not_new_n1020__5;
  wire new_n4619_;
  wire new_n8995_;
  wire new_n6512_;
  wire not_new_n991__0;
  wire not_new_n8602_;
  wire new_n6324_;
  wire new_n10317_;
  wire not_new_n601__5;
  wire new_n2705_;
  wire new_n2304_;
  wire not_new_n3824_;
  wire not_new_n627__16284135979104490;
  wire not_new_n8845__2;
  wire new_n1664_;
  wire not_new_n7601_;
  wire not_new_n4772__0;
  wire not_new_n598__3430;
  wire not_new_n587__797922662976120010;
  wire not_new_n7445_;
  wire not_new_n8504_;
  wire new_n5381_;
  wire not_new_n7670__0;
  wire not_new_n4748__0;
  wire po191;
  wire new_n1637_;
  wire not_new_n10146_;
  wire new_n9126_;
  wire not_new_n3375__1;
  wire new_n7188_;
  wire not_new_n6717_;
  wire new_n8363_;
  wire not_new_n5433__0;
  wire not_new_n5470__0;
  wire new_n8135_;
  wire not_new_n609__9;
  wire not_new_n589__185621159210175743024531636712070;
  wire not_new_n5572_;
  wire not_new_n4107_;
  wire new_n4837_;
  wire new_n2197_;
  wire not_new_n1534__6;
  wire po242;
  wire not_new_n6868_;
  wire new_n9006_;
  wire not_new_n4948_;
  wire new_n2829_;
  wire not_new_n1963_;
  wire not_new_n7006_;
  wire or_not_new_n1406__not_new_n1407_;
  wire not_new_n3569_;
  wire new_n1829_;
  wire not_new_n768_;
  wire new_n3652_;
  wire new_n1242_;
  wire new_n2778_;
  wire not_new_n3923_;
  wire not_new_n9967__0;
  wire not_new_n8285__0;
  wire po289;
  wire new_n8042_;
  wire not_pi179_4;
  wire not_new_n3315__2824752490;
  wire new_n9420_;
  wire not_new_n6538__1;
  wire new_n3956_;
  wire new_n8025_;
  wire new_n3261_;
  wire not_new_n9684_;
  wire new_n6715_;
  wire new_n10115_;
  wire not_new_n9819_;
  wire not_new_n6502__0;
  wire new_n2636_;
  wire not_po296_367033682172941254412302110320336601888010;
  wire new_n9552_;
  wire not_new_n595__57648010;
  wire new_n4596_;
  wire new_n2048_;
  wire not_new_n4792__0;
  wire not_new_n638__5585458640832840070;
  wire not_pi009_0;
  wire new_n1807_;
  wire new_n7726_;
  wire not_new_n5135_;
  wire not_new_n626__1;
  wire not_new_n1159__0;
  wire new_n7444_;
  wire not_new_n9159_;
  wire not_new_n6413_;
  wire new_n4688_;
  wire not_new_n5147_;
  wire not_new_n4797_;
  wire not_new_n647__138412872010;
  wire key_gate_110;
  wire new_n4928_;
  wire not_pi056_2;
  wire new_n6097_;
  wire not_pi033_5;
  wire not_new_n3115_;
  wire not_new_n3274_;
  wire not_new_n1061__1;
  wire new_n6751_;
  wire new_n4696_;
  wire not_pi259;
  wire new_n7130_;
  wire not_new_n644__4;
  wire new_n5459_;
  wire new_n1244_;
  wire not_new_n1904_;
  wire new_n1632_;
  wire new_n7490_;
  wire new_n3476_;
  wire not_pi257_2;
  wire new_n10101_;
  wire new_n6012_;
  wire not_new_n9741_;
  wire not_new_n9576_;
  wire new_n2529_;
  wire new_n10085_;
  wire new_n1304_;
  wire not_new_n7197_;
  wire new_n7491_;
  wire new_n9715_;
  wire new_n9696_;
  wire not_new_n1212_;
  wire new_n7586_;
  wire new_n9721_;
  wire new_n2993_;
  wire or_not_new_n2964__not_new_n2967_;
  wire not_new_n584__0;
  wire not_new_n1168__0;
  wire not_new_n2959_;
  wire not_new_n589__332329305696010;
  wire new_n8584_;
  wire not_new_n4015_;
  wire not_new_n687_;
  wire not_new_n586__968890104070;
  wire not_new_n10042__0;
  wire new_n2278_;
  wire not_pi055_1;
  wire not_new_n4999__0;
  wire new_n6351_;
  wire not_new_n599__138412872010;
  wire not_new_n3690_;
  wire new_n3149_;
  wire new_n6034_;
  wire new_n9713_;
  wire not_new_n1583__8;
  wire new_n3039_;
  wire not_new_n3683_;
  wire not_new_n1037__70;
  wire not_new_n1440_;
  wire or_or_not_new_n2189__not_new_n2186__not_new_n2187_;
  wire not_new_n9108_;
  wire new_n7280_;
  wire not_new_n8800_;
  wire not_new_n5084__2;
  wire not_new_n6504__0;
  wire new_n9528_;
  wire new_n6322_;
  wire not_new_n8065_;
  wire not_new_n646__2326305139872070;
  wire not_new_n7396_;
  wire not_new_n1041__5;
  wire new_n636_;
  wire not_new_n8471_;
  wire not_new_n1213_;
  wire not_new_n1065__39098210485829880490;
  wire not_new_n3235_;
  wire not_new_n642__5;
  wire and_new_n1217__new_n1218_;
  wire new_n6065_;
  wire not_new_n4807__0;
  wire and_new_n2992__new_n998_;
  wire new_n9435_;
  wire not_new_n2611_;
  wire new_n7702_;
  wire not_new_n8191_;
  wire not_new_n3785_;
  wire not_new_n4424_;
  wire not_new_n4596_;
  wire new_n6936_;
  wire not_new_n2091_;
  wire not_new_n1041__6;
  wire new_n6389_;
  wire not_new_n5341_;
  wire new_n8896_;
  wire not_new_n1597__968890104070;
  wire not_new_n1035__24010;
  wire new_n10321_;
  wire new_n9109_;
  wire not_new_n7303_;
  wire not_new_n1049__0;
  wire not_new_n10218_;
  wire new_n6365_;
  wire not_new_n1613__113988951853731430;
  wire new_n4767_;
  wire not_new_n7642__0;
  wire not_new_n4715_;
  wire new_n2270_;
  wire new_n1179_;
  wire not_pi059_2;
  wire new_n7554_;
  wire not_new_n9889_;
  wire not_new_n1413_;
  wire not_new_n3148_;
  wire and_not_pi040_3_not_pi041_2;
  wire new_n6769_;
  wire not_new_n607__4;
  wire not_new_n8294_;
  wire not_new_n1588__6782230728490;
  wire new_n4313_;
  wire not_new_n639__39098210485829880490;
  wire new_n3727_;
  wire new_n3086_;
  wire new_n9903_;
  wire new_n1487_;
  wire not_new_n7146_;
  wire new_n8230_;
  wire not_new_n950_;
  wire not_new_n610__24010;
  wire not_new_n626__47475615099430;
  wire not_new_n3368_;
  wire not_new_n633__968890104070;
  wire not_new_n9636_;
  wire new_n6827_;
  wire not_new_n5116_;
  wire not_new_n647__332329305696010;
  wire not_new_n8992_;
  wire not_new_n4451_;
  wire not_new_n8225_;
  wire not_new_n7759_;
  wire not_new_n1830_;
  wire new_n2104_;
  wire or_not_new_n10219__not_new_n10220_;
  wire new_n6850_;
  wire not_new_n1031__70;
  wire not_new_n9934_;
  wire not_new_n1591__7;
  wire not_new_n6457_;
  wire not_new_n2653_;
  wire or_not_new_n2980__not_new_n2979_;
  wire not_new_n599__16284135979104490;
  wire new_n5337_;
  wire new_n4731_;
  wire not_new_n1603__403536070;
  wire new_n7053_;
  wire not_new_n1604__6782230728490;
  wire new_n4780_;
  wire new_n8106_;
  wire new_n8911_;
  wire not_new_n7124_;
  wire not_new_n648__7;
  wire not_new_n1027__39098210485829880490;
  wire not_new_n5183_;
  wire not_new_n628__8;
  wire new_n5273_;
  wire not_new_n5452_;
  wire not_pi176_3;
  wire not_new_n3387_;
  wire new_n7985_;
  wire not_new_n1599__19773267430;
  wire not_new_n3661_;
  wire not_pi154;
  wire new_n5917_;
  wire not_new_n1611__2824752490;
  wire new_n8922_;
  wire not_new_n629__70;
  wire not_new_n2757_;
  wire not_new_n8333_;
  wire not_new_n1377_;
  wire not_new_n6663_;
  wire not_new_n5066__0;
  wire not_new_n7020__0;
  wire new_n4453_;
  wire not_new_n9972__0;
  wire not_new_n7721_;
  wire not_new_n1067__19773267430;
  wire new_n8724_;
  wire new_n4880_;
  wire new_n5508_;
  wire not_new_n1604_;
  wire new_n2647_;
  wire not_new_n9816_;
  wire not_new_n5741__2;
  wire not_new_n7004__0;
  wire not_new_n699_;
  wire not_new_n928__2824752490;
  wire or_not_new_n2747__not_new_n2746_;
  wire not_new_n4983_;
  wire new_n5695_;
  wire new_n1002_;
  wire new_n6711_;
  wire new_n7159_;
  wire new_n9354_;
  wire new_n4291_;
  wire new_n3133_;
  wire not_new_n2586_;
  wire and_and_new_n2707__new_n2708__new_n3822_;
  wire new_n7594_;
  wire not_new_n6075_;
  wire not_new_n1631_;
  wire not_new_n6068__0;
  wire new_n3446_;
  wire new_n6980_;
  wire not_new_n4124__2;
  wire new_n1782_;
  wire new_n6630_;
  wire new_n6363_;
  wire not_new_n1175_;
  wire not_new_n3488_;
  wire not_new_n7907_;
  wire new_n3767_;
  wire not_new_n3105_;
  wire not_new_n3928__0;
  wire not_pi059_1;
  wire new_n8543_;
  wire not_new_n7620__1;
  wire not_new_n9225_;
  wire not_new_n8119_;
  wire not_new_n3816_;
  wire new_n1378_;
  wire not_new_n2563_;
  wire not_new_n5597__1;
  wire not_new_n591__7;
  wire new_n3111_;
  wire not_new_n1055__490;
  wire po237;
  wire not_new_n625__657123623635342801395430;
  wire new_n5190_;
  wire new_n9403_;
  wire new_n6115_;
  wire new_n10122_;
  wire new_n8825_;
  wire not_new_n7594_;
  wire new_n5439_;
  wire new_n3796_;
  wire new_n954_;
  wire not_pi221;
  wire not_new_n8048_;
  wire not_new_n1584__2824752490;
  wire new_n5245_;
  wire not_new_n992_;
  wire not_new_n5706_;
  wire new_n3117_;
  wire new_n9910_;
  wire not_new_n7912_;
  wire not_new_n5093_;
  wire not_po296_9095436801298611408202050198891430;
  wire not_new_n4946__0;
  wire new_n5940_;
  wire new_n8805_;
  wire new_n9969_;
  wire not_new_n2920_;
  wire not_new_n8650_;
  wire or_not_new_n7906__not_new_n7780_;
  wire po188;
  wire or_not_new_n8448__not_new_n8419_;
  wire new_n7093_;
  wire new_n3343_;
  wire new_n7090_;
  wire not_new_n598__113988951853731430;
  wire new_n1561_;
  wire not_new_n6245_;
  wire not_new_n1069__10;
  wire new_n2663_;
  wire new_n604_;
  wire new_n1642_;
  wire not_new_n5412_;
  wire and_new_n2276__new_n2279_;
  wire new_n7543_;
  wire not_new_n8854_;
  wire not_new_n7162_;
  wire new_n6045_;
  wire new_n4758_;
  wire new_n10326_;
  wire new_n5255_;
  wire new_n5028_;
  wire new_n1681_;
  wire not_new_n8368_;
  wire not_new_n4089_;
  wire new_n7078_;
  wire not_new_n8082_;
  wire not_new_n4926_;
  wire new_n6687_;
  wire not_new_n7432_;
  wire not_new_n5800_;
  wire not_new_n5975_;
  wire new_n6468_;
  wire new_n8900_;
  wire not_new_n7244_;
  wire not_new_n8351_;
  wire not_new_n4232_;
  wire new_n1475_;
  wire not_new_n4802__0;
  wire new_n2294_;
  wire new_n7757_;
  wire not_new_n6671_;
  wire not_pi136_3;
  wire not_new_n9645_;
  wire new_n2469_;
  wire new_n1249_;
  wire not_new_n9854__2;
  wire not_new_n8201_;
  wire not_new_n8426_;
  wire not_new_n3185__7;
  wire new_n1973_;
  wire not_new_n1041__3430;
  wire new_n3040_;
  wire new_n9920_;
  wire new_n9214_;
  wire or_or_not_new_n2946__not_new_n2949__not_new_n2948_;
  wire not_new_n644__332329305696010;
  wire new_n5825_;
  wire new_n8548_;
  wire not_new_n9725_;
  wire not_new_n631__2824752490;
  wire not_new_n1441_;
  wire not_new_n1015__2;
  wire not_new_n5380_;
  wire new_n4473_;
  wire not_new_n640__113988951853731430;
  wire not_pi261_1;
  wire not_new_n3919__0;
  wire not_new_n4663_;
  wire new_n3211_;
  wire po079;
  wire not_new_n9537_;
  wire new_n8731_;
  wire and_new_n2200__new_n2203_;
  wire new_n5559_;
  wire not_new_n7049_;
  wire not_new_n2074_;
  wire not_new_n2553_;
  wire new_n8309_;
  wire not_new_n647__70;
  wire new_n8355_;
  wire or_not_new_n6373__not_new_n6413_;
  wire not_new_n8883_;
  wire not_new_n4934_;
  wire not_new_n7607_;
  wire and_new_n1858__new_n1861_;
  wire new_n3447_;
  wire new_n8507_;
  wire not_new_n8271_;
  wire new_n4646_;
  wire not_pi224;
  wire not_new_n7329_;
  wire not_new_n1053__47475615099430;
  wire not_new_n8139__0;
  wire not_new_n1596__16284135979104490;
  wire not_new_n4031_;
  wire not_new_n628__657123623635342801395430;
  wire not_new_n1602__2;
  wire new_n4620_;
  wire not_new_n3372__5;
  wire not_new_n3162_;
  wire not_new_n4619_;
  wire not_new_n1247_;
  wire not_pi095;
  wire new_n6374_;
  wire not_new_n1437_;
  wire or_not_new_n2497__not_new_n1568_;
  wire not_new_n4123_;
  wire new_n3640_;
  wire not_new_n1248_;
  wire not_new_n7644__0;
  wire new_n1391_;
  wire and_new_n1801__new_n1804_;
  wire not_new_n1576__9;
  wire new_n7502_;
  wire not_new_n6373__4;
  wire not_new_n1037__6782230728490;
  wire new_n3007_;
  wire new_n4571_;
  wire new_n6178_;
  wire not_new_n2676_;
  wire new_n8981_;
  wire not_new_n7470_;
  wire not_new_n5460_;
  wire not_new_n3667_;
  wire not_new_n585__490;
  wire not_new_n4168_;
  wire not_new_n1601__24010;
  wire not_new_n1538__3;
  wire or_or_not_new_n1331__not_new_n1329__not_new_n2268_;
  wire not_new_n9318_;
  wire not_new_n8177_;
  wire not_new_n600__1;
  wire new_n8605_;
  wire not_new_n643__70;
  wire not_new_n5425_;
  wire not_new_n7007__0;
  wire not_new_n6918_;
  wire not_new_n2887_;
  wire new_n8473_;
  wire not_new_n1611__0;
  wire not_new_n9540_;
  wire new_n8895_;
  wire not_new_n7367_;
  wire new_n4730_;
  wire not_new_n1531_;
  wire or_not_new_n4835__not_new_n4777_;
  wire not_new_n4780__0;
  wire not_new_n2605_;
  wire not_new_n7906_;
  wire new_n3890_;
  wire new_n5742_;
  wire not_new_n3976__0;
  wire not_new_n6577_;
  wire new_n5975_;
  wire not_new_n1613__2326305139872070;
  wire new_n2640_;
  wire new_n8052_;
  wire not_new_n9403_;
  wire not_new_n6737__1;
  wire new_n5965_;
  wire new_n2129_;
  wire not_new_n7651__2;
  wire not_new_n10041__0;
  wire new_n2076_;
  wire new_n10248_;
  wire new_n6256_;
  wire not_new_n630__8235430;
  wire new_n3374_;
  wire new_n6159_;
  wire new_n6986_;
  wire not_new_n4930_;
  wire not_new_n1598__3;
  wire new_n8757_;
  wire new_n5554_;
  wire not_new_n594__1;
  wire new_n4049_;
  wire not_new_n4802_;
  wire not_new_n5210_;
  wire new_n4201_;
  wire new_n2364_;
  wire not_new_n1921_;
  wire not_new_n618__19773267430;
  wire new_n5392_;
  wire new_n4078_;
  wire new_n3547_;
  wire new_n2366_;
  wire not_new_n3216_;
  wire new_n1686_;
  wire not_new_n581__0;
  wire not_pi268;
  wire new_n4034_;
  wire not_new_n3035_;
  wire not_new_n9351_;
  wire not_new_n8897__0;
  wire not_new_n5196_;
  wire not_new_n640__5;
  wire new_n5168_;
  wire po152;
  wire new_n6010_;
  wire new_n6304_;
  wire po124;
  wire not_new_n1041__0;
  wire not_new_n607__0;
  wire not_new_n1416_;
  wire not_new_n4115_;
  wire not_new_n9523_;
  wire new_n5692_;
  wire not_new_n1055__57648010;
  wire not_new_n8064_;
  wire not_new_n5199_;
  wire new_n1880_;
  wire not_new_n6452_;
  wire not_new_n5889_;
  wire not_new_n3677_;
  wire po108;
  wire not_new_n6146_;
  wire new_n9842_;
  wire or_not_new_n9612__not_new_n9611_;
  wire not_new_n9987_;
  wire new_n3302_;
  wire not_pi109;
  wire new_n5446_;
  wire not_new_n999__1;
  wire not_new_n1065_;
  wire not_pi250_2;
  wire not_new_n5108_;
  wire not_new_n1598__7;
  wire new_n4598_;
  wire or_not_new_n2695__not_new_n2694_;
  wire new_n3988_;
  wire not_new_n7996_;
  wire not_new_n7890_;
  wire new_n2287_;
  wire or_not_new_n3091__not_new_n3090_;
  wire po218;
  wire not_new_n9894_;
  wire new_n2036_;
  wire not_new_n6544_;
  wire new_n8684_;
  wire new_n9048_;
  wire not_pi031_0;
  wire not_new_n1764_;
  wire new_n2318_;
  wire not_new_n4484_;
  wire new_n4720_;
  wire not_new_n8963__1;
  wire new_n4771_;
  wire not_new_n645__19773267430;
  wire not_new_n2931_;
  wire not_new_n5527_;
  wire new_n2623_;
  wire not_new_n6051_;
  wire not_new_n3374_;
  wire new_n7753_;
  wire new_n1864_;
  wire not_new_n622__2326305139872070;
  wire new_n8749_;
  wire new_n6338_;
  wire or_not_new_n3110__not_new_n3109_;
  wire not_new_n1187_;
  wire not_pi215;
  wire not_pi016;
  wire new_n923_;
  wire not_new_n758_;
  wire key_gate_76;
  wire new_n3156_;
  wire new_n8075_;
  wire new_n2295_;
  wire not_new_n9635_;
  wire not_new_n1445_;
  wire new_n9674_;
  wire new_n2615_;
  wire new_n6613_;
  wire not_new_n1605__1;
  wire not_new_n4683_;
  wire new_n1497_;
  wire po142;
  wire and_new_n1238__new_n1837_;
  wire new_n5816_;
  wire new_n6492_;
  wire new_n3841_;
  wire not_new_n4431__0;
  wire new_n8549_;
  wire not_new_n9550_;
  wire not_new_n611__5;
  wire not_new_n602__19773267430;
  wire new_n5924_;
  wire not_pi123;
  wire not_new_n3282_;
  wire new_n6189_;
  wire not_new_n7328_;
  wire and_new_n2105__new_n2108_;
  wire not_new_n622__168070;
  wire not_new_n1601__3;
  wire not_new_n8596__3;
  wire new_n1017_;
  wire new_n7864_;
  wire new_n8212_;
  wire not_new_n4975__0;
  wire not_new_n6541_;
  wire not_new_n1819_;
  wire new_n7403_;
  wire po178;
  wire not_new_n1045__47475615099430;
  wire not_new_n1611__24010;
  wire new_n9117_;
  wire not_new_n1403_;
  wire new_n9350_;
  wire not_new_n5039_;
  wire new_n8372_;
  wire new_n4158_;
  wire new_n3971_;
  wire not_new_n8278__0;
  wire not_new_n5482__0;
  wire not_pi171_1;
  wire new_n2745_;
  wire not_new_n1919__0;
  wire not_new_n5427__0;
  wire not_pi169_3;
  wire new_n9363_;
  wire not_new_n6537_;
  wire new_n3768_;
  wire not_new_n7443_;
  wire not_new_n1069__4;
  wire not_new_n4776__0;
  wire not_new_n9362_;
  wire new_n5403_;
  wire not_new_n1576__8235430;
  wire new_n6792_;
  wire new_n1578_;
  wire new_n6190_;
  wire not_po296_21838143759917965991093122527538323430;
  wire new_n5410_;
  wire not_new_n6634_;
  wire new_n1201_;
  wire and_new_n1242__new_n1856_;
  wire not_new_n5924_;
  wire not_new_n621__332329305696010;
  wire not_new_n3510_;
  wire not_new_n1055_;
  wire not_new_n5111__0;
  wire not_new_n581__1176490;
  wire not_new_n8446_;
  wire new_n8777_;
  wire not_new_n5841_;
  wire not_new_n5479_;
  wire new_n9648_;
  wire not_new_n3331_;
  wire new_n9502_;
  wire not_new_n2946_;
  wire not_new_n5463_;
  wire new_n8618_;
  wire not_new_n6761__0;
  wire new_n6791_;
  wire new_n8102_;
  wire not_new_n4188_;
  wire not_new_n7110_;
  wire and_new_n933__new_n935_;
  wire not_new_n617__3430;
  wire not_new_n9616_;
  wire new_n8865_;
  wire not_new_n3315__2326305139872070;
  wire new_n6437_;
  wire not_new_n7703_;
  wire new_n2472_;
  wire new_n7077_;
  wire not_new_n4898__1;
  wire not_new_n4468__0;
  wire not_new_n1253_;
  wire not_new_n4843__1;
  wire not_new_n1205_;
  wire new_n10150_;
  wire new_n1256_;
  wire or_not_new_n2727__not_new_n2730_;
  wire not_new_n8801_;
  wire not_new_n7304_;
  wire new_n6135_;
  wire not_new_n10127_;
  wire new_n5871_;
  wire not_pi162_0;
  wire not_po296_332329305696010;
  wire new_n9609_;
  wire new_n10233_;
  wire new_n1739_;
  wire new_n4093_;
  wire not_pi167_1;
  wire new_n4335_;
  wire new_n7604_;
  wire new_n7647_;
  wire new_n8615_;
  wire not_new_n2885_;
  wire not_new_n5354_;
  wire not_new_n7628__0;
  wire not_new_n4739_;
  wire new_n1953_;
  wire or_not_new_n2776__not_new_n2779_;
  wire new_n4754_;
  wire new_n4934_;
  wire not_new_n1041__1176490;
  wire not_new_n7261_;
  wire new_n6768_;
  wire new_n5976_;
  wire not_new_n10006_;
  wire new_n1310_;
  wire not_new_n2033__0;
  wire not_new_n4582_;
  wire not_new_n9852_;
  wire not_new_n6595_;
  wire new_n4802_;
  wire not_new_n8127_;
  wire not_new_n588__0;
  wire not_new_n740__1;
  wire not_new_n4393_;
  wire key_gate_105;
  wire key_gate_20;
  wire and_and_not_pi060_1_not_pi059_1_not_pi058_1;
  wire not_new_n589__445676403263631959001900459745680070;
  wire not_new_n589__490;
  wire new_n4503_;
  wire not_new_n7818_;
  wire not_new_n9944_;
  wire not_new_n3867_;
  wire new_n7037_;
  wire not_new_n3190_;
  wire not_new_n6691__0;
  wire not_new_n5381_;
  wire or_or_not_new_n6239__not_new_n6350__not_new_n6232__3;
  wire new_n8918_;
  wire new_n9058_;
  wire not_new_n1043__19773267430;
  wire not_new_n3577_;
  wire or_or_not_new_n2865__not_new_n2868__not_new_n2867_;
  wire not_new_n3934__0;
  wire not_new_n7420_;
  wire not_new_n8549_;
  wire po089;
  wire not_new_n6160_;
  wire not_new_n3372__7;
  wire not_new_n9215_;
  wire not_new_n600__168070;
  wire not_new_n9788_;
  wire not_new_n1027__1;
  wire not_new_n1600__8;
  wire not_new_n9926_;
  wire not_new_n4829__1;
  wire new_n1443_;
  wire new_n3124_;
  wire new_n6797_;
  wire not_new_n8579_;
  wire not_new_n596__5;
  wire new_n8444_;
  wire new_n6348_;
  wire new_n1212_;
  wire not_new_n587__490;
  wire not_new_n1603__1;
  wire new_n6001_;
  wire new_n6962_;
  wire not_new_n642__24010;
  wire new_n3413_;
  wire new_n3864_;
  wire not_new_n621__797922662976120010;
  wire new_n3525_;
  wire not_new_n1055__19773267430;
  wire not_new_n7031__1;
  wire and_new_n1298__new_n2122_;
  wire not_new_n7267_;
  wire not_new_n4432_;
  wire not_new_n6414_;
  wire new_n8423_;
  wire not_new_n626__4;
  wire new_n4354_;
  wire not_new_n3315__138412872010;
  wire not_new_n8936_;
  wire not_new_n1611_;
  wire new_n9974_;
  wire new_n2818_;
  wire or_not_new_n1024__2_not_new_n1028__3;
  wire new_n7882_;
  wire not_new_n9403__0;
  wire new_n4843_;
  wire not_new_n749_;
  wire new_n9345_;
  wire new_n4694_;
  wire not_new_n7872_;
  wire new_n7054_;
  wire not_new_n6839_;
  wire new_n5896_;
  wire new_n8462_;
  wire not_new_n9800_;
  wire not_new_n6181_;
  wire new_n3799_;
  wire new_n10289_;
  wire not_new_n5820_;
  wire not_new_n6982__2;
  wire new_n10227_;
  wire not_new_n4203_;
  wire new_n6955_;
  wire not_new_n6020_;
  wire not_new_n1027__403536070;
  wire not_new_n2982_;
  wire not_new_n2593_;
  wire not_new_n9198_;
  wire not_new_n10200_;
  wire not_new_n2858_;
  wire not_new_n6588_;
  wire not_new_n7234_;
  wire not_new_n623__4;
  wire not_new_n1009__2;
  wire not_new_n619__490;
  wire not_new_n6373__2;
  wire new_n6050_;
  wire not_new_n586__24010;
  wire not_po296_3430;
  wire new_n4765_;
  wire not_new_n6974__968890104070;
  wire new_n1285_;
  wire not_new_n605__168070;
  wire not_new_n617__93874803376477543056490;
  wire po193;
  wire not_new_n8281_;
  wire not_new_n591__9;
  wire not_new_n3706_;
  wire not_new_n6636__0;
  wire new_n3026_;
  wire new_n10311_;
  wire not_new_n4620_;
  wire not_new_n1005_;
  wire new_n2959_;
  wire new_n4202_;
  wire not_new_n1520_;
  wire new_n5048_;
  wire new_n9705_;
  wire new_n2727_;
  wire not_new_n9875_;
  wire not_new_n10193_;
  wire new_n7245_;
  wire new_n3641_;
  wire not_new_n1589__8;
  wire not_new_n645__4;
  wire new_n2298_;
  wire not_new_n9685_;
  wire not_new_n619__24010;
  wire new_n5007_;
  wire new_n5514_;
  wire new_n8227_;
  wire not_new_n6508__0;
  wire new_n9457_;
  wire new_n5324_;
  wire new_n1602_;
  wire not_new_n647__1176490;
  wire not_new_n6150_;
  wire new_n4946_;
  wire not_new_n3535_;
  wire not_new_n1581__403536070;
  wire new_n5085_;
  wire not_pi035_1;
  wire new_n7777_;
  wire new_n9810_;
  wire new_n9362_;
  wire new_n3222_;
  wire not_new_n3860_;
  wire not_new_n2801_;
  wire not_new_n4416__0;
  wire not_new_n1596__57648010;
  wire not_new_n634__5;
  wire not_new_n4092_;
  wire not_new_n8507_;
  wire new_n9921_;
  wire not_new_n8455_;
  wire not_pi160_0;
  wire new_n9442_;
  wire not_new_n4528_;
  wire not_new_n618__16284135979104490;
  wire not_new_n10062_;
  wire new_n6695_;
  wire not_new_n6035_;
  wire not_new_n6946_;
  wire not_new_n5774__0;
  wire not_new_n3955_;
  wire new_n8535_;
  wire key_gate_18;
  wire new_n3585_;
  wire not_new_n635__4;
  wire new_n2525_;
  wire not_new_n742__1;
  wire not_new_n1580__490;
  wire not_new_n6140_;
  wire new_n7008_;
  wire not_new_n647__47475615099430;
  wire not_new_n4753_;
  wire new_n2887_;
  wire not_new_n4716_;
  wire not_pi119_0;
  wire not_new_n7363_;
  wire new_n6258_;
  wire new_n7155_;
  wire new_n6478_;
  wire not_new_n5478_;
  wire not_new_n8047_;
  wire not_new_n9242_;
  wire not_new_n644_;
  wire not_new_n8256__0;
  wire new_n3977_;
  wire not_new_n7718_;
  wire not_pi108;
  wire new_n2543_;
  wire new_n4878_;
  wire new_n9081_;
  wire or_not_new_n1958__not_new_n1959_;
  wire new_n1649_;
  wire not_new_n2171_;
  wire new_n667_;
  wire not_new_n634__2824752490;
  wire not_new_n7435_;
  wire new_n1617_;
  wire new_n1895_;
  wire not_new_n8787_;
  wire new_n4569_;
  wire new_n4537_;
  wire new_n5075_;
  wire or_not_new_n1570__not_new_n2502_;
  wire new_n4865_;
  wire new_n8320_;
  wire not_new_n9600_;
  wire new_n1897_;
  wire not_new_n4135__1;
  wire new_n7758_;
  wire new_n3424_;
  wire not_new_n4771_;
  wire not_new_n9401_;
  wire new_n1363_;
  wire new_n9141_;
  wire new_n7241_;
  wire not_new_n1583__0;
  wire not_new_n3315__5;
  wire not_new_n5186__0;
  wire new_n3050_;
  wire not_new_n7658__0;
  wire not_new_n5686__1;
  wire new_n5533_;
  wire new_n6654_;
  wire new_n10333_;
  wire not_new_n8994_;
  wire new_n2903_;
  wire not_new_n6373__7;
  wire not_new_n4161_;
  wire not_new_n8976_;
  wire new_n7651_;
  wire not_new_n9147_;
  wire not_new_n2911_;
  wire not_new_n3829_;
  wire not_new_n5295_;
  wire not_new_n4988__0;
  wire new_n9076_;
  wire not_new_n4444__0;
  wire new_n6618_;
  wire not_new_n622__5;
  wire not_new_n595__968890104070;
  wire not_new_n638__332329305696010;
  wire not_new_n626__797922662976120010;
  wire new_n4490_;
  wire not_new_n630__10;
  wire not_new_n3184__24010;
  wire new_n6830_;
  wire not_pi142_2;
  wire not_new_n5188_;
  wire not_new_n4757_;
  wire not_new_n620__4;
  wire new_n2189_;
  wire new_n4909_;
  wire new_n1818_;
  wire not_new_n633__113988951853731430;
  wire new_n2134_;
  wire new_n10164_;
  wire or_not_new_n3170__not_new_n3169_;
  wire not_new_n9361__0;
  wire not_new_n9951__0;
  wire not_new_n1728__332329305696010;
  wire not_new_n7069_;
  wire not_new_n8147_;
  wire not_new_n1595_;
  wire not_new_n2624_;
  wire new_n6985_;
  wire new_n5318_;
  wire not_po296_7;
  wire not_new_n7204_;
  wire not_new_n1583__168070;
  wire new_n8970_;
  wire not_new_n7653_;
  wire and_and_new_n2143__new_n2146__new_n2144_;
  wire new_n2265_;
  wire not_new_n8702_;
  wire new_n5397_;
  wire not_new_n775__490;
  wire new_n9625_;
  wire new_n10318_;
  wire new_n2115_;
  wire not_new_n7153__0;
  wire not_new_n3973_;
  wire not_new_n989_;
  wire not_new_n1580__9;
  wire not_new_n593__3430;
  wire not_new_n6373__0;
  wire not_new_n618__273687473400809163430;
  wire new_n5759_;
  wire not_new_n2034_;
  wire new_n7739_;
  wire not_new_n5441_;
  wire new_n2353_;
  wire not_new_n960_;
  wire not_new_n4451__0;
  wire not_new_n3315__10;
  wire new_n3018_;
  wire not_new_n603__2;
  wire not_new_n2306_;
  wire new_n2942_;
  wire new_n3917_;
  wire new_n9896_;
  wire not_new_n5956__0;
  wire not_new_n9716_;
  wire new_n8496_;
  wire new_n4328_;
  wire new_n6254_;
  wire new_n6590_;
  wire not_new_n8506_;
  wire new_n2592_;
  wire not_new_n1588__3;
  wire key_gate_83;
  wire not_new_n2344_;
  wire new_n6528_;
  wire not_new_n8172_;
  wire new_n3364_;
  wire and_new_n1839__new_n1842_;
  wire not_pi037_3;
  wire new_n1544_;
  wire new_n8442_;
  wire new_n7809_;
  wire not_new_n6611_;
  wire not_new_n4818__1;
  wire not_new_n7809__0;
  wire new_n9243_;
  wire not_new_n637__70;
  wire new_n8621_;
  wire not_new_n6499_;
  wire not_pi017_0;
  wire not_new_n1063__47475615099430;
  wire not_new_n617__3;
  wire not_pi255;
  wire not_new_n3450_;
  wire not_new_n642__8235430;
  wire not_new_n2958_;
  wire not_new_n9284_;
  wire not_new_n6475__1;
  wire not_new_n6685_;
  wire not_new_n6474_;
  wire not_new_n7321__0;
  wire new_n706_;
  wire new_n5994_;
  wire not_new_n4718__0;
  wire not_new_n3215_;
  wire new_n8177_;
  wire not_new_n1597__8;
  wire not_new_n6053_;
  wire not_new_n1962_;
  wire not_new_n7528_;
  wire new_n9028_;
  wire not_new_n7692_;
  wire not_new_n7900_;
  wire new_n8469_;
  wire not_new_n5005_;
  wire not_new_n5137_;
  wire new_n2432_;
  wire not_new_n7010_;
  wire not_new_n9226_;
  wire not_pi153_0;
  wire not_new_n646__0;
  wire not_new_n4264_;
  wire not_new_n6546__0;
  wire not_new_n7667_;
  wire new_n9957_;
  wire not_new_n5050_;
  wire new_n8375_;
  wire new_n5478_;
  wire not_new_n632__5585458640832840070;
  wire not_new_n1585__3;
  wire not_new_n9062_;
  wire new_n1215_;
  wire not_new_n2799_;
  wire new_n5681_;
  wire not_new_n7439__2;
  wire new_n7943_;
  wire new_n8828_;
  wire not_new_n1051__2824752490;
  wire not_new_n1611__8235430;
  wire new_n3709_;
  wire not_new_n5674__0;
  wire not_new_n1597__47475615099430;
  wire new_n7303_;
  wire not_new_n4535_;
  wire new_n1936_;
  wire not_new_n635__24010;
  wire new_n7042_;
  wire new_n723_;
  wire new_n4866_;
  wire not_new_n1035__168070;
  wire new_n4984_;
  wire not_new_n8745_;
  wire not_pi053_3;
  wire not_new_n1584__403536070;
  wire not_new_n7269_;
  wire not_pi129_2;
  wire not_new_n9508_;
  wire new_n4225_;
  wire not_new_n10224_;
  wire not_new_n7556_;
  wire new_n6780_;
  wire new_n2031_;
  wire new_n9865_;
  wire not_new_n1583__1176490;
  wire not_new_n5476_;
  wire not_new_n7607__0;
  wire not_new_n4475_;
  wire and_and_and_new_n1463__new_n1465__new_n1464__new_n3720_;
  wire po297;
  wire new_n9657_;
  wire new_n3560_;
  wire new_n9360_;
  wire new_n7863_;
  wire not_new_n747_;
  wire not_new_n603__5;
  wire not_new_n775__968890104070;
  wire not_new_n723__1;
  wire not_new_n2783_;
  wire not_new_n1053__1;
  wire not_new_n7101_;
  wire not_new_n9298_;
  wire not_new_n4569_;
  wire not_new_n643__3430;
  wire not_new_n1149__0;
  wire new_n7007_;
  wire not_new_n8963_;
  wire and_and_new_n1972__new_n1975__new_n1973_;
  wire new_n7195_;
  wire new_n1408_;
  wire new_n10108_;
  wire not_new_n4922_;
  wire not_new_n4132__0;
  wire new_n8261_;
  wire not_new_n1601__2;
  wire not_new_n6159_;
  wire not_new_n621__1176490;
  wire not_new_n9394_;
  wire not_new_n10041_;
  wire new_n8128_;
  wire new_n5417_;
  wire or_not_new_n3097__not_new_n3096_;
  wire not_new_n1585__9;
  wire new_n10070_;
  wire new_n9828_;
  wire not_pi140_1;
  wire not_new_n8595__6;
  wire not_pi174_1;
  wire not_new_n610__2;
  wire not_new_n1011__5;
  wire not_new_n4526_;
  wire new_n4980_;
  wire not_new_n8822_;
  wire new_n4481_;
  wire new_n1348_;
  wire not_new_n7436__1;
  wire or_not_new_n929__not_new_n931_;
  wire new_n10116_;
  wire not_new_n5601_;
  wire new_n643_;
  wire not_new_n8946_;
  wire not_new_n7330_;
  wire not_new_n8963__0;
  wire not_new_n5465__0;
  wire not_new_n1031__7;
  wire or_not_new_n6363__not_new_n6358_;
  wire not_new_n7034__1;
  wire new_n8241_;
  wire new_n9449_;
  wire new_n4189_;
  wire new_n5699_;
  wire po115;
  wire not_new_n615_;
  wire not_new_n3551_;
  wire new_n6676_;
  wire new_n1339_;
  wire not_new_n5074_;
  wire not_new_n4496_;
  wire new_n2087_;
  wire new_n8864_;
  wire new_n8647_;
  wire not_new_n1312_;
  wire not_new_n6772_;
  wire new_n3716_;
  wire not_pi061_0;
  wire not_new_n1581__24010;
  wire and_new_n7597__new_n7953_;
  wire not_new_n581__47475615099430;
  wire not_new_n740__0;
  wire not_new_n2187_;
  wire not_pi169_1;
  wire not_new_n8713_;
  wire new_n6161_;
  wire key_gate_115;
  wire new_n9129_;
  wire new_n5120_;
  wire or_not_new_n2034__not_new_n2035_;
  wire not_new_n1027__3430;
  wire not_new_n618__0;
  wire not_new_n3184__3430;
  wire new_n6224_;
  wire new_n9845_;
  wire new_n9302_;
  wire not_new_n3883_;
  wire not_new_n6165_;
  wire new_n8954_;
  wire new_n6160_;
  wire new_n8322_;
  wire and_new_n1754__new_n1755_;
  wire not_new_n5427_;
  wire not_po296_4;
  wire new_n3823_;
  wire not_new_n1534__7;
  wire not_new_n1051__10;
  wire new_n5084_;
  wire new_n5625_;
  wire new_n5619_;
  wire not_new_n9414__0;
  wire not_new_n598__70;
  wire new_n6317_;
  wire new_n5451_;
  wire new_n10271_;
  wire not_new_n591__968890104070;
  wire new_n7747_;
  wire not_new_n8798__2;
  wire new_n5039_;
  wire not_new_n4218_;
  wire or_not_new_n2545__not_new_n2544_;
  wire not_new_n6242__3;
  wire new_n4662_;
  wire not_new_n1728__0;
  wire or_not_new_n2547__not_new_n2551_;
  wire not_new_n6640__2;
  wire new_n8832_;
  wire not_new_n9217_;
  wire and_new_n8753__new_n8754_;
  wire not_new_n628__968890104070;
  wire not_new_n9900_;
  wire not_new_n638__47475615099430;
  wire not_new_n3977_;
  wire not_new_n8320_;
  wire not_new_n5442_;
  wire new_n6436_;
  wire not_new_n1165_;
  wire not_new_n2800_;
  wire new_n581_;
  wire not_new_n4600_;
  wire not_new_n596__8;
  wire new_n1750_;
  wire not_new_n5742_;
  wire not_new_n1047__490;
  wire new_n9538_;
  wire not_new_n9598_;
  wire new_n3701_;
  wire new_n9766_;
  wire not_new_n9721_;
  wire not_new_n5658_;
  wire not_new_n7555_;
  wire not_new_n1506_;
  wire not_pi273_1;
  wire new_n4479_;
  wire new_n6035_;
  wire new_n9253_;
  wire not_new_n7632__0;
  wire new_n7501_;
  wire new_n6210_;
  wire or_or_not_new_n3944__not_new_n3914__1_not_new_n4014__4;
  wire not_new_n3209_;
  wire not_new_n7094_;
  wire new_n9423_;
  wire not_new_n1510_;
  wire not_new_n9855__0;
  wire not_new_n9880__0;
  wire not_new_n6676_;
  wire not_new_n5481__0;
  wire not_new_n609__490;
  wire new_n5033_;
  wire not_new_n3695_;
  wire or_or_or_not_new_n2847__not_new_n2850__not_new_n2849__not_new_n2851_;
  wire not_new_n628__39098210485829880490;
  wire new_n5895_;
  wire new_n2250_;
  wire not_new_n9966__0;
  wire new_n8770_;
  wire or_not_new_n1319__not_new_n1317_;
  wire new_n5626_;
  wire not_new_n4511_;
  wire not_new_n8686_;
  wire not_new_n6958_;
  wire new_n3338_;
  wire new_n2579_;
  wire not_new_n7598__1;
  wire not_new_n10260_;
  wire not_new_n5643_;
  wire not_new_n1535_;
  wire not_new_n633__5;
  wire new_n3213_;
  wire new_n5972_;
  wire not_new_n2764_;
  wire new_n4417_;
  wire and_and_new_n2010__new_n2013__new_n2011_;
  wire new_n6312_;
  wire new_n8458_;
  wire not_new_n4284_;
  wire not_new_n1597__4;
  wire new_n1648_;
  wire not_new_n8590_;
  wire not_new_n3129_;
  wire new_n9111_;
  wire new_n7152_;
  wire not_new_n1580__24010;
  wire not_new_n1061__0;
  wire not_new_n7516_;
  wire new_n3148_;
  wire not_new_n594__47475615099430;
  wire new_n5650_;
  wire not_new_n4130__1;
  wire not_pi253_0;
  wire not_new_n6808_;
  wire not_new_n8541_;
  wire not_new_n625__4;
  wire new_n10204_;
  wire new_n4583_;
  wire new_n3660_;
  wire not_new_n9663_;
  wire new_n10088_;
  wire new_n7673_;
  wire new_n9410_;
  wire not_new_n4635_;
  wire not_new_n6978__1;
  wire not_new_n6630_;
  wire not_new_n1351_;
  wire new_n759_;
  wire new_n6125_;
  wire or_or_not_new_n1863__not_new_n1864__not_new_n1866_;
  wire new_n3221_;
  wire not_new_n1049__2326305139872070;
  wire not_new_n4471_;
  wire not_new_n7580_;
  wire not_new_n9161_;
  wire not_new_n9899_;
  wire new_n6694_;
  wire new_n10036_;
  wire not_new_n628__138412872010;
  wire new_n6087_;
  wire new_n5018_;
  wire not_new_n600__70;
  wire not_new_n3364_;
  wire not_new_n633__47475615099430;
  wire new_n1628_;
  wire new_n4992_;
  wire not_new_n7663__2;
  wire not_new_n630__2326305139872070;
  wire new_n6243_;
  wire not_new_n595__3430;
  wire new_n7296_;
  wire or_not_new_n2265__not_new_n2262_;
  wire not_new_n2346_;
  wire not_new_n6394_;
  wire new_n4499_;
  wire not_new_n9418_;
  wire new_n9396_;
  wire new_n8617_;
  wire new_n2943_;
  wire not_new_n587__19773267430;
  wire new_n6965_;
  wire not_new_n8901_;
  wire new_n4467_;
  wire or_or_or_not_new_n2946__not_new_n2949__not_new_n2948__not_new_n2950_;
  wire po081;
  wire not_pi026_0;
  wire new_n7136_;
  wire not_new_n7768_;
  wire and_new_n1326__new_n2255_;
  wire new_n5289_;
  wire not_new_n9842_;
  wire new_n1654_;
  wire new_n5546_;
  wire not_new_n6242_;
  wire not_new_n3185__19773267430;
  wire not_new_n4122__2;
  wire not_new_n6475_;
  wire not_pi258_1;
  wire not_new_n4000__0;
  wire not_new_n745__0;
  wire new_n9664_;
  wire or_or_not_new_n2547__not_new_n2551__not_new_n1425_;
  wire new_n5450_;
  wire not_po296_1742514982336908143055105517947102601079450420187483430;
  wire not_new_n1576__3;
  wire not_new_n8181_;
  wire not_new_n1602__2824752490;
  wire not_new_n621__968890104070;
  wire new_n7459_;
  wire not_new_n4425__0;
  wire key_gate_54;
  wire new_n970_;
  wire new_n10279_;
  wire new_n3049_;
  wire not_new_n989__70;
  wire not_new_n4156_;
  wire po245;
  wire new_n2335_;
  wire new_n4887_;
  wire new_n2207_;
  wire not_new_n9815_;
  wire new_n4553_;
  wire not_new_n3998_;
  wire not_new_n1018__7;
  wire or_not_new_n2655__not_new_n2654_;
  wire not_new_n3107_;
  wire new_n7320_;
  wire or_or_not_new_n1977__not_new_n1978__not_new_n1980_;
  wire not_new_n4209_;
  wire not_new_n611__9;
  wire not_pi262;
  wire new_n2238_;
  wire new_n8308_;
  wire new_n5837_;
  wire not_new_n7629_;
  wire not_new_n7515_;
  wire not_new_n1585__490;
  wire not_new_n3482_;
  wire not_new_n2693_;
  wire new_n6031_;
  wire not_new_n3144_;
  wire not_new_n4500__0;
  wire not_new_n1028__10;
  wire new_n4237_;
  wire new_n8946_;
  wire not_pi193;
  wire new_n5325_;
  wire not_new_n586__6;
  wire new_n9284_;
  wire new_n9531_;
  wire new_n4071_;
  wire new_n7539_;
  wire not_new_n4686_;
  wire new_n7196_;
  wire not_new_n8913_;
  wire new_n5395_;
  wire not_new_n775__1;
  wire and_new_n1338__new_n2312_;
  wire new_n1620_;
  wire new_n6199_;
  wire or_or_or_not_new_n2776__not_new_n2779__not_new_n2778__not_new_n2780_;
  wire not_new_n600__5;
  wire new_n5440_;
  wire new_n1265_;
  wire not_new_n4137__1;
  wire not_new_n1534__797922662976120010;
  wire not_new_n647__5;
  wire and_and_new_n1053__new_n6232__new_n6395_;
  wire not_new_n6631__1;
  wire not_new_n1045__2;
  wire new_n3681_;
  wire not_new_n1061__3;
  wire key_gate_86;
  wire new_n1498_;
  wire not_new_n4257_;
  wire not_new_n7380_;
  wire not_new_n1028__4;
  wire not_new_n4285_;
  wire new_n10114_;
  wire not_new_n7554_;
  wire not_new_n2975_;
  wire not_new_n581__445676403263631959001900459745680070;
  wire not_new_n1006__4;
  wire not_new_n984__490;
  wire not_new_n6093_;
  wire new_n9757_;
  wire new_n10332_;
  wire new_n3625_;
  wire new_n4829_;
  wire not_new_n9929__0;
  wire new_n5375_;
  wire new_n7317_;
  wire new_n8400_;
  wire new_n6878_;
  wire not_new_n10005_;
  wire new_n6988_;
  wire not_new_n9934__0;
  wire not_new_n1537__1176490;
  wire new_n8847_;
  wire or_not_new_n2615__not_new_n2614_;
  wire not_new_n600__3430;
  wire new_n9978_;
  wire new_n6453_;
  wire not_new_n598__138412872010;
  wire new_n9189_;
  wire not_new_n8875_;
  wire new_n2879_;
  wire new_n3132_;
  wire new_n3618_;
  wire not_new_n7739__2;
  wire po045;
  wire not_new_n4084_;
  wire new_n1937_;
  wire not_new_n7115__0;
  wire not_po296;
  wire not_new_n9552_;
  wire new_n3062_;
  wire not_new_n8357_;
  wire not_new_n6242__1;
  wire new_n6366_;
  wire not_new_n765_;
  wire new_n625_;
  wire not_new_n591__8235430;
  wire not_new_n6354_;
  wire new_n8465_;
  wire and_new_n2314__new_n2317_;
  wire not_new_n1027__13410686196639649008070;
  wire not_po296_5585458640832840070;
  wire not_new_n3462_;
  wire not_new_n1018__6;
  wire not_new_n3399_;
  wire not_new_n645__1;
  wire new_n7984_;
  wire new_n10023_;
  wire new_n7398_;
  wire new_n4514_;
  wire not_new_n677_;
  wire not_new_n605__24010;
  wire not_new_n581__9;
  wire key_gate_102;
  wire not_new_n1479_;
  wire new_n7620_;
  wire not_new_n1601__93874803376477543056490;
  wire not_new_n638__2824752490;
  wire new_n3356_;
  wire not_new_n9935_;
  wire not_new_n1537__797922662976120010;
  wire new_n5511_;
  wire not_new_n4946_;
  wire not_new_n1581__168070;
  wire not_new_n8167_;
  wire new_n5379_;
  wire new_n9007_;
  wire new_n3515_;
  wire new_n602_;
  wire new_n3458_;
  wire new_n4306_;
  wire new_n1763_;
  wire new_n8607_;
  wire not_new_n3530_;
  wire not_new_n6963_;
  wire new_n1956_;
  wire not_pi260_3;
  wire po256;
  wire new_n7475_;
  wire not_new_n7143__0;
  wire not_new_n4223_;
  wire not_new_n10122_;
  wire not_new_n989__24010;
  wire po043;
  wire not_new_n9038_;
  wire not_new_n6233_;
  wire or_or_not_new_n2577__not_new_n2581__not_new_n1431_;
  wire or_not_new_n1553__not_new_n1376_;
  wire not_new_n4098_;
  wire not_new_n6090_;
  wire new_n7458_;
  wire not_new_n775__2824752490;
  wire new_n6564_;
  wire new_n5082_;
  wire not_new_n3272_;
  wire new_n8853_;
  wire not_new_n7610_;
  wire not_new_n3210_;
  wire new_n5997_;
  wire new_n8134_;
  wire new_n4011_;
  wire not_new_n2916_;
  wire not_pi021;
  wire not_pi139_1;
  wire not_new_n5096_;
  wire new_n6113_;
  wire not_po296_3788186922656647816827176259430;
  wire not_pi064_0;
  wire not_new_n4965_;
  wire new_n10226_;
  wire not_new_n9382__0;
  wire not_new_n1597__10;
  wire new_n2405_;
  wire new_n3328_;
  wire not_new_n1614_;
  wire not_new_n2734_;
  wire new_n2696_;
  wire not_new_n9118__0;
  wire new_n5722_;
  wire new_n4883_;
  wire not_new_n1881__0;
  wire new_n8247_;
  wire not_new_n645__2;
  wire new_n7678_;
  wire po253;
  wire or_or_or_not_new_n6226__0_not_new_n6336__not_new_n6373__5_not_new_n6242__2;
  wire not_new_n594__0;
  wire not_new_n3901_;
  wire new_n9401_;
  wire not_new_n9406_;
  wire not_new_n10029__0;
  wire not_new_n8966_;
  wire not_new_n6979__0;
  wire not_new_n3497_;
  wire new_n1328_;
  wire new_n1321_;
  wire new_n9299_;
  wire new_n8699_;
  wire not_new_n6443__6;
  wire new_n7256_;
  wire new_n5529_;
  wire not_new_n7627__2;
  wire new_n8887_;
  wire not_new_n724__0;
  wire po086;
  wire not_new_n586__490;
  wire not_new_n1602__19773267430;
  wire new_n7044_;
  wire new_n2527_;
  wire not_new_n5916__0;
  wire not_new_n1013__3;
  wire not_new_n2502_;
  wire new_n7585_;
  wire not_new_n3481_;
  wire new_n3642_;
  wire not_new_n5322_;
  wire not_new_n1585__138412872010;
  wire not_new_n4179_;
  wire not_new_n1232_;
  wire new_n4705_;
  wire new_n3745_;
  wire new_n3675_;
  wire new_n1342_;
  wire new_n4316_;
  wire not_pi263_1;
  wire not_new_n5752_;
  wire not_new_n1039__113988951853731430;
  wire not_new_n5408_;
  wire not_new_n2591_;
  wire not_new_n5782_;
  wire not_new_n9667_;
  wire not_new_n9914_;
  wire not_new_n7091_;
  wire not_new_n8216_;
  wire not_new_n7611_;
  wire not_new_n3130_;
  wire new_n5346_;
  wire not_new_n9854__1;
  wire not_new_n688_;
  wire new_n4768_;
  wire not_new_n4110_;
  wire not_new_n1589__403536070;
  wire not_new_n4996_;
  wire new_n1331_;
  wire new_n9158_;
  wire new_n10068_;
  wire new_n4103_;
  wire new_n10052_;
  wire not_new_n5443_;
  wire new_n8302_;
  wire new_n10111_;
  wire not_new_n8898_;
  wire not_new_n589__4;
  wire new_n2580_;
  wire new_n6567_;
  wire new_n8794_;
  wire not_po296_8235430;
  wire not_new_n4316_;
  wire new_n4898_;
  wire new_n4957_;
  wire not_new_n7664__0;
  wire new_n4528_;
  wire not_new_n3781_;
  wire new_n10143_;
  wire not_new_n1024__0;
  wire new_n679_;
  wire not_new_n7904_;
  wire new_n6725_;
  wire new_n6896_;
  wire new_n4444_;
  wire or_not_new_n1323__not_new_n1321_;
  wire not_new_n4676_;
  wire new_n8787_;
  wire not_new_n1596__19773267430;
  wire not_new_n6332_;
  wire not_new_n610__5;
  wire new_n6301_;
  wire not_new_n2342_;
  wire not_new_n1055__1176490;
  wire new_n3020_;
  wire not_new_n606__70;
  wire not_new_n2167_;
  wire not_new_n4135__0;
  wire new_n9516_;
  wire not_new_n6303_;
  wire not_new_n611__8;
  wire not_new_n588__9;
  wire not_new_n8515_;
  wire new_n6346_;
  wire not_new_n1580__332329305696010;
  wire not_new_n5894_;
  wire not_new_n8275_;
  wire new_n3262_;
  wire new_n4044_;
  wire not_new_n8658_;
  wire not_new_n5193_;
  wire new_n7212_;
  wire not_new_n9339_;
  wire new_n9286_;
  wire new_n2399_;
  wire not_new_n1199_;
  wire not_new_n6777_;
  wire new_n8063_;
  wire new_n1298_;
  wire not_new_n2247_;
  wire new_n9444_;
  wire new_n7692_;
  wire not_new_n1045__1;
  wire not_new_n4170__0;
  wire new_n5796_;
  wire not_new_n2795_;
  wire new_n6822_;
  wire new_n1772_;
  wire not_new_n1576__3430;
  wire new_n9261_;
  wire not_new_n2634_;
  wire new_n3619_;
  wire not_new_n8884_;
  wire not_pi097_0;
  wire not_new_n631__2;
  wire new_n6306_;
  wire not_new_n5377_;
  wire new_n1980_;
  wire not_new_n3940_;
  wire new_n9779_;
  wire new_n2861_;
  wire not_new_n1585__0;
  wire not_new_n4445__0;
  wire new_n9169_;
  wire new_n7926_;
  wire not_new_n5581_;
  wire not_new_n629__0;
  wire not_new_n8870_;
  wire not_new_n9015_;
  wire not_new_n4122_;
  wire new_n1701_;
  wire new_n3406_;
  wire new_n3519_;
  wire new_n7359_;
  wire new_n3097_;
  wire not_pi176_1;
  wire new_n9716_;
  wire and_new_n3804__new_n3807_;
  wire not_new_n10248_;
  wire not_new_n1323_;
  wire not_new_n1621_;
  wire not_new_n637_;
  wire new_n5470_;
  wire new_n6296_;
  wire and_new_n2517__new_n2518_;
  wire not_new_n1576__57648010;
  wire new_n6891_;
  wire not_new_n4713_;
  wire new_n4655_;
  wire not_new_n4993__0;
  wire new_n8448_;
  wire or_not_new_n1158__0_not_new_n8713__1;
  wire not_new_n4842_;
  wire not_new_n1583__70;
  wire new_n659_;
  wire not_new_n1341_;
  wire not_new_n4245_;
  wire not_new_n1071__138412872010;
  wire new_n3534_;
  wire not_new_n3959_;
  wire new_n6136_;
  wire not_new_n9079_;
  wire not_new_n626__332329305696010;
  wire not_new_n764_;
  wire new_n7171_;
  wire new_n7583_;
  wire new_n5925_;
  wire new_n4440_;
  wire not_new_n8849_;
  wire not_new_n6126_;
  wire not_new_n7620__0;
  wire or_not_new_n10045__1_not_new_n9855__1;
  wire new_n3083_;
  wire not_new_n628__3430;
  wire new_n8143_;
  wire new_n2277_;
  wire new_n7402_;
  wire not_new_n1535__0;
  wire new_n3509_;
  wire new_n4431_;
  wire not_new_n2134_;
  wire not_new_n7448__0;
  wire not_new_n5769_;
  wire not_new_n1020__7;
  wire not_new_n643__6782230728490;
  wire new_n7763_;
  wire not_new_n10083_;
  wire not_new_n1491_;
  wire not_new_n622__7;
  wire not_new_n647__0;
  wire new_n6424_;
  wire key_gate_38;
  wire not_new_n3925_;
  wire new_n9722_;
  wire not_new_n1730__0;
  wire not_new_n7019_;
  wire not_new_n10329_;
  wire po280;
  wire not_new_n4779__0;
  wire new_n1945_;
  wire not_new_n9866_;
  wire new_n7725_;
  wire new_n3430_;
  wire not_new_n4226_;
  wire not_new_n4835_;
  wire not_new_n8235_;
  wire not_new_n5681_;
  wire not_new_n1043__8235430;
  wire po266;
  wire not_new_n1059__4;
  wire not_new_n3372__39098210485829880490;
  wire not_new_n3185__3;
  wire new_n5698_;
  wire new_n7298_;
  wire not_pi165_0;
  wire or_not_new_n6897__not_new_n6798_;
  wire new_n2795_;
  wire not_new_n7427__0;
  wire new_n1337_;
  wire and_new_n1043__new_n6232_;
  wire new_n3813_;
  wire not_new_n1591__3;
  wire not_new_n5920__0;
  wire new_n5372_;
  wire not_new_n644__2824752490;
  wire or_or_or_not_new_n2874__not_new_n2877__not_new_n2876__not_new_n2878_;
  wire not_new_n5078_;
  wire not_new_n7781__0;
  wire new_n8406_;
  wire not_new_n634__0;
  wire not_new_n4200_;
  wire not_new_n664_;
  wire not_new_n1069__968890104070;
  wire not_new_n6709_;
  wire new_n2143_;
  wire new_n4175_;
  wire new_n7358_;
  wire not_new_n9248_;
  wire new_n9309_;
  wire new_n7665_;
  wire new_n6977_;
  wire not_new_n6000_;
  wire not_new_n6607_;
  wire new_n10031_;
  wire new_n2899_;
  wire not_new_n595__5;
  wire not_new_n1159_;
  wire not_new_n10198_;
  wire not_new_n4265_;
  wire not_new_n922__1;
  wire new_n2517_;
  wire not_new_n9761_;
  wire new_n9908_;
  wire not_new_n7773_;
  wire new_n2991_;
  wire and_new_n2697__new_n2698_;
  wire new_n9729_;
  wire not_new_n606__5;
  wire new_n6105_;
  wire new_n2659_;
  wire not_new_n585__2326305139872070;
  wire new_n4281_;
  wire new_n4565_;
  wire not_new_n5704_;
  wire not_new_n2888_;
  wire new_n7474_;
  wire new_n8491_;
  wire not_new_n928__7;
  wire new_n3987_;
  wire not_new_n7152__0;
  wire or_not_new_n5203__not_new_n5087__0;
  wire new_n8057_;
  wire new_n3571_;
  wire new_n4607_;
  wire not_new_n3397_;
  wire new_n6151_;
  wire not_pi144_2;
  wire new_n3329_;
  wire not_new_n6479_;
  wire not_new_n610__70;
  wire not_new_n5200_;
  wire not_new_n610__8235430;
  wire not_new_n989__19773267430;
  wire not_new_n8660_;
  wire not_new_n4158_;
  wire not_new_n5595_;
  wire new_n4033_;
  wire not_new_n3214_;
  wire not_new_n10177_;
  wire new_n7001_;
  wire new_n5647_;
  wire new_n4585_;
  wire not_new_n9381_;
  wire not_new_n7167_;
  wire new_n2747_;
  wire not_new_n644__16284135979104490;
  wire not_new_n4113_;
  wire not_new_n597__8;
  wire new_n9244_;
  wire not_new_n734__0;
  wire new_n1979_;
  wire not_new_n3011_;
  wire not_new_n618__10;
  wire not_new_n617__138412872010;
  wire and_and_not_pi048_2_not_pi047_2_not_pi050_2;
  wire new_n5803_;
  wire new_n2535_;
  wire not_new_n9013__0;
  wire new_n5911_;
  wire new_n4466_;
  wire not_new_n7445__1;
  wire new_n2753_;
  wire not_new_n1368_;
  wire not_new_n3474_;
  wire new_n7080_;
  wire new_n3852_;
  wire not_new_n775__332329305696010;
  wire new_n8502_;
  wire or_not_new_n1307__not_new_n1305_;
  wire not_new_n3737_;
  wire not_new_n8246_;
  wire new_n10161_;
  wire new_n3718_;
  wire not_new_n6299_;
  wire new_n5365_;
  wire new_n6009_;
  wire not_new_n1537__19773267430;
  wire new_n9876_;
  wire not_new_n1296_;
  wire not_new_n2643_;
  wire new_n10174_;
  wire not_new_n4999__1;
  wire key_gate_107;
  wire not_new_n1031__8;
  wire not_new_n1782_;
  wire not_new_n5663_;
  wire not_new_n629__47475615099430;
  wire not_new_n1616__968890104070;
  wire not_new_n8043_;
  wire new_n9164_;
  wire new_n10090_;
  wire not_new_n6238_;
  wire po206;
  wire key_gate_44;
  wire not_new_n1512_;
  wire not_new_n6443__3430;
  wire new_n6790_;
  wire new_n2463_;
  wire new_n3404_;
  wire and_and_new_n2086__new_n2089__new_n2087_;
  wire not_new_n9478_;
  wire not_new_n7778_;
  wire not_new_n3123_;
  wire new_n6542_;
  wire not_new_n2644_;
  wire not_new_n4240_;
  wire new_n1562_;
  wire new_n5209_;
  wire new_n3306_;
  wire new_n5845_;
  wire not_new_n631__13410686196639649008070;
  wire not_new_n9900__0;
  wire not_new_n1039__8235430;
  wire not_new_n9005_;
  wire not_new_n2810_;
  wire not_new_n3290_;
  wire new_n7776_;
  wire not_pi078;
  wire or_pi033_pi035;
  wire new_n696_;
  wire not_new_n1581__5;
  wire not_new_n9436_;
  wire not_new_n4913_;
  wire new_n4671_;
  wire not_new_n4155_;
  wire new_n7376_;
  wire not_new_n994__138412872010;
  wire not_new_n10148_;
  wire not_new_n7018__1;
  wire not_new_n1049__3;
  wire not_new_n6621_;
  wire not_new_n5114_;
  wire new_n9650_;
  wire not_new_n3556_;
  wire new_n9834_;
  wire or_not_new_n1596__403536070_not_new_n7586_;
  wire not_new_n7749_;
  wire not_new_n5057_;
  wire or_or_not_new_n6226__0_not_new_n6336__not_new_n6373__5;
  wire not_new_n1591__47475615099430;
  wire not_new_n5791__1;
  wire not_new_n602__138412872010;
  wire not_new_n642__19773267430;
  wire not_new_n1409_;
  wire new_n3436_;
  wire not_new_n5656_;
  wire not_new_n6661_;
  wire not_new_n594__8235430;
  wire not_new_n621__5585458640832840070;
  wire new_n7602_;
  wire new_n1214_;
  wire not_new_n3300_;
  wire not_new_n6593_;
  wire new_n3485_;
  wire new_n6398_;
  wire not_new_n628__4;
  wire not_new_n8420_;
  wire new_n8785_;
  wire new_n6974_;
  wire new_n6138_;
  wire not_new_n9670_;
  wire not_new_n4761__0;
  wire new_n1268_;
  wire new_n4960_;
  wire new_n2341_;
  wire new_n8881_;
  wire not_new_n1594__0;
  wire new_n8122_;
  wire not_new_n9871_;
  wire not_new_n1611__6;
  wire not_new_n6272_;
  wire not_new_n2076_;
  wire new_n6641_;
  wire new_n10325_;
  wire new_n5868_;
  wire new_n7846_;
  wire new_n5057_;
  wire new_n5838_;
  wire new_n8341_;
  wire not_new_n7142_;
  wire new_n8723_;
  wire new_n5409_;
  wire new_n5665_;
  wire not_new_n1027__9;
  wire new_n4121_;
  wire not_new_n624__8;
  wire not_new_n5750_;
  wire not_new_n7876_;
  wire not_new_n5037_;
  wire new_n8180_;
  wire not_new_n5336_;
  wire new_n1419_;
  wire new_n4245_;
  wire or_not_new_n6780__not_new_n6662_;
  wire not_new_n6046_;
  wire new_n5184_;
  wire not_new_n1585__2824752490;
  wire or_not_new_n6073__not_new_n6048_;
  wire not_new_n2967_;
  wire new_n10337_;
  wire new_n6098_;
  wire not_new_n723__0;
  wire not_new_n1014__6;
  wire new_n3010_;
  wire new_n7005_;
  wire not_new_n3850_;
  wire new_n2162_;
  wire new_n4434_;
  wire new_n5066_;
  wire not_new_n6173_;
  wire new_n4433_;
  wire new_n8840_;
  wire new_n2675_;
  wire not_new_n3318__0;
  wire not_new_n4317_;
  wire not_new_n9138_;
  wire not_new_n6059_;
  wire new_n6150_;
  wire po064;
  wire new_n2900_;
  wire new_n1933_;
  wire new_n3037_;
  wire not_new_n1589__3430;
  wire not_new_n1580__47475615099430;
  wire new_n6053_;
  wire not_new_n1150_;
  wire not_new_n6270_;
  wire not_new_n639__3430;
  wire new_n3699_;
  wire not_new_n641__8;
  wire new_n1629_;
  wire not_new_n6524__2;
  wire new_n8138_;
  wire new_n1707_;
  wire new_n3738_;
  wire new_n6605_;
  wire not_new_n1182_;
  wire not_new_n7883_;
  wire not_new_n1037__47475615099430;
  wire new_n9863_;
  wire not_new_n4512_;
  wire not_new_n1071__3;
  wire new_n4910_;
  wire po219;
  wire not_new_n608__8;
  wire new_n2211_;
  wire po263;
  wire not_new_n3800_;
  wire new_n7929_;
  wire new_n7119_;
  wire not_new_n7632_;
  wire not_new_n3531_;
  wire new_n6286_;
  wire not_new_n1631__168070;
  wire not_new_n5290_;
  wire new_n5887_;
  wire not_po296_19773267430;
  wire new_n4847_;
  wire new_n8619_;
  wire not_new_n617__9;
  wire not_new_n645__6782230728490;
  wire new_n9150_;
  wire not_new_n5825_;
  wire not_new_n8983_;
  wire new_n1835_;
  wire not_new_n586__0;
  wire not_new_n3184__9;
  wire new_n8054_;
  wire not_new_n1631__2326305139872070;
  wire new_n9361_;
  wire new_n3837_;
  wire not_new_n775__10;
  wire not_new_n1251_;
  wire not_new_n1016__2;
  wire po068;
  wire new_n7914_;
  wire not_new_n3241_;
  wire new_n8165_;
  wire not_new_n8183_;
  wire or_not_new_n6337__not_new_n6373__6;
  wire new_n2708_;
  wire not_new_n4458__0;
  wire not_new_n8897_;
  wire not_new_n2168_;
  wire not_new_n7808_;
  wire not_pi195;
  wire not_new_n6765_;
  wire not_new_n5182_;
  wire not_new_n2348__0;
  wire not_new_n8261_;
  wire not_new_n1538__16284135979104490;
  wire new_n584_;
  wire not_new_n9029_;
  wire new_n3691_;
  wire not_new_n6443__1176490;
  wire not_new_n9082_;
  wire not_new_n8340_;
  wire not_new_n4613_;
  wire not_pi045_1;
  wire not_new_n645_;
  wire new_n2061_;
  wire new_n6625_;
  wire not_new_n1612__70;
  wire new_n10126_;
  wire new_n6870_;
  wire not_new_n626__657123623635342801395430;
  wire not_new_n8174_;
  wire new_n1203_;
  wire new_n8921_;
  wire new_n7356_;
  wire not_new_n3309_;
  wire not_new_n6235_;
  wire not_new_n9028__0;
  wire not_new_n6339_;
  wire not_new_n10046__0;
  wire not_new_n593__968890104070;
  wire not_pi274_2;
  wire not_new_n1429_;
  wire not_new_n1069__2824752490;
  wire new_n1944_;
  wire not_new_n3315__16284135979104490;
  wire new_n1553_;
  wire not_new_n5890_;
  wire or_not_new_n3152__not_new_n3151_;
  wire new_n6167_;
  wire new_n4051_;
  wire not_new_n2789_;
  wire not_new_n4764_;
  wire not_new_n1536__5;
  wire not_new_n1041__19773267430;
  wire new_n5253_;
  wire new_n2242_;
  wire new_n2973_;
  wire new_n1317_;
  wire not_new_n4402_;
  wire po207;
  wire new_n5163_;
  wire new_n8166_;
  wire not_new_n6718_;
  wire not_pi140;
  wire new_n5046_;
  wire new_n4087_;
  wire new_n3386_;
  wire new_n2329_;
  wire not_new_n1631__16284135979104490;
  wire not_new_n9768_;
  wire not_pi272_2;
  wire not_new_n1176__0;
  wire new_n6499_;
  wire new_n3179_;
  wire new_n10166_;
  wire not_new_n8722_;
  wire not_new_n8135_;
  wire new_n10141_;
  wire not_new_n612__0;
  wire not_new_n5742__1;
  wire not_pi269_0;
  wire not_new_n1982_;
  wire not_new_n9199_;
  wire new_n8467_;
  wire not_new_n1057__70;
  wire not_new_n4801_;
  wire not_new_n984__2824752490;
  wire new_n9107_;
  wire new_n4806_;
  wire not_new_n8521_;
  wire not_new_n8123_;
  wire new_n6240_;
  wire not_new_n1063__5;
  wire not_new_n3296_;
  wire not_new_n9387__0;
  wire new_n3559_;
  wire new_n1535_;
  wire not_new_n589__6782230728490;
  wire not_new_n7028__0;
  wire not_new_n638__5;
  wire not_new_n6498__0;
  wire not_new_n1024__1;
  wire new_n7263_;
  wire not_pi064_2326305139872070;
  wire new_n4527_;
  wire new_n692_;
  wire new_n7617_;
  wire and_new_n2508__new_n2510_;
  wire not_new_n8150_;
  wire new_n649_;
  wire not_new_n1059__403536070;
  wire or_not_new_n1901__not_new_n1902_;
  wire new_n3978_;
  wire or_not_new_n2971__not_new_n2970_;
  wire not_pi146_3;
  wire new_n8223_;
  wire not_new_n1537_;
  wire not_new_n3739_;
  wire new_n2731_;
  wire not_new_n8419_;
  wire not_new_n6527_;
  wire new_n5217_;
  wire new_n6919_;
  wire not_new_n8453_;
  wire not_new_n9101_;
  wire and_new_n3780__new_n3783_;
  wire new_n1157_;
  wire not_new_n5368_;
  wire new_n9448_;
  wire new_n1883_;
  wire new_n3831_;
  wire not_new_n3930_;
  wire not_new_n9878_;
  wire new_n7830_;
  wire not_new_n3195_;
  wire new_n6587_;
  wire not_new_n8189_;
  wire not_new_n603__0;
  wire not_new_n5952_;
  wire new_n7192_;
  wire not_new_n5084__1;
  wire not_new_n589__152867006319425761937651857692768264010;
  wire not_new_n8518_;
  wire not_new_n9614_;
  wire and_new_n1286__new_n2065_;
  wire not_new_n732_;
  wire not_new_n8155__2;
  wire not_new_n594__16284135979104490;
  wire new_n3783_;
  wire not_new_n7612_;
  wire not_new_n625__9;
  wire not_new_n9769_;
  wire new_n4945_;
  wire not_new_n4309_;
  wire not_new_n1565_;
  wire not_new_n7333_;
  wire new_n6388_;
  wire new_n5219_;
  wire not_new_n4845_;
  wire not_new_n6974__8;
  wire not_new_n624__0;
  wire new_n3479_;
  wire not_new_n5906_;
  wire not_new_n8596_;
  wire new_n6117_;
  wire new_n3456_;
  wire new_n3327_;
  wire new_n5725_;
  wire new_n631_;
  wire or_not_new_n7715__not_new_n7714_;
  wire not_new_n1616__4;
  wire not_new_n5786__1;
  wire not_new_n5792__0;
  wire new_n984_;
  wire not_new_n7212__0;
  wire not_new_n6634__0;
  wire not_new_n6071_;
  wire new_n2465_;
  wire not_new_n1631__3;
  wire and_new_n2513__new_n2512_;
  wire not_new_n636__8;
  wire not_new_n618__2824752490;
  wire new_n8515_;
  wire new_n4625_;
  wire not_new_n6642_;
  wire not_new_n6145_;
  wire not_new_n2018_;
  wire not_new_n7131_;
  wire not_new_n6177_;
  wire and_and_new_n2200__new_n2203__new_n2201_;
  wire not_new_n10249_;
  wire new_n1392_;
  wire new_n7770_;
  wire not_new_n5640_;
  wire not_new_n4593_;
  wire not_new_n4237_;
  wire po278;
  wire new_n1441_;
  wire not_new_n595__2824752490;
  wire new_n4971_;
  wire not_new_n1598__2326305139872070;
  wire not_new_n10245_;
  wire and_new_n3306__new_n3305_;
  wire not_new_n694_;
  wire not_new_n619__1;
  wire not_new_n5566_;
  wire not_new_n2749_;
  wire new_n5092_;
  wire new_n2067_;
  wire not_new_n3562_;
  wire not_new_n4939_;
  wire new_n1423_;
  wire new_n2443_;
  wire new_n3084_;
  wire new_n3425_;
  wire not_new_n2794_;
  wire not_new_n4381_;
  wire not_pi260_2;
  wire not_new_n636__5;
  wire or_not_new_n1339__not_new_n1337_;
  wire not_new_n581__6168735096280623662907561568153897267931784070;
  wire new_n10119_;
  wire new_n7923_;
  wire new_n6899_;
  wire not_pi179;
  wire not_new_n5095__0;
  wire or_not_new_n4240__not_new_n4343_;
  wire new_n7598_;
  wire new_n6106_;
  wire new_n4168_;
  wire new_n7189_;
  wire new_n1361_;
  wire not_new_n7896_;
  wire not_new_n7724_;
  wire not_new_n602__8235430;
  wire new_n6347_;
  wire not_new_n7670_;
  wire new_n743_;
  wire new_n4540_;
  wire not_new_n8850_;
  wire not_new_n7649__0;
  wire not_new_n9099__0;
  wire new_n9439_;
  wire not_new_n4426_;
  wire not_new_n3245_;
  wire not_new_n8113_;
  wire not_new_n9956__0;
  wire not_new_n3101_;
  wire or_not_new_n6353__not_new_n6232__5;
  wire new_n6280_;
  wire not_new_n9557_;
  wire not_new_n8106__0;
  wire not_new_n4612_;
  wire new_n4002_;
  wire not_new_n5884__0;
  wire not_po296_2;
  wire not_new_n6528_;
  wire not_new_n10171_;
  wire not_new_n2543_;
  wire not_new_n8348_;
  wire not_new_n10046_;
  wire not_new_n632__332329305696010;
  wire new_n8624_;
  wire not_new_n4163__1;
  wire not_new_n1602__24010;
  wire not_new_n3471_;
  wire not_new_n595__2;
  wire new_n8977_;
  wire not_new_n5444__0;
  wire or_or_not_new_n1263__not_new_n1261__not_new_n1945_;
  wire new_n3214_;
  wire not_new_n7138__0;
  wire not_new_n8265__2;
  wire not_new_n10154_;
  wire not_new_n6660_;
  wire not_new_n1381_;
  wire not_new_n633__3430;
  wire not_new_n647__3;
  wire not_new_n5959_;
  wire not_new_n1061__9;
  wire not_new_n8441_;
  wire new_n6003_;
  wire new_n5740_;
  wire not_new_n7044__0;
  wire not_new_n775__403536070;
  wire not_new_n6030_;
  wire not_new_n604__6782230728490;
  wire not_new_n7164_;
  wire not_new_n7856_;
  wire not_new_n4992__0;
  wire not_new_n7148_;
  wire not_new_n5393_;
  wire new_n3765_;
  wire new_n4280_;
  wire new_n9912_;
  wire not_new_n9584_;
  wire not_pi090;
  wire not_pi175_3;
  wire new_n10055_;
  wire new_n4975_;
  wire new_n1975_;
  wire new_n9631_;
  wire not_new_n7132_;
  wire and_new_n8828__new_n9210_;
  wire not_new_n8058_;
  wire new_n6536_;
  wire new_n9297_;
  wire not_new_n1613__57648010;
  wire not_new_n647__2326305139872070;
  wire new_n1428_;
  wire new_n2330_;
  wire not_new_n6350_;
  wire not_new_n1006__1;
  wire not_pi184;
  wire not_new_n1007__6;
  wire not_new_n1063__16284135979104490;
  wire not_new_n6195_;
  wire not_new_n8344_;
  wire not_new_n3882_;
  wire new_n10184_;
  wire not_new_n9433_;
  wire not_new_n4677_;
  wire new_n3756_;
  wire new_n4679_;
  wire new_n8726_;
  wire new_n9249_;
  wire new_n4513_;
  wire new_n3685_;
  wire not_pi223;
  wire not_new_n940__0;
  wire new_n6183_;
  wire new_n4210_;
  wire new_n6166_;
  wire new_n4068_;
  wire new_n8366_;
  wire not_new_n586__113988951853731430;
  wire not_new_n4119__1;
  wire not_new_n4816__0;
  wire not_pi161;
  wire not_new_n5599_;
  wire new_n640_;
  wire new_n4761_;
  wire not_new_n1061__138412872010;
  wire not_new_n1045__332329305696010;
  wire new_n6902_;
  wire not_new_n3184__168070;
  wire or_not_new_n4816__not_new_n4751_;
  wire new_n5811_;
  wire new_n4988_;
  wire new_n5265_;
  wire not_new_n7578_;
  wire new_n3112_;
  wire new_n6667_;
  wire not_new_n4987_;
  wire not_new_n2526_;
  wire not_new_n2245_;
  wire not_new_n7479_;
  wire and_and_new_n2162__new_n2165__new_n2163_;
  wire not_new_n6976_;
  wire new_n10284_;
  wire not_new_n6446_;
  wire or_or_not_new_n2838__not_new_n2841__not_new_n2840_;
  wire not_new_n1580__1;
  wire new_n6154_;
  wire not_new_n611__1176490;
  wire not_new_n2741_;
  wire new_n6129_;
  wire new_n7216_;
  wire not_new_n1603__2824752490;
  wire new_n1245_;
  wire new_n8059_;
  wire not_new_n589__16284135979104490;
  wire new_n6295_;
  wire not_new_n5621_;
  wire not_new_n2758_;
  wire not_new_n2161_;
  wire new_n4010_;
  wire new_n9923_;
  wire or_or_not_new_n1473__not_new_n2722__not_new_n2723_;
  wire new_n9380_;
  wire new_n3914_;
  wire new_n1756_;
  wire new_n1621_;
  wire not_new_n607_;
  wire not_new_n1065__57648010;
  wire not_new_n7645_;
  wire not_new_n8522_;
  wire not_new_n1063__19773267430;
  wire not_new_n3273_;
  wire po267;
  wire not_new_n3767_;
  wire not_new_n617__2326305139872070;
  wire not_new_n6010_;
  wire not_new_n5262_;
  wire new_n7793_;
  wire not_new_n4340_;
  wire new_n4594_;
  wire not_pi073;
  wire new_n7194_;
  wire new_n6976_;
  wire not_new_n594__1176490;
  wire new_n1515_;
  wire not_new_n7662__0;
  wire new_n4423_;
  wire not_new_n6761_;
  wire new_n7348_;
  wire not_new_n1581__8;
  wire new_n1525_;
  wire not_new_n6133_;
  wire new_n3795_;
  wire new_n3291_;
  wire not_new_n4118_;
  wire not_new_n8886_;
  wire not_new_n9554_;
  wire not_new_n10157_;
  wire new_n8092_;
  wire not_new_n640__1176490;
  wire new_n7405_;
  wire not_new_n5056__0;
  wire new_n2949_;
  wire not_new_n3981_;
  wire not_new_n8595_;
  wire not_new_n7589_;
  wire not_new_n610__7;
  wire new_n2992_;
  wire new_n1154_;
  wire new_n8692_;
  wire not_new_n6697_;
  wire new_n3648_;
  wire not_new_n3982__0;
  wire not_new_n1067__7;
  wire not_new_n588__24010;
  wire not_new_n1583__490;
  wire not_new_n1581__2824752490;
  wire new_n9359_;
  wire not_new_n7077_;
  wire not_new_n3340_;
  wire not_new_n3248_;
  wire not_new_n989__6;
  wire new_n5488_;
  wire new_n6855_;
  wire new_n10341_;
  wire not_new_n4072__0;
  wire not_new_n7481_;
  wire not_pi265_3;
  wire new_n1805_;
  wire not_new_n9585_;
  wire new_n1815_;
  wire not_new_n1977_;
  wire new_n2483_;
  wire key_gate_1;
  wire not_new_n8074_;
  wire new_n4242_;
  wire new_n8457_;
  wire not_new_n589__225393402906922580878632490;
  wire po241;
  wire not_new_n586__9;
  wire new_n8137_;
  wire not_new_n4669_;
  wire new_n4912_;
  wire new_n1405_;
  wire or_not_new_n1159__0_not_new_n8794__0;
  wire not_new_n6613__3;
  wire new_n8251_;
  wire not_new_n7489_;
  wire not_new_n6937_;
  wire not_new_n6540__1;
  wire not_new_n2348_;
  wire new_n7026_;
  wire not_new_n10010_;
  wire key_gate_84;
  wire not_pi034_2;
  wire new_n9952_;
  wire new_n5405_;
  wire not_new_n9477_;
  wire new_n7965_;
  wire not_new_n4846_;
  wire not_new_n6906_;
  wire new_n4572_;
  wire not_new_n731_;
  wire not_new_n3929__0;
  wire and_new_n4405__new_n4330_;
  wire new_n4004_;
  wire new_n2306_;
  wire not_new_n10239_;
  wire new_n1184_;
  wire new_n3949_;
  wire not_new_n604__10;
  wire not_new_n9606_;
  wire new_n7759_;
  wire new_n3089_;
  wire not_new_n1398_;
  wire not_new_n4227_;
  wire not_new_n1208_;
  wire not_new_n4955_;
  wire not_new_n646__4;
  wire new_n4100_;
  wire new_n3092_;
  wire new_n6415_;
  wire new_n5476_;
  wire new_n6041_;
  wire not_new_n7648__2;
  wire new_n2871_;
  wire new_n6274_;
  wire new_n952_;
  wire new_n1755_;
  wire not_new_n6300_;
  wire new_n7013_;
  wire not_new_n7930_;
  wire not_new_n3856_;
  wire po222;
  wire new_n2246_;
  wire new_n6872_;
  wire not_new_n622__70;
  wire new_n8053_;
  wire new_n7622_;
  wire not_new_n4898__0;
  wire not_new_n8908_;
  wire not_new_n7113__2;
  wire new_n1346_;
  wire not_new_n1027__968890104070;
  wire new_n9045_;
  wire not_new_n6531__1;
  wire not_pi264_0;
  wire new_n3005_;
  wire and_and_new_n2325__new_n2332__new_n2333_;
  wire new_n7608_;
  wire not_new_n3383_;
  wire not_new_n8217_;
  wire new_n5210_;
  wire po295;
  wire not_new_n7752_;
  wire new_n8501_;
  wire po056;
  wire new_n4450_;
  wire not_new_n1601__797922662976120010;
  wire and_new_n2143__new_n2146_;
  wire new_n3680_;
  wire not_new_n3776_;
  wire not_new_n599__8;
  wire new_n6939_;
  wire not_new_n1037__113988951853731430;
  wire not_new_n4452_;
  wire not_new_n8296_;
  wire new_n2447_;
  wire not_new_n7830_;
  wire new_n5799_;
  wire new_n6743_;
  wire new_n8284_;
  wire not_new_n7230_;
  wire not_new_n7382_;
  wire new_n6052_;
  wire po122;
  wire not_new_n1728__3;
  wire new_n5532_;
  wire not_new_n1672_;
  wire not_new_n6248_;
  wire not_new_n1041__24010;
  wire new_n3078_;
  wire not_new_n5293_;
  wire new_n2673_;
  wire not_new_n1617_;
  wire not_new_n1047__403536070;
  wire new_n6238_;
  wire not_new_n5744_;
  wire not_pi166_1;
  wire not_new_n989__8235430;
  wire not_po298_10;
  wire not_new_n6443__1;
  wire not_new_n5559_;
  wire new_n2939_;
  wire new_n8569_;
  wire new_n3819_;
  wire not_new_n7679_;
  wire or_not_new_n1055__168070_not_new_n6325_;
  wire not_new_n3315__6;
  wire not_po298_9;
  wire or_or_or_not_pi269_1_not_pi260_1_not_pi257_1_not_pi248_1;
  wire new_n4348_;
  wire not_new_n581__16284135979104490;
  wire not_new_n607__5;
  wire not_new_n3946_;
  wire not_new_n629__403536070;
  wire new_n2072_;
  wire new_n9653_;
  wire new_n3095_;
  wire or_or_not_new_n2284__not_new_n2281__not_new_n2282_;
  wire new_n7690_;
  wire new_n4904_;
  wire new_n9257_;
  wire new_n1859_;
  wire new_n2217_;
  wire not_new_n5764__0;
  wire not_new_n3334_;
  wire not_new_n1554_;
  wire not_new_n1599__10;
  wire not_new_n1591_;
  wire not_new_n5662_;
  wire new_n7084_;
  wire not_new_n5426_;
  wire not_new_n1616__9;
  wire new_n2108_;
  wire not_new_n2842_;
  wire new_n5601_;
  wire not_po296_43181145673964365640352930977077280875522488490;
  wire new_n2096_;
  wire not_new_n4838_;
  wire not_new_n7342_;
  wire new_n3510_;
  wire new_n6880_;
  wire not_new_n7005__0;
  wire not_new_n5000__0;
  wire new_n6774_;
  wire not_new_n1598__10;
  wire not_new_n1067__24010;
  wire not_new_n9782_;
  wire new_n5956_;
  wire not_new_n8877_;
  wire or_not_new_n1555__not_new_n2434_;
  wire not_new_n617__403536070;
  wire new_n2039_;
  wire new_n2398_;
  wire or_not_new_n6340__not_new_n6341_;
  wire new_n6597_;
  wire new_n1908_;
  wire not_new_n5446_;
  wire not_new_n8340__0;
  wire new_n2032_;
  wire not_new_n1378_;
  wire new_n3817_;
  wire new_n947_;
  wire not_new_n8826_;
  wire new_n3631_;
  wire key_gate_98;
  wire not_new_n1551_;
  wire new_n6320_;
  wire not_new_n4914_;
  wire not_new_n7013__1;
  wire not_new_n4426__0;
  wire new_n8858_;
  wire not_new_n2072_;
  wire not_new_n8442_;
  wire new_n8354_;
  wire not_new_n5706__1;
  wire not_pi208;
  wire new_n7132_;
  wire not_new_n6193_;
  wire new_n6491_;
  wire not_new_n1010__0;
  wire new_n5657_;
  wire new_n3623_;
  wire not_new_n1037__8235430;
  wire or_or_not_new_n1271__not_new_n1269__not_new_n1983_;
  wire new_n10022_;
  wire new_n3102_;
  wire new_n2528_;
  wire new_n3620_;
  wire new_n8978_;
  wire or_or_not_new_n2091__not_new_n2092__not_new_n2094_;
  wire not_new_n1767_;
  wire not_new_n1580_;
  wire not_new_n8032_;
  wire not_new_n9282_;
  wire new_n1325_;
  wire new_n7161_;
  wire not_new_n6601_;
  wire not_new_n1605__2;
  wire not_new_n4165_;
  wire not_new_n6916_;
  wire new_n10032_;
  wire not_new_n589__168070;
  wire not_new_n3382_;
  wire not_new_n631__490;
  wire new_n4755_;
  wire new_n9749_;
  wire not_new_n4176_;
  wire not_new_n1018_;
  wire not_new_n10176_;
  wire new_n6758_;
  wire not_new_n5596_;
  wire new_n3590_;
  wire not_pi182_0;
  wire not_new_n3054_;
  wire new_n4769_;
  wire or_not_new_n2170__not_new_n2167_;
  wire new_n1526_;
  wire new_n6599_;
  wire new_n4959_;
  wire not_new_n3702_;
  wire new_n4611_;
  wire new_n9238_;
  wire new_n2131_;
  wire not_new_n1154_;
  wire new_n3460_;
  wire not_new_n1039__2326305139872070;
  wire not_new_n4827__1;
  wire not_new_n3956_;
  wire not_new_n8145_;
  wire new_n4795_;
  wire not_new_n581__6782230728490;
  wire new_n5830_;
  wire new_n2723_;
  wire not_po298_2;
  wire not_new_n3372__16284135979104490;
  wire or_or_not_new_n1787__not_new_n1788__not_new_n1790_;
  wire not_new_n4116__2;
  wire new_n3835_;
  wire new_n2853_;
  wire not_new_n8837__0;
  wire new_n1694_;
  wire new_n4458_;
  wire not_new_n8655_;
  wire not_new_n7702_;
  wire not_new_n1537__968890104070;
  wire not_new_n3310__6;
  wire not_new_n9964__0;
  wire key_gate_116;
  wire not_po296_1577753820348458066150427430;
  wire not_new_n4670_;
  wire not_new_n7574_;
  wire not_pi226;
  wire not_new_n8508_;
  wire new_n746_;
  wire not_new_n7440_;
  wire not_new_n5276_;
  wire not_new_n629__9;
  wire not_new_n3081_;
  wire not_new_n1065__8235430;
  wire new_n7870_;
  wire new_n4239_;
  wire not_new_n5365_;
  wire new_n5251_;
  wire not_new_n581__3119734822845423713013303218219760490;
  wire new_n8736_;
  wire not_new_n928__10;
  wire not_new_n629__5;
  wire not_new_n647__10;
  wire not_new_n1536__3;
  wire not_new_n1612_;
  wire not_new_n7638_;
  wire or_not_new_n3155__not_new_n3154_;
  wire not_new_n5813__0;
  wire not_new_n7895_;
  wire not_new_n602__0;
  wire new_n8929_;
  wire new_n5538_;
  wire new_n4962_;
  wire not_new_n993_;
  wire po180;
  wire not_new_n724_;
  wire not_new_n9969__0;
  wire new_n6535_;
  wire not_new_n609__0;
  wire not_new_n4330_;
  wire new_n3394_;
  wire new_n3391_;
  wire not_new_n8606_;
  wire new_n1536_;
  wire not_new_n6521_;
  wire not_new_n1037__3;
  wire not_po296_125892552985318850263419623839875454447587430;
  wire not_new_n632__10;
  wire not_new_n8545_;
  wire new_n9336_;
  wire not_new_n1043__57648010;
  wire new_n8580_;
  wire not_new_n7451__1;
  wire not_new_n9454_;
  wire not_new_n6616_;
  wire not_new_n4260_;
  wire new_n4109_;
  wire not_new_n9059__0;
  wire not_new_n1622_;
  wire not_new_n5078__1;
  wire not_new_n4343_;
  wire not_new_n639__47475615099430;
  wire not_new_n7358_;
  wire new_n4925_;
  wire not_pi133_0;
  wire new_n1297_;
  wire new_n7242_;
  wire not_new_n4987__0;
  wire not_new_n5568_;
  wire not_new_n6984__0;
  wire not_new_n6633__1;
  wire not_new_n5701_;
  wire new_n6714_;
  wire not_new_n1023_;
  wire not_new_n10110_;
  wire not_new_n3232_;
  wire new_n2201_;
  wire new_n10117_;
  wire not_pi064_5;
  wire not_new_n3361_;
  wire not_new_n9906__0;
  wire not_new_n8233_;
  wire not_new_n9124_;
  wire not_new_n1714_;
  wire not_new_n1615__0;
  wire not_new_n3985_;
  wire not_new_n9344_;
  wire new_n5982_;
  wire not_new_n6187_;
  wire new_n6665_;
  wire not_new_n5189_;
  wire not_new_n7936_;
  wire new_n7379_;
  wire not_new_n994__19773267430;
  wire not_new_n4902_;
  wire and_new_n4974__new_n5376_;
  wire not_new_n9544_;
  wire new_n9758_;
  wire not_new_n598__0;
  wire not_new_n5000_;
  wire new_n4302_;
  wire new_n8967_;
  wire not_new_n4692_;
  wire not_new_n10208_;
  wire new_n1382_;
  wire new_n5277_;
  wire new_n6571_;
  wire not_new_n630__57648010;
  wire new_n5469_;
  wire not_new_n7606_;
  wire new_n4606_;
  wire new_n6007_;
  wire not_new_n3311__0;
  wire not_new_n7035__0;
  wire po074;
  wire new_n7134_;
  wire not_new_n1045__0;
  wire new_n4319_;
  wire not_new_n7013_;
  wire new_n6450_;
  wire not_new_n9811_;
  wire not_new_n775__2;
  wire key_gate_11;
  wire not_new_n4106_;
  wire not_new_n7940_;
  wire new_n727_;
  wire or_or_or_not_new_n2497__not_new_n1568__not_new_n2498__not_new_n2500_;
  wire new_n5996_;
  wire new_n3729_;
  wire new_n7221_;
  wire not_new_n10273_;
  wire not_pi024;
  wire not_new_n1069__57648010;
  wire not_new_n630__332329305696010;
  wire new_n7031_;
  wire not_new_n10071_;
  wire not_new_n2835_;
  wire not_new_n7106_;
  wire new_n8420_;
  wire new_n3478_;
  wire not_new_n7422_;
  wire new_n8871_;
  wire not_new_n625__490;
  wire new_n6457_;
  wire not_new_n7320_;
  wire new_n6396_;
  wire not_new_n4126__1;
  wire new_n5738_;
  wire not_new_n6631_;
  wire new_n2839_;
  wire new_n2261_;
  wire new_n7041_;
  wire not_new_n610__1176490;
  wire new_n8890_;
  wire new_n7478_;
  wire po262;
  wire new_n9964_;
  wire not_new_n4810_;
  wire new_n3614_;
  wire not_new_n593__6;
  wire new_n2641_;
  wire new_n9295_;
  wire and_new_n2067__new_n2070_;
  wire new_n5553_;
  wire new_n9826_;
  wire not_new_n6698_;
  wire new_n7532_;
  wire po137;
  wire not_new_n1601__273687473400809163430;
  wire not_new_n6458_;
  wire not_new_n2936_;
  wire new_n1941_;
  wire new_n4019_;
  wire po158;
  wire new_n6175_;
  wire not_new_n1436_;
  wire not_new_n10129_;
  wire new_n6628_;
  wire new_n5384_;
  wire new_n1677_;
  wire not_pi157;
  wire new_n4067_;
  wire not_new_n1611__47475615099430;
  wire new_n9656_;
  wire not_new_n641__138412872010;
  wire not_new_n8130_;
  wire new_n2009_;
  wire new_n1744_;
  wire not_new_n10234_;
  wire not_new_n10043_;
  wire not_new_n8844_;
  wire not_new_n3942_;
  wire not_new_n6974__2326305139872070;
  wire not_pi018;
  wire not_new_n9443_;
  wire not_new_n1603__6;
  wire not_new_n2613_;
  wire not_pi064_2824752490;
  wire not_new_n1057__2824752490;
  wire new_n8815_;
  wire new_n1789_;
  wire not_new_n1563_;
  wire new_n8870_;
  wire not_new_n6206_;
  wire not_new_n1390_;
  wire not_new_n1014_;
  wire new_n3935_;
  wire not_new_n2788_;
  wire not_new_n1596__8235430;
  wire not_new_n607__3;
  wire po296;
  wire not_new_n8781_;
  wire new_n4097_;
  wire po038;
  wire not_new_n9085_;
  wire not_new_n4461__0;
  wire new_n5792_;
  wire not_new_n6346_;
  wire new_n2946_;
  wire new_n9469_;
  wire not_new_n9028_;
  wire new_n6814_;
  wire new_n5107_;
  wire not_new_n8154__0;
  wire not_pi250_1;
  wire new_n10188_;
  wire new_n3219_;
  wire new_n2411_;
  wire new_n6417_;
  wire not_new_n9888__0;
  wire new_n3325_;
  wire new_n5228_;
  wire or_or_not_new_n9893__not_new_n9890__0_not_new_n10266_;
  wire not_new_n9964_;
  wire not_new_n644__8235430;
  wire new_n9751_;
  wire new_n3162_;
  wire not_new_n7650_;
  wire new_n7815_;
  wire not_new_n1158__1;
  wire not_new_n949_;
  wire not_new_n596__490;
  wire not_new_n1538__113988951853731430;
  wire new_n6229_;
  wire not_new_n5562_;
  wire not_new_n8999_;
  wire not_new_n9687_;
  wire not_new_n1216_;
  wire not_new_n5748_;
  wire not_new_n1291_;
  wire new_n7133_;
  wire new_n1678_;
  wire new_n7891_;
  wire new_n5185_;
  wire not_new_n7536_;
  wire new_n1210_;
  wire not_pi036_2;
  wire new_n9961_;
  wire new_n2071_;
  wire po091;
  wire not_new_n7640_;
  wire new_n8630_;
  wire new_n9273_;
  wire new_n5302_;
  wire not_new_n1055__24010;
  wire new_n3388_;
  wire not_new_n10219_;
  wire new_n5789_;
  wire new_n3992_;
  wire not_new_n4467__0;
  wire not_new_n6613_;
  wire not_new_n3681_;
  wire not_new_n1002__1;
  wire not_new_n994_;
  wire not_new_n6232__2;
  wire not_new_n586__8235430;
  wire not_new_n4133__1;
  wire and_new_n3315__new_n923_;
  wire new_n10222_;
  wire new_n9115_;
  wire po140;
  wire not_new_n606__168070;
  wire not_new_n1069__8;
  wire new_n2688_;
  wire not_new_n1615_;
  wire or_or_or_not_new_n6226__not_new_n6323__not_new_n6324__not_new_n6242_;
  wire not_new_n1536__70;
  wire new_n3942_;
  wire not_new_n1018__2;
  wire new_n8333_;
  wire not_new_n1061__4;
  wire not_new_n5416_;
  wire not_new_n6633__0;
  wire not_new_n7000_;
  wire not_new_n7645__0;
  wire not_new_n1063__332329305696010;
  wire not_new_n5195__0;
  wire not_new_n8561_;
  wire not_new_n2785_;
  wire new_n2817_;
  wire not_new_n8924_;
  wire new_n8418_;
  wire not_new_n628__5;
  wire not_new_n3437_;
  wire new_n8742_;
  wire not_new_n9963__0;
  wire not_new_n9193_;
  wire new_n3931_;
  wire not_new_n3579_;
  wire new_n2963_;
  wire or_or_not_new_n2776__not_new_n2779__not_new_n2778_;
  wire new_n1573_;
  wire not_pi177_2;
  wire new_n1438_;
  wire not_new_n607__6;
  wire po040;
  wire new_n9490_;
  wire new_n6775_;
  wire not_new_n7112_;
  wire new_n2676_;
  wire not_new_n7669_;
  wire new_n1266_;
  wire new_n5229_;
  wire not_new_n600__968890104070;
  wire new_n6494_;
  wire new_n8833_;
  wire not_new_n598__403536070;
  wire not_new_n1862_;
  wire new_n4581_;
  wire new_n4117_;
  wire key_gate_39;
  wire new_n1773_;
  wire new_n7626_;
  wire not_new_n1293_;
  wire not_pi158;
  wire new_n2301_;
  wire not_po298_6;
  wire new_n1592_;
  wire not_new_n638__10;
  wire not_new_n4071__0;
  wire new_n9376_;
  wire new_n6578_;
  wire not_new_n586__70;
  wire new_n6483_;
  wire not_pi014_0;
  wire new_n2985_;
  wire not_new_n4447__0;
  wire not_new_n4001_;
  wire not_new_n9024_;
  wire not_new_n6135_;
  wire not_new_n10317_;
  wire not_new_n1602__6;
  wire not_new_n946_;
  wire not_new_n5750__0;
  wire not_new_n4161__1;
  wire not_new_n1613_;
  wire not_new_n9983_;
  wire new_n3378_;
  wire not_new_n7387_;
  wire not_new_n7588_;
  wire not_new_n4216_;
  wire not_new_n598__2326305139872070;
  wire not_new_n10191_;
  wire po272;
  wire not_new_n6974__3;
  wire not_new_n581__70;
  wire not_new_n1047__8235430;
  wire new_n4415_;
  wire and_new_n1745__new_n1744_;
  wire not_new_n6486_;
  wire not_new_n593__8;
  wire po287;
  wire new_n8255_;
  wire not_new_n8819_;
  wire not_new_n5449_;
  wire not_new_n4469_;
  wire new_n8932_;
  wire new_n6316_;
  wire new_n10139_;
  wire not_new_n631__8;
  wire new_n9886_;
  wire new_n4552_;
  wire new_n9236_;
  wire not_new_n1536__138412872010;
  wire or_not_new_n1546__not_new_n1362_;
  wire not_pi269_2;
  wire not_new_n1391_;
  wire not_new_n639__7;
  wire new_n2391_;
  wire not_new_n6566_;
  wire new_n8819_;
  wire not_new_n3199_;
  wire new_n1767_;
  wire not_new_n3185__168070;
  wire new_n6600_;
  wire not_new_n8811_;
  wire new_n5465_;
  wire not_new_n1596__6782230728490;
  wire new_n4180_;
  wire not_new_n9683_;
  wire new_n6551_;
  wire not_new_n621__1;
  wire new_n2412_;
  wire key_gate_25;
  wire not_new_n629_;
  wire not_new_n5668_;
  wire new_n3415_;
  wire not_new_n3974_;
  wire not_new_n6443__7;
  wire new_n6640_;
  wire not_new_n8473_;
  wire not_new_n3332_;
  wire new_n10293_;
  wire not_new_n583_;
  wire not_new_n10147_;
  wire new_n8472_;
  wire not_new_n8162__2;
  wire new_n5015_;
  wire new_n4261_;
  wire new_n6152_;
  wire new_n6314_;
  wire new_n3584_;
  wire new_n4726_;
  wire not_new_n8596__2;
  wire not_new_n3384__0;
  wire new_n6197_;
  wire not_new_n6804_;
  wire not_new_n9500_;
  wire not_new_n8213_;
  wire not_new_n8659_;
  wire not_new_n8322_;
  wire new_n6722_;
  wire not_new_n1039__9;
  wire not_new_n636__70;
  wire not_new_n3565_;
  wire not_new_n8981_;
  wire not_new_n5454_;
  wire not_new_n4699_;
  wire new_n7843_;
  wire not_new_n9630_;
  wire new_n3976_;
  wire new_n10120_;
  wire not_new_n1631__8235430;
  wire new_n7683_;
  wire not_new_n7627__0;
  wire new_n4677_;
  wire new_n3337_;
  wire new_n7270_;
  wire not_new_n1059__968890104070;
  wire not_new_n7897_;
  wire new_n9020_;
  wire or_not_new_n2091__not_new_n2092_;
  wire new_n6699_;
  wire new_n5132_;
  wire and_new_n2627__new_n2628_;
  wire po055;
  wire not_new_n9594__0;
  wire not_new_n3736_;
  wire new_n2728_;
  wire new_n4931_;
  wire not_new_n4443__0;
  wire new_n9924_;
  wire not_new_n8376__0;
  wire not_pi112_0;
  wire not_new_n4994_;
  wire new_n2558_;
  wire new_n4404_;
  wire new_n3224_;
  wire new_n10076_;
  wire new_n935_;
  wire new_n1569_;
  wire not_new_n4228_;
  wire new_n8161_;
  wire not_new_n4812_;
  wire not_new_n9771_;
  wire not_new_n8583_;
  wire not_new_n1063__1;
  wire not_new_n4465_;
  wire not_new_n9931_;
  wire new_n1506_;
  wire not_new_n611_;
  wire new_n3339_;
  wire not_new_n640__1;
  wire not_new_n5753__0;
  wire not_new_n5928__0;
  wire not_new_n4985__0;
  wire not_new_n6755_;
  wire not_new_n1327_;
  wire not_new_n4984__1;
  wire new_n8533_;
  wire new_n3238_;
  wire new_n4508_;
  wire not_new_n6415_;
  wire not_new_n4197_;
  wire not_new_n1039__2824752490;
  wire new_n4817_;
  wire not_new_n8089_;
  wire not_new_n3878_;
  wire not_new_n3928_;
  wire or_or_not_new_n6240__not_new_n6330__not_new_n6331_;
  wire not_new_n6443__9;
  wire not_new_n7010__0;
  wire not_new_n1061__70;
  wire new_n5639_;
  wire not_new_n7614__0;
  wire new_n6785_;
  wire new_n4534_;
  wire new_n3875_;
  wire not_new_n8965_;
  wire not_new_n8392_;
  wire new_n2872_;
  wire not_new_n1037__138412872010;
  wire new_n5098_;
  wire not_new_n999_;
  wire not_new_n5802_;
  wire new_n8198_;
  wire not_pi034_1;
  wire not_new_n628__1176490;
  wire new_n664_;
  wire not_pi162;
  wire new_n6682_;
  wire not_new_n2035_;
  wire not_new_n775__7;
  wire new_n3340_;
  wire new_n6710_;
  wire not_new_n7139__0;
  wire new_n6395_;
  wire new_n2867_;
  wire not_new_n2494_;
  wire new_n7766_;
  wire not_new_n3691_;
  wire new_n2955_;
  wire not_new_n8930_;
  wire not_new_n9383_;
  wire not_new_n8288_;
  wire not_new_n589__7490483309651862334944941026945644936490;
  wire not_new_n7715_;
  wire key_gate_48;
  wire not_new_n5479__0;
  wire not_new_n1013__7;
  wire not_new_n602__168070;
  wire new_n3921_;
  wire not_new_n1588__3430;
  wire not_new_n1588__8235430;
  wire not_new_n1612__403536070;
  wire new_n9544_;
  wire not_new_n1397_;
  wire not_new_n1589__2;
  wire new_n3067_;
  wire not_new_n922__0;
  wire new_n4699_;
  wire not_new_n9056__0;
  wire new_n5416_;
  wire not_new_n3819_;
  wire new_n7148_;
  wire not_new_n8499_;
  wire new_n8702_;
  wire not_new_n984__168070;
  wire new_n2054_;
  wire new_n4775_;
  wire not_new_n3087_;
  wire not_new_n9216_;
  wire new_n9797_;
  wire not_new_n9965__0;
  wire not_new_n8423_;
  wire not_new_n631__138412872010;
  wire new_n8868_;
  wire not_new_n5280_;
  wire new_n3897_;
  wire not_new_n5269_;
  wire not_po296_2326305139872070;
  wire not_new_n586__797922662976120010;
  wire not_new_n9926__0;
  wire new_n9471_;
  wire not_pi250_3;
  wire not_new_n8141__0;
  wire not_new_n6615_;
  wire new_n4651_;
  wire not_new_n1612__8;
  wire not_new_n3185__403536070;
  wire not_new_n7754__3;
  wire not_new_n9982_;
  wire new_n5278_;
  wire new_n8623_;
  wire not_new_n1065__6;
  wire not_new_n1432_;
  wire not_new_n2825_;
  wire new_n7434_;
  wire new_n8653_;
  wire new_n1167_;
  wire new_n4885_;
  wire new_n8604_;
  wire not_new_n7663__1;
  wire new_n1161_;
  wire not_new_n7643_;
  wire not_new_n2185__0;
  wire not_new_n968_;
  wire not_pi020_0;
  wire new_n8594_;
  wire not_new_n6499__0;
  wire new_n5191_;
  wire not_new_n635__968890104070;
  wire not_new_n6689_;
  wire not_new_n1787_;
  wire not_new_n7845_;
  wire not_new_n626__13410686196639649008070;
  wire not_new_n7678_;
  wire not_new_n10257_;
  wire not_new_n7020_;
  wire not_new_n8134_;
  wire not_new_n3918_;
  wire not_new_n9754_;
  wire or_or_not_new_n1283__not_new_n1281__not_new_n2040_;
  wire new_n4252_;
  wire not_new_n5767__2;
  wire not_new_n645__70;
  wire new_n4264_;
  wire new_n1668_;
  wire not_new_n3321_;
  wire not_new_n4829__0;
  wire not_new_n7074_;
  wire not_new_n10003_;
  wire po291;
  wire new_n5370_;
  wire new_n4295_;
  wire not_new_n589__1299348114471230201171721456984490;
  wire new_n3762_;
  wire not_new_n5791__2;
  wire new_n6946_;
  wire not_new_n1009__0;
  wire or_or_not_new_n2740__not_new_n2743__not_new_n2742_;
  wire or_not_new_n5266__not_new_n5206_;
  wire new_n7992_;
  wire not_new_n5862_;
  wire not_new_n3678_;
  wire not_new_n1536__9;
  wire not_new_n596__0;
  wire not_new_n1396_;
  wire not_new_n4705_;
  wire not_new_n9106_;
  wire new_n8012_;
  wire not_new_n1612__2326305139872070;
  wire not_new_n1041__1;
  wire not_new_n4119_;
  wire or_or_not_new_n1939__not_new_n1940__not_new_n1942_;
  wire not_new_n4128__1;
  wire not_new_n5702_;
  wire new_n8061_;
  wire not_new_n1035__1176490;
  wire new_n8242_;
  wire not_new_n624__1;
  wire not_new_n1534__10;
  wire not_new_n1069__138412872010;
  wire new_n7879_;
  wire new_n3586_;
  wire not_new_n594__8;
  wire not_new_n2300_;
  wire new_n5186_;
  wire not_new_n7080_;
  wire new_n6251_;
  wire not_new_n7009_;
  wire and_new_n2404__new_n2403_;
  wire not_new_n8481_;
  wire not_new_n775__3430;
  wire and_new_n1460__new_n1466_;
  wire not_new_n4427__0;
  wire not_new_n7339_;
  wire not_new_n1583__9;
  wire not_new_n9141_;
  wire not_new_n7771_;
  wire not_new_n1943_;
  wire not_new_n6531__0;
  wire not_new_n602__3430;
  wire new_n7749_;
  wire not_new_n2128__0;
  wire not_new_n8182_;
  wire new_n6187_;
  wire new_n9534_;
  wire not_new_n1591__9;
  wire not_new_n5301_;
  wire key_gate_97;
  wire not_new_n3553_;
  wire new_n4936_;
  wire new_n5927_;
  wire not_new_n8985_;
  wire new_n5363_;
  wire new_n6042_;
  wire new_n4487_;
  wire not_new_n596__47475615099430;
  wire not_new_n8355_;
  wire not_new_n7357__0;
  wire not_new_n9385__0;
  wire new_n2002_;
  wire new_n10157_;
  wire not_new_n10018__0;
  wire not_new_n3315__3430;
  wire new_n7076_;
  wire not_new_n1600__332329305696010;
  wire not_new_n4789_;
  wire new_n3470_;
  wire new_n3915_;
  wire not_po296_12197604876358357001385738625629718207556152941312384010;
  wire new_n5970_;
  wire new_n2984_;
  wire not_new_n7126_;
  wire not_new_n9129_;
  wire not_new_n1043__2824752490;
  wire new_n1531_;
  wire new_n2452_;
  wire new_n3495_;
  wire new_n1840_;
  wire new_n9301_;
  wire not_new_n8242_;
  wire new_n3621_;
  wire not_new_n2847_;
  wire not_new_n10165_;
  wire not_new_n5206_;
  wire not_new_n618__47475615099430;
  wire not_pi167_2;
  wire not_pi061_2;
  wire new_n3816_;
  wire not_new_n1055__6782230728490;
  wire new_n3646_;
  wire new_n2862_;
  wire not_new_n643__3;
  wire not_new_n1604__3;
  wire not_new_n3679_;
  wire po002;
  wire not_new_n625__797922662976120010;
  wire not_new_n4656_;
  wire not_new_n1049__1;
  wire not_new_n1049__968890104070;
  wire not_new_n632__2326305139872070;
  wire not_new_n4121__0;
  wire new_n8866_;
  wire new_n8817_;
  wire not_new_n631__5585458640832840070;
  wire not_new_n9455_;
  wire not_new_n4979__0;
  wire not_new_n2893_;
  wire not_new_n2711_;
  wire new_n8789_;
  wire not_pi064_19773267430;
  wire not_new_n9543_;
  wire new_n7810_;
  wire not_new_n9475_;
  wire not_new_n5794__0;
  wire not_new_n9425_;
  wire not_pi248_0;
  wire new_n4916_;
  wire not_new_n9691_;
  wire not_pi064_4;
  wire not_new_n1043__4;
  wire not_new_n6232__5;
  wire new_n8661_;
  wire not_new_n2939_;
  wire not_new_n622__8235430;
  wire not_new_n1421_;
  wire po234;
  wire not_new_n628__6;
  wire new_n9215_;
  wire not_new_n8872_;
  wire not_new_n6232__4;
  wire new_n4515_;
  wire not_new_n6825_;
  wire not_new_n8864_;
  wire new_n4728_;
  wire not_new_n7638__0;
  wire new_n3818_;
  wire new_n5525_;
  wire new_n2843_;
  wire new_n6652_;
  wire not_new_n645__10;
  wire not_new_n5456__0;
  wire new_n9438_;
  wire not_new_n7797_;
  wire not_new_n638_;
  wire new_n4877_;
  wire not_new_n1862__0;
  wire po113;
  wire new_n734_;
  wire new_n6700_;
  wire new_n4562_;
  wire not_new_n4210_;
  wire not_new_n10044_;
  wire not_new_n10242_;
  wire new_n6960_;
  wire not_new_n4577_;
  wire not_new_n4956_;
  wire new_n5937_;
  wire not_pi053_2;
  wire not_new_n3178_;
  wire not_new_n5458__0;
  wire not_new_n10318_;
  wire not_new_n3917_;
  wire new_n2865_;
  wire not_new_n1883_;
  wire new_n1658_;
  wire not_new_n2351_;
  wire new_n8964_;
  wire new_n9434_;
  wire not_new_n6798_;
  wire not_new_n1039__10;
  wire not_pi262_0;
  wire not_new_n1037__5;
  wire new_n8897_;
  wire new_n3801_;
  wire new_n1413_;
  wire new_n2981_;
  wire not_new_n1613__7;
  wire not_new_n3787_;
  wire new_n4053_;
  wire not_pi178_0;
  wire not_po298;
  wire not_new_n9082__0;
  wire not_new_n3925__0;
  wire not_new_n9612_;
  wire not_pi129_0;
  wire not_pi121_0;
  wire not_new_n9512__2;
  wire not_new_n1536__403536070;
  wire not_new_n5749__2;
  wire not_new_n8595__1;
  wire not_new_n1538__4;
  wire not_new_n7789_;
  wire new_n5315_;
  wire not_new_n3895_;
  wire new_n8345_;
  wire not_new_n599__6782230728490;
  wire not_new_n648__3;
  wire not_new_n1624_;
  wire not_new_n619__8;
  wire new_n3202_;
  wire not_pi135_2;
  wire not_new_n6473__1;
  wire not_new_n9269_;
  wire new_n1309_;
  wire new_n2297_;
  wire not_new_n8954_;
  wire not_pi171_3;
  wire new_n7635_;
  wire new_n9897_;
  wire new_n8401_;
  wire and_and_not_pi056_1_not_pi055_1_not_pi054_1;
  wire not_pi042_0;
  wire not_new_n1537__168070;
  wire not_new_n1055__2824752490;
  wire not_new_n6476_;
  wire not_new_n8107_;
  wire not_new_n7569_;
  wire new_n4896_;
  wire not_new_n1534__5;
  wire new_n1938_;
  wire not_new_n9087_;
  wire not_new_n8689_;
  wire not_new_n6286_;
  wire po150;
  wire not_new_n3131_;
  wire new_n938_;
  wire not_new_n8502_;
  wire not_new_n7675_;
  wire not_new_n1053__3430;
  wire not_po296_85383234134508499009700170379408027452893070589186688070;
  wire not_new_n6620__0;
  wire po251;
  wire not_pi071;
  wire new_n10146_;
  wire not_new_n3840_;
  wire not_new_n8552_;
  wire not_new_n726__0;
  wire new_n1358_;
  wire not_new_n4509_;
  wire not_new_n635__3;
  wire not_new_n9379_;
  wire not_new_n928__332329305696010;
  wire not_new_n1888_;
  wire not_new_n1061__6782230728490;
  wire not_new_n7691_;
  wire new_n4738_;
  wire not_new_n1012__4;
  wire new_n2119_;
  wire not_new_n1061__47475615099430;
  wire not_new_n10192_;
  wire not_new_n7648__1;
  wire not_po296_52433383167563036344614587188619514555430;
  wire not_new_n8879_;
  wire not_new_n7288_;
  wire new_n7663_;
  wire new_n6839_;
  wire new_n2367_;
  wire new_n6479_;
  wire not_new_n7938_;
  wire not_new_n1599__6;
  wire not_new_n1606__4;
  wire new_n5222_;
  wire not_new_n631__93874803376477543056490;
  wire new_n7822_;
  wire new_n8049_;
  wire new_n3883_;
  wire not_new_n3475_;
  wire new_n8718_;
  wire not_new_n2615_;
  wire new_n3499_;
  wire not_new_n4102_;
  wire not_pi259_0;
  wire not_new_n638__225393402906922580878632490;
  wire not_new_n7362_;
  wire po298;
  wire not_new_n4827__0;
  wire new_n2660_;
  wire new_n3913_;
  wire not_new_n4957__0;
  wire new_n8557_;
  wire not_new_n627__7;
  wire new_n3794_;
  wire not_new_n6497__0;
  wire not_new_n636__7;
  wire new_n4509_;
  wire not_new_n1728__10;
  wire new_n4920_;
  wire not_new_n7827__0;
  wire not_new_n1317_;
  wire not_new_n3791_;
  wire new_n5807_;
  wire new_n3318_;
  wire not_pi255_3;
  wire not_new_n1903_;
  wire not_new_n600__2;
  wire not_new_n6641_;
  wire not_new_n7990_;
  wire not_new_n6974__3430;
  wire not_new_n7831_;
  wire not_new_n612__2;
  wire not_new_n8910_;
  wire not_new_n9243_;
  wire and_new_n6977__new_n7377_;
  wire not_new_n3286_;
  wire new_n8290_;
  wire not_new_n9862_;
  wire not_new_n8916_;
  wire new_n3674_;
  wire not_new_n1585__16284135979104490;
  wire not_new_n775__6782230728490;
  wire not_new_n9955__0;
  wire new_n6612_;
  wire not_new_n9422_;
  wire not_new_n593__47475615099430;
  wire not_pi037_1;
  wire not_new_n4959__0;
  wire not_new_n8151_;
  wire not_new_n5686__0;
  wire new_n5354_;
  wire new_n8710_;
  wire not_new_n628__273687473400809163430;
  wire not_new_n4990_;
  wire not_new_n4841__1;
  wire new_n741_;
  wire not_new_n4728_;
  wire new_n6671_;
  wire not_new_n5876_;
  wire not_new_n2988_;
  wire not_new_n8239_;
  wire not_pi135_1;
  wire not_new_n602__57648010;
  wire not_new_n1536__4;
  wire not_new_n3185__968890104070;
  wire new_n8403_;
  wire not_new_n4932_;
  wire not_new_n6635__4;
  wire not_new_n5316_;
  wire new_n5580_;
  wire not_new_n633__7;
  wire not_new_n742_;
  wire not_new_n6448_;
  wire new_n1634_;
  wire not_new_n9415_;
  wire new_n8373_;
  wire new_n9953_;
  wire not_new_n5480_;
  wire not_new_n634__57648010;
  wire new_n7229_;
  wire not_pi011;
  wire new_n5169_;
  wire not_new_n5826_;
  wire not_new_n10032_;
  wire new_n9352_;
  wire not_new_n7775_;
  wire new_n4461_;
  wire not_new_n3253_;
  wire not_new_n8276_;
  wire new_n2876_;
  wire not_new_n3186_;
  wire not_new_n983_;
  wire not_new_n599__1;
  wire not_new_n588__5;
  wire new_n2637_;
  wire new_n7127_;
  wire new_n2495_;
  wire not_new_n603__4;
  wire not_new_n10135_;
  wire not_new_n6981__0;
  wire not_new_n8012_;
  wire not_pi251;
  wire not_new_n1768__0;
  wire new_n7205_;
  wire not_new_n9406__0;
  wire key_gate_82;
  wire not_new_n3745_;
  wire new_n5083_;
  wire and_new_n2998__new_n998_;
  wire new_n8908_;
  wire new_n7588_;
  wire new_n748_;
  wire new_n4873_;
  wire not_new_n1069__7;
  wire new_n7473_;
  wire new_n5307_;
  wire not_new_n9302_;
  wire not_new_n643__8;
  wire new_n5907_;
  wire new_n4251_;
  wire not_new_n7754__0;
  wire and_new_n8104__new_n8464_;
  wire not_new_n8436_;
  wire not_new_n6483_;
  wire not_new_n5132_;
  wire new_n1771_;
  wire not_new_n3092_;
  wire not_new_n9541__0;
  wire or_not_new_n4410__not_new_n609_;
  wire not_new_n7694_;
  wire and_new_n5082__new_n5423_;
  wire new_n1819_;
  wire not_new_n3268_;
  wire not_new_n5974__0;
  wire not_new_n8292_;
  wire not_new_n1583__403536070;
  wire not_new_n4463__0;
  wire new_n7342_;
  wire new_n8837_;
  wire not_new_n4474_;
  wire new_n2697_;
  wire not_new_n1534__3;
  wire new_n8460_;
  wire new_n2866_;
  wire new_n3548_;
  wire not_pi256_1;
  wire new_n7259_;
  wire not_new_n3329_;
  wire new_n2112_;
  wire and_new_n6373__new_n6254_;
  wire new_n2312_;
  wire not_new_n594__9;
  wire new_n9040_;
  wire new_n7947_;
  wire not_new_n9105_;
  wire not_new_n7596_;
  wire not_new_n4126_;
  wire new_n1871_;
  wire not_new_n9461_;
  wire not_new_n2942_;
  wire new_n3930_;
  wire not_new_n6474__0;
  wire not_new_n1584__47475615099430;
  wire not_new_n5113__0;
  wire new_n9626_;
  wire or_not_new_n1243__not_new_n1241_;
  wire new_n7974_;
  wire new_n2010_;
  wire not_new_n625__4599865365447399609768010;
  wire new_n5074_;
  wire not_new_n1071__9;
  wire not_new_n3369__0;
  wire not_new_n597__2326305139872070;
  wire not_new_n1728__113988951853731430;
  wire new_n2947_;
  wire not_pi134;
  wire not_new_n2751_;
  wire not_new_n5739_;
  wire new_n6172_;
  wire not_new_n4997_;
  wire not_new_n10259_;
  wire new_n1326_;
  wire not_new_n4016_;
  wire or_not_new_n1267__not_new_n1265_;
  wire not_new_n3367_;
  wire new_n9418_;
  wire not_new_n9904_;
  wire not_new_n8094_;
  wire not_new_n7109__1;
  wire not_new_n3182__0;
  wire not_new_n6895_;
  wire not_new_n4633_;
  wire not_new_n4122__1;
  wire not_new_n648__490;
  wire new_n9563_;
  wire not_new_n1594__490;
  wire not_new_n2242__0;
  wire not_new_n595__4;
  wire not_new_n7146__1;
  wire new_n3997_;
  wire not_new_n5608_;
  wire not_new_n10225_;
  wire not_new_n4231_;
  wire new_n4140_;
  wire not_pi239;
  wire new_n703_;
  wire new_n9082_;
  wire not_new_n3489_;
  wire not_new_n2664_;
  wire not_new_n957_;
  wire new_n2249_;
  wire not_pi142_0;
  wire not_new_n4014__2;
  wire not_new_n9882_;
  wire new_n1277_;
  wire not_new_n9188_;
  wire not_new_n730_;
  wire new_n6621_;
  wire not_new_n3311__4;
  wire not_new_n1631__47475615099430;
  wire new_n2429_;
  wire not_new_n9610__0;
  wire new_n5561_;
  wire not_new_n1604__490;
  wire not_new_n631__225393402906922580878632490;
  wire not_new_n1584__5;
  wire not_new_n9430_;
  wire new_n9874_;
  wire new_n3710_;
  wire not_new_n643__968890104070;
  wire not_new_n5306_;
  wire not_new_n1003_;
  wire not_new_n6541__1;
  wire and_and_not_pi044_1_not_pi043_1_not_pi046_1;
  wire new_n5804_;
  wire not_new_n1580__4;
  wire new_n8906_;
  wire not_new_n7433__0;
  wire or_not_new_n5441__not_new_n5617__1;
  wire new_n4077_;
  wire not_new_n4456_;
  wire not_new_n1013__6;
  wire not_new_n7945_;
  wire not_new_n585__7;
  wire new_n6911_;
  wire not_new_n6469_;
  wire not_new_n7185_;
  wire new_n9675_;
  wire not_new_n6217_;
  wire or_not_new_n649__0_not_new_n4287_;
  wire not_new_n628__7;
  wire new_n5172_;
  wire not_new_n1069__6782230728490;
  wire new_n1630_;
  wire not_new_n3394_;
  wire not_pi085;
  wire not_new_n7600_;
  wire not_new_n9343_;
  wire po257;
  wire not_new_n6211_;
  wire not_new_n600__7;
  wire not_new_n1004__3;
  wire new_n1492_;
  wire new_n2755_;
  wire not_pi174_3;
  wire not_new_n4272_;
  wire new_n3360_;
  wire not_new_n6500_;
  wire not_new_n4546_;
  wire new_n7954_;
  wire not_new_n5350_;
  wire not_new_n1239_;
  wire new_n3513_;
  wire not_new_n7656__0;
  wire new_n4323_;
  wire new_n6575_;
  wire new_n6787_;
  wire not_new_n4287_;
  wire not_new_n6999__0;
  wire new_n1362_;
  wire not_new_n984__47475615099430;
  wire not_new_n928__3430;
  wire not_new_n596__332329305696010;
  wire not_new_n8842_;
  wire not_po298_968890104070;
  wire not_new_n9010_;
  wire new_n4756_;
  wire new_n2896_;
  wire not_new_n7429_;
  wire not_new_n627__8;
  wire not_new_n3582_;
  wire new_n8541_;
  wire and_new_n1322__new_n2236_;
  wire new_n2164_;
  wire not_new_n7427_;
  wire not_new_n7024__0;
  wire not_new_n4498_;
  wire not_new_n8123__0;
  wire not_new_n3491_;
  wire new_n1690_;
  wire not_pi098;
  wire new_n8294_;
  wire new_n4390_;
  wire new_n7383_;
  wire new_n8901_;
  wire new_n9122_;
  wire not_new_n4412_;
  wire new_n9217_;
  wire not_new_n1049__1176490;
  wire new_n5145_;
  wire not_pi113;
  wire not_new_n4135_;
  wire not_pi125;
  wire not_new_n7184_;
  wire new_n7579_;
  wire not_new_n5570_;
  wire not_new_n1616__24010;
  wire not_new_n9986_;
  wire new_n4398_;
  wire not_new_n2865_;
  wire not_new_n7476_;
  wire not_new_n5197__0;
  wire new_n2533_;
  wire not_new_n7602__0;
  wire new_n10238_;
  wire new_n2927_;
  wire new_n3905_;
  wire new_n7614_;
  wire not_new_n7707_;
  wire not_new_n1581__16284135979104490;
  wire not_pi064_3430;
  wire new_n2247_;
  wire not_new_n1537__70;
  wire new_n8277_;
  wire not_new_n8823_;
  wire not_new_n589__1070069044235980333563563003849377848070;
  wire not_new_n5828_;
  wire not_new_n1045__968890104070;
  wire not_new_n3372__2824752490;
  wire or_not_new_n4461__not_new_n609__0;
  wire new_n6701_;
  wire not_pi126;
  wire or_or_not_new_n6226__not_new_n6323__not_new_n6324_;
  wire po239;
  wire not_new_n7609_;
  wire not_new_n6518__0;
  wire new_n4634_;
  wire new_n8916_;
  wire not_new_n5936_;
  wire not_new_n621__3430;
  wire not_new_n1603__9;
  wire new_n2386_;
  wire new_n1280_;
  wire not_new_n4433_;
  wire not_new_n1009__6;
  wire not_new_n1061__403536070;
  wire or_not_new_n3118__not_new_n3119_;
  wire not_new_n3184__403536070;
  wire not_new_n1023__0;
  wire not_new_n597__24010;
  wire not_new_n646__16284135979104490;
  wire not_new_n3183_;
  wire new_n8342_;
  wire not_new_n5343_;
  wire not_new_n8928_;
  wire new_n2511_;
  wire new_n5203_;
  wire new_n10080_;
  wire not_new_n5008_;
  wire new_n5041_;
  wire new_n4536_;
  wire not_new_n6503__0;
  wire not_new_n5107_;
  wire not_new_n6533_;
  wire new_n2607_;
  wire not_new_n8613_;
  wire not_new_n2566_;
  wire new_n8107_;
  wire not_new_n8865_;
  wire new_n1394_;
  wire not_new_n630__5;
  wire not_new_n6405_;
  wire not_new_n6952_;
  wire new_n10315_;
  wire new_n1893_;
  wire new_n4118_;
  wire not_new_n8120_;
  wire new_n3070_;
  wire not_new_n5313_;
  wire new_n4271_;
  wire new_n9881_;
  wire new_n1708_;
  wire not_new_n4104_;
  wire new_n3760_;
  wire not_new_n9267_;
  wire not_new_n4013_;
  wire new_n5596_;
  wire new_n8239_;
  wire new_n10218_;
  wire not_new_n1013__2;
  wire not_pi064_24010;
  wire new_n6903_;
  wire and_new_n3064__new_n998_;
  wire new_n5043_;
  wire not_new_n627__2824752490;
  wire new_n3599_;
  wire not_new_n4283_;
  wire new_n4743_;
  wire not_new_n8799_;
  wire new_n6433_;
  wire new_n2136_;
  wire not_new_n3988_;
  wire not_new_n6196_;
  wire new_n3118_;
  wire new_n8376_;
  wire new_n1700_;
  wire not_new_n9494__0;
  wire new_n6305_;
  wire not_new_n7857_;
  wire not_new_n5013_;
  wire not_new_n1580__3;
  wire new_n4352_;
  wire not_new_n994__4;
  wire not_new_n1055__10;
  wire not_new_n2244_;
  wire not_new_n4118__2;
  wire not_new_n728_;
  wire new_n7973_;
  wire not_new_n3060_;
  wire not_new_n1604__968890104070;
  wire new_n7679_;
  wire not_new_n2623_;
  wire not_new_n8905_;
  wire new_n2892_;
  wire new_n5758_;
  wire new_n8109_;
  wire new_n4963_;
  wire new_n1043_;
  wire not_new_n8169_;
  wire not_new_n3733_;
  wire new_n8412_;
  wire not_new_n7381_;
  wire new_n5668_;
  wire new_n8318_;
  wire new_n6709_;
  wire new_n1318_;
  wire or_not_new_n2953__not_new_n2952_;
  wire new_n4231_;
  wire new_n9906_;
  wire not_new_n5769__0;
  wire not_new_n5242_;
  wire new_n8711_;
  wire new_n4602_;
  wire not_new_n9421_;
  wire not_new_n3983_;
  wire not_new_n5392_;
  wire new_n9518_;
  wire not_new_n8851_;
  wire not_new_n5407_;
  wire not_new_n9932_;
  wire not_new_n3992__0;
  wire not_new_n1599__968890104070;
  wire new_n2840_;
  wire not_new_n3189_;
  wire new_n8694_;
  wire not_new_n5505_;
  wire or_or_not_new_n2557__not_new_n2561__not_new_n1427_;
  wire and_and_new_n3792__new_n3795__new_n3801_;
  wire new_n3192_;
  wire new_n7893_;
  wire not_new_n1594__8235430;
  wire not_new_n2803_;
  wire not_new_n6041_;
  wire new_n8680_;
  wire not_new_n632__2;
  wire or_not_new_n6590__not_new_n6589_;
  wire not_new_n994__16284135979104490;
  wire new_n1194_;
  wire new_n4478_;
  wire new_n3622_;
  wire not_new_n5443__0;
  wire and_new_n6365__new_n6439_;
  wire new_n589_;
  wire not_new_n4303_;
  wire not_new_n9331_;
  wire or_not_pi269_2_not_pi248_2;
  wire new_n661_;
  wire new_n5598_;
  wire new_n9744_;
  wire not_new_n3198_;
  wire new_n10074_;
  wire not_new_n1031__0;
  wire not_new_n9919_;
  wire new_n5669_;
  wire new_n4891_;
  wire not_new_n6806_;
  wire not_new_n6638_;
  wire not_pi001;
  wire not_new_n7610__1;
  wire or_not_new_n4812__not_new_n4736_;
  wire new_n8421_;
  wire new_n2732_;
  wire new_n6088_;
  wire not_new_n1905_;
  wire new_n2051_;
  wire not_new_n4286_;
  wire not_new_n2971_;
  wire not_new_n3185__9;
  wire not_new_n608__10;
  wire new_n6022_;
  wire not_new_n6510_;
  wire new_n9491_;
  wire new_n1581_;
  wire not_new_n7514_;
  wire new_n4005_;
  wire not_new_n6835_;
  wire not_new_n634__8;
  wire new_n8018_;
  wire not_new_n9950__1;
  wire not_new_n3823_;
  wire new_n2350_;
  wire not_new_n8855_;
  wire not_new_n8256__1;
  wire not_new_n8112__1;
  wire new_n9075_;
  wire new_n3555_;
  wire not_new_n644__3;
  wire not_pi184_0;
  wire not_new_n5720__0;
  wire new_n5211_;
  wire not_new_n630__19773267430;
  wire new_n9143_;
  wire not_new_n1597__9;
  wire not_new_n1600__70;
  wire not_new_n610__57648010;
  wire not_new_n9740_;
  wire not_new_n2052_;
  wire not_new_n1055__2;
  wire not_new_n4476_;
  wire po015;
  wire new_n3116_;
  wire not_new_n2567_;
  wire not_new_n8720__0;
  wire and_new_n6388__new_n6313_;
  wire new_n7436_;
  wire new_n2273_;
  wire not_new_n3072_;
  wire new_n2128_;
  wire not_new_n7754_;
  wire new_n9871_;
  wire new_n7318_;
  wire new_n6770_;
  wire new_n7211_;
  wire new_n8100_;
  wire not_new_n607__1;
  wire not_pi146_0;
  wire new_n2980_;
  wire not_new_n7671__0;
  wire not_new_n5156_;
  wire and_new_n4295__new_n4334_;
  wire not_new_n1055__8;
  wire not_new_n1051__490;
  wire new_n5503_;
  wire not_new_n719_;
  wire not_new_n6954_;
  wire not_new_n1053__5;
  wire not_new_n621__19773267430;
  wire new_n5155_;
  wire not_new_n9315_;
  wire new_n10298_;
  wire not_new_n4124_;
  wire not_new_n6368_;
  wire or_or_not_new_n2072__not_new_n2073__not_new_n2075_;
  wire not_new_n591__2824752490;
  wire new_n6200_;
  wire not_new_n3317_;
  wire new_n10203_;
  wire not_new_n4807__1;
  wire not_new_n6925_;
  wire new_n8752_;
  wire new_n3848_;
  wire not_new_n8371_;
  wire not_new_n4219_;
  wire new_n7447_;
  wire new_n8273_;
  wire new_n5915_;
  wire not_new_n4942_;
  wire new_n1811_;
  wire not_new_n8558_;
  wire new_n9228_;
  wire not_new_n8434_;
  wire po157;
  wire not_new_n989__403536070;
  wire key_gate_118;
  wire not_new_n9981_;
  wire not_new_n635__113988951853731430;
  wire not_new_n642__332329305696010;
  wire new_n5877_;
  wire new_n8282_;
  wire not_new_n9901_;
  wire new_n3257_;
  wire not_new_n5452__0;
  wire new_n9975_;
  wire not_new_n7544_;
  wire not_new_n10126_;
  wire new_n8727_;
  wire new_n2192_;
  wire not_pi064_1;
  wire not_new_n9140_;
  wire new_n1196_;
  wire new_n6928_;
  wire not_new_n9930__0;
  wire new_n9266_;
  wire new_n3063_;
  wire new_n10113_;
  wire new_n7902_;
  wire not_new_n1538__5;
  wire not_pi064_70;
  wire not_new_n3375__5;
  wire not_new_n3372__4;
  wire new_n4064_;
  wire new_n9315_;
  wire new_n2219_;
  wire not_new_n7031_;
  wire new_n5481_;
  wire new_n7336_;
  wire not_new_n5052_;
  wire new_n3265_;
  wire not_new_n7143_;
  wire new_n8067_;
  wire new_n1774_;
  wire not_pi104_0;
  wire and_new_n1543__new_n2376_;
  wire not_new_n7603_;
  wire not_new_n4662_;
  wire new_n7963_;
  wire not_new_n7759__1;
  wire not_new_n6859_;
  wire not_new_n5972_;
  wire not_new_n2862_;
  wire po195;
  wire new_n6355_;
  wire new_n6144_;
  wire new_n1962_;
  wire not_new_n8633_;
  wire new_n8036_;
  wire new_n4272_;
  wire not_new_n6307_;
  wire new_n7096_;
  wire not_new_n2303_;
  wire new_n8511_;
  wire new_n4311_;
  wire not_new_n6047_;
  wire not_new_n589__3;
  wire new_n7025_;
  wire new_n1059_;
  wire not_new_n4597_;
  wire new_n3516_;
  wire not_new_n1538__2824752490;
  wire not_new_n8207_;
  wire not_pi138_1;
  wire new_n728_;
  wire not_new_n2535_;
  wire not_new_n10158_;
  wire not_new_n1602__403536070;
  wire not_pi114;
  wire not_new_n1868_;
  wire new_n1259_;
  wire not_new_n1612__7;
  wire new_n7568_;
  wire new_n7323_;
  wire new_n3981_;
  wire not_new_n8258_;
  wire not_new_n5799_;
  wire not_new_n1028__490;
  wire new_n1397_;
  wire new_n7277_;
  wire new_n985_;
  wire and_and_new_n1043__new_n6232__new_n6229_;
  wire not_new_n1600__47475615099430;
  wire new_n1024_;
  wire not_new_n609__7;
  wire new_n7010_;
  wire not_new_n640__24010;
  wire new_n10209_;
  wire po175;
  wire not_new_n4434_;
  wire new_n5852_;
  wire not_new_n1687_;
  wire new_n2975_;
  wire not_new_n7454__0;
  wire not_new_n1728__9;
  wire new_n4353_;
  wire not_new_n8427_;
  wire or_not_new_n8833__not_new_n8830__0;
  wire new_n7945_;
  wire not_pi047_3;
  wire new_n1234_;
  wire not_new_n603__19773267430;
  wire not_new_n6673_;
  wire new_n7185_;
  wire not_new_n7342__0;
  wire new_n6252_;
  wire not_new_n647__19773267430;
  wire new_n5813_;
  wire not_new_n4828_;
  wire new_n4345_;
  wire not_new_n5620_;
  wire not_new_n4417__0;
  wire new_n7066_;
  wire new_n10137_;
  wire not_new_n6625_;
  wire new_n4675_;
  wire not_new_n984__1;
  wire not_new_n5914_;
  wire not_new_n9854__0;
  wire not_new_n1049__7;
  wire new_n8205_;
  wire new_n5495_;
  wire not_new_n627__6;
  wire new_n4798_;
  wire new_n7214_;
  wire new_n6407_;
  wire new_n9748_;
  wire new_n2998_;
  wire or_or_not_new_n2227__not_new_n2224__not_new_n2225_;
  wire new_n5593_;
  wire new_n9259_;
  wire new_n3107_;
  wire not_new_n5531_;
  wire new_n5111_;
  wire not_pi244;
  wire new_n9917_;
  wire new_n5719_;
  wire not_new_n8520_;
  wire not_new_n3837_;
  wire not_pi015;
  wire new_n2383_;
  wire not_new_n4126__0;
  wire not_new_n8595__3;
  wire not_new_n9536_;
  wire not_new_n5140_;
  wire new_n3721_;
  wire not_new_n3032_;
  wire not_new_n2614_;
  wire new_n1692_;
  wire new_n2643_;
  wire or_or_not_new_n4246__not_new_n4350__not_new_n669_;
  wire not_new_n1995__0;
  wire po210;
  wire new_n3155_;
  wire new_n7904_;
  wire not_new_n3921__0;
  wire not_pi183_0;
  wire not_new_n1037__968890104070;
  wire not_new_n589__8235430;
  wire not_new_n5033_;
  wire or_or_not_new_n6337__not_new_n6373__6_not_new_n6338_;
  wire new_n4760_;
  wire new_n590_;
  wire new_n7483_;
  wire not_new_n1051__138412872010;
  wire po292;
  wire not_new_n8303_;
  wire new_n6562_;
  wire new_n1680_;
  wire new_n3749_;
  wire new_n6520_;
  wire not_new_n1057__47475615099430;
  wire and_new_n8304__new_n8299_;
  wire new_n9688_;
  wire new_n6824_;
  wire new_n9305_;
  wire not_po296_77309937197074445241370944070;
  wire not_new_n1613__3430;
  wire not_new_n1051__70;
  wire new_n1974_;
  wire not_new_n7424__0;
  wire new_n3240_;
  wire new_n2396_;
  wire not_new_n6613__1;
  wire not_new_n5746__0;
  wire new_n6761_;
  wire not_new_n634__9;
  wire not_new_n5781_;
  wire not_new_n10204_;
  wire new_n7328_;
  wire new_n8306_;
  wire not_new_n4322__0;
  wire new_n8889_;
  wire not_new_n3516_;
  wire not_new_n5733__0;
  wire not_new_n9083_;
  wire not_new_n1598__1;
  wire not_new_n5550_;
  wire new_n3285_;
  wire new_n5891_;
  wire new_n1627_;
  wire not_new_n6517_;
  wire not_pi133_3;
  wire not_new_n3463_;
  wire not_new_n7753_;
  wire not_new_n1057__6;
  wire not_new_n9873_;
  wire not_new_n7599_;
  wire not_new_n5808__1;
  wire not_new_n1231_;
  wire not_new_n9373__1;
  wire not_new_n6443__16284135979104490;
  wire new_n6122_;
  wire new_n7687_;
  wire new_n5521_;
  wire not_new_n3897_;
  wire not_new_n4963_;
  wire not_new_n6994__0;
  wire not_new_n6580_;
  wire new_n1270_;
  wire not_new_n605__3;
  wire not_new_n637__1;
  wire not_new_n655_;
  wire not_new_n3120_;
  wire new_n4325_;
  wire po248;
  wire not_new_n3416_;
  wire new_n1481_;
  wire not_new_n5474__0;
  wire new_n8508_;
  wire not_new_n3654_;
  wire not_new_n4129__1;
  wire new_n2078_;
  wire new_n3603_;
  wire new_n2672_;
  wire not_new_n1597__1;
  wire not_new_n7960_;
  wire not_new_n602__5;
  wire not_new_n1013__5;
  wire not_new_n5335_;
  wire new_n4083_;
  wire not_new_n7629__0;
  wire new_n5963_;
  wire not_pi058_3;
  wire not_new_n646__10;
  wire new_n8009_;
  wire new_n8888_;
  wire not_pi255_0;
  wire not_new_n1583__6;
  wire not_new_n3311__3;
  wire new_n1402_;
  wire not_new_n8711_;
  wire not_new_n8206_;
  wire new_n2276_;
  wire not_new_n739__0;
  wire new_n1473_;
  wire new_n2557_;
  wire new_n4256_;
  wire new_n7824_;
  wire not_new_n9411_;
  wire not_new_n1039__6;
  wire new_n6968_;
  wire not_po298_403536070;
  wire new_n1963_;
  wire or_not_new_n2890__not_new_n2889_;
  wire not_new_n3570_;
  wire not_new_n9848_;
  wire not_new_n1581__1176490;
  wire not_new_n1602__138412872010;
  wire new_n8633_;
  wire new_n9356_;
  wire new_n8276_;
  wire new_n3389_;
  wire not_new_n7211_;
  wire new_n4820_;
  wire not_new_n9489_;
  wire new_n8512_;
  wire not_new_n3428_;
  wire not_new_n5493_;
  wire not_new_n3879_;
  wire new_n4037_;
  wire not_new_n9399_;
  wire not_new_n1597__2824752490;
  wire not_new_n7913_;
  wire new_n3843_;
  wire new_n3311_;
  wire new_n2055_;
  wire not_new_n8271__2;
  wire not_new_n6608_;
  wire new_n4009_;
  wire new_n9855_;
  wire new_n8208_;
  wire not_new_n9280_;
  wire new_n7204_;
  wire new_n5751_;
  wire not_new_n2263_;
  wire new_n8678_;
  wire not_new_n5905__2;
  wire not_new_n1009__4;
  wire new_n8746_;
  wire new_n10079_;
  wire not_new_n3185__47475615099430;
  wire new_n7487_;
  wire not_new_n3826_;
  wire new_n5729_;
  wire new_n5801_;
  wire not_pi018_0;
  wire and_new_n8874__new_n9276_;
  wire not_new_n8808_;
  wire not_new_n3803_;
  wire new_n5471_;
  wire not_new_n2903_;
  wire new_n4616_;
  wire new_n4208_;
  wire not_new_n644__113988951853731430;
  wire not_new_n599__7;
  wire not_new_n3439_;
  wire not_new_n10015_;
  wire not_new_n3427_;
  wire new_n3530_;
  wire new_n1985_;
  wire new_n5342_;
  wire new_n9707_;
  wire not_new_n587__332329305696010;
  wire not_new_n1594__7;
  wire not_new_n642__70;
  wire not_new_n1589__57648010;
  wire not_new_n1589__968890104070;
  wire not_new_n1163_;
  wire not_new_n6530_;
  wire new_n3579_;
  wire not_new_n1295_;
  wire new_n3061_;
  wire not_new_n8244__2;
  wire not_new_n663_;
  wire not_new_n3657_;
  wire not_new_n624__70;
  wire new_n4032_;
  wire po114;
  wire not_new_n3298_;
  wire not_new_n1588__7;
  wire new_n9986_;
  wire not_new_n635__332329305696010;
  wire new_n9349_;
  wire not_new_n2509__8;
  wire not_new_n8653_;
  wire not_new_n4769_;
  wire not_new_n648__5;
  wire not_new_n6883_;
  wire new_n7523_;
  wire new_n2047_;
  wire new_n980_;
  wire new_n7597_;
  wire new_n6406_;
  wire not_new_n4807_;
  wire not_new_n1599__3;
  wire new_n2300_;
  wire new_n4364_;
  wire not_new_n7403_;
  wire not_pi127_0;
  wire not_pi076;
  wire new_n3184_;
  wire or_or_not_new_n6327__not_new_n6373__2_not_new_n1051__490;
  wire not_new_n8929_;
  wire not_new_n8738_;
  wire new_n3336_;
  wire not_new_n744_;
  wire not_new_n3269_;
  wire not_new_n3680_;
  wire new_n7476_;
  wire new_n2221_;
  wire not_new_n6373__6;
  wire not_new_n601__3430;
  wire new_n4358_;
  wire new_n5564_;
  wire and_new_n8884__new_n9290_;
  wire not_new_n7488_;
  wire new_n1296_;
  wire not_new_n1049__57648010;
  wire new_n3805_;
  wire not_new_n4725_;
  wire new_n7465_;
  wire not_new_n9757_;
  wire not_new_n6175_;
  wire not_new_n8101_;
  wire new_n9857_;
  wire not_new_n1601__13410686196639649008070;
  wire new_n4682_;
  wire new_n5070_;
  wire not_new_n4745_;
  wire new_n992_;
  wire new_n1781_;
  wire new_n6158_;
  wire not_new_n1041__7;
  wire not_new_n4510__0;
  wire not_new_n4837__0;
  wire not_new_n1553_;
  wire not_new_n2541_;
  wire not_new_n4192_;
  wire new_n5659_;
  wire new_n9680_;
  wire not_new_n5547_;
  wire new_n3181_;
  wire new_n2224_;
  wire not_new_n1938_;
  wire new_n925_;
  wire new_n2563_;
  wire not_new_n8255_;
  wire new_n6244_;
  wire not_new_n7180_;
  wire new_n4362_;
  wire and_new_n1330__new_n2274_;
  wire new_n8305_;
  wire and_and_and_new_n1460__new_n1466__new_n1458__new_n1459_;
  wire not_new_n4446__0;
  wire new_n2370_;
  wire not_new_n926_;
  wire not_new_n9959_;
  wire new_n7267_;
  wire not_new_n6117_;
  wire new_n5753_;
  wire not_new_n6977__0;
  wire not_new_n1059_;
  wire new_n3342_;
  wire new_n3688_;
  wire new_n7555_;
  wire not_new_n9966_;
  wire new_n7637_;
  wire not_new_n636__47475615099430;
  wire new_n8081_;
  wire not_new_n3458_;
  wire not_new_n7653__0;
  wire not_new_n3936_;
  wire new_n7377_;
  wire not_new_n10185_;
  wire not_new_n7146__0;
  wire not_new_n8899__0;
  wire not_new_n4759__0;
  wire new_n3939_;
  wire new_n9220_;
  wire not_new_n8080_;
  wire new_n2902_;
  wire new_n7979_;
  wire not_new_n4144_;
  wire new_n9736_;
  wire new_n5151_;
  wire not_new_n10029__2;
  wire not_new_n7602_;
  wire not_new_n626__968890104070;
  wire not_new_n1597__16284135979104490;
  wire new_n8010_;
  wire new_n6163_;
  wire not_new_n1045__9;
  wire not_new_n2186_;
  wire not_new_n647__9;
  wire new_n2174_;
  wire new_n6268_;
  wire new_n2972_;
  wire new_n9717_;
  wire new_n2413_;
  wire not_new_n1605_;
  wire not_new_n5851_;
  wire not_new_n6482__1;
  wire new_n2804_;
  wire new_n2739_;
  wire not_new_n6875_;
  wire not_new_n4507_;
  wire new_n4031_;
  wire new_n9031_;
  wire new_n9949_;
  wire new_n2144_;
  wire new_n7645_;
  wire po294;
  wire not_new_n8330_;
  wire new_n10338_;
  wire not_new_n3136_;
  wire new_n3290_;
  wire new_n1902_;
  wire new_n6221_;
  wire new_n7708_;
  wire not_new_n6488_;
  wire or_or_not_new_n2617__not_new_n2621__not_new_n1439_;
  wire not_new_n6235__0;
  wire new_n6553_;
  wire new_n2785_;
  wire new_n3842_;
  wire new_n4570_;
  wire not_new_n9885_;
  wire new_n9087_;
  wire not_new_n9421__0;
  wire new_n8629_;
  wire not_new_n5812_;
  wire new_n2833_;
  wire not_new_n4735__0;
  wire not_pi043_3;
  wire new_n9178_;
  wire new_n5656_;
  wire not_new_n609__1;
  wire not_new_n4726__0;
  wire new_n1746_;
  wire new_n4322_;
  wire new_n3715_;
  wire new_n9745_;
  wire not_new_n10276_;
  wire not_new_n6983_;
  wire new_n8226_;
  wire not_new_n1488_;
  wire not_new_n6200_;
  wire new_n5311_;
  wire new_n5402_;
  wire not_new_n8376_;
  wire not_new_n6513_;
  wire new_n5462_;
  wire new_n6192_;
  wire not_new_n967_;
  wire new_n1619_;
  wire not_new_n9326__1;
  wire not_new_n642__1176490;
  wire not_new_n1534__2;
  wire not_new_n8980_;
  wire not_new_n6740_;
  wire not_new_n1576__47475615099430;
  wire new_n10186_;
  wire not_new_n6017_;
  wire not_new_n3991__0;
  wire not_new_n7513_;
  wire not_new_n5976_;
  wire not_new_n6993__1;
  wire not_new_n4563_;
  wire not_new_n8222_;
  wire not_new_n3916__0;
  wire not_new_n5551_;
  wire or_not_new_n8941__not_new_n8811_;
  wire new_n8254_;
  wire not_new_n9512__0;
  wire not_new_n3862_;
  wire and_new_n6369__new_n6320_;
  wire new_n7735_;
  wire new_n3231_;
  wire not_new_n587__968890104070;
  wire new_n3368_;
  wire not_new_n10121_;
  wire not_new_n6264_;
  wire new_n5865_;
  wire new_n1282_;
  wire not_new_n5317_;
  wire new_n6721_;
  wire not_new_n602__332329305696010;
  wire po166;
  wire new_n4645_;
  wire new_n2512_;
  wire not_new_n8503_;
  wire not_new_n3310__70;
  wire new_n3227_;
  wire not_new_n4351_;
  wire new_n8159_;
  wire not_new_n1071__57648010;
  wire not_new_n1045__5585458640832840070;
  wire new_n7669_;
  wire not_new_n1428_;
  wire new_n1858_;
  wire not_new_n5898__0;
  wire not_new_n597__138412872010;
  wire new_n8186_;
  wire not_new_n6945_;
  wire not_pi004_0;
  wire new_n7145_;
  wire new_n8019_;
  wire not_new_n6534_;
  wire not_new_n604__19773267430;
  wire not_new_n625__57648010;
  wire new_n5810_;
  wire not_new_n9373_;
  wire new_n1954_;
  wire not_new_n1534__1176490;
  wire new_n2482_;
  wire new_n1955_;
  wire not_new_n2778_;
  wire new_n7903_;
  wire new_n5282_;
  wire not_new_n1585__2;
  wire not_new_n641_;
  wire not_new_n602__7;
  wire new_n2027_;
  wire not_new_n5794__2;
  wire not_new_n3184__7;
  wire new_n2103_;
  wire new_n1922_;
  wire new_n6016_;
  wire po050;
  wire not_new_n5286__0;
  wire new_n2303_;
  wire not_pi157_0;
  wire not_new_n1015__0;
  wire new_n7467_;
  wire not_new_n3185__2326305139872070;
  wire not_new_n9495_;
  wire new_n3541_;
  wire not_new_n10036_;
  wire not_new_n6683__0;
  wire new_n7528_;
  wire new_n3486_;
  wire not_new_n7286_;
  wire not_new_n643__8235430;
  wire not_new_n4733__0;
  wire new_n9300_;
  wire new_n4389_;
  wire new_n2768_;
  wire not_new_n1585__3430;
  wire new_n9370_;
  wire new_n6992_;
  wire new_n3300_;
  wire not_new_n3784_;
  wire and_new_n1334__new_n2293_;
  wire new_n9498_;
  wire not_new_n8001_;
  wire new_n7207_;
  wire new_n4947_;
  wire not_new_n2768_;
  wire not_new_n3749_;
  wire not_new_n5353_;
  wire not_new_n928__16284135979104490;
  wire new_n9395_;
  wire not_new_n630__1;
  wire not_new_n1604__19773267430;
  wire not_new_n7196_;
  wire not_new_n7630__0;
  wire not_new_n4552_;
  wire not_new_n9844_;
  wire new_n3438_;
  wire new_n4169_;
  wire new_n5704_;
  wire not_new_n8856_;
  wire not_new_n4780_;
  wire not_new_n4117__1;
  wire new_n6297_;
  wire not_new_n9954__0;
  wire not_new_n1013__1;
  wire new_n5499_;
  wire new_n1542_;
  wire not_new_n599__403536070;
  wire not_new_n5679_;
  wire not_new_n3656_;
  wire new_n8311_;
  wire not_new_n7043__0;
  wire new_n8952_;
  wire not_pi143_2;
  wire not_new_n10313_;
  wire not_new_n1043__138412872010;
  wire not_new_n10034__0;
  wire not_new_n1576__8;
  wire new_n5892_;
  wire not_new_n1600__0;
  wire not_new_n7029__0;
  wire new_n3549_;
  wire and_new_n1540__new_n2361_;
  wire not_new_n1576__10;
  wire not_new_n7604__0;
  wire and_new_n8982__new_n9323_;
  wire new_n5192_;
  wire not_new_n589__39098210485829880490;
  wire not_new_n6882_;
  wire not_new_n640__7;
  wire new_n6434_;
  wire new_n7246_;
  wire key_gate_16;
  wire new_n4855_;
  wire new_n1876_;
  wire and_and_new_n6385__new_n6386__new_n6241_;
  wire not_new_n3372__93874803376477543056490;
  wire new_n9966_;
  wire new_n1442_;
  wire not_new_n1013__4;
  wire new_n5377_;
  wire new_n3980_;
  wire new_n4940_;
  wire new_n2587_;
  wire not_pi174_2;
  wire new_n10185_;
  wire new_n9023_;
  wire new_n9104_;
  wire not_new_n1584__3430;
  wire not_new_n6827_;
  wire po047;
  wire not_pi247_0;
  wire not_new_n8005_;
  wire new_n3041_;
  wire not_new_n1168_;
  wire not_new_n8710_;
  wire not_new_n4221_;
  wire new_n9844_;
  wire not_new_n6157_;
  wire new_n7235_;
  wire not_new_n7663_;
  wire not_new_n7169_;
  wire new_n2177_;
  wire not_new_n587__7;
  wire new_n4549_;
  wire not_new_n8185_;
  wire not_new_n1616__8;
  wire not_new_n8887__0;
  wire not_new_n5469__0;
  wire new_n7027_;
  wire not_new_n928__6;
  wire not_new_n617__19773267430;
  wire not_new_n5903_;
  wire not_new_n1380_;
  wire po187;
  wire not_new_n9970_;
  wire not_new_n618__13410686196639649008070;
  wire not_new_n5044_;
  wire not_new_n8291_;
  wire new_n6266_;
  wire not_new_n1585__2326305139872070;
  wire not_new_n6258_;
  wire not_new_n8377_;
  wire not_new_n9379__0;
  wire not_new_n3196_;
  wire not_new_n4083_;
  wire not_new_n1613__490;
  wire not_pi025_0;
  wire not_new_n1726_;
  wire new_n8002_;
  wire not_new_n4929_;
  wire new_n2827_;
  wire new_n675_;
  wire not_new_n5683_;
  wire not_new_n585__4;
  wire not_new_n2227_;
  wire new_n6455_;
  wire new_n2781_;
  wire new_n9946_;
  wire new_n4772_;
  wire new_n2475_;
  wire new_n4211_;
  wire not_new_n1536__10;
  wire new_n4426_;
  wire new_n3908_;
  wire new_n1412_;
  wire not_new_n1631__6782230728490;
  wire new_n4554_;
  wire not_new_n4189_;
  wire new_n1364_;
  wire new_n8698_;
  wire new_n5954_;
  wire not_new_n1602__16284135979104490;
  wire not_new_n4723_;
  wire not_new_n9712_;
  wire new_n5893_;
  wire not_new_n609__5;
  wire po131;
  wire not_new_n1583__47475615099430;
  wire not_new_n1067__332329305696010;
  wire not_new_n1537__2326305139872070;
  wire new_n1596_;
  wire new_n7394_;
  wire not_new_n6975_;
  wire not_new_n9240_;
  wire not_new_n2854_;
  wire or_not_new_n2625__not_new_n2624_;
  wire not_new_n7133_;
  wire not_new_n3472_;
  wire not_new_n1580__10;
  wire not_new_n1881_;
  wire new_n4013_;
  wire not_new_n632__24010;
  wire not_new_n7550_;
  wire new_n7498_;
  wire new_n4454_;
  wire not_new_n4831__1;
  wire not_new_n5664_;
  wire new_n3199_;
  wire not_pi200;
  wire new_n5327_;
  wire not_new_n5015_;
  wire not_new_n1053__0;
  wire not_new_n1536_;
  wire new_n1641_;
  wire new_n3604_;
  wire not_new_n9870_;
  wire new_n7577_;
  wire new_n1827_;
  wire new_n9123_;
  wire new_n1457_;
  wire new_n4739_;
  wire not_new_n10009_;
  wire new_n5283_;
  wire not_po296_3;
  wire not_new_n6561_;
  wire not_new_n2340_;
  wire not_new_n9386_;
  wire new_n9755_;
  wire not_new_n637__2;
  wire not_new_n3685_;
  wire not_new_n8277_;
  wire not_new_n5318_;
  wire not_new_n5211_;
  wire not_new_n10138_;
  wire new_n3757_;
  wire new_n6771_;
  wire not_new_n5919__0;
  wire not_new_n589__26517308458596534717790233816010;
  wire not_new_n586__16284135979104490;
  wire not_new_n2784_;
  wire or_not_new_n9103__not_new_n8987__0;
  wire new_n9394_;
  wire new_n2035_;
  wire new_n1460_;
  wire not_new_n2696_;
  wire not_new_n1602__490;
  wire not_new_n1002__6;
  wire not_new_n1576__168070;
  wire not_new_n1596__2824752490;
  wire not_new_n5597__0;
  wire not_new_n7867_;
  wire new_n1053_;
  wire not_new_n1642_;
  wire new_n3610_;
  wire not_new_n4424__0;
  wire not_new_n4749_;
  wire not_new_n7995_;
  wire not_new_n10283_;
  wire new_n3538_;
  wire new_n2935_;
  wire not_new_n6885_;
  wire not_new_n1053__490;
  wire not_new_n10186_;
  wire not_new_n6872_;
  wire not_new_n8140__0;
  wire new_n2135_;
  wire new_n3626_;
  wire new_n5732_;
  wire not_new_n593__9;
  wire not_new_n989__9;
  wire and_and_new_n2048__new_n2051__new_n2049_;
  wire new_n9258_;
  wire not_pi040;
  wire not_new_n633__39098210485829880490;
  wire not_new_n1616__332329305696010;
  wire not_new_n3438_;
  wire not_new_n10007_;
  wire not_new_n8828_;
  wire new_n8883_;
  wire new_n7667_;
  wire not_new_n638__138412872010;
  wire new_n5921_;
  wire not_new_n8244__3;
  wire new_n1468_;
  wire new_n10234_;
  wire and_new_n3768__new_n3771_;
  wire not_new_n587__8;
  wire new_n6759_;
  wire not_new_n8799__1;
  wire new_n10006_;
  wire new_n8307_;
  wire new_n2968_;
  wire new_n3297_;
  wire not_new_n5231_;
  wire not_new_n7004__1;
  wire not_new_n701_;
  wire not_new_n1004__6;
  wire new_n2589_;
  wire new_n10274_;
  wire not_new_n3718_;
  wire not_new_n4748_;
  wire not_new_n603__10;
  wire new_n4610_;
  wire new_n7237_;
  wire new_n8117_;
  wire new_n9690_;
  wire not_new_n3975_;
  wire new_n4186_;
  wire new_n700_;
  wire new_n9051_;
  wire not_new_n1600__4;
  wire not_new_n4175_;
  wire not_new_n3372__3;
  wire not_new_n8338_;
  wire not_new_n1594__10;
  wire not_new_n7657__0;
  wire not_new_n1012__2;
  wire not_new_n6498_;
  wire not_new_n7683_;
  wire new_n1359_;
  wire not_new_n7475_;
  wire not_new_n629__8235430;
  wire new_n3598_;
  wire not_new_n630__403536070;
  wire new_n8612_;
  wire not_new_n8830__1;
  wire not_new_n9390_;
  wire not_new_n1600__1;
  wire not_new_n3931__0;
  wire not_new_n1601__57648010;
  wire not_new_n3250_;
  wire new_n7955_;
  wire new_n9889_;
  wire not_new_n8410_;
  wire not_new_n1580__403536070;
  wire new_n1432_;
  wire not_new_n5746__1;
  wire and_new_n2379__new_n2378_;
  wire not_new_n6995__1;
  wire new_n3344_;
  wire not_pi132_2;
  wire not_new_n2275_;
  wire new_n2340_;
  wire new_n10009_;
  wire not_new_n1158_;
  wire new_n7101_;
  wire new_n9190_;
  wire new_n8365_;
  wire not_new_n5491__0;
  wire not_new_n5796__0;
  wire not_new_n581__2824752490;
  wire or_not_new_n1295__not_new_n1293_;
  wire or_or_not_new_n6334__not_new_n6232__0_not_new_n6235__0;
  wire not_new_n7480_;
  wire not_new_n8835_;
  wire not_new_n9347_;
  wire not_new_n8107__0;
  wire not_new_n1426_;
  wire not_new_n3779_;
  wire not_new_n3372__24010;
  wire new_n2146_;
  wire not_new_n3884_;
  wire new_n5863_;
  wire not_new_n9846_;
  wire not_new_n1538__138412872010;
  wire not_new_n7203_;
  wire not_new_n638__4599865365447399609768010;
  wire not_new_n2504_;
  wire key_gate_126;
  wire not_new_n3185__332329305696010;
  wire not_new_n10145_;
  wire new_n3420_;
  wire new_n4830_;
  wire new_n4198_;
  wire not_new_n628__2326305139872070;
  wire new_n1260_;
  wire not_new_n587__403536070;
  wire new_n4419_;
  wire not_new_n7108_;
  wire new_n1519_;
  wire not_new_n648__332329305696010;
  wire not_new_n3725_;
  wire new_n4561_;
  wire new_n3289_;
  wire not_new_n6496__1;
  wire and_new_n9905__new_n10320_;
  wire new_n6456_;
  wire not_new_n617__1176490;
  wire new_n1891_;
  wire not_new_n10336_;
  wire new_n1501_;
  wire new_n9572_;
  wire new_n9321_;
  wire new_n9340_;
  wire not_pi003;
  wire not_new_n6814_;
  wire not_new_n6774_;
  wire not_new_n631__2326305139872070;
  wire new_n5200_;
  wire not_new_n9923_;
  wire not_new_n1607__5;
  wire not_new_n633__403536070;
  wire new_n5292_;
  wire new_n8164_;
  wire new_n2439_;
  wire not_new_n9556_;
  wire not_new_n631__19773267430;
  wire not_new_n8114_;
  wire not_new_n4485__0;
  wire new_n10246_;
  wire not_new_n630__6;
  wire not_new_n5885_;
  wire not_new_n8290_;
  wire new_n4056_;
  wire new_n9027_;
  wire not_new_n622__1;
  wire new_n10263_;
  wire not_new_n2056_;
  wire not_pi253_1;
  wire not_new_n1071__0;
  wire new_n1213_;
  wire not_new_n8424_;
  wire not_new_n648__39098210485829880490;
  wire new_n8029_;
  wire not_new_n1055__0;
  wire and_new_n2707__new_n2708_;
  wire not_new_n1063__0;
  wire or_or_not_new_n1882__not_new_n1883__not_new_n1885_;
  wire not_new_n5947_;
  wire not_new_n586__2824752490;
  wire not_pi177;
  wire not_new_n3853_;
  wire new_n9034_;
  wire not_new_n638__2326305139872070;
  wire not_new_n581__21838143759917965991093122527538323430;
  wire new_n5179_;
  wire new_n2546_;
  wire not_new_n2419_;
  wire not_pi270;
  wire or_not_new_n2827__not_new_n2826_;
  wire new_n5969_;
  wire new_n1008_;
  wire not_new_n1071__7;
  wire new_n8463_;
  wire not_new_n6976__1;
  wire not_new_n6994__1;
  wire new_n8834_;
  wire new_n7773_;
  wire po156;
  wire new_n582_;
  wire new_n7504_;
  wire new_n6298_;
  wire not_new_n1631__5;
  wire not_new_n7040__1;
  wire not_pi006_0;
  wire new_n7817_;
  wire new_n8069_;
  wire new_n8195_;
  wire new_n9909_;
  wire new_n3461_;
  wire not_new_n7454__1;
  wire not_new_n1589__9;
  wire not_new_n9707_;
  wire new_n4854_;
  wire and_new_n2086__new_n2089_;
  wire new_n8343_;
  wire not_new_n646__1;
  wire not_new_n7415__0;
  wire not_new_n589__13410686196639649008070;
  wire not_new_n4460_;
  wire new_n3746_;
  wire new_n5590_;
  wire new_n6563_;
  wire or_not_new_n3397__not_new_n3398_;
  wire po003;
  wire new_n2453_;
  wire new_n1289_;
  wire not_pi126_0;
  wire new_n9400_;
  wire new_n1286_;
  wire new_n8784_;
  wire new_n5177_;
  wire new_n3119_;
  wire new_n5573_;
  wire new_n4394_;
  wire not_new_n8796_;
  wire new_n6550_;
  wire new_n1513_;
  wire key_gate_30;
  wire not_new_n1067__6;
  wire not_new_n3548_;
  wire po136;
  wire not_new_n4800_;
  wire not_new_n609__6;
  wire and_and_new_n6227__new_n6232__new_n6229_;
  wire not_new_n10002_;
  wire new_n7181_;
  wire not_new_n4129_;
  wire not_new_n4607_;
  wire not_new_n6519_;
  wire not_new_n1536__8;
  wire new_n7755_;
  wire new_n4840_;
  wire not_new_n7656_;
  wire not_new_n1990_;
  wire not_new_n5308_;
  wire not_new_n4933_;
  wire new_n4438_;
  wire not_new_n1922_;
  wire not_new_n6067_;
  wire new_n10313_;
  wire new_n1312_;
  wire not_new_n3414_;
  wire not_new_n3574_;
  wire not_pi121;
  wire new_n7721_;
  wire new_n9724_;
  wire new_n962_;
  wire not_new_n638__6;
  wire not_new_n6691_;
  wire not_new_n8597_;
  wire not_new_n7801__0;
  wire new_n7803_;
  wire not_new_n3876_;
  wire new_n3138_;
  wire or_not_new_n9893__not_new_n9890__0;
  wire not_new_n7825_;
  wire not_new_n1059__47475615099430;
  wire not_new_n8023_;
  wire not_new_n8063_;
  wire not_new_n7312_;
  wire new_n622_;
  wire new_n5815_;
  wire new_n2873_;
  wire not_new_n2439_;
  wire not_new_n9371_;
  wire not_new_n6223__0;
  wire new_n4691_;
  wire or_or_not_new_n1247__not_new_n1245__not_new_n1869_;
  wire or_not_new_n6348__not_new_n6232__2;
  wire not_pi183;
  wire new_n9955_;
  wire or_or_not_new_n1239__not_new_n1237__not_new_n1831_;
  wire not_new_n7928_;
  wire not_new_n4155__0;
  wire not_pi062_0;
  wire not_new_n7315_;
  wire new_n10190_;
  wire not_new_n1043__7;
  wire not_new_n638__19773267430;
  wire new_n4982_;
  wire not_new_n1914_;
  wire new_n4591_;
  wire not_pi035_2;
  wire not_new_n6478__0;
  wire new_n5586_;
  wire new_n2812_;
  wire not_new_n8168_;
  wire new_n9603_;
  wire not_new_n4215_;
  wire and_new_n10034__new_n10289_;
  wire not_new_n7372_;
  wire not_new_n6089_;
  wire not_new_n3387__0;
  wire not_new_n9305_;
  wire new_n3539_;
  wire not_new_n9801_;
  wire not_new_n2318__0;
  wire new_n9888_;
  wire not_pi190;
  wire not_new_n3310__1;
  wire new_n3260_;
  wire not_new_n3422_;
  wire not_new_n640__2;
  wire new_n1186_;
  wire not_new_n8386_;
  wire not_new_n2850_;
  wire not_new_n1016__4;
  wire not_new_n8477_;
  wire not_new_n9652_;
  wire not_new_n8593_;
  wire new_n9324_;
  wire new_n7551_;
  wire new_n4609_;
  wire not_pi147;
  wire not_new_n3512_;
  wire new_n672_;
  wire not_new_n776_;
  wire not_new_n589__47475615099430;
  wire not_new_n7326_;
  wire not_new_n7634__0;
  wire not_new_n6865_;
  wire new_n3264_;
  wire new_n10046_;
  wire not_new_n1602__0;
  wire not_new_n1053__3;
  wire not_new_n8896_;
  wire not_new_n8746_;
  wire not_pi166_0;
  wire not_new_n7641_;
  wire not_new_n1027__138412872010;
  wire not_new_n928__24010;
  wire and_and_new_n1820__new_n1823__new_n1821_;
  wire new_n1607_;
  wire new_n2365_;
  wire not_new_n587__3430;
  wire not_new_n3372__70;
  wire new_n4344_;
  wire not_new_n9952__0;
  wire not_new_n582_;
  wire not_new_n10134_;
  wire new_n9269_;
  wire not_po296_6;
  wire not_new_n3705_;
  wire new_n9464_;
  wire new_n6402_;
  wire new_n2813_;
  wire not_new_n1340_;
  wire and_new_n1731__new_n1732_;
  wire new_n8561_;
  wire not_new_n633__24010;
  wire not_new_n5004_;
  wire new_n4723_;
  wire not_new_n1598_;
  wire not_new_n8105_;
  wire not_new_n4962_;
  wire not_new_n4124__0;
  wire new_n7977_;
  wire new_n2322_;
  wire not_new_n1472_;
  wire new_n7308_;
  wire not_pi263;
  wire not_new_n9492_;
  wire new_n7894_;
  wire not_new_n626__24010;
  wire not_new_n9448_;
  wire new_n6289_;
  wire not_new_n608__70;
  wire new_n5701_;
  wire not_new_n5844_;
  wire not_new_n3666_;
  wire not_new_n4530_;
  wire not_new_n1581__490;
  wire new_n8272_;
  wire not_new_n3184__19773267430;
  wire new_n9089_;
  wire new_n8151_;
  wire not_new_n9915__1;
  wire new_n2820_;
  wire new_n7552_;
  wire not_new_n2805_;
  wire new_n10051_;
  wire new_n8371_;
  wire not_new_n1597__19773267430;
  wire not_new_n2128_;
  wire not_new_n610__10;
  wire not_new_n1009_;
  wire not_new_n7884_;
  wire not_new_n1240_;
  wire new_n8732_;
  wire new_n1723_;
  wire not_new_n1001_;
  wire not_new_n5850_;
  wire not_new_n1043__5;
  wire not_new_n3869_;
  wire not_new_n4920_;
  wire not_new_n7125_;
  wire and_new_n6481__new_n6853_;
  wire not_new_n3686_;
  wire not_new_n1602__113988951853731430;
  wire not_new_n596_;
  wire not_new_n6182_;
  wire not_new_n8156__0;
  wire not_new_n1591__5;
  wire not_new_n4009_;
  wire not_new_n630__2824752490;
  wire new_n2156_;
  wire new_n5356_;
  wire new_n7437_;
  wire new_n5017_;
  wire not_new_n8699_;
  wire not_new_n8798__0;
  wire not_new_n1603__47475615099430;
  wire not_new_n8373_;
  wire new_n10302_;
  wire not_new_n4844_;
  wire new_n9275_;
  wire not_new_n1249_;
  wire new_n1793_;
  wire po213;
  wire not_new_n619__57648010;
  wire not_new_n8813_;
  wire not_new_n5806_;
  wire not_new_n10120_;
  wire not_new_n1049__403536070;
  wire or_not_new_n6250__not_new_n6371_;
  wire not_new_n581__332329305696010;
  wire new_n3736_;
  wire new_n2422_;
  wire not_new_n5326_;
  wire not_new_n4181_;
  wire new_n3682_;
  wire not_new_n5762__0;
  wire new_n7838_;
  wire new_n7925_;
  wire not_new_n8978_;
  wire not_new_n581__2569235775210588780886114772242356213216070;
  wire not_new_n8957_;
  wire not_new_n9227_;
  wire not_new_n4945__1;
  wire not_new_n737_;
  wire new_n1384_;
  wire not_new_n633__797922662976120010;
  wire new_n8843_;
  wire new_n3491_;
  wire new_n5026_;
  wire not_new_n6720_;
  wire not_new_n8725_;
  wire new_n2928_;
  wire not_new_n1591__8235430;
  wire new_n8187_;
  wire new_n10047_;
  wire not_new_n6063_;
  wire not_new_n4827_;
  wire not_new_n8580_;
  wire not_new_n6656__0;
  wire new_n9770_;
  wire new_n6272_;
  wire new_n6404_;
  wire not_new_n581__8;
  wire not_new_n6679_;
  wire not_new_n1043__8;
  wire not_new_n4113__1;
  wire new_n4566_;
  wire not_new_n6559_;
  wire not_new_n8996__0;
  wire new_n9536_;
  wire new_n4150_;
  wire not_new_n6443__2824752490;
  wire not_new_n1536__3430;
  wire not_new_n5277_;
  wire new_n5331_;
  wire new_n628_;
  wire new_n1844_;
  wire new_n5651_;
  wire not_new_n4792__1;
  wire new_n3027_;
  wire not_new_n8067_;
  wire not_new_n644__7;
  wire not_new_n9130_;
  wire not_new_n1584__968890104070;
  wire not_new_n599__1176490;
  wire not_new_n9620_;
  wire not_new_n1063_;
  wire not_new_n2994_;
  wire new_n2790_;
  wire new_n3793_;
  wire not_new_n1012__5;
  wire new_n2034_;
  wire not_new_n9542_;
  wire not_new_n4119__0;
  wire and_new_n6983__new_n7398_;
  wire not_new_n8200_;
  wire not_new_n7622_;
  wire not_new_n1017_;
  wire not_new_n4808_;
  wire not_new_n7701_;
  wire not_new_n1537__490;
  wire new_n9458_;
  wire new_n6807_;
  wire new_n2285_;
  wire not_po296_103677930763188441902487387275962551382129494864490;
  wire not_new_n3360_;
  wire and_new_n1991__new_n1994_;
  wire not_new_n1065__2;
  wire not_new_n619__2824752490;
  wire not_new_n636__10;
  wire not_new_n4744_;
  wire key_gate_4;
  wire not_new_n613__4;
  wire not_new_n9251_;
  wire new_n3873_;
  wire not_pi163;
  wire new_n2664_;
  wire new_n7808_;
  wire not_new_n5552_;
  wire not_new_n593__1176490;
  wire not_new_n8266__0;
  wire not_new_n617__1;
  wire not_new_n1063__168070;
  wire not_new_n2147_;
  wire not_new_n2133_;
  wire not_new_n6727_;
  wire new_n9829_;
  wire new_n8716_;
  wire not_new_n621__4;
  wire not_new_n3168_;
  wire new_n8738_;
  wire new_n3514_;
  wire not_new_n3423_;
  wire new_n7505_;
  wire not_new_n10166_;
  wire not_new_n7033__1;
  wire not_new_n646__7;
  wire new_n1898_;
  wire new_n1802_;
  wire not_new_n1580__5;
  wire and_and_new_n2029__new_n2032__new_n2030_;
  wire not_new_n4527_;
  wire not_new_n4291_;
  wire new_n4927_;
  wire not_new_n7661__0;
  wire not_new_n5061_;
  wire not_new_n3279_;
  wire not_new_n8525_;
  wire not_new_n9607_;
  wire not_new_n3275_;
  wire not_new_n4784_;
  wire not_new_n1037__0;
  wire not_new_n3417_;
  wire not_pi108_0;
  wire new_n2626_;
  wire not_new_n6087_;
  wire and_not_pi040_1_not_pi039_1;
  wire not_new_n9353_;
  wire new_n4043_;
  wire new_n8032_;
  wire not_new_n629__2;
  wire new_n3568_;
  wire not_new_n5557_;
  wire not_new_n4627_;
  wire not_new_n5043_;
  wire not_new_n3384__1;
  wire new_n2467_;
  wire not_new_n622__490;
  wire not_new_n5782__0;
  wire not_new_n581__797922662976120010;
  wire not_new_n9601_;
  wire not_new_n1598__8;
  wire not_new_n3217_;
  wire not_new_n1591__6782230728490;
  wire new_n7144_;
  wire not_new_n4146_;
  wire new_n3322_;
  wire new_n8779_;
  wire new_n1808_;
  wire new_n7424_;
  wire new_n1251_;
  wire new_n4296_;
  wire not_new_n4529_;
  wire not_new_n7911_;
  wire not_new_n611__57648010;
  wire new_n7847_;
  wire new_n2848_;
  wire not_new_n6919_;
  wire not_new_n7835_;
  wire new_n9576_;
  wire not_new_n637__8235430;
  wire not_new_n928__70;
  wire new_n6514_;
  wire not_new_n7128_;
  wire or_or_or_not_new_n2727__not_new_n2730__not_new_n2729__not_new_n2731_;
  wire new_n7048_;
  wire new_n6910_;
  wire new_n1806_;
  wire new_n9242_;
  wire new_n729_;
  wire not_new_n8175_;
  wire new_n5237_;
  wire not_new_n1626_;
  wire not_new_n9509_;
  wire new_n1741_;
  wire new_n1625_;
  wire not_new_n625__2;
  wire not_new_n5532_;
  wire new_n9296_;
  wire not_new_n1805_;
  wire not_new_n634__4;
  wire and_and_new_n1739__new_n1740__new_n1742_;
  wire not_new_n3808_;
  wire new_n8072_;
  wire new_n1977_;
  wire not_new_n6841_;
  wire not_new_n5498__0;
  wire new_n2491_;
  wire new_n5993_;
  wire not_new_n9338_;
  wire new_n10050_;
  wire not_new_n7364_;
  wire new_n5600_;
  wire new_n3206_;
  wire not_new_n7671_;
  wire new_n4653_;
  wire not_new_n1584__6;
  wire new_n5262_;
  wire new_n8213_;
  wire not_new_n3308_;
  wire not_new_n1607__1176490;
  wire new_n10165_;
  wire not_new_n6726_;
  wire new_n2690_;
  wire not_new_n1027__2326305139872070;
  wire new_n4460_;
  wire new_n5449_;
  wire not_new_n1007_;
  wire not_pi102;
  wire not_new_n7919_;
  wire new_n7102_;
  wire not_new_n6514__0;
  wire not_new_n9962__0;
  wire not_new_n10125_;
  wire not_new_n6677__0;
  wire not_new_n9991_;
  wire new_n2773_;
  wire new_n8755_;
  wire new_n3576_;
  wire not_new_n3457_;
  wire not_new_n2564_;
  wire not_new_n4982_;
  wire not_new_n1607__8235430;
  wire new_n9235_;
  wire not_new_n4818_;
  wire new_n1354_;
  wire not_new_n3406_;
  wire not_new_n9733_;
  wire not_new_n5786__2;
  wire or_not_new_n9327__0_not_new_n9524__0;
  wire not_new_n737__0;
  wire not_new_n4454_;
  wire new_n8088_;
  wire new_n9655_;
  wire not_new_n9507_;
  wire not_new_n1055__47475615099430;
  wire not_new_n1616__47475615099430;
  wire not_pi064_1176490;
  wire not_new_n2556_;
  wire not_new_n1031__3430;
  wire not_new_n603__9;
  wire not_new_n648__57648010;
  wire not_pi231;
  wire not_new_n4806_;
  wire not_new_n7433_;
  wire not_new_n1045__24010;
  wire new_n8324_;
  wire not_new_n741__1;
  wire new_n7610_;
  wire new_n3624_;
  wire not_new_n4540_;
  wire new_n7457_;
  wire or_not_new_n1563__not_new_n2474_;
  wire not_new_n647__403536070;
  wire not_new_n1789_;
  wire new_n2245_;
  wire new_n5897_;
  wire not_new_n1444_;
  wire new_n2554_;
  wire not_new_n1619_;
  wire new_n7413_;
  wire new_n9237_;
  wire new_n1924_;
  wire not_new_n2807_;
  wire new_n1761_;
  wire not_new_n5577_;
  wire not_new_n1599__2;
  wire not_pi177_0;
  wire not_new_n9211_;
  wire not_new_n7577_;
  wire new_n3331_;
  wire not_new_n2831_;
  wire new_n5005_;
  wire new_n2616_;
  wire not_new_n9100_;
  wire not_new_n638__8;
  wire not_new_n1468_;
  wire new_n5526_;
  wire not_pi064_138412872010;
  wire new_n5617_;
  wire not_new_n632__39098210485829880490;
  wire new_n5139_;
  wire new_n7411_;
  wire not_new_n588__8235430;
  wire not_new_n4813_;
  wire new_n9460_;
  wire not_new_n612__3;
  wire not_new_n8858_;
  wire not_new_n10031_;
  wire not_new_n984__2326305139872070;
  wire new_n4893_;
  wire not_new_n775__57648010;
  wire new_n4250_;
  wire not_new_n646__2824752490;
  wire new_n724_;
  wire new_n3072_;
  wire not_new_n6507_;
  wire not_new_n7045__2;
  wire new_n3901_;
  wire not_new_n9350_;
  wire new_n6104_;
  wire not_new_n10024_;
  wire new_n1822_;
  wire not_new_n10184_;
  wire new_n1969_;
  wire new_n3991_;
  wire not_new_n593__24010;
  wire not_new_n5339_;
  wire not_new_n974_;
  wire new_n4623_;
  wire not_pi052_1;
  wire not_new_n4501_;
  wire not_new_n4172__0;
  wire not_pi131_2;
  wire not_pi191;
  wire new_n8495_;
  wire new_n8155_;
  wire new_n7596_;
  wire new_n2198_;
  wire not_new_n2509__168070;
  wire not_new_n8671_;
  wire not_new_n7457_;
  wire new_n3068_;
  wire not_new_n1589__332329305696010;
  wire new_n4955_;
  wire not_new_n2663_;
  wire not_new_n6123_;
  wire new_n6510_;
  wire not_new_n704_;
  wire not_new_n5988_;
  wire not_new_n1328_;
  wire new_n6863_;
  wire new_n5435_;
  wire not_new_n5240_;
  wire not_new_n643__9;
  wire not_new_n617__13410686196639649008070;
  wire new_n7203_;
  wire not_new_n1047__9;
  wire not_new_n2626_;
  wire not_new_n647__57648010;
  wire not_new_n602__2326305139872070;
  wire not_new_n641__1;
  wire not_new_n1344_;
  wire not_new_n591__797922662976120010;
  wire not_new_n7027__0;
  wire new_n9044_;
  wire not_new_n1017__4;
  wire new_n4618_;
  wire new_n8748_;
  wire new_n4278_;
  wire or_or_not_new_n2749__not_new_n2752__not_new_n2751_;
  wire new_n6427_;
  wire not_new_n5473__0;
  wire not_new_n8076_;
  wire not_new_n1601__16284135979104490;
  wire not_new_n1588_;
  wire new_n635_;
  wire not_po296_63668057609090279857414351392240010;
  wire and_new_n6244__new_n6372_;
  wire not_new_n633__4;
  wire not_new_n9300_;
  wire new_n4445_;
  wire not_new_n648__3430;
  wire new_n5424_;
  wire not_new_n1581__3430;
  wire not_new_n5548_;
  wire new_n4888_;
  wire not_new_n9368_;
  wire not_new_n642__3;
  wire not_new_n7662_;
  wire not_new_n1636_;
  wire new_n9930_;
  wire not_new_n5689_;
  wire not_new_n9609_;
  wire new_n2401_;
  wire or_or_not_new_n2607__not_new_n2611__not_new_n1437_;
  wire not_new_n604__0;
  wire new_n9116_;
  wire new_n939_;
  wire not_new_n2970_;
  wire new_n3591_;
  wire not_new_n638__7;
  wire not_new_n9699_;
  wire new_n7658_;
  wire not_new_n8450_;
  wire not_new_n7421_;
  wire not_new_n5502_;
  wire not_new_n7729_;
  wire new_n8347_;
  wire not_new_n1602__3430;
  wire new_n6431_;
  wire not_new_n1039__138412872010;
  wire not_new_n9940__0;
  wire not_new_n4510_;
  wire not_pi049_1;
  wire not_new_n1604__1;
  wire not_new_n9144_;
  wire not_new_n5591_;
  wire po001;
  wire new_n4901_;
  wire not_new_n4554_;
  wire new_n1507_;
  wire new_n7884_;
  wire new_n7595_;
  wire not_new_n1599__8;
  wire po147;
  wire not_new_n3772_;
  wire not_new_n5261_;
  wire not_new_n6184_;
  wire not_new_n1569__0;
  wire new_n4683_;
  wire new_n3906_;
  wire new_n1393_;
  wire new_n2130_;
  wire not_new_n10137_;
  wire not_new_n3167_;
  wire new_n2714_;
  wire not_new_n775__138412872010;
  wire not_new_n3655_;
  wire new_n738_;
  wire new_n9899_;
  wire not_new_n7005_;
  wire new_n1371_;
  wire or_not_new_n1549__not_new_n1368_;
  wire new_n2691_;
  wire new_n8201_;
  wire new_n7581_;
  wire not_new_n639__1176490;
  wire new_n2933_;
  wire not_new_n2747_;
  wire not_new_n1027__2;
  wire not_new_n5401_;
  wire not_new_n4002_;
  wire not_new_n7100_;
  wire new_n1728_;
  wire not_new_n989__3430;
  wire not_new_n7613_;
  wire new_n5104_;
  wire new_n6675_;
  wire not_new_n1538__70;
  wire not_new_n1603__24010;
  wire not_new_n6034_;
  wire not_new_n740_;
  wire not_new_n8360_;
  wire new_n3254_;
  wire new_n1031_;
  wire new_n3376_;
  wire not_new_n9917_;
  wire not_new_n4970_;
  wire not_new_n720__0;
  wire not_new_n1067__4;
  wire new_n4637_;
  wire new_n2226_;
  wire new_n6278_;
  wire new_n1067_;
  wire new_n7966_;
  wire not_new_n8845_;
  wire not_new_n5502__0;
  wire new_n8790_;
  wire new_n3237_;
  wire not_new_n1588__113988951853731430;
  wire not_new_n647_;
  wire new_n5295_;
  wire not_new_n7971_;
  wire not_new_n8307_;
  wire new_n2262_;
  wire not_pi048_0;
  wire new_n3178_;
  wire not_new_n9666_;
  wire new_n10049_;
  wire new_n4492_;
  wire not_new_n3349_;
  wire new_n3605_;
  wire not_new_n2730_;
  wire not_new_n4548_;
  wire not_new_n624__9;
  wire not_pi178_3;
  wire new_n3454_;
  wire not_new_n1514_;
  wire new_n5081_;
  wire not_new_n6012_;
  wire new_n5113_;
  wire and_and_new_n1754__new_n1755__new_n1757_;
  wire new_n6288_;
  wire new_n6067_;
  wire not_new_n1039__332329305696010;
  wire new_n7258_;
  wire new_n1721_;
  wire new_n2894_;
  wire not_new_n8081_;
  wire not_new_n8894_;
  wire not_new_n597__70;
  wire not_new_n5890__2;
  wire not_new_n6985__0;
  wire new_n3986_;
  wire not_new_n7780_;
  wire new_n8786_;
  wire new_n9175_;
  wire not_new_n6991_;
  wire not_new_n8173_;
  wire not_new_n626__2;
  wire not_new_n2817_;
  wire not_new_n618__7;
  wire not_new_n7038__0;
  wire new_n5773_;
  wire new_n3909_;
  wire not_new_n2976_;
  wire not_new_n603__6;
  wire not_po296_445676403263631959001900459745680070;
  wire new_n9059_;
  wire not_new_n647__1;
  wire not_new_n8577_;
  wire not_pi254_0;
  wire new_n7625_;
  wire new_n4942_;
  wire not_new_n9088_;
  wire or_or_not_new_n6335__not_new_n6373__4_not_new_n1071__490;
  wire not_new_n3976_;
  wire new_n2772_;
  wire new_n4022_;
  wire new_n6893_;
  wire not_new_n627_;
  wire not_new_n10015__0;
  wire not_new_n5619_;
  wire not_new_n4030__0;
  wire new_n8756_;
  wire or_or_or_not_new_n2919__not_new_n2922__not_new_n2921__not_new_n2923_;
  wire new_n8359_;
  wire not_new_n617__332329305696010;
  wire new_n2786_;
  wire new_n7462_;
  wire new_n2988_;
  wire new_n6651_;
  wire not_new_n1021__0;
  wire not_new_n4314_;
  wire not_new_n7631__2;
  wire new_n4305_;
  wire new_n7631_;
  wire new_n2634_;
  wire new_n1663_;
  wire new_n3243_;
  wire new_n2406_;
  wire not_new_n1864_;
  wire new_n8470_;
  wire not_new_n5282_;
  wire not_pi252_0;
  wire new_n5524_;
  wire new_n2835_;
  wire not_new_n4814__0;
  wire not_pi136_0;
  wire not_new_n9593_;
  wire new_n6092_;
  wire not_new_n4242_;
  wire new_n3190_;
  wire not_new_n625__19773267430;
  wire po028;
  wire not_new_n7406__2;
  wire not_new_n9266_;
  wire new_n5285_;
  wire or_or_or_not_new_n6897__not_new_n6798__not_new_n6826__not_new_n6827_;
  wire not_new_n1043__2;
  wire new_n7868_;
  wire not_new_n2742_;
  wire not_pi229;
  wire not_new_n721__0;
  wire new_n7866_;
  wire not_new_n6366_;
  wire new_n7472_;
  wire not_new_n1057__2;
  wire not_new_n1456_;
  wire new_n7715_;
  wire not_new_n5485_;
  wire new_n3888_;
  wire not_new_n7665__0;
  wire not_new_n1598__138412872010;
  wire new_n1906_;
  wire not_new_n2722_;
  wire not_new_n8328_;
  wire new_n9377_;
  wire not_new_n9507__0;
  wire new_n4535_;
  wire not_new_n8853_;
  wire new_n4612_;
  wire not_new_n7918_;
  wire new_n5515_;
  wire not_new_n581__7490483309651862334944941026945644936490;
  wire new_n4304_;
  wire not_new_n617__797922662976120010;
  wire new_n2573_;
  wire new_n1729_;
  wire new_n5072_;
  wire new_n8705_;
  wire new_n10171_;
  wire not_new_n7021__0;
  wire or_or_or_not_new_n2758__not_new_n2761__not_new_n2760__not_new_n2762_;
  wire not_new_n9977_;
  wire not_new_n6788_;
  wire new_n8404_;
  wire not_new_n9994_;
  wire not_new_n5818_;
  wire not_new_n8248__2;
  wire not_new_n3584_;
  wire not_new_n5543_;
  wire not_new_n1273_;
  wire new_n10048_;
  wire not_new_n6768_;
  wire not_new_n3887_;
  wire not_new_n5482_;
  wire not_new_n5881_;
  wire new_n7744_;
  wire new_n8005_;
  wire new_n3918_;
  wire not_new_n598__5;
  wire not_new_n2154_;
  wire not_new_n5712_;
  wire not_new_n5166_;
  wire not_new_n1773_;
  wire not_new_n2509__9;
  wire new_n5309_;
  wire new_n9038_;
  wire new_n4605_;
  wire new_n3387_;
  wire not_new_n1631__0;
  wire not_new_n10240_;
  wire not_new_n5908_;
  wire not_new_n3710_;
  wire new_n5522_;
  wire new_n5894_;
  wire or_not_new_n680__not_new_n4322_;
  wire not_new_n1613__332329305696010;
  wire not_new_n7725_;
  wire new_n5246_;
  wire new_n2791_;
  wire not_new_n8084_;
  wire new_n7876_;
  wire not_new_n1067__1;
  wire new_n1653_;
  wire or_or_not_new_n1158__0_not_new_n8713__1_not_new_n8785_;
  wire not_new_n7648__0;
  wire not_new_n4153_;
  wire not_new_n9954_;
  wire not_new_n8153_;
  wire not_new_n608__24010;
  wire not_new_n5600_;
  wire and_new_n1278__new_n2027_;
  wire not_new_n1039__5585458640832840070;
  wire not_new_n5406_;
  wire new_n6330_;
  wire new_n9064_;
  wire not_new_n1601__0;
  wire not_new_n4503_;
  wire and_and_new_n1877__new_n1880__new_n1878_;
  wire not_new_n601__168070;
  wire new_n7319_;
  wire new_n2012_;
  wire new_n2886_;
  wire not_new_n3184__70;
  wire new_n3700_;
  wire new_n7779_;
  wire new_n3249_;
  wire new_n2382_;
  wire new_n9840_;
  wire not_new_n1584__8;
  wire new_n9248_;
  wire not_new_n4040_;
  wire new_n8084_;
  wire not_new_n7666_;
  wire new_n711_;
  wire new_n9106_;
  wire not_new_n10110__0;
  wire new_n2720_;
  wire not_pi064_7;
  wire not_new_n4815_;
  wire not_new_n618__4599865365447399609768010;
  wire not_new_n7114_;
  wire and_new_n1318__new_n2217_;
  wire not_new_n5208_;
  wire not_new_n994__10;
  wire not_new_n1017__3;
  wire not_new_n636__138412872010;
  wire new_n3131_;
  wire not_new_n1281_;
  wire not_new_n775__4;
  wire new_n7961_;
  wire not_new_n1588__2326305139872070;
  wire not_new_n3929_;
  wire new_n9145_;
  wire new_n9364_;
  wire not_new_n9023_;
  wire not_new_n1728__8235430;
  wire not_new_n4794__0;
  wire not_new_n7001_;
  wire not_new_n1824_;
  wire new_n4685_;
  wire not_new_n7022__0;
  wire not_new_n5455__0;
  wire not_new_n5815_;
  wire not_new_n9383__0;
  wire not_new_n8912_;
  wire not_new_n5519__0;
  wire new_n5786_;
  wire new_n2702_;
  wire not_new_n10295_;
  wire not_new_n1580__0;
  wire not_new_n5402_;
  wire and_new_n1314__new_n2198_;
  wire not_new_n7774__0;
  wire not_new_n9192_;
  wire new_n6595_;
  wire not_new_n7415_;
  wire new_n3662_;
  wire not_new_n2925_;
  wire not_new_n1051__3430;
  wire not_new_n6932_;
  wire new_n4212_;
  wire new_n2748_;
  wire not_new_n618__32199057558131797268376070;
  wire new_n3416_;
  wire not_new_n10328_;
  wire new_n7354_;
  wire not_new_n6592_;
  wire not_new_n1015__3;
  wire not_pi064_168070;
  wire new_n6319_;
  wire po224;
  wire new_n6821_;
  wire not_pi139_3;
  wire not_new_n5614_;
  wire not_new_n637__7;
  wire not_po298_19773267430;
  wire not_new_n8030_;
  wire new_n4951_;
  wire not_new_n4120_;
  wire new_n8934_;
  wire not_new_n3098_;
  wire new_n9970_;
  wire not_new_n3880_;
  wire new_n4969_;
  wire new_n1896_;
  wire new_n1595_;
  wire not_new_n4502_;
  wire not_new_n3658_;
  wire new_n6799_;
  wire not_new_n638__1;
  wire not_new_n3138_;
  wire new_n3188_;
  wire new_n5912_;
  wire not_new_n3978__0;
  wire and_new_n2409__new_n2408_;
  wire new_n4411_;
  wire not_new_n8114__0;
  wire new_n1847_;
  wire not_new_n624__10;
  wire not_new_n1576__70;
  wire new_n8667_;
  wire not_new_n9855__1;
  wire not_new_n9221_;
  wire new_n9589_;
  wire or_or_not_new_n1275__not_new_n1273__not_new_n2002_;
  wire not_new_n6524__1;
  wire new_n4642_;
  wire new_n7032_;
  wire new_n8758_;
  wire new_n9487_;
  wire new_n4939_;
  wire not_new_n7052_;
  wire new_n3742_;
  wire not_new_n7455_;
  wire new_n3058_;
  wire not_new_n9366_;
  wire not_new_n9095__0;
  wire not_new_n10128__0;
  wire not_new_n6019_;
  wire not_new_n627__24010;
  wire not_new_n6820_;
  wire new_n4397_;
  wire not_new_n9327__0;
  wire not_new_n1065__1176490;
  wire new_n936_;
  wire new_n1843_;
  wire new_n9928_;
  wire not_new_n10237_;
  wire new_n3558_;
  wire new_n7392_;
  wire not_new_n619__10;
  wire not_new_n3160_;
  wire new_n9866_;
  wire new_n4342_;
  wire not_pi051;
  wire new_n2094_;
  wire not_new_n7138_;
  wire new_n9484_;
  wire or_not_new_n9631__not_new_n9515__0;
  wire not_new_n722__1;
  wire not_new_n7412__0;
  wire new_n9389_;
  wire not_pi047_4;
  wire new_n9661_;
  wire new_n8693_;
  wire not_new_n5960_;
  wire not_new_n750_;
  wire new_n5774_;
  wire not_new_n5684_;
  wire not_new_n775__6;
  wire not_new_n10020__0;
  wire new_n1758_;
  wire not_new_n929_;
  wire new_n7547_;
  wire not_new_n639__5585458640832840070;
  wire new_n4080_;
  wire not_new_n5001_;
  wire not_new_n8956__0;
  wire not_new_n630__138412872010;
  wire not_new_n621__2824752490;
  wire new_n4069_;
  wire new_n8614_;
  wire not_new_n8485_;
  wire not_new_n646__1176490;
  wire not_new_n2759_;
  wire new_n8131_;
  wire new_n941_;
  wire not_new_n3157_;
  wire not_new_n1597__3430;
  wire not_new_n5017_;
  wire new_n3965_;
  wire new_n9809_;
  wire po020;
  wire new_n5064_;
  wire not_new_n5788_;
  wire new_n6837_;
  wire new_n6943_;
  wire not_new_n984__0;
  wire not_new_n5795__0;
  wire not_pi043_2;
  wire new_n10191_;
  wire new_n7934_;
  wire not_new_n6793_;
  wire not_new_n10170_;
  wire new_n2562_;
  wire new_n6898_;
  wire not_new_n9219_;
  wire not_new_n9360_;
  wire not_new_n602_;
  wire not_new_n8317_;
  wire key_gate_100;
  wire not_po296_168070;
  wire not_new_n1576_;
  wire not_new_n5743__0;
  wire not_new_n9468_;
  wire not_new_n669_;
  wire not_new_n4430__0;
  wire not_new_n596__2326305139872070;
  wire not_new_n2449_;
  wire not_new_n586__57648010;
  wire new_n3004_;
  wire not_new_n5192__0;
  wire new_n8985_;
  wire new_n983_;
  wire not_new_n7030__0;
  wire new_n2088_;
  wire not_new_n3409_;
  wire not_new_n3442_;
  wire not_new_n1717_;
  wire new_n1892_;
  wire not_new_n601__332329305696010;
  wire not_new_n1602__5;
  wire new_n1272_;
  wire new_n5226_;
  wire new_n2384_;
  wire new_n5112_;
  wire new_n8121_;
  wire new_n976_;
  wire not_new_n8251_;
  wire not_new_n1607__19773267430;
  wire new_n3055_;
  wire new_n6690_;
  wire not_new_n1043__16284135979104490;
  wire new_n4937_;
  wire not_new_n1347_;
  wire not_new_n625__403536070;
  wire not_new_n9314_;
  wire new_n2906_;
  wire not_new_n597__2824752490;
  wire not_new_n7424__1;
  wire not_new_n6787_;
  wire not_pi089;
  wire not_new_n4125_;
  wire not_new_n6533__0;
  wire not_new_n1061__7;
  wire new_n6704_;
  wire not_new_n7148__0;
  wire new_n2438_;
  wire new_n9735_;
  wire not_new_n4760_;
  wire po007;
  wire new_n2521_;
  wire new_n9561_;
  wire new_n2780_;
  wire new_n5505_;
  wire not_new_n3260_;
  wire or_not_new_n2527__not_new_n2531_;
  wire not_new_n6097_;
  wire not_new_n2531_;
  wire new_n2281_;
  wire new_n3000_;
  wire new_n8332_;
  wire not_new_n8838_;
  wire not_new_n1370_;
  wire not_new_n7807_;
  wire new_n3521_;
  wire not_new_n5430__0;
  wire not_new_n5899__0;
  wire not_new_n8407_;
  wire not_new_n7616__0;
  wire new_n3984_;
  wire not_pi275_2;
  wire not_new_n8180_;
  wire new_n5746_;
  wire not_new_n9688_;
  wire new_n7507_;
  wire new_n2859_;
  wire not_pi046_0;
  wire new_n2931_;
  wire new_n8499_;
  wire not_new_n5328_;
  wire new_n8646_;
  wire not_new_n8569_;
  wire new_n5428_;
  wire not_new_n9920_;
  wire new_n7417_;
  wire not_new_n632__403536070;
  wire not_new_n9373__0;
  wire and_and_new_n6251__new_n6371__new_n1597_;
  wire not_new_n632__8235430;
  wire not_new_n9190_;
  wire not_new_n4442_;
  wire not_new_n7829_;
  wire not_new_n7837_;
  wire or_not_new_n3122__not_new_n3121_;
  wire not_new_n4415_;
  wire not_new_n2949_;
  wire not_new_n4525_;
  wire new_n5175_;
  wire not_new_n3263_;
  wire not_new_n6475__2;
  wire not_new_n636__8235430;
  wire new_n1823_;
  wire not_new_n1588__19773267430;
  wire new_n629_;
  wire not_new_n589__2;
  wire not_new_n7598__2;
  wire new_n1529_;
  wire not_new_n3185__1176490;
  wire not_new_n602__968890104070;
  wire new_n6206_;
  wire not_new_n630__16284135979104490;
  wire new_n4240_;
  wire new_n3704_;
  wire not_new_n7661_;
  wire po032;
  wire new_n3128_;
  wire new_n3276_;
  wire not_new_n4300_;
  wire new_n10225_;
  wire not_new_n1047__6782230728490;
  wire new_n9551_;
  wire not_new_n1037__168070;
  wire new_n8505_;
  wire not_new_n2704_;
  wire not_new_n6617__2;
  wire or_not_new_n2129__not_new_n2130_;
  wire new_n1867_;
  wire new_n6184_;
  wire new_n5574_;
  wire or_or_not_new_n6339__not_new_n6232__1_not_new_n6242__3;
  wire new_n5394_;
  wire not_new_n7046_;
  wire not_pi116_0;
  wire not_new_n1596__168070;
  wire not_new_n6826_;
  wire not_new_n5490_;
  wire new_n6626_;
  wire not_new_n1534__4;
  wire not_new_n1631__113988951853731430;
  wire new_n8487_;
  wire key_gate_85;
  wire not_new_n3312_;
  wire not_po298_3;
  wire new_n7989_;
  wire not_new_n954_;
  wire new_n3862_;
  wire or_or_not_new_n1295__not_new_n1293__not_new_n2097_;
  wire not_new_n8984__2;
  wire new_n5820_;
  wire not_new_n8500_;
  wire new_n2089_;
  wire new_n5215_;
  wire new_n6465_;
  wire not_new_n7402_;
  wire not_new_n5680__0;
  wire new_n9868_;
  wire new_n6226_;
  wire not_new_n7212_;
  wire new_n1449_;
  wire not_new_n928__2326305139872070;
  wire po282;
  wire or_not_new_n1558__not_new_n2449_;
  wire new_n3948_;
  wire not_new_n648__4;
  wire not_new_n1612__10;
  wire new_n1175_;
  wire not_new_n8150__2;
  wire new_n3532_;
  wire new_n9061_;
  wire new_n10133_;
  wire key_gate_93;
  wire not_new_n1031__10;
  wire not_new_n8353_;
  wire not_new_n9896_;
  wire not_new_n8119__0;
  wire not_pi144_0;
  wire not_new_n9482_;
  wire not_new_n706_;
  wire not_new_n2870_;
  wire new_n4996_;
  wire new_n2538_;
  wire not_new_n4767__0;
  wire new_n4517_;
  wire not_pi148_0;
  wire not_new_n9657_;
  wire not_new_n7039__0;
  wire new_n1862_;
  wire not_po296_968890104070;
  wire new_n3526_;
  wire not_new_n594__6;
  wire new_n2194_;
  wire new_n10310_;
  wire not_new_n5230_;
  wire not_new_n8876_;
  wire not_new_n775__5;
  wire not_new_n8829_;
  wire new_n6294_;
  wire new_n3453_;
  wire new_n6681_;
  wire new_n4040_;
  wire new_n6636_;
  wire not_new_n3470_;
  wire new_n5314_;
  wire new_n7964_;
  wire and_new_n9510__new_n9851_;
  wire new_n2970_;
  wire not_new_n2112_;
  wire not_new_n6996__0;
  wire new_n5597_;
  wire not_new_n6650__0;
  wire new_n2490_;
  wire new_n7028_;
  wire not_pi273;
  wire not_new_n3979_;
  wire new_n7508_;
  wire not_new_n9984_;
  wire not_new_n8598_;
  wire new_n5943_;
  wire new_n2229_;
  wire new_n5513_;
  wire not_new_n4132__1;
  wire new_n6971_;
  wire new_n9720_;
  wire not_new_n5513_;
  wire not_pi180;
  wire not_new_n6658_;
  wire not_new_n626__4599865365447399609768010;
  wire new_n2548_;
  wire new_n9574_;
  wire not_new_n628__113988951853731430;
  wire new_n3861_;
  wire not_new_n1597__0;
  wire not_new_n3665_;
  wire new_n7752_;
  wire new_n10092_;
  wire new_n5683_;
  wire new_n5427_;
  wire new_n3808_;
  wire po174;
  wire po110;
  wire not_pi180_0;
  wire new_n4979_;
  wire not_new_n6507__1;
  wire new_n5602_;
  wire not_new_n617__70;
  wire new_n2825_;
  wire not_new_n9563_;
  wire not_new_n1352_;
  wire new_n6223_;
  wire not_new_n984__3;
  wire new_n2595_;
  wire new_n4377_;
  wire not_new_n5470_;
  wire not_pi047_2;
  wire new_n2816_;
  wire not_new_n603__70;
  wire not_new_n5731_;
  wire new_n5260_;
  wire not_new_n10269_;
  wire new_n9590_;
  wire new_n5587_;
  wire new_n5605_;
  wire not_new_n7955_;
  wire not_new_n5058__0;
  wire new_n4600_;
  wire not_new_n5387_;
  wire new_n5149_;
  wire not_new_n6684_;
  wire not_new_n6447_;
  wire not_new_n4988_;
  wire not_new_n8830__0;
  wire not_new_n6363_;
  wire not_new_n5209__0;
  wire new_n1964_;
  wire not_new_n6511_;
  wire new_n10173_;
  wire not_new_n9157_;
  wire or_or_not_new_n2758__not_new_n2761__not_new_n2760_;
  wire new_n8682_;
  wire new_n2267_;
  wire not_new_n9538_;
  wire not_new_n6736_;
  wire not_new_n10061_;
  wire not_new_n9239_;
  wire not_pi048_1;
  wire new_n2316_;
  wire not_new_n1009__1;
  wire or_not_new_n3363__not_new_n583__0;
  wire new_n2718_;
  wire not_new_n4481_;
  wire not_new_n7693_;
  wire not_new_n644__490;
  wire not_new_n4804__0;
  wire new_n4406_;
  wire not_new_n8199_;
  wire new_n2995_;
  wire new_n9673_;
  wire new_n3789_;
  wire not_new_n7758_;
  wire not_new_n1037__7;
  wire not_new_n632_;
  wire not_new_n1538__1;
  wire new_n2161_;
  wire new_n6485_;
  wire not_new_n9988_;
  wire new_n5761_;
  wire new_n4273_;
  wire not_new_n3003_;
  wire not_new_n5471__0;
  wire not_new_n594__2;
  wire new_n9911_;
  wire new_n4763_;
  wire not_new_n7305_;
  wire not_new_n1019__4;
  wire not_new_n5111_;
  wire not_new_n589__19773267430;
  wire new_n1338_;
  wire not_new_n3711_;
  wire new_n7453_;
  wire not_new_n589__0;
  wire new_n7695_;
  wire new_n2042_;
  wire not_new_n3820_;
  wire new_n6871_;
  wire new_n3803_;
  wire not_new_n3325_;
  wire new_n2433_;
  wire not_new_n7115_;
  wire new_n9285_;
  wire new_n7164_;
  wire not_new_n7412_;
  wire not_new_n10258_;
  wire not_new_n1151_;
  wire not_new_n7066_;
  wire not_new_n645__6;
  wire new_n5890_;
  wire not_new_n9377__0;
  wire new_n7549_;
  wire not_new_n6370__1;
  wire not_new_n3132_;
  wire not_new_n5716_;
  wire not_new_n1053__2326305139872070;
  wire not_new_n7882_;
  wire not_pi053;
  wire not_new_n8986_;
  wire not_new_n6975__1;
  wire new_n4387_;
  wire not_new_n4460__0;
  wire new_n5207_;
  wire key_gate_122;
  wire not_new_n7410_;
  wire not_new_n619__8235430;
  wire new_n5201_;
  wire new_n7538_;
  wire not_new_n3069_;
  wire not_new_n585__6;
  wire new_n2945_;
  wire not_new_n9319_;
  wire new_n6103_;
  wire not_new_n4169__0;
  wire new_n5223_;
  wire not_new_n2015_;
  wire new_n9431_;
  wire not_new_n4440__0;
  wire not_pi065;
  wire not_new_n4449__0;
  wire not_new_n3372__8235430;
  wire new_n5672_;
  wire not_new_n5352_;
  wire new_n3108_;
  wire new_n8408_;
  wire new_n7674_;
  wire not_new_n8907_;
  wire not_new_n6493__0;
  wire not_pi266;
  wire not_pi057_0;
  wire new_n6593_;
  wire new_n2658_;
  wire new_n9386_;
  wire new_n10178_;
  wire new_n3733_;
  wire not_new_n2776_;
  wire not_new_n7529_;
  wire not_new_n6792_;
  wire new_n1638_;
  wire not_new_n8314__0;
  wire new_n9047_;
  wire not_new_n7860_;
  wire not_pi034;
  wire not_new_n1612__332329305696010;
  wire new_n5095_;
  wire new_n8769_;
  wire not_po296_11044276742439206463052992010;
  wire not_new_n5729_;
  wire new_n8783_;
  wire new_n5000_;
  wire new_n3807_;
  wire new_n2145_;
  wire not_new_n1584__70;
  wire not_new_n4533_;
  wire new_n8157_;
  wire or_not_new_n1315__not_new_n1313_;
  wire not_new_n585__2;
  wire not_new_n2090__0;
  wire not_new_n5284_;
  wire or_not_new_n1239__not_new_n1237_;
  wire not_po298_2824752490;
  wire not_new_n9879__1;
  wire new_n4416_;
  wire not_new_n8308__0;
  wire new_n1765_;
  wire not_new_n980_;
  wire not_new_n596__7;
  wire new_n4933_;
  wire not_new_n589__3119734822845423713013303218219760490;
  wire new_n7676_;
  wire not_new_n1031__138412872010;
  wire new_n6929_;
  wire not_new_n6134_;
  wire not_new_n9099_;
  wire not_new_n4054_;
  wire not_new_n7038__1;
  wire new_n9328_;
  wire not_new_n7719_;
  wire and_and_new_n8723__new_n1174__new_n8719_;
  wire not_new_n6978_;
  wire new_n2395_;
  wire not_new_n589__273687473400809163430;
  wire new_n4672_;
  wire not_new_n1041__70;
  wire not_new_n598__6;
  wire not_new_n9861_;
  wire not_new_n1585__70;
  wire not_new_n6491_;
  wire new_n8022_;
  wire not_new_n1599__6782230728490;
  wire not_new_n737__1;
  wire new_n4681_;
  wire or_or_not_new_n2874__not_new_n2877__not_new_n2876_;
  wire not_new_n3659_;
  wire not_new_n984__19773267430;
  wire new_n2775_;
  wire not_new_n3310__2;
  wire not_new_n9428__0;
  wire not_new_n3797_;
  wire new_n4732_;
  wire not_new_n5742__2;
  wire not_new_n6462_;
  wire new_n6809_;
  wire not_new_n9053_;
  wire not_new_n636__9;
  wire not_new_n1448_;
  wire new_n5709_;
  wire new_n10025_;
  wire new_n8433_;
  wire not_new_n5695_;
  wire po132;
  wire new_n8532_;
  wire not_new_n6443__47475615099430;
  wire new_n2763_;
  wire not_new_n8931_;
  wire not_new_n1071__2;
  wire new_n6670_;
  wire not_new_n641__0;
  wire not_new_n7768__0;
  wire not_new_n1607__2824752490;
  wire not_new_n1022_;
  wire not_new_n3084_;
  wire not_new_n7394_;
  wire new_n8163_;
  wire key_gate_114;
  wire not_new_n3145_;
  wire not_new_n586__403536070;
  wire not_new_n638__797922662976120010;
  wire not_new_n3833_;
  wire new_n9714_;
  wire not_new_n6535_;
  wire new_n7011_;
  wire or_not_new_n2575__not_new_n2574_;
  wire not_new_n645__168070;
  wire new_n8153_;
  wire not_new_n604__24010;
  wire new_n2190_;
  wire not_new_n6554_;
  wire new_n6213_;
  wire not_new_n1012__1;
  wire new_n8656_;
  wire new_n9638_;
  wire new_n3253_;
  wire new_n7855_;
  wire not_new_n5680_;
  wire new_n4218_;
  wire new_n5584_;
  wire new_n3175_;
  wire not_new_n5078__2;
  wire not_new_n1047__6;
  wire not_new_n8846_;
  wire not_new_n7754__2;
  wire and_new_n10032__new_n580_;
  wire new_n9554_;
  wire not_new_n6763_;
  wire not_new_n631__403536070;
  wire new_n9282_;
  wire not_new_n9943_;
  wire not_new_n5426__0;
  wire new_n8428_;
  wire new_n2066_;
  wire new_n6645_;
  wire not_new_n7113__1;
  wire new_n9289_;
  wire not_new_n608__4;
  wire not_new_n7044_;
  wire new_n8668_;
  wire not_new_n5400_;
  wire and_and_new_n8724__new_n8726__new_n8728_;
  wire not_new_n1009__5;
  wire new_n8966_;
  wire not_new_n2147__0;
  wire new_n3417_;
  wire not_new_n8329_;
  wire not_new_n618__8;
  wire not_new_n613__5;
  wire not_new_n6450_;
  wire and_new_n1446__new_n2659_;
  wire not_new_n627__968890104070;
  wire not_new_n10123_;
  wire not_new_n641__7;
  wire new_n6746_;
  wire and_and_new_n4298__new_n4341__new_n4345_;
  wire new_n5399_;
  wire not_new_n9726_;
  wire or_or_not_new_n8528__not_new_n8429__not_new_n8457_;
  wire new_n9131_;
  wire not_new_n4966_;
  wire not_new_n1202_;
  wire not_new_n8054_;
  wire not_new_n3075_;
  wire not_new_n1604__7;
  wire not_new_n645__9;
  wire new_n9905_;
  wire not_new_n3200_;
  wire po105;
  wire new_n9737_;
  wire new_n933_;
  wire not_new_n9058_;
  wire not_new_n4568_;
  wire new_n3048_;
  wire not_new_n8573_;
  wire new_n8080_;
  wire not_new_n3519_;
  wire not_new_n1534__403536070;
  wire not_new_n1045__5;
  wire not_new_n1161__0;
  wire new_n1013_;
  wire not_new_n611__403536070;
  wire new_n4578_;
  wire not_new_n5495_;
  wire not_new_n7347_;
  wire new_n657_;
  wire new_n8014_;
  wire new_n8936_;
  wire new_n5274_;
  wire not_new_n3576_;
  wire not_new_n6745__0;
  wire not_new_n9979_;
  wire and_and_new_n6369__new_n6320__new_n6230_;
  wire new_n1246_;
  wire new_n3212_;
  wire or_or_not_new_n1773__not_new_n1213__not_new_n1214_;
  wire not_new_n1599__403536070;
  wire not_new_n9424_;
  wire not_new_n8159_;
  wire not_new_n4791_;
  wire new_n4500_;
  wire not_new_n9644_;
  wire not_new_n3372__797922662976120010;
  wire new_n8356_;
  wire not_new_n1065__47475615099430;
  wire not_new_n630__24010;
  wire not_new_n8104__0;
  wire new_n3785_;
  wire not_new_n1548_;
  wire new_n6367_;
  wire not_new_n6908_;
  wire new_n6698_;
  wire new_n2686_;
  wire not_new_n1071__3430;
  wire new_n7668_;
  wire not_new_n3560_;
  wire not_new_n7007_;
  wire not_new_n6057_;
  wire not_new_n8653__0;
  wire not_new_n626__57648010;
  wire new_n3023_;
  wire not_pi257_3;
  wire new_n2926_;
  wire not_new_n4275_;
  wire not_new_n3802_;
  wire new_n1550_;
  wire not_new_n612__7;
  wire not_new_n2772_;
  wire new_n1486_;
  wire not_new_n1065__168070;
  wire not_new_n4319__0;
  wire not_new_n1538__168070;
  wire or_not_pi245_0_not_new_n1625_;
  wire not_new_n4282_;
  wire new_n8192_;
  wire not_new_n2284_;
  wire new_n2974_;
  wire not_new_n10004_;
  wire new_n1590_;
  wire not_new_n600__10;
  wire not_new_n6575_;
  wire not_new_n8685_;
  wire not_new_n3388_;
  wire not_new_n603__7;
  wire not_new_n4936_;
  wire new_n8651_;
  wire new_n5434_;
  wire new_n7355_;
  wire new_n5840_;
  wire not_new_n5798__0;
  wire not_new_n3663_;
  wire new_n7174_;
  wire new_n9176_;
  wire not_new_n8271__1;
  wire new_n678_;
  wire not_new_n4673_;
  wire not_new_n1588__39098210485829880490;
  wire not_new_n8859_;
  wire new_n8434_;
  wire not_pi210;
  wire not_new_n1604__113988951853731430;
  wire not_new_n3125_;
  wire new_n4258_;
  wire not_new_n594__138412872010;
  wire new_n9485_;
  wire new_n1011_;
  wire new_n7915_;
  wire new_n5520_;
  wire or_or_or_not_new_n2820__not_new_n2823__not_new_n2822__not_new_n2824_;
  wire new_n6307_;
  wire not_new_n2718_;
  wire new_n4421_;
  wire not_new_n618__9;
  wire not_new_n1591__1;
  wire new_n2657_;
  wire not_new_n1775_;
  wire not_new_n7366__1;
  wire new_n6344_;
  wire not_new_n1406_;
  wire not_new_n10027_;
  wire not_new_n5511_;
  wire not_new_n6212_;
  wire not_new_n8097_;
  wire not_new_n5459_;
  wire not_new_n6526_;
  wire new_n6958_;
  wire not_new_n5079_;
  wire not_new_n9829_;
  wire not_new_n4112_;
  wire new_n7030_;
  wire not_new_n1431_;
  wire not_new_n8869_;
  wire not_new_n8816_;
  wire not_new_n594__3;
  wire and_and_new_n1801__new_n1804__new_n1802_;
  wire not_new_n1604__332329305696010;
  wire new_n658_;
  wire not_new_n637__6;
  wire or_not_new_n1564__not_new_n2479_;
  wire new_n5782_;
  wire not_new_n648__797922662976120010;
  wire and_new_n2424__new_n2423_;
  wire not_new_n601__3;
  wire new_n993_;
  wire not_new_n10075_;
  wire not_new_n611__19773267430;
  wire new_n9685_;
  wire not_pi275_3;
  wire po036;
  wire not_new_n1043__1176490;
  wire not_new_n8934_;
  wire not_new_n7454_;
  wire new_n3323_;
  wire not_new_n7728_;
  wire new_n3966_;
  wire not_new_n7129_;
  wire not_new_n9835_;
  wire not_pi238;
  wire new_n6448_;
  wire new_n9416_;
  wire or_not_new_n5430__0_not_pi130_2;
  wire not_pi116;
  wire key_gate_15;
  wire new_n3186_;
  wire po048;
  wire new_n4370_;
  wire new_n9627_;
  wire new_n4746_;
  wire not_new_n581_;
  wire not_new_n7024_;
  wire or_not_new_n2617__not_new_n2621_;
  wire new_n10152_;
  wire not_new_n4125__0;
  wire not_new_n643__113988951853731430;
  wire po268;
  wire not_new_n9487__0;
  wire new_n6466_;
  wire not_new_n984__6;
  wire not_new_n624__57648010;
  wire or_not_new_n2765__not_new_n2764_;
  wire not_new_n6639_;
  wire not_new_n5759_;
  wire not_new_n2264_;
  wire new_n1915_;
  wire not_new_n630__6782230728490;
  wire not_new_n6529_;
  wire new_n9587_;
  wire new_n9711_;
  wire new_n4977_;
  wire new_n4902_;
  wire not_new_n7008__1;
  wire new_n6865_;
  wire new_n3583_;
  wire not_new_n7067_;
  wire not_new_n7887_;
  wire not_new_n3949_;
  wire not_new_n8618_;
  wire new_n8768_;
  wire new_n3578_;
  wire not_new_n8854__0;
  wire not_new_n1438_;
  wire not_new_n8572_;
  wire new_n8062_;
  wire new_n3414_;
  wire po144;
  wire not_new_n2684_;
  wire not_new_n621__24010;
  wire not_new_n5734_;
  wire not_pi247;
  wire not_new_n589__70;
  wire not_new_n581__1915812313805664144010;
  wire not_new_n1067__490;
  wire not_pi054_0;
  wire not_new_n5508_;
  wire not_new_n636__1;
  wire not_new_n6586_;
  wire new_n2427_;
  wire new_n7703_;
  wire not_new_n6983__1;
  wire not_new_n9900__1;
  wire not_new_n4989_;
  wire not_new_n9506__2;
  wire new_n7407_;
  wire new_n9186_;
  wire not_new_n2945_;
  wire not_new_n8848__0;
  wire new_n610_;
  wire not_new_n4448_;
  wire not_new_n639__273687473400809163430;
  wire new_n5359_;
  wire not_new_n8177__0;
  wire new_n3198_;
  wire not_new_n594__2326305139872070;
  wire new_n4120_;
  wire not_new_n7600__0;
  wire not_new_n4756_;
  wire new_n8211_;
  wire not_new_n3372__273687473400809163430;
  wire new_n5376_;
  wire not_new_n2484_;
  wire new_n3492_;
  wire not_new_n6309_;
  wire new_n10288_;
  wire not_pi164;
  wire not_new_n5192_;
  wire new_n6359_;
  wire not_new_n6341_;
  wire not_new_n5995_;
  wire new_n4892_;
  wire new_n9067_;
  wire not_new_n1604__403536070;
  wire not_po298_138412872010;
  wire not_new_n634__332329305696010;
  wire not_new_n621__490;
  wire not_new_n1537__57648010;
  wire new_n7442_;
  wire not_new_n648__1176490;
  wire new_n5947_;
  wire not_new_n2636_;
  wire not_new_n604__403536070;
  wire not_new_n4506_;
  wire not_new_n622__138412872010;
  wire new_n8861_;
  wire not_new_n1051__0;
  wire new_n5100_;
  wire not_new_n604__3;
  wire not_new_n4877_;
  wire not_new_n581__1;
  wire not_new_n732__1;
  wire not_new_n5799__0;
  wire new_n1150_;
  wire not_pi062;
  wire not_new_n6158_;
  wire not_new_n3448_;
  wire new_n10267_;
  wire not_new_n5539_;
  wire new_n7710_;
  wire not_new_n8536_;
  wire new_n5099_;
  wire not_new_n4809__0;
  wire not_new_n1065__138412872010;
  wire new_n3393_;
  wire not_new_n2334_;
  wire or_not_new_n3094__not_new_n3093_;
  wire new_n7865_;
  wire new_n1736_;
  wire new_n3283_;
  wire not_new_n5537_;
  wire new_n6165_;
  wire not_new_n2338_;
  wire not_new_n5478__0;
  wire not_new_n5510_;
  wire new_n7927_;
  wire not_pi094;
  wire new_n2445_;
  wire new_n9581_;
  wire not_new_n625__138412872010;
  wire not_new_n5615_;
  wire new_n9398_;
  wire not_new_n9970__0;
  wire not_new_n4296_;
  wire not_new_n2246_;
  wire new_n7002_;
  wire not_new_n9171_;
  wire not_new_n8681_;
  wire not_pi138;
  wire new_n9187_;
  wire not_new_n3184__5;
  wire not_new_n648__0;
  wire not_new_n1365_;
  wire not_new_n6492__0;
  wire not_new_n632__1176490;
  wire po139;
  wire new_n1575_;
  wire not_new_n625__113988951853731430;
  wire not_new_n8713__1;
  wire not_new_n5513__0;
  wire not_new_n1536__5585458640832840070;
  wire new_n8023_;
  wire not_new_n5278_;
  wire new_n5749_;
  wire not_new_n4191_;
  wire not_new_n8845__0;
  wire not_new_n3528_;
  wire key_gate_49;
  wire not_new_n7951_;
  wire not_new_n639__19773267430;
  wire not_pi169;
  wire not_new_n693_;
  wire not_new_n8958__0;
  wire not_new_n4028_;
  wire not_new_n3185__6782230728490;
  wire new_n4871_;
  wire new_n3601_;
  wire new_n10087_;
  wire new_n8007_;
  wire not_new_n9693_;
  wire new_n3854_;
  wire not_po298_57648010;
  wire not_new_n1041__4;
  wire new_n3189_;
  wire new_n9584_;
  wire not_new_n3041_;
  wire not_new_n7801_;
  wire not_new_n1053__10;
  wire not_new_n8267_;
  wire new_n4889_;
  wire new_n9731_;
  wire not_new_n5773_;
  wire not_new_n5372_;
  wire not_new_n4468_;
  wire new_n4852_;
  wire new_n4485_;
  wire new_n1388_;
  wire new_n6447_;
  wire not_new_n6094_;
  wire not_new_n4410__0;
  wire new_n6015_;
  wire not_new_n3311__8235430;
  wire not_new_n4930__1;
  wire not_new_n4431_;
  wire new_n8383_;
  wire not_new_n1027__7;
  wire new_n7248_;
  wire new_n1672_;
  wire not_new_n9365__0;
  wire not_new_n1604__10;
  wire new_n7696_;
  wire not_new_n7250_;
  wire not_new_n3915__0;
  wire not_new_n6232_;
  wire new_n9870_;
  wire not_new_n1419_;
  wire not_new_n7929_;
  wire or_or_or_not_new_n1773__not_new_n1213__not_new_n1214__not_new_n1775_;
  wire not_new_n632__2824752490;
  wire not_new_n928__6782230728490;
  wire not_new_n1071__8;
  wire new_n6353_;
  wire not_new_n4131_;
  wire new_n9323_;
  wire new_n4221_;
  wire not_new_n10081_;
  wire not_new_n7626__0;
  wire not_new_n7592_;
  wire not_new_n1055__9;
  wire new_n2359_;
  wire not_new_n6505_;
  wire new_n4412_;
  wire not_new_n3763_;
  wire new_n4706_;
  wire new_n1720_;
  wire new_n2291_;
  wire new_n2470_;
  wire new_n6386_;
  wire not_new_n626__3430;
  wire not_new_n1045__273687473400809163430;
  wire new_n1851_;
  wire new_n3402_;
  wire new_n6688_;
  wire new_n9802_;
  wire new_n9030_;
  wire new_n7998_;
  wire new_n8836_;
  wire not_new_n3255_;
  wire not_new_n702_;
  wire new_n7599_;
  wire not_new_n609__10;
  wire new_n1618_;
  wire not_new_n1581__6782230728490;
  wire not_new_n2824_;
  wire new_n3928_;
  wire and_new_n6395__new_n6396_;
  wire new_n5775_;
  wire not_new_n5767__1;
  wire not_new_n1613__19773267430;
  wire not_new_n4843__0;
  wire not_new_n7154_;
  wire not_new_n9729_;
  wire new_n10042_;
  wire new_n2996_;
  wire or_not_new_n7046__not_new_n7265_;
  wire not_new_n3372__47475615099430;
  wire new_n997_;
  wire not_new_n8836_;
  wire not_new_n5677_;
  wire not_new_n631__10;
  wire new_n3804_;
  wire or_not_new_n5041__not_new_n4911_;
  wire not_new_n7617_;
  wire new_n5581_;
  wire po281;
  wire not_new_n8656_;
  wire new_n8579_;
  wire not_new_n6870_;
  wire not_new_n596__10;
  wire not_new_n6687_;
  wire not_new_n7842_;
  wire new_n8931_;
  wire new_n2233_;
  wire new_n3208_;
  wire not_new_n6539_;
  wire not_new_n5756__0;
  wire not_new_n1028__3;
  wire new_n1959_;
  wire not_new_n1043__9;
  wire not_new_n1002_;
  wire not_new_n5500_;
  wire new_n5582_;
  wire not_new_n627__332329305696010;
  wire or_or_not_new_n1299__not_new_n1297__not_new_n2116_;
  wire not_new_n4487__0;
  wire not_new_n1584__0;
  wire not_new_n10144__0;
  wire key_gate_91;
  wire new_n9317_;
  wire new_n5710_;
  wire not_new_n618__70;
  wire not_new_n5564_;
  wire not_new_n7777_;
  wire not_new_n1383_;
  wire not_new_n4330__0;
  wire new_n8891_;
  wire new_n10144_;
  wire new_n3087_;
  wire new_n4638_;
  wire new_n9203_;
  wire new_n7261_;
  wire not_new_n1607__6;
  wire new_n1407_;
  wire not_new_n4751__0;
  wire not_new_n1589__138412872010;
  wire not_new_n10294_;
  wire new_n2577_;
  wire not_new_n3941_;
  wire not_new_n638__6782230728490;
  wire not_new_n635__7;
  wire not_new_n646__968890104070;
  wire not_pi132_0;
  wire new_n6509_;
  wire new_n7682_;
  wire new_n3459_;
  wire not_new_n3430_;
  wire not_new_n581__19773267430;
  wire not_new_n1939_;
  wire or_not_new_n2675__not_new_n2674_;
  wire not_new_n4719_;
  wire new_n2526_;
  wire not_new_n8396_;
  wire not_new_n4911_;
  wire new_n6413_;
  wire new_n3170_;
  wire new_n7463_;
  wire new_n9357_;
  wire not_new_n625__7;
  wire not_new_n5270_;
  wire new_n2017_;
  wire not_new_n3372__57648010;
  wire po269;
  wire not_new_n631__1;
  wire new_n2369_;
  wire new_n9391_;
  wire new_n2163_;
  wire not_new_n2304_;
  wire new_n7705_;
  wire po024;
  wire not_new_n4014__4;
  wire new_n7574_;
  wire not_new_n6007_;
  wire new_n1601_;
  wire not_new_n10278_;
  wire new_n6410_;
  wire new_n6867_;
  wire not_new_n3315__70;
  wire not_new_n8952_;
  wire new_n1688_;
  wire not_pi006;
  wire new_n6740_;
  wire new_n3713_;
  wire not_new_n9391_;
  wire not_new_n625__3430;
  wire new_n2178_;
  wire new_n5087_;
  wire not_new_n2607_;
  wire new_n4710_;
  wire new_n5339_;
  wire new_n6343_;
  wire new_n6991_;
  wire not_new_n9169_;
  wire not_new_n4502__0;
  wire new_n6440_;
  wire and_and_and_not_pi051_1_not_pi050_1_not_pi049_1_not_pi048_1;
  wire new_n1458_;
  wire not_new_n3206_;
  wire not_new_n5430_;
  wire not_new_n2036_;
  wire not_pi117;
  wire or_or_not_pi269_1_not_pi260_1_not_pi257_1;
  wire new_n4523_;
  wire new_n5293_;
  wire new_n2172_;
  wire new_n3508_;
  wire not_new_n8701_;
  wire new_n591_;
  wire new_n5294_;
  wire new_n3812_;
  wire not_pi058;
  wire new_n2484_;
  wire new_n5204_;
  wire new_n2124_;
  wire not_new_n4707_;
  wire not_new_n6539__1;
  wire not_new_n619__968890104070;
  wire new_n5124_;
  wire not_new_n5041_;
  wire new_n6733_;
  wire or_or_not_new_n6160__not_new_n6161__not_new_n6090_;
  wire not_new_n4805_;
  wire new_n4639_;
  wire new_n5347_;
  wire not_new_n5760_;
  wire not_new_n6993__0;
  wire new_n737_;
  wire not_new_n1006__6;
  wire not_new_n621__3;
  wire not_new_n4575_;
  wire new_n9440_;
  wire new_n5641_;
  wire or_or_not_new_n1251__not_new_n1249__not_new_n1888_;
  wire new_n1759_;
  wire not_new_n1581__19773267430;
  wire not_new_n1063__968890104070;
  wire not_new_n9959__0;
  wire new_n1695_;
  wire new_n7842_;
  wire new_n6046_;
  wire not_new_n3310__10;
  wire not_new_n626__225393402906922580878632490;
  wire new_n1240_;
  wire new_n8631_;
  wire new_n6706_;
  wire not_new_n1826_;
  wire new_n4082_;
  wire not_new_n6038_;
  wire not_new_n3193_;
  wire not_new_n8713__0;
  wire not_new_n9484_;
  wire new_n4197_;
  wire not_new_n6039_;
  wire not_new_n5882__1;
  wire not_new_n4905_;
  wire not_new_n5112_;
  wire new_n5995_;
  wire new_n8041_;
  wire new_n3711_;
  wire not_new_n1597__6782230728490;
  wire not_new_n1067_;
  wire not_new_n1065__70;
  wire new_n6017_;
  wire not_new_n739_;
  wire not_new_n4238_;
  wire not_new_n648_;
  wire new_n5135_;
  wire po164;
  wire new_n6261_;
  wire not_new_n8158__0;
  wire not_new_n1063__1176490;
  wire not_new_n647__24010;
  wire and_new_n1250__new_n1894_;
  wire not_new_n625__3;
  wire and_new_n5268__new_n5267_;
  wire new_n5444_;
  wire new_n8640_;
  wire not_new_n7894_;
  wire new_n3567_;
  wire not_pi064_5585458640832840070;
  wire new_n7202_;
  wire not_new_n8139__1;
  wire not_new_n1569_;
  wire not_new_n8662_;
  wire new_n8196_;
  wire not_new_n3947_;
  wire new_n3441_;
  wire not_new_n7444_;
  wire not_new_n591__8;
  wire new_n5004_;
  wire not_new_n3960_;
  wire po208;
  wire new_n4199_;
  wire not_new_n731__1;
  wire new_n9130_;
  wire new_n3400_;
  wire not_new_n1596__10;
  wire new_n6570_;
  wire new_n9084_;
  wire new_n2522_;
  wire not_new_n3924_;
  wire new_n7609_;
  wire new_n1191_;
  wire not_new_n1504_;
  wire not_new_n603__8;
  wire not_new_n7385_;
  wire not_new_n1267_;
  wire not_new_n741_;
  wire not_new_n596__1176490;
  wire not_new_n633__16284135979104490;
  wire new_n1253_;
  wire not_new_n9402__0;
  wire not_new_n3890_;
  wire not_new_n591__0;
  wire not_new_n642__9;
  wire not_new_n7975_;
  wire not_new_n5846_;
  wire new_n8829_;
  wire not_new_n639__70;
  wire not_new_n1069__0;
  wire new_n2632_;
  wire not_pi135_3;
  wire new_n6146_;
  wire new_n6508_;
  wire new_n3705_;
  wire not_new_n3805_;
  wire not_new_n628__9;
  wire not_new_n1564_;
  wire and_new_n6417__new_n6418_;
  wire not_new_n1596__1915812313805664144010;
  wire not_new_n1613__6782230728490;
  wire new_n7038_;
  wire not_new_n5555_;
  wire not_new_n1567_;
  wire not_new_n5519_;
  wire new_n8297_;
  wire new_n6072_;
  wire not_new_n1538__24010;
  wire new_n10223_;
  wire new_n2090_;
  wire new_n9800_;
  wire new_n5764_;
  wire new_n4042_;
  wire or_not_new_n7316__not_new_n7186_;
  wire not_new_n638__0;
  wire new_n8271_;
  wire not_new_n5724_;
  wire new_n7480_;
  wire not_new_n1611__490;
  wire not_new_n9876_;
  wire not_new_n5477__0;
  wire new_n8060_;
  wire not_new_n4835__1;
  wire not_new_n598__2;
  wire not_new_n989__8;
  wire new_n1704_;
  wire not_new_n754_;
  wire new_n7110_;
  wire not_pi165_1;
  wire new_n8525_;
  wire not_new_n3672_;
  wire not_new_n4462__0;
  wire not_new_n1616__70;
  wire new_n7313_;
  wire new_n8449_;
  wire not_pi176_0;
  wire not_new_n1028__9;
  wire not_new_n9874_;
  wire not_new_n8322__0;
  wire not_new_n7735__2;
  wire new_n7135_;
  wire new_n8686_;
  wire new_n1832_;
  wire not_new_n613__3;
  wire not_pi039_4;
  wire new_n10260_;
  wire or_not_new_n9084__not_new_n9083_;
  wire not_new_n5475__0;
  wire not_new_n2123_;
  wire not_new_n634__24010;
  wire not_pi101_0;
  wire not_new_n8629_;
  wire or_or_or_not_new_n2955__not_new_n2958__not_new_n2957__not_new_n2959_;
  wire new_n5126_;
  wire new_n2151_;
  wire not_new_n7139__1;
  wire not_new_n3315__4;
  wire new_n9046_;
  wire new_n6603_;
  wire new_n5794_;
  wire not_new_n1031__168070;
  wire new_n4558_;
  wire not_new_n7564_;
  wire not_new_n5743_;
  wire not_new_n6476__0;
  wire new_n7593_;
  wire not_new_n7699_;
  wire not_new_n1010__1;
  wire new_n8011_;
  wire new_n7040_;
  wire new_n1512_;
  wire not_new_n728__1;
  wire not_new_n1999_;
  wire not_new_n4097_;
  wire not_new_n9292_;
  wire not_new_n1808_;
  wire new_n8824_;
  wire not_new_n1616__6;
  wire not_new_n607__10;
  wire not_new_n4906_;
  wire not_new_n2876_;
  wire not_po296_0;
  wire not_po296_13410686196639649008070;
  wire not_new_n604__332329305696010;
  wire new_n2407_;
  wire new_n3505_;
  wire not_new_n675_;
  wire not_new_n922_;
  wire new_n662_;
  wire not_new_n7026_;
  wire new_n8562_;
  wire not_new_n9084_;
  wire not_new_n6644__0;
  wire new_n1679_;
  wire not_new_n2748_;
  wire not_new_n621__8235430;
  wire new_n1661_;
  wire new_n3973_;
  wire new_n5051_;
  wire and_new_n6375__new_n6382_;
  wire not_new_n4162_;
  wire new_n1206_;
  wire new_n927_;
  wire or_not_new_n2567__not_new_n2571_;
  wire not_new_n7497_;
  wire new_n5141_;
  wire new_n9159_;
  wire new_n4604_;
  wire and_new_n1542__new_n2371_;
  wire not_new_n9661_;
  wire not_new_n1192_;
  wire not_pi249_2;
  wire new_n8976_;
  wire not_new_n1047__47475615099430;
  wire new_n2908_;
  wire not_new_n4090_;
  wire not_pi057_1;
  wire not_new_n4435__0;
  wire not_new_n6509__0;
  wire or_or_not_new_n2820__not_new_n2823__not_new_n2822_;
  wire new_n9147_;
  wire or_not_new_n2973__not_new_n2976_;
  wire not_new_n7170__0;
  wire not_pi052;
  wire not_new_n6033_;
  wire not_new_n631__39098210485829880490;
  wire new_n4446_;
  wire not_new_n8009_;
  wire not_new_n4276_;
  wire new_n6202_;
  wire not_new_n9065_;
  wire not_new_n609__24010;
  wire not_new_n8595__4;
  wire not_new_n9513_;
  wire new_n8807_;
  wire new_n1872_;
  wire new_n5280_;
  wire not_new_n9714_;
  wire not_new_n596__24010;
  wire not_new_n6659_;
  wire not_new_n627__168070;
  wire new_n6803_;
  wire new_n8685_;
  wire not_new_n581__490;
  wire not_new_n3436_;
  wire new_n5407_;
  wire new_n5080_;
  wire not_new_n8632_;
  wire new_n3573_;
  wire not_new_n1603__5;
  wire not_new_n5304_;
  wire not_new_n4136__0;
  wire new_n6435_;
  wire not_new_n6331_;
  wire new_n7509_;
  wire not_new_n4271_;
  wire not_new_n7409__0;
  wire not_new_n1728__403536070;
  wire new_n1454_;
  wire not_new_n6950_;
  wire not_new_n2166__0;
  wire new_n8436_;
  wire new_n4489_;
  wire not_new_n5457_;
  wire not_new_n10324_;
  wire not_new_n10173_;
  wire not_new_n2732_;
  wire new_n8202_;
  wire new_n4641_;
  wire not_new_n5626_;
  wire new_n5290_;
  wire not_new_n9821_;
  wire new_n6659_;
  wire not_new_n628__5585458640832840070;
  wire not_new_n7449_;
  wire new_n9973_;
  wire not_new_n1600__2;
  wire new_n7468_;
  wire new_n8191_;
  wire new_n4429_;
  wire not_new_n8104__1;
  wire new_n9041_;
  wire not_new_n6375_;
  wire not_pi007_0;
  wire not_new_n1774_;
  wire not_new_n2075_;
  wire not_new_n638__1176490;
  wire new_n3281_;
  wire new_n7942_;
  wire not_new_n10073__0;
  wire or_not_new_n4839__not_new_n4767_;
  wire not_po296_35561530251773635572553173835655155124070416738520070;
  wire new_n2394_;
  wire new_n3955_;
  wire new_n3433_;
  wire new_n8909_;
  wire not_new_n597__4;
  wire not_new_n4638_;
  wire new_n3223_;
  wire not_new_n1781_;
  wire not_new_n628__16284135979104490;
  wire not_new_n1957_;
  wire not_new_n1200_;
  wire not_new_n7002_;
  wire not_new_n7433__1;
  wire not_new_n9050_;
  wire not_new_n7103_;
  wire not_new_n8959_;
  wire new_n1604_;
  wire not_new_n4456__0;
  wire new_n8304_;
  wire new_n9501_;
  wire not_new_n597__57648010;
  wire new_n3296_;
  wire not_new_n1537__16284135979104490;
  wire not_new_n7089_;
  wire not_new_n5754__2;
  wire not_new_n2830_;
  wire not_new_n3918__0;
  wire new_n3866_;
  wire not_new_n639__6782230728490;
  wire new_n2195_;
  wire not_new_n1153__0;
  wire not_new_n7155__1;
  wire new_n9982_;
  wire new_n2147_;
  wire new_n4379_;
  wire new_n7730_;
  wire not_new_n1039__2;
  wire new_n945_;
  wire new_n6405_;
  wire new_n3570_;
  wire new_n5714_;
  wire new_n5233_;
  wire new_n7310_;
  wire not_new_n1585__6782230728490;
  wire not_new_n3529_;
  wire not_new_n3986__0;
  wire not_new_n9942_;
  wire not_new_n1047__3430;
  wire po154;
  wire new_n6170_;
  wire not_new_n3378_;
  wire not_new_n8108__0;
  wire not_new_n9408__0;
  wire po042;
  wire not_pi055_2;
  wire not_new_n8163_;
  wire not_new_n2319_;
  wire new_n6978_;
  wire not_new_n1580__8235430;
  wire not_new_n7447_;
  wire not_new_n1061__16284135979104490;
  wire new_n9639_;
  wire not_new_n1594__4;
  wire new_n6901_;
  wire not_new_n4755_;
  wire not_new_n8413_;
  wire not_new_n599__968890104070;
  wire not_new_n5300_;
  wire not_new_n8422_;
  wire new_n4403_;
  wire new_n6245_;
  wire not_new_n3097_;
  wire not_new_n6325_;
  wire not_pi122;
  wire new_n1029_;
  wire not_new_n1538__0;
  wire new_n7464_;
  wire not_new_n4839_;
  wire not_new_n5006_;
  wire not_new_n646__24010;
  wire or_not_new_n6782__not_new_n6621_;
  wire not_pi254;
  wire new_n7406_;
  wire new_n10043_;
  wire new_n3468_;
  wire new_n9915_;
  wire new_n3712_;
  wire not_new_n9417_;
  wire not_new_n1019__5;
  wire not_new_n635__5;
  wire not_new_n595__2326305139872070;
  wire new_n4577_;
  wire new_n8636_;
  wire new_n9509_;
  wire not_new_n1611__19773267430;
  wire new_n5144_;
  wire not_new_n5742__0;
  wire not_new_n1790_;
  wire not_new_n7534_;
  wire not_new_n3938_;
  wire new_n3412_;
  wire not_new_n735_;
  wire not_new_n1376_;
  wire key_gate_50;
  wire new_n1673_;
  wire or_not_new_n1554__not_new_n2429_;
  wire new_n4670_;
  wire not_new_n10018_;
  wire not_new_n642__403536070;
  wire new_n9134_;
  wire not_pi091;
  wire not_new_n6185_;
  wire new_n1041_;
  wire new_n2006_;
  wire new_n6048_;
  wire not_new_n618__968890104070;
  wire not_new_n1031__9;
  wire new_n937_;
  wire not_new_n7405_;
  wire not_new_n1611__3;
  wire new_n5636_;
  wire not_new_n8688_;
  wire not_new_n9833_;
  wire not_new_n633__57648010;
  wire not_new_n759_;
  wire not_new_n5405_;
  wire new_n8108_;
  wire not_new_n4190_;
  wire not_new_n6977__1;
  wire new_n2049_;
  wire new_n2321_;
  wire new_n6207_;
  wire not_new_n4422__0;
  wire not_new_n1319_;
  wire not_new_n638__3430;
  wire not_new_n5438__0;
  wire not_new_n3172_;
  wire new_n9972_;
  wire not_new_n5915_;
  wire new_n3788_;
  wire new_n6293_;
  wire not_new_n8368__1;
  wire new_n1659_;
  wire not_new_n1043__2326305139872070;
  wire new_n8169_;
  wire not_new_n581__367033682172941254412302110320336601888010;
  wire not_new_n9313_;
  wire not_new_n5717_;
  wire not_new_n10293_;
  wire new_n4179_;
  wire not_new_n1944_;
  wire not_new_n3742_;
  wire not_new_n589__541169560379521116689596608490;
  wire not_new_n723_;
  wire new_n6198_;
  wire not_new_n1035__5;
  wire not_new_n8917_;
  wire or_not_new_n6239__not_new_n6350_;
  wire not_new_n1612__57648010;
  wire not_new_n1602__1176490;
  wire not_new_n3237_;
  wire new_n6661_;
  wire not_new_n4230_;
  wire or_not_new_n3140__not_new_n3139_;
  wire new_n2541_;
  wire new_n6913_;
  wire new_n5463_;
  wire or_not_new_n934__not_new_n933__0;
  wire new_n944_;
  wire not_new_n7931_;
  wire not_new_n4121__1;
  wire new_n3656_;
  wire or_not_new_n1562__not_new_n2469_;
  wire new_n1307_;
  wire new_n4223_;
  wire not_new_n5817_;
  wire not_new_n8869__0;
  wire new_n600_;
  wire new_n5035_;
  wire not_pi099;
  wire not_new_n619__9;
  wire not_new_n7097_;
  wire not_new_n8635_;
  wire not_new_n3573_;
  wire new_n5734_;
  wire new_n1023_;
  wire new_n1357_;
  wire not_new_n8286_;
  wire new_n7912_;
  wire not_new_n1556_;
  wire not_new_n1063__6;
  wire new_n3411_;
  wire new_n7361_;
  wire not_new_n8400_;
  wire new_n3419_;
  wire not_new_n8625_;
  wire new_n9637_;
  wire not_new_n6603_;
  wire not_new_n6479__1;
  wire new_n1565_;
  wire not_new_n5494_;
  wire new_n1554_;
  wire not_new_n1599__2824752490;
  wire new_n9206_;
  wire not_new_n3318_;
  wire not_new_n684_;
  wire not_new_n589__403536070;
  wire not_new_n4770_;
  wire new_n3457_;
  wire not_new_n6538__0;
  wire not_new_n1585__8;
  wire not_new_n4698_;
  wire new_n1999_;
  wire new_n6339_;
  wire not_new_n622__968890104070;
  wire not_new_n635__2;
  wire new_n6689_;
  wire not_new_n640__490;
  wire not_new_n3185__1;
  wire new_n7416_;
  wire new_n4047_;
  wire new_n1284_;
  wire new_n10201_;
  wire not_new_n5496__0;
  wire not_new_n1067__2;
  wire new_n6228_;
  wire not_new_n5593_;
  wire not_new_n7452_;
  wire not_po296_1;
  wire not_new_n4735_;
  wire not_new_n5694_;
  wire new_n8174_;
  wire new_n651_;
  wire not_new_n5891_;
  wire not_new_n7722_;
  wire not_new_n646__138412872010;
  wire new_n2966_;
  wire not_new_n973_;
  wire new_n1935_;
  wire not_new_n3670_;
  wire new_n9585_;
  wire not_new_n8937_;
  wire not_new_n594__7;
  wire new_n7166_;
  wire new_n1754_;
  wire not_new_n7753__0;
  wire not_new_n8553_;
  wire new_n8456_;
  wire not_new_n7041_;
  wire new_n7534_;
  wire not_new_n2890_;
  wire not_new_n9940_;
  wire new_n7184_;
  wire not_new_n3372__113988951853731430;
  wire new_n7049_;
  wire not_new_n9958__0;
  wire new_n1381_;
  wire new_n7697_;
  wire new_n9890_;
  wire new_n8235_;
  wire not_new_n4214_;
  wire new_n4148_;
  wire not_new_n9742_;
  wire new_n6140_;
  wire not_new_n10032__0;
  wire new_n10066_;
  wire not_new_n2851_;
  wire not_new_n9566_;
  wire not_new_n7345__1;
  wire new_n6124_;
  wire not_new_n4134__0;
  wire not_new_n10017_;
  wire new_n9597_;
  wire not_new_n9957__0;
  wire new_n5188_;
  wire not_new_n620__0;
  wire not_new_n9345_;
  wire not_new_n4566_;
  wire new_n8038_;
  wire not_new_n3446_;
  wire new_n9615_;
  wire not_new_n9880_;
  wire new_n8238_;
  wire new_n4777_;
  wire not_pi194;
  wire new_n8089_;
  wire not_new_n5148_;
  wire not_new_n1702_;
  wire not_new_n610__3430;
  wire new_n9959_;
  wire not_new_n1599__490;
  wire not_new_n3814_;
  wire not_new_n1049__332329305696010;
  wire not_new_n3834_;
  wire new_n1372_;
  wire not_new_n1039__6782230728490;
  wire not_new_n639__8235430;
  wire new_n8231_;
  wire not_new_n591__57648010;
  wire new_n3975_;
  wire not_new_n2286_;
  wire new_n5916_;
  wire new_n5760_;
  wire not_new_n10216_;
  wire new_n8248_;
  wire new_n7874_;
  wire new_n6959_;
  wire new_n9616_;
  wire not_new_n10205_;
  wire new_n9950_;
  wire not_new_n3511_;
  wire not_pi060_2;
  wire not_new_n1027__16284135979104490;
  wire new_n8337_;
  wire new_n8476_;
  wire not_new_n1264_;
  wire not_new_n9708_;
  wire po271;
  wire new_n4378_;
  wire new_n9873_;
  wire not_new_n9694_;
  wire not_new_n2963_;
  wire new_n2346_;
  wire not_new_n8841_;
  wire not_new_n9333_;
  wire not_new_n634__1176490;
  wire not_new_n3919_;
  wire not_new_n9195_;
  wire not_pi041;
  wire new_n4108_;
  wire not_new_n1613__4;
  wire and_new_n2414__new_n2413_;
  wire new_n5160_;
  wire not_new_n642__8;
  wire new_n3437_;
  wire new_n770_;
  wire or_or_not_new_n1335__not_new_n1333__not_new_n2287_;
  wire new_n2749_;
  wire not_new_n4201_;
  wire new_n4443_;
  wire not_new_n1355_;
  wire not_new_n5816_;
  wire new_n4999_;
  wire not_new_n627__1;
  wire new_n3979_;
  wire not_new_n5431__0;
  wire not_new_n8959__0;
  wire not_new_n3757_;
  wire not_new_n3443_;
  wire new_n1733_;
  wire not_new_n1051__168070;
  wire not_new_n593__403536070;
  wire not_new_n1260_;
  wire new_n4176_;
  wire not_new_n5092_;
  wire new_n2059_;
  wire new_n5187_;
  wire not_new_n1599__1176490;
  wire not_new_n1581__9;
  wire not_new_n638__273687473400809163430;
  wire not_new_n1579_;
  wire not_new_n6762_;
  wire not_new_n627__6782230728490;
  wire new_n932_;
  wire not_new_n6979__1;
  wire new_n2223_;
  wire new_n8559_;
  wire not_new_n7553_;
  wire not_new_n9080_;
  wire not_new_n9744_;
  wire not_new_n4565_;
  wire new_n7684_;
  wire new_n9255_;
  wire not_new_n1599__3430;
  wire new_n4930_;
  wire not_new_n7053_;
  wire not_new_n1041__8235430;
  wire not_new_n3558_;
  wire not_new_n5045_;
  wire not_new_n6702_;
  wire new_n7333_;
  wire not_new_n9584__0;
  wire not_new_n4065_;
  wire new_n6502_;
  wire new_n1769_;
  wire and_new_n6326__new_n6241_;
  wire not_new_n2714_;
  wire new_n3312_;
  wire not_new_n3372__168070;
  wire new_n9948_;
  wire not_new_n8039_;
  wire not_new_n6728_;
  wire new_n9922_;
  wire not_new_n7512_;
  wire not_new_n5009_;
  wire or_or_not_new_n1555__not_new_n2434__not_new_n1379_;
  wire not_new_n3295_;
  wire new_n5182_;
  wire new_n2264_;
  wire new_n5334_;
  wire new_n5712_;
  wire new_n8270_;
  wire new_n5472_;
  wire not_new_n8472_;
  wire new_n6944_;
  wire not_new_n6999_;
  wire not_new_n6297_;
  wire new_n5875_;
  wire new_n2263_;
  wire not_new_n746_;
  wire new_n5344_;
  wire new_n2919_;
  wire not_new_n644__3430;
  wire not_new_n637__8;
  wire not_new_n9358_;
  wire not_new_n1976__0;
  wire not_new_n635__6;
  wire not_new_n1561_;
  wire not_new_n7002__0;
  wire not_new_n2581_;
  wire new_n5512_;
  wire not_new_n10105_;
  wire not_new_n6110_;
  wire new_n4524_;
  wire not_new_n4116__1;
  wire new_n3972_;
  wire not_new_n9947_;
  wire key_gate_109;
  wire new_n5127_;
  wire not_new_n7468_;
  wire new_n3431_;
  wire new_n5238_;
  wire not_new_n7879_;
  wire new_n6650_;
  wire not_new_n2769_;
  wire new_n5106_;
  wire new_n10281_;
  wire not_new_n6992__1;
  wire not_new_n597__168070;
  wire po035;
  wire new_n8471_;
  wire not_new_n5682_;
  wire new_n2052_;
  wire new_n4575_;
  wire new_n7691_;
  wire not_new_n588__6;
  wire not_new_n5848_;
  wire not_new_n637__2824752490;
  wire not_new_n7538_;
  wire not_new_n2880_;
  wire not_new_n7352_;
  wire new_n6877_;
  wire new_n8744_;
  wire new_n6638_;
  wire not_new_n5649_;
  wire new_n7137_;
  wire not_new_n1057__24010;
  wire not_new_n7824_;
  wire new_n6764_;
  wire new_n3054_;
  wire new_n9904_;
  wire new_n4061_;
  wire not_new_n1538__6;
  wire new_n8425_;
  wire not_new_n7925_;
  wire po214;
  wire not_new_n1069__5;
  wire new_n7686_;
  wire not_new_n10024__0;
  wire not_pi152_0;
  wire not_new_n3126_;
  wire not_new_n6373__3;
  wire not_new_n1941_;
  wire new_n1949_;
  wire not_new_n5641_;
  wire new_n10250_;
  wire new_n1477_;
  wire new_n3282_;
  wire not_new_n1602__4;
  wire new_n9592_;
  wire new_n6833_;
  wire new_n5599_;
  wire new_n7575_;
  wire new_n2631_;
  wire new_n9891_;
  wire not_pi161_1;
  wire not_pi218;
  wire not_pi019;
  wire not_new_n8411_;
  wire new_n7878_;
  wire not_new_n1611__3430;
  wire not_pi055;
  wire not_new_n632__6;
  wire not_new_n10136_;
  wire not_new_n6873_;
  wire not_new_n3538_;
  wire not_new_n7598__0;
  wire not_new_n2040_;
  wire not_new_n8154_;
  wire not_new_n6449_;
  wire new_n1009_;
  wire new_n6950_;
  wire not_new_n8721_;
  wire not_new_n7043_;
  wire new_n8534_;
  wire not_new_n2204_;
  wire new_n1589_;
  wire not_new_n7153_;
  wire not_new_n1605__4;
  wire not_new_n1071_;
  wire not_new_n8248__0;
  wire not_new_n4113__2;
  wire not_new_n6131_;
  wire not_new_n8176_;
  wire not_new_n8085_;
  wire not_new_n6226_;
  wire new_n7112_;
  wire not_new_n625__16284135979104490;
  wire not_new_n4933__0;
  wire not_new_n1596__6;
  wire new_n6778_;
  wire not_new_n8205_;
  wire not_new_n2207_;
  wire not_new_n1309_;
  wire new_n5979_;
  wire not_new_n4114__1;
  wire not_new_n2792_;
  wire new_n6753_;
  wire not_new_n8188_;
  wire not_new_n627__70;
  wire not_new_n593__8235430;
  wire not_new_n5431__1;
  wire not_new_n6483__0;
  wire not_new_n6967_;
  wire new_n608_;
  wire not_new_n7155__0;
  wire new_n4112_;
  wire new_n4326_;
  wire new_n5329_;
  wire new_n5181_;
  wire new_n1582_;
  wire not_new_n8366_;
  wire not_new_n7462_;
  wire not_new_n3405_;
  wire new_n4451_;
  wire and_and_and_new_n6227__new_n6232__new_n6229__new_n6317_;
  wire not_new_n8265__1;
  wire not_new_n9549_;
  wire new_n4027_;
  wire new_n6927_;
  wire not_new_n6649_;
  wire not_new_n4841_;
  wire not_new_n591_;
  wire or_or_not_new_n2587__not_new_n2591__not_new_n1433_;
  wire not_new_n3372__490;
  wire not_new_n3841_;
  wire not_new_n630__39098210485829880490;
  wire new_n8572_;
  wire not_new_n1031__5;
  wire not_new_n5399_;
  wire not_new_n4969_;
  wire new_n8364_;
  wire not_new_n4494_;
  wire not_new_n5451__0;
  wire not_pi124_0;
  wire not_new_n2498_;
  wire not_new_n6739_;
  wire not_pi054_1;
  wire not_new_n1071__70;
  wire new_n10008_;
  wire not_new_n2028_;
  wire not_new_n8860_;
  wire key_gate_78;
  wire not_new_n4433__0;
  wire not_new_n5785_;
  wire new_n3347_;
  wire not_new_n760_;
  wire new_n9937_;
  wire not_new_n5558_;
  wire or_not_new_n5917__not_new_n5719__0;
  wire new_n1022_;
  wire not_new_n10115_;
  wire not_new_n624__5;
  wire new_n3247_;
  wire not_new_n6519__1;
  wire new_n6505_;
  wire not_new_n2955_;
  wire new_n4521_;
  wire po145;
  wire new_n4385_;
  wire new_n2187_;
  wire not_new_n6531__2;
  wire new_n8001_;
  wire not_new_n3855_;
  wire not_new_n6984__1;
  wire new_n9021_;
  wire new_n2602_;
  wire new_n9348_;
  wire new_n4324_;
  wire not_new_n10008_;
  wire not_new_n1047__19773267430;
  wire new_n3220_;
  wire not_new_n9139_;
  wire new_n9337_;
  wire new_n7737_;
  wire new_n8417_;
  wire not_new_n2791_;
  wire new_n3056_;
  wire not_new_n2454_;
  wire not_new_n628_;
  wire new_n5244_;
  wire new_n3047_;
  wire new_n2978_;
  wire new_n7780_;
  wire not_new_n1580__6;
  wire not_new_n606__57648010;
  wire not_new_n1602__70;
  wire not_new_n600__1176490;
  wire new_n6473_;
  wire not_new_n989__1176490;
  wire new_n9864_;
  wire not_new_n9207_;
  wire not_new_n8393_;
  wire not_new_n3434_;
  wire not_new_n9470_;
  wire not_pi249;
  wire not_new_n3185__2824752490;
  wire not_new_n3372__138412872010;
  wire not_new_n3391_;
  wire not_new_n9622_;
  wire not_new_n1602_;
  wire new_n4935_;
  wire not_new_n4469__0;
  wire not_new_n1024__2;
  wire not_new_n7414_;
  wire and_new_n1254__new_n1913_;
  wire not_new_n7151_;
  wire new_n9004_;
  wire not_new_n644__6782230728490;
  wire not_new_n3315__8;
  wire new_n6464_;
  wire new_n4818_;
  wire new_n7281_;
  wire not_new_n648__24010;
  wire new_n5708_;
  wire new_n9140_;
  wire not_new_n4014_;
  wire not_new_n7406_;
  wire not_new_n3999_;
  wire new_n9846_;
  wire not_new_n9511__0;
  wire new_n1171_;
  wire not_new_n1011__8;
  wire key_gate_10;
  wire not_new_n9590_;
  wire not_pi137_0;
  wire new_n6376_;
  wire new_n2206_;
  wire not_new_n4003_;
  wire po000;
  wire not_new_n1065__968890104070;
  wire not_new_n6951_;
  wire new_n4139_;
  wire new_n10182_;
  wire new_n10290_;
  wire new_n9582_;
  wire new_n2588_;
  wire new_n6107_;
  wire not_new_n8265__0;
  wire not_new_n4081_;
  wire not_new_n588__968890104070;
  wire new_n2188_;
  wire not_new_n591__2326305139872070;
  wire new_n9925_;
  wire new_n2736_;
  wire not_new_n637__10;
  wire not_new_n7792_;
  wire not_new_n5507__0;
  wire not_new_n6191_;
  wire not_new_n8134__1;
  wire new_n4477_;
  wire new_n9397_;
  wire not_new_n7603__1;
  wire new_n7400_;
  wire new_n8439_;
  wire not_new_n7626_;
  wire not_new_n7008_;
  wire or_or_not_new_n2597__not_new_n2601__not_new_n1435_;
  wire not_new_n3184__2824752490;
  wire new_n4900_;
  wire not_new_n6459_;
  wire not_new_n5523_;
  wire not_new_n7325_;
  wire new_n8176_;
  wire new_n2105_;
  wire new_n5413_;
  wire not_new_n7950_;
  wire new_n6766_;
  wire or_or_not_new_n2919__not_new_n2922__not_new_n2921_;
  wire new_n9618_;
  wire new_n5348_;
  wire new_n6664_;
  wire new_n6840_;
  wire new_n623_;
  wire new_n3673_;
  wire not_new_n3093_;
  wire not_pi052_0;
  wire new_n5899_;
  wire not_new_n3254_;
  wire new_n5833_;
  wire not_new_n642__7;
  wire not_new_n6986_;
  wire not_new_n7706_;
  wire new_n3995_;
  wire not_po298_1176490;
  wire new_n9694_;
  wire not_new_n9229_;
  wire not_new_n8142_;
  wire not_new_n598__9;
  wire new_n4092_;
  wire not_new_n3525_;
  wire new_n1702_;
  wire and_new_n2124__new_n2127_;
  wire not_new_n1067__2824752490;
  wire not_new_n9336_;
  wire not_new_n635__490;
  wire new_n1598_;
  wire and_new_n2642__new_n2641_;
  wire not_new_n598__1176490;
  wire not_new_n5068_;
  wire new_n9594_;
  wire not_pi145;
  wire new_n10130_;
  wire not_new_n5819_;
  wire new_n1909_;
  wire new_n1770_;
  wire new_n969_;
  wire new_n7222_;
  wire not_new_n3197_;
  wire not_new_n1919_;
  wire not_new_n9893__0;
  wire not_new_n7723_;
  wire new_n7513_;
  wire not_new_n9235_;
  wire not_new_n3962_;
  wire not_new_n1598__968890104070;
  wire new_n722_;
  wire not_new_n9690_;
  wire new_n6116_;
  wire new_n3210_;
  wire new_n5974_;
  wire not_new_n2242_;
  wire new_n1655_;
  wire new_n3429_;
  wire not_new_n10124_;
  wire not_new_n5202_;
  wire or_not_new_n2284__not_new_n2281_;
  wire not_new_n3044_;
  wire not_new_n9602_;
  wire not_new_n736_;
  wire not_new_n6974__4;
  wire not_new_n3806_;
  wire new_n7510_;
  wire new_n4669_;
  wire new_n1842_;
  wire not_new_n1297_;
  wire not_new_n10306_;
  wire new_n3036_;
  wire not_new_n2185_;
  wire not_new_n7331_;
  wire not_new_n7585_;
  wire not_new_n6479__0;
  wire not_new_n9380_;
  wire not_new_n10327_;
  wire new_n2895_;
  wire not_new_n928__47475615099430;
  wire not_new_n6298_;
  wire new_n9318_;
  wire not_new_n1580__2326305139872070;
  wire not_new_n8266__4;
  wire not_new_n10101_;
  wire not_new_n8803_;
  wire new_n8513_;
  wire new_n6942_;
  wire new_n6615_;
  wire new_n9462_;
  wire not_new_n8248_;
  wire new_n7393_;
  wire new_n5638_;
  wire new_n3434_;
  wire not_new_n3927__0;
  wire not_new_n1039__490;
  wire not_new_n1027__4;
  wire not_new_n634__1;
  wire not_new_n1008__3;
  wire new_n9445_;
  wire not_new_n2109__0;
  wire new_n2314_;
  wire not_new_n7257_;
  wire not_new_n4071__3;
  wire new_n10285_;
  wire not_new_n4117__0;
  wire not_new_n588__19773267430;
  wire not_new_n1768__1;
  wire not_new_n599__47475615099430;
  wire not_new_n8417_;
  wire not_new_n6242__4;
  wire new_n2921_;
  wire new_n943_;
  wire new_n2782_;
  wire new_n2920_;
  wire or_not_new_n1557__not_new_n2444_;
  wire new_n9271_;
  wire not_new_n6993_;
  wire not_new_n622__57648010;
  wire new_n673_;
  wire not_new_n6959_;
  wire key_gate_14;
  wire new_n1917_;
  wire new_n1991_;
  wire new_n9804_;
  wire not_new_n3515_;
  wire new_n10276_;
  wire new_n1532_;
  wire not_new_n9901__0;
  wire not_new_n984__3430;
  wire not_new_n6349_;
  wire new_n5914_;
  wire new_n5258_;
  wire not_new_n5690_;
  wire new_n4119_;
  wire not_new_n5031_;
  wire not_new_n9917__0;
  wire not_new_n6477__0;
  wire not_new_n3541_;
  wire new_n8450_;
  wire new_n5176_;
  wire new_n4111_;
  wire not_new_n1588__70;
  wire not_new_n8644_;
  wire new_n4248_;
  wire not_new_n4177_;
  wire not_new_n1485_;
  wire new_n1828_;
  wire or_not_new_n5448__not_new_n5597__1;
  wire not_new_n1007__4;
  wire not_new_n6358_;
  wire new_n4427_;
  wire new_n7390_;
  wire not_new_n1614__0;
  wire not_new_n5912_;
  wire not_new_n1591__57648010;
  wire new_n6090_;
  wire not_new_n594__968890104070;
  wire not_pi033_0;
  wire not_new_n6490_;
  wire not_new_n3724_;
  wire new_n1037_;
  wire not_new_n7242_;
  wire new_n3409_;
  wire not_pi250;
  wire and_and_new_n2257__new_n2260__new_n2258_;
  wire not_new_n6464_;
  wire new_n6914_;
  wire new_n7952_;
  wire not_new_n10063_;
  wire not_new_n3912_;
  wire not_new_n1848_;
  wire not_new_n5379_;
  wire not_new_n6170_;
  wire not_new_n9414_;
  wire not_pi026;
  wire not_new_n591__5585458640832840070;
  wire not_new_n2534_;
  wire not_new_n9910__0;
  wire new_n3501_;
  wire not_new_n608__490;
  wire not_new_n5958_;
  wire not_new_n9412_;
  wire or_not_pi257_3_not_pi260_3;
  wire not_pi014;
  wire not_new_n5787_;
  wire new_n5721_;
  wire new_n6051_;
  wire not_new_n6240_;
  wire not_new_n979_;
  wire new_n10020_;
  wire new_n3911_;
  wire or_not_new_n1024__0_not_new_n3384__2;
  wire not_new_n1793_;
  wire new_n6055_;
  wire not_new_n1546_;
  wire new_n4254_;
  wire not_new_n6583_;
  wire not_new_n8144_;
  wire not_new_n8162__1;
  wire new_n5864_;
  wire not_new_n8713__2;
  wire not_new_n594_;
  wire or_or_not_new_n1557__not_new_n2444__not_new_n1383_;
  wire not_new_n3684_;
  wire new_n8600_;
  wire new_n6729_;
  wire not_new_n2320_;
  wire not_new_n8208_;
  wire not_new_n1537__2;
  wire not_new_n3517_;
  wire not_new_n5805__0;
  wire new_n7750_;
  wire not_new_n2917_;
  wire not_new_n4217_;
  wire not_new_n3500_;
  wire not_pi173_2;
  wire not_new_n1045__16284135979104490;
  wire or_not_new_n5893__0_not_new_n6159__0;
  wire not_new_n581__881247870897231951843937366879128181133112010;
  wire new_n8588_;
  wire new_n6476_;
  wire not_new_n738__0;
  wire new_n9768_;
  wire new_n3215_;
  wire not_new_n5594_;
  wire new_n4041_;
  wire not_new_n609__3430;
  wire new_n4243_;
  wire not_new_n5793__0;
  wire not_new_n6999__1;
  wire not_new_n5737_;
  wire new_n8112_;
  wire or_or_not_new_n6349__not_new_n6373__7_not_new_n1041__490;
  wire new_n2741_;
  wire not_new_n1596__2;
  wire not_new_n3311_;
  wire not_po296_93874803376477543056490;
  wire not_pi260_4;
  wire not_new_n4473__0;
  wire not_new_n9519_;
  wire new_n9227_;
  wire not_new_n6694_;
  wire not_new_n7189_;
  wire not_new_n9679_;
  wire new_n3589_;
  wire new_n4872_;
  wire not_new_n10016_;
  wire not_new_n604__1;
  wire new_n4658_;
  wire not_new_n631__4;
  wire new_n8142_;
  wire not_new_n6168_;
  wire not_new_n1907_;
  wire and_new_n2995__new_n998_;
  wire not_new_n5579_;
  wire not_new_n2808_;
  wire not_new_n4786_;
  wire not_new_n2096_;
  wire new_n6257_;
  wire not_new_n7272_;
  wire not_new_n1065__3;
  wire po095;
  wire not_new_n7732_;
  wire new_n9404_;
  wire new_n2989_;
  wire not_new_n8293_;
  wire or_not_new_n1342__not_new_n1343_;
  wire or_not_new_n2926__not_new_n2925_;
  wire new_n7098_;
  wire not_new_n3734_;
  wire not_new_n8799__0;
  wire new_n4697_;
  wire not_new_n5749__0;
  wire not_new_n680_;
  wire new_n8119_;
  wire new_n7548_;
  wire new_n9014_;
  wire new_n2292_;
  wire not_new_n2923_;
  wire not_new_n6665_;
  wire new_n6377_;
  wire new_n9601_;
  wire not_new_n4133__2;
  wire not_new_n7974_;
  wire not_new_n3778_;
  wire new_n3348_;
  wire new_n994_;
  wire new_n8910_;
  wire new_n1446_;
  wire new_n2331_;
  wire not_new_n4253_;
  wire new_n6449_;
  wire new_n9492_;
  wire new_n2857_;
  wire new_n8759_;
  wire new_n8709_;
  wire new_n5312_;
  wire not_new_n1057__3430;
  wire new_n3527_;
  wire not_new_n5060_;
  wire not_new_n586__1;
  wire not_new_n622__0;
  wire new_n4483_;
  wire not_new_n603__1176490;
  wire new_n6849_;
  wire key_gate_79;
  wire po090;
  wire new_n599_;
  wire new_n6619_;
  wire new_n2448_;
  wire not_new_n1588__4;
  wire not_new_n8532_;
  wire new_n6470_;
  wire new_n8563_;
  wire not_new_n643__332329305696010;
  wire not_new_n7650__0;
  wire not_new_n634__490;
  wire or_not_new_n6508__1_not_new_n6600_;
  wire new_n1021_;
  wire not_new_n8574_;
  wire new_n5671_;
  wire new_n2651_;
  wire not_new_n8219_;
  wire new_n9012_;
  wire not_new_n3669_;
  wire not_new_n7747_;
  wire new_n1202_;
  wire new_n6493_;
  wire new_n1925_;
  wire not_new_n7781_;
  wire not_new_n10107_;
  wire not_new_n5078__3;
  wire new_n8129_;
  wire not_new_n6780_;
  wire not_new_n2509__1176490;
  wire new_n4614_;
  wire not_new_n640__2326305139872070;
  wire po058;
  wire new_n3384_;
  wire not_new_n5275_;
  wire not_pi051_0;
  wire not_new_n1069__6;
  wire not_new_n6723_;
  wire not_new_n1534__490;
  wire not_new_n4113__0;
  wire not_new_n8108_;
  wire not_new_n1053__8;
  wire not_new_n1766_;
  wire not_new_n4809_;
  wire and_new_n1972__new_n1975_;
  wire new_n9600_;
  wire not_new_n9011_;
  wire new_n2286_;
  wire new_n7791_;
  wire new_n9837_;
  wire new_n2576_;
  wire not_new_n751_;
  wire not_new_n8369_;
  wire not_new_n9587_;
  wire not_new_n6124_;
  wire not_new_n5492__0;
  wire not_pi265_1;
  wire not_new_n4233_;
  wire po109;
  wire not_new_n4726_;
  wire not_new_n6526__0;
  wire not_new_n10309_;
  wire new_n5374_;
  wire not_new_n591__2;
  wire not_new_n4515_;
  wire not_new_n6478_;
  wire not_new_n644__47475615099430;
  wire new_n5330_;
  wire not_new_n5496_;
  wire not_new_n4691_;
  wire not_new_n1607__24010;
  wire not_new_n1039__1;
  wire not_new_n7635__0;
  wire not_new_n622__47475615099430;
  wire not_new_n6487__2;
  wire not_new_n1374_;
  wire new_n7344_;
  wire new_n7589_;
  wire not_new_n8098_;
  wire not_new_n1053__403536070;
  wire not_new_n4025_;
  wire new_n6069_;
  wire and_new_n6373__new_n6389_;
  wire not_new_n600__0;
  wire and_new_n6451__new_n6799_;
  wire new_n5640_;
  wire not_new_n1538__403536070;
  wire new_n5016_;
  wire new_n7649_;
  wire new_n3615_;
  wire new_n3830_;
  wire not_new_n9539__0;
  wire new_n2822_;
  wire new_n3677_;
  wire new_n9231_;
  wire not_new_n4664_;
  wire not_new_n10141_;
  wire new_n9054_;
  wire not_new_n3096_;
  wire not_new_n8041_;
  wire not_new_n8788_;
  wire not_new_n6179_;
  wire new_n1414_;
  wire not_new_n1228_;
  wire new_n3059_;
  wire not_new_n600__403536070;
  wire not_new_n5012_;
  wire new_n2456_;
  wire new_n3410_;
  wire not_new_n2899_;
  wire new_n5281_;
  wire new_n6579_;
  wire new_n5170_;
  wire new_n5686_;
  wire new_n4447_;
  wire not_new_n7611__2;
  wire not_new_n9365_;
  wire not_new_n5982_;
  wire not_new_n1576__24010;
  wire not_new_n5395_;
  wire new_n9995_;
  wire not_new_n595__6;
  wire not_new_n603__47475615099430;
  wire new_n9382_;
  wire new_n1854_;
  wire not_new_n3194_;
  wire not_new_n1693_;
  wire new_n2584_;
  wire new_n4668_;
  wire new_n3399_;
  wire new_n8574_;
  wire new_n3279_;
  wire new_n2259_;
  wire not_new_n2115_;
  wire not_new_n7572_;
  wire not_new_n606__1;
  wire new_n6823_;
  wire new_n3273_;
  wire not_new_n1585__1176490;
  wire not_new_n9335_;
  wire not_new_n7917_;
  wire new_n7786_;
  wire not_new_n4459_;
  wire not_new_n4604_;
  wire not_pi147_2;
  wire not_new_n5435__1;
  wire not_new_n2985_;
  wire not_new_n9633_;
  wire new_n4964_;
  wire not_new_n2726_;
  wire new_n9313_;
  wire not_new_n6564_;
  wire not_new_n7648_;
  wire new_n1208_;
  wire not_new_n9036_;
  wire new_n2050_;
  wire new_n8570_;
  wire not_new_n8249_;
  wire not_new_n611__7;
  wire new_n7118_;
  wire new_n5818_;
  wire new_n10224_;
  wire not_new_n3432_;
  wire not_new_n1536__2;
  wire new_n8690_;
  wire not_new_n1558_;
  wire new_n7428_;
  wire new_n1299_;
  wire not_new_n640__70;
  wire new_n4476_;
  wire not_pi257_5;
  wire not_new_n9720_;
  wire not_new_n581__968890104070;
  wire new_n2711_;
  wire not_new_n7284_;
  wire new_n6573_;
  wire new_n7371_;
  wire new_n9170_;
  wire not_new_n1013__0;
  wire not_new_n4779_;
  wire not_new_n7624__0;
  wire not_new_n1607__2;
  wire new_n2519_;
  wire new_n749_;
  wire not_new_n6643_;
  wire not_new_n1594__2;
  wire new_n687_;
  wire not_new_n2294_;
  wire new_n7239_;
  wire new_n3134_;
  wire po285;
  wire not_new_n6576_;
  wire not_new_n7343_;
  wire new_n4430_;
  wire not_new_n8164_;
  wire not_new_n1069__24010;
  wire new_n2752_;
  wire not_new_n4538_;
  wire not_new_n7840_;
  wire not_new_n8833__0;
  wire not_new_n3342_;
  wire new_n5987_;
  wire not_new_n9078_;
  wire not_pi083;
  wire new_n3751_;
  wire not_new_n8805_;
  wire new_n10320_;
  wire not_new_n1607__7;
  wire new_n1197_;
  wire new_n4151_;
  wire not_new_n6635__2;
  wire not_new_n1028_;
  wire not_new_n6712_;
  wire new_n4836_;
  wire not_new_n2796_;
  wire not_new_n1583__57648010;
  wire not_new_n1045__7;
  wire not_new_n597__332329305696010;
  wire new_n9102_;
  wire not_new_n2149_;
  wire new_n2649_;
  wire new_n2098_;
  wire not_new_n2777_;
  wire not_new_n928__5;
  wire not_new_n1631__3430;
  wire po014;
  wire not_new_n6898_;
  wire not_new_n8088_;
  wire new_n8017_;
  wire and_new_n10033__new_n3902_;
  wire not_new_n1589__3;
  wire not_new_n1612__4;
  wire not_new_n3372__1915812313805664144010;
  wire not_new_n2709_;
  wire new_n4029_;
  wire new_n9049_;
  wire not_new_n7277_;
  wire new_n5369_;
  wire not_new_n1043__24010;
  wire new_n8928_;
  wire not_new_n7293_;
  wire new_n4629_;
  wire not_new_n2979_;
  wire not_new_n8113__2;
  wire new_n2620_;
  wire not_new_n8223_;
  wire or_not_new_n2072__not_new_n2073_;
  wire not_new_n6488__0;
  wire not_new_n9589_;
  wire new_n7493_;
  wire or_not_new_n2208__not_new_n2205_;
  wire new_n4436_;
  wire not_new_n9523__1;
  wire not_new_n9097_;
  wire not_new_n1059__7;
  wire not_new_n7739__1;
  wire new_n10098_;
  wire new_n6522_;
  wire new_n2476_;
  wire not_new_n1594__3430;
  wire not_new_n596__968890104070;
  wire not_new_n618__332329305696010;
  wire not_new_n7192_;
  wire not_new_n634__8235430;
  wire not_new_n5928_;
  wire new_n3012_;
  wire new_n7275_;
  wire new_n2073_;
  wire not_new_n1601__5;
  wire not_new_n1170_;
  wire not_new_n3315__57648010;
  wire not_new_n4239_;
  wire not_pi011_0;
  wire not_new_n1039__968890104070;
  wire new_n6421_;
  wire not_new_n5795_;
  wire not_pi119;
  wire not_new_n1537__10;
  wire not_new_n2497_;
  wire not_new_n8132_;
  wire new_n5303_;
  wire not_new_n7458_;
  wire not_new_n1067__2326305139872070;
  wire new_n9686_;
  wire not_new_n1945_;
  wire not_new_n587__16284135979104490;
  wire new_n9610_;
  wire key_gate_96;
  wire not_new_n9410_;
  wire po069;
  wire new_n3927_;
  wire not_new_n4411__0;
  wire or_or_not_new_n1559__not_new_n2454__not_new_n1387_;
  wire new_n7970_;
  wire not_new_n1720_;
  wire new_n8635_;
  wire not_new_n953_;
  wire not_new_n680__0;
  wire new_n2496_;
  wire not_new_n7597__1;
  wire not_new_n5629_;
  wire not_new_n1049__2;
  wire new_n2794_;
  wire not_new_n2966_;
  wire not_new_n7680_;
  wire not_new_n9867__0;
  wire new_n2881_;
  wire new_n1153_;
  wire not_new_n4115__1;
  wire not_new_n1067__168070;
  wire new_n5823_;
  wire new_n5821_;
  wire new_n5557_;
  wire not_new_n7170_;
  wire new_n2834_;
  wire not_new_n5790_;
  wire not_new_n6083_;
  wire not_new_n1596__13410686196639649008070;
  wire new_n3493_;
  wire new_n3707_;
  wire new_n7765_;
  wire not_new_n6709__0;
  wire new_n9291_;
  wire not_new_n9056_;
  wire not_new_n3927_;
  wire not_new_n4001__1;
  wire not_new_n3827_;
  wire new_n10056_;
  wire or_not_new_n2577__not_new_n2581_;
  wire new_n2308_;
  wire or_not_new_n1763__not_new_n1764_;
  wire new_n7896_;
  wire new_n7948_;
  wire not_new_n611__4;
  wire new_n9163_;
  wire not_new_n2479_;
  wire not_new_n2719_;
  wire not_new_n626__8235430;
  wire new_n4365_;
  wire not_new_n8046_;
  wire not_new_n5984__0;
  wire new_n2215_;
  wire not_new_n4154_;
  wire new_n3574_;
  wire new_n10255_;
  wire new_n2116_;
  wire or_not_new_n9694__not_new_n9634_;
  wire not_new_n2078_;
  wire not_new_n642__2326305139872070;
  wire not_new_n6731_;
  wire not_new_n588__797922662976120010;
  wire po049;
  wire new_n10109_;
  wire not_new_n10109_;
  wire not_new_n6161_;
  wire not_pi044_1;
  wire not_new_n4950__0;
  wire not_new_n7388_;
  wire not_new_n646__490;
  wire new_n8729_;
  wire new_n9883_;
  wire not_new_n1576__7;
  wire not_new_n640__168070;
  wire new_n3304_;
  wire not_new_n4470_;
  wire not_new_n5739__0;
  wire new_n3958_;
  wire not_new_n4974__0;
  wire not_new_n1265_;
  wire or_not_new_n2605__not_new_n2604_;
  wire new_n1374_;
  wire new_n3293_;
  wire new_n7087_;
  wire new_n3684_;
  wire not_new_n1537__332329305696010;
  wire new_n4747_;
  wire new_n9372_;
  wire not_new_n638__1915812313805664144010;
  wire not_new_n7179_;
  wire new_n6926_;
  wire new_n2449_;
  wire new_n7257_;
  wire not_new_n4757__0;
  wire not_new_n640__968890104070;
  wire not_new_n2740_;
  wire new_n1302_;
  wire not_new_n689_;
  wire new_n8803_;
  wire not_pi061_1;
  wire new_n10306_;
  wire new_n3130_;
  wire new_n1353_;
  wire new_n7871_;
  wire not_new_n3311__168070;
  wire not_new_n5710_;
  wire not_new_n9624_;
  wire not_new_n7252_;
  wire not_new_n4072_;
  wire not_new_n1329_;
  wire new_n9367_;
  wire not_new_n4204_;
  wire new_n8854_;
  wire new_n2916_;
  wire not_new_n2710_;
  wire not_new_n7716_;
  wire not_new_n3480_;
  wire not_new_n2054_;
  wire not_new_n6233__0;
  wire not_new_n1612__2;
  wire not_new_n5833_;
  wire new_n7086_;
  wire new_n6173_;
  wire new_n10012_;
  wire po138;
  wire new_n9327_;
  wire not_new_n6443__403536070;
  wire new_n3017_;
  wire new_n7191_;
  wire new_n8489_;
  wire new_n4545_;
  wire new_n708_;
  wire not_new_n1597__403536070;
  wire new_n4831_;
  wire new_n7772_;
  wire not_pi170_1;
  wire not_new_n7216_;
  wire not_new_n5823_;
  wire new_n7321_;
  wire not_new_n6104_;
  wire new_n3357_;
  wire new_n5687_;
  wire new_n9250_;
  wire new_n10296_;
  wire not_new_n8271__0;
  wire not_new_n8230_;
  wire not_new_n5514_;
  wire not_new_n7543_;
  wire new_n2473_;
  wire new_n5660_;
  wire new_n9999_;
  wire not_new_n3327_;
  wire new_n5886_;
  wire not_new_n4305_;
  wire new_n1691_;
  wire not_new_n1847_;
  wire not_new_n1611__6782230728490;
  wire new_n3954_;
  wire not_new_n4928_;
  wire new_n2097_;
  wire new_n4246_;
  wire not_new_n9637_;
  wire new_n3014_;
  wire not_new_n2717_;
  wire not_new_n3287_;
  wire not_new_n589__77309937197074445241370944070;
  wire not_new_n1455_;
  wire new_n9983_;
  wire new_n2915_;
  wire not_new_n1425_;
  wire new_n8873_;
  wire not_pi230;
  wire not_new_n603_;
  wire new_n5827_;
  wire and_new_n5938__new_n5933_;
  wire not_new_n632__16284135979104490;
  wire not_new_n8287__0;
  wire not_new_n6008_;
  wire new_n6810_;
  wire not_new_n3384__3;
  wire not_new_n5063__1;
  wire new_n5941_;
  wire not_new_n1728__16284135979104490;
  wire not_new_n596__168070;
  wire new_n5874_;
  wire not_new_n2765_;
  wire not_new_n645__1176490;
  wire not_new_n4292_;
  wire not_new_n4775__0;
  wire not_new_n7321_;
  wire not_new_n8316_;
  wire not_new_n6620_;
  wire new_n1603_;
  wire new_n5230_;
  wire new_n5903_;
  wire new_n9329_;
  wire new_n5741_;
  wire new_n3798_;
  wire new_n7530_;
  wire new_n3820_;
  wire new_n10314_;
  wire not_pi270_0;
  wire not_new_n610__6;
  wire new_n2831_;
  wire new_n4283_;
  wire not_new_n604__6;
  wire new_n4597_;
  wire not_new_n6486__0;
  wire not_new_n4928__0;
  wire new_n10266_;
  wire not_new_n1583__5;
  wire not_new_n603__2824752490;
  wire not_new_n6114_;
  wire po255;
  wire not_new_n8196_;
  wire and_new_n9412__new_n9818_;
  wire not_new_n1018__3;
  wire not_new_n2969_;
  wire not_new_n3931_;
  wire not_new_n601__7;
  wire not_new_n3913__0;
  wire new_n7299_;
  wire new_n5549_;
  wire new_n8394_;
  wire new_n9678_;
  wire new_n9247_;
  wire not_new_n589__1176490;
  wire not_new_n1049__138412872010;
  wire or_not_new_n2847__not_new_n2850_;
  wire not_new_n2190_;
  wire not_new_n5644_;
  wire not_new_n2509__2;
  wire not_new_n1272_;
  wire not_new_n8150__1;
  wire not_new_n591__6;
  wire not_new_n6631__0;
  wire not_new_n3184__8;
  wire not_new_n4157__0;
  wire not_new_n6373_;
  wire not_new_n1596__797922662976120010;
  wire not_new_n2957_;
  wire not_pi023;
  wire new_n7363_;
  wire not_pi260_0;
  wire new_n5498_;
  wire not_new_n3675_;
  wire not_new_n5687_;
  wire not_new_n3310__7;
  wire not_new_n1011__3;
  wire new_n2628_;
  wire new_n4544_;
  wire not_new_n3184__57648010;
  wire not_new_n4293_;
  wire new_n4012_;
  wire new_n6290_;
  wire new_n8430_;
  wire not_new_n8231_;
  wire new_n5523_;
  wire not_new_n2037_;
  wire not_new_n7618__0;
  wire new_n9168_;
  wire not_new_n591__168070;
  wire not_new_n948_;
  wire not_new_n4984_;
  wire not_new_n4441_;
  wire not_new_n8871_;
  wire not_new_n6443__24010;
  wire new_n5420_;
  wire new_n1950_;
  wire not_new_n3932_;
  wire not_new_n9814_;
  wire not_new_n994__1;
  wire new_n3792_;
  wire not_new_n10073_;
  wire not_new_n5733_;
  wire not_new_n8490_;
  wire not_new_n1004__2;
  wire not_new_n1589__70;
  wire new_n6684_;
  wire new_n6909_;
  wire not_new_n7436_;
  wire new_n666_;
  wire not_new_n625__5;
  wire not_new_n591__70;
  wire new_n7295_;
  wire not_new_n5458_;
  wire not_new_n4793__0;
  wire not_pi048_4;
  wire not_new_n600__57648010;
  wire not_pi258;
  wire not_new_n6651_;
  wire not_new_n9447_;
  wire not_new_n4261_;
  wire not_new_n9900__2;
  wire new_n2110_;
  wire not_new_n2225_;
  wire not_new_n7943_;
  wire not_new_n8991__0;
  wire not_new_n2536_;
  wire new_n2936_;
  wire not_new_n1588__403536070;
  wire not_pi142;
  wire not_new_n1920_;
  wire not_new_n9374_;
  wire not_pi132_1;
  wire new_n1410_;
  wire new_n9644_;
  wire new_n8571_;
  wire not_new_n3384__6;
  wire not_new_n6974__70;
  wire not_pi143_1;
  wire new_n1340_;
  wire not_new_n7735_;
  wire not_new_n7713_;
  wire new_n8381_;
  wire po104;
  wire not_new_n1059__0;
  wire and_new_n7662__new_n7994_;
  wire not_new_n8546_;
  wire not_new_n7064_;
  wire not_new_n8596__1;
  wire new_n4814_;
  wire new_n8194_;
  wire not_new_n1728__3430;
  wire not_pi164_2;
  wire new_n8813_;
  wire or_or_not_new_n4240__not_new_n4343__not_new_n704_;
  wire new_n4206_;
  wire not_new_n1584__3;
  wire not_new_n626__39098210485829880490;
  wire not_new_n4825_;
  wire not_new_n7849_;
  wire new_n2868_;
  wire new_n4105_;
  wire not_new_n1051__7;
  wire not_new_n587__3;
  wire new_n714_;
  wire new_n10344_;
  wire not_new_n1008__1;
  wire not_new_n4572_;
  wire not_new_n1611__7;
  wire new_n1199_;
  wire new_n9526_;
  wire new_n9066_;
  wire not_new_n8279_;
  wire not_new_n1018__0;
  wire not_pi118;
  wire new_n8395_;
  wire not_new_n2855_;
  wire not_new_n6154_;
  wire new_n4356_;
  wire new_n1787_;
  wire not_new_n2755_;
  wire not_new_n8129__0;
  wire not_new_n1690_;
  wire not_new_n7947_;
  wire not_new_n4174__0;
  wire new_n8203_;
  wire new_n7043_;
  wire new_n8528_;
  wire not_new_n8630_;
  wire not_new_n4017__0;
  wire new_n2800_;
  wire not_new_n744__0;
  wire new_n1809_;
  wire not_new_n652_;
  wire not_new_n8899__3;
  wire new_n3483_;
  wire new_n2735_;
  wire new_n2796_;
  wire not_new_n8599_;
  wire not_new_n8098__0;
  wire not_new_n9133_;
  wire new_n6079_;
  wire not_new_n1037__57648010;
  wire not_new_n1584__4;
  wire new_n9304_;
  wire new_n8409_;
  wire not_new_n1470_;
  wire not_new_n5445_;
  wire not_new_n6974__8235430;
  wire new_n3269_;
  wire new_n9408_;
  wire not_new_n3926_;
  wire new_n7362_;
  wire not_new_n8109_;
  wire not_new_n8092_;
  wire new_n1931_;
  wire new_n7286_;
  wire new_n1264_;
  wire not_new_n1063__2326305139872070;
  wire not_new_n1530_;
  wire not_pi086;
  wire new_n4788_;
  wire not_new_n604__138412872010;
  wire not_new_n690_;
  wire new_n3477_;
  wire new_n10134_;
  wire not_new_n1161_;
  wire new_n5944_;
  wire new_n8455_;
  wire not_new_n4366_;
  wire not_new_n599__168070;
  wire not_new_n4583_;
  wire not_pi175_2;
  wire new_n9000_;
  wire new_n1960_;
  wire not_new_n9892_;
  wire new_n6300_;
  wire not_new_n1047__70;
  wire not_new_n10183_;
  wire new_n4516_;
  wire not_new_n594__19773267430;
  wire not_new_n4935_;
  wire new_n4200_;
  wire new_n3250_;
  wire not_new_n5774_;
  wire not_new_n6171_;
  wire new_n10100_;
  wire new_n8438_;
  wire new_n9319_;
  wire new_n9971_;
  wire not_new_n6525_;
  wire and_new_n6016__new_n5855_;
  wire not_new_n3362_;
  wire not_new_n1039__5;
  wire new_n7307_;
  wire not_new_n633__168070;
  wire not_new_n1287_;
  wire not_new_n10235_;
  wire not_new_n619__403536070;
  wire new_n9108_;
  wire not_new_n1537__7;
  wire not_new_n627__0;
  wire new_n4425_;
  wire new_n9811_;
  wire not_new_n2109_;
  wire not_new_n626__10;
  wire not_new_n588__490;
  wire new_n6825_;
  wire not_new_n5162_;
  wire not_new_n5686_;
  wire new_n6820_;
  wire new_n8994_;
  wire not_new_n1051__1;
  wire not_new_n7646_;
  wire not_new_n2902_;
  wire new_n3140_;
  wire not_new_n1057__8235430;
  wire not_pi134_0;
  wire not_new_n928__3;
  wire new_n9799_;
  wire not_new_n627__9;
  wire not_new_n5696_;
  wire not_new_n3709_;
  wire not_new_n928__403536070;
  wire new_n10118_;
  wire new_n2852_;
  wire new_n7232_;
  wire new_n5939_;
  wire new_n5613_;
  wire not_new_n617__273687473400809163430;
  wire new_n5988_;
  wire new_n9702_;
  wire not_new_n5199__0;
  wire not_new_n635__6782230728490;
  wire not_new_n10026_;
  wire or_or_not_new_n4933__not_new_n4930__0_not_new_n5322_;
  wire new_n6292_;
  wire not_new_n5978_;
  wire new_n3683_;
  wire not_new_n1583__19773267430;
  wire not_new_n10199_;
  wire not_new_n6893_;
  wire new_n5362_;
  wire not_new_n601__2;
  wire new_n3153_;
  wire not_new_n4159__1;
  wire not_new_n630__7;
  wire new_n3180_;
  wire not_new_n4457_;
  wire or_not_new_n2607__not_new_n2611_;
  wire new_n1788_;
  wire new_n9994_;
  wire not_new_n7446_;
  wire new_n1482_;
  wire not_new_n8370_;
  wire new_n6925_;
  wire not_new_n1601__168070;
  wire new_n9179_;
  wire new_n9691_;
  wire new_n3504_;
  wire new_n758_;
  wire new_n5068_;
  wire not_new_n1536__2326305139872070;
  wire not_new_n3572_;
  wire not_new_n4455__0;
  wire new_n1484_;
  wire not_new_n596__1;
  wire new_n7439_;
  wire not_new_n630__1176490;
  wire not_new_n5654_;
  wire new_n5429_;
  wire new_n9417_;
  wire not_new_n8137__0;
  wire not_new_n6018_;
  wire new_n6186_;
  wire not_new_n8202_;
  wire not_new_n4438_;
  wire not_new_n6328_;
  wire not_pi168;
  wire new_n8762_;
  wire key_gate_63;
  wire not_new_n8595__5;
  wire not_new_n670_;
  wire or_or_not_new_n6363__not_new_n6358__not_new_n6361_;
  wire new_n4719_;
  wire not_new_n9491_;
  wire not_new_n7748_;
  wire or_not_new_n6318__not_new_n6373__0;
  wire not_new_n631__332329305696010;
  wire not_new_n641__9;
  wire not_new_n1590_;
  wire not_new_n642__968890104070;
  wire not_new_n3280_;
  wire not_new_n8875__0;
  wire not_new_n3310__5;
  wire new_n4388_;
  wire new_n1406_;
  wire new_n2841_;
  wire new_n4700_;
  wire not_new_n7735__0;
  wire not_new_n5084__0;
  wire new_n6748_;
  wire not_new_n4082_;
  wire new_n6390_;
  wire not_new_n4534_;
  wire not_new_n1666_;
  wire new_n9316_;
  wire not_new_n5719__0;
  wire not_new_n1708_;
  wire not_new_n4797__1;
  wire new_n7820_;
  wire not_new_n3176_;
  wire new_n9730_;
  wire new_n4207_;
  wire and_new_n8984__new_n9245_;
  wire new_n9307_;
  wire new_n6354_;
  wire not_new_n8158__2;
  wire not_new_n989__332329305696010;
  wire new_n4826_;
  wire not_new_n4136_;
  wire not_new_n1059__57648010;
  wire po189;
  wire new_n776_;
  wire not_new_n5374_;
  wire new_n7578_;
  wire not_new_n5534_;
  wire not_new_n3466_;
  wire not_new_n8134__0;
  wire not_new_n7874_;
  wire new_n8632_;
  wire new_n8077_;
  wire not_new_n3426_;
  wire not_new_n1783_;
  wire not_new_n598__10;
  wire not_pi151;
  wire not_new_n588_;
  wire not_new_n4921_;
  wire not_new_n5424_;
  wire not_new_n628__70;
  wire new_n958_;
  wire new_n10207_;
  wire new_n2810_;
  wire not_new_n4544_;
  wire not_new_n1594__70;
  wire new_n9820_;
  wire new_n9387_;
  wire new_n6411_;
  wire po250;
  wire not_new_n3020_;
  wire or_not_new_n3965__not_new_n3966_;
  wire not_new_n4455_;
  wire not_new_n3177_;
  wire not_new_n6769_;
  wire not_new_n9946__0;
  wire new_n10176_;
  wire new_n9441_;
  wire not_new_n6635_;
  wire new_n1341_;
  wire new_n7940_;
  wire or_not_new_n2903__not_new_n1483_;
  wire new_n3195_;
  wire new_n4632_;
  wire po120;
  wire new_n4526_;
  wire and_new_n1915__new_n1918_;
  wire not_new_n6040_;
  wire or_not_new_n2872__not_new_n2871_;
  wire new_n9468_;
  wire new_n2912_;
  wire new_n735_;
  wire not_new_n6964_;
  wire new_n3511_;
  wire new_n9569_;
  wire key_gate_62;
  wire not_new_n8538_;
  wire new_n9311_;
  wire not_new_n9337_;
  wire not_new_n4310_;
  wire not_new_n4117_;
  wire not_new_n4414__0;
  wire new_n5948_;
  wire new_n4235_;
  wire new_n5216_;
  wire not_new_n5238_;
  wire not_new_n6974__168070;
  wire not_new_n9173_;
  wire new_n8393_;
  wire not_new_n6465_;
  wire not_pi172_2;
  wire not_new_n648__2;
  wire not_new_n4765__0;
  wire new_n5383_;
  wire new_n5853_;
  wire not_new_n1067__6782230728490;
  wire new_n2805_;
  wire new_n2693_;
  wire not_new_n1600__7;
  wire new_n8818_;
  wire new_n2053_;
  wire new_n4259_;
  wire new_n5980_;
  wire not_new_n646__57648010;
  wire new_n9505_;
  wire not_new_n636__3;
  wire not_new_n5229_;
  wire new_n2389_;
  wire not_new_n4464_;
  wire new_n7064_;
  wire new_n5953_;
  wire not_new_n587__138412872010;
  wire new_n10343_;
  wire new_n8772_;
  wire not_new_n1631__797922662976120010;
  wire not_new_n647__7;
  wire not_new_n5631_;
  wire new_n7288_;
  wire new_n8149_;
  wire new_n7741_;
  wire new_n10029_;
  wire not_new_n9845_;
  wire not_new_n8984__0;
  wire not_new_n1049_;
  wire not_new_n616_;
  wire not_new_n1529_;
  wire new_n3668_;
  wire not_new_n619__6;
  wire not_new_n1063__24010;
  wire new_n2196_;
  wire not_new_n4951__0;
  wire new_n6544_;
  wire not_new_n5083__0;
  wire not_new_n5868_;
  wire new_n5161_;
  wire not_new_n1607__3430;
  wire new_n5527_;
  wire new_n9383_;
  wire not_new_n644__19773267430;
  wire new_n10160_;
  wire not_new_n3799_;
  wire new_n8095_;
  wire not_new_n4898_;
  wire new_n3983_;
  wire not_new_n6290_;
  wire new_n7619_;
  wire new_n8087_;
  wire new_n7335_;
  wire new_n5023_;
  wire not_pi033_4;
  wire not_new_n1011__4;
  wire new_n8237_;
  wire not_new_n4964_;
  wire not_new_n7360_;
  wire new_n1834_;
  wire new_n7500_;
  wire not_new_n7932__0;
  wire not_new_n2345__0;
  wire key_gate_19;
  wire new_n4574_;
  wire or_not_new_n4843__not_new_n4757_;
  wire not_new_n5285_;
  wire not_new_n5803__0;
  wire not_new_n1534__0;
  wire not_new_n4723__0;
  wire not_new_n6337_;
  wire new_n9094_;
  wire not_pi162_1;
  wire new_n3326_;
  wire new_n5059_;
  wire new_n4187_;
  wire new_n7875_;
  wire not_new_n7240_;
  wire new_n9195_;
  wire not_new_n7056_;
  wire not_pi106_0;
  wire not_new_n8564_;
  wire new_n1683_;
  wire new_n1555_;
  wire new_n4314_;
  wire new_n9602_;
  wire new_n7326_;
  wire new_n7541_;
  wire not_new_n3413_;
  wire new_n8218_;
  wire new_n8590_;
  wire not_new_n4427_;
  wire not_new_n1595__0;
  wire not_new_n1612__47475615099430;
  wire new_n5371_;
  wire not_new_n617__6782230728490;
  wire new_n6054_;
  wire new_n3109_;
  wire new_n1860_;
  wire new_n4244_;
  wire not_new_n624__4;
  wire not_new_n587__57648010;
  wire not_new_n9967_;
  wire new_n9188_;
  wire new_n762_;
  wire new_n3644_;
  wire new_n1149_;
  wire not_new_n6840_;
  wire not_pi065_0;
  wire not_pi249_1;
  wire not_new_n8321_;
  wire new_n2754_;
  wire not_new_n775__168070;
  wire not_new_n1603__2;
  wire not_new_n643__1;
  wire not_new_n6896_;
  wire new_n3602_;
  wire not_new_n1728__57648010;
  wire not_pi165_2;
  wire not_new_n631__3430;
  wire new_n6876_;
  wire not_new_n4994__0;
  wire or_not_new_n6817__not_new_n6788_;
  wire new_n4703_;
  wire not_new_n1027_;
  wire po093;
  wire not_new_n643__797922662976120010;
  wire not_new_n601__403536070;
  wire not_new_n4680_;
  wire new_n9234_;
  wire new_n5071_;
  wire not_new_n1057__490;
  wire new_n1424_;
  wire new_n4396_;
  wire new_n2479_;
  wire not_new_n604_;
  wire new_n3002_;
  wire new_n5928_;
  wire or_not_new_n1255__not_new_n1253_;
  wire not_new_n6555_;
  wire new_n1863_;
  wire new_n3542_;
  wire new_n7641_;
  wire po030;
  wire not_pi173_3;
  wire not_new_n691_;
  wire new_n7527_;
  wire not_new_n6541__0;
  wire new_n5718_;
  wire key_gate_77;
  wire not_new_n5447__0;
  wire not_new_n8528_;
  wire not_new_n1053__16284135979104490;
  wire not_new_n5807__1;
  wire new_n7612_;
  wire new_n9793_;
  wire not_new_n3310__3;
  wire not_new_n4166_;
  wire new_n6452_;
  wire not_new_n633__6;
  wire new_n9533_;
  wire new_n8048_;
  wire new_n8296_;
  wire not_new_n1051__2;
  wire new_n7627_;
  wire new_n9432_;
  wire new_n4308_;
  wire not_new_n5456_;
  wire or_or_not_new_n2785__not_new_n2788__not_new_n2787_;
  wire new_n2957_;
  wire new_n7172_;
  wire new_n3473_;
  wire not_new_n6923_;
  wire not_new_n6636_;
  wire new_n613_;
  wire not_new_n1601__138412872010;
  wire not_new_n2861_;
  wire new_n7564_;
  wire not_new_n4824_;
  wire not_new_n1300_;
  wire not_new_n585__968890104070;
  wire not_new_n8086_;
  wire new_n8477_;
  wire not_new_n588__2824752490;
  wire and_new_n3055__new_n998_;
  wire not_new_n3240_;
  wire not_new_n3121_;
  wire not_new_n9201_;
  wire new_n1866_;
  wire new_n2309_;
  wire new_n5486_;
  wire not_new_n624__2;
  wire new_n10034_;
  wire not_new_n1041__138412872010;
  wire new_n6972_;
  wire not_new_n3398_;
  wire and_new_n2394__new_n2393_;
  wire not_new_n3425_;
  wire new_n652_;
  wire new_n6838_;
  wire not_new_n1537__47475615099430;
  wire not_new_n1257_;
  wire new_n2460_;
  wire not_new_n9968__0;
  wire not_pi058_1;
  wire not_new_n8289__0;
  wire not_new_n726_;
  wire new_n1927_;
  wire not_new_n6850_;
  wire not_new_n612__4;
  wire new_n3065_;
  wire not_new_n1071__2824752490;
  wire new_n1651_;
  wire new_n10172_;
  wire not_new_n984__138412872010;
  wire not_new_n631__4599865365447399609768010;
  wire not_new_n3185__3430;
  wire not_new_n6054_;
  wire new_n5055_;
  wire new_n6907_;
  wire new_n5197_;
  wire not_new_n3103_;
  wire not_new_n4413_;
  wire new_n9652_;
  wire new_n4172_;
  wire not_new_n6021_;
  wire new_n3502_;
  wire not_new_n5775_;
  wire not_new_n7450_;
  wire not_new_n1585__5;
  wire not_new_n2575_;
  wire not_new_n4754_;
  wire not_new_n9072_;
  wire not_new_n1160__0;
  wire not_new_n1589__2326305139872070;
  wire new_n9128_;
  wire not_new_n628__13410686196639649008070;
  wire or_not_new_n1561__not_new_n2464_;
  wire new_n1015_;
  wire not_new_n9587__0;
  wire not_new_n1035__7;
  wire new_n1932_;
  wire po100;
  wire new_n5545_;
  wire not_new_n3230_;
  wire not_pi252_1;
  wire not_po298_1;
  wire new_n718_;
  wire not_new_n8639_;
  wire not_new_n6443_;
  wire new_n3369_;
  wire new_n6765_;
  wire not_new_n7841_;
  wire new_n4810_;
  wire new_n4091_;
  wire or_or_not_new_n2034__not_new_n2035__not_new_n2037_;
  wire not_new_n8737_;
  wire new_n4586_;
  wire new_n9741_;
  wire new_n1156_;
  wire new_n8666_;
  wire new_n5881_;
  wire not_new_n598__4;
  wire not_new_n4148_;
  wire new_n2608_;
  wire not_new_n7366__0;
  wire not_new_n9599_;
  wire new_n8778_;
  wire new_n3372_;
  wire new_n5908_;
  wire not_new_n5447__1;
  wire not_pi048_3;
  wire not_pi135_0;
  wire not_new_n8873_;
  wire not_new_n1583__8235430;
  wire and_and_new_n8692__new_n8691__new_n8695_;
  wire new_n2685_;
  wire not_new_n951_;
  wire not_new_n3239_;
  wire new_n5461_;
  wire new_n2269_;
  wire not_new_n657_;
  wire new_n10062_;
  wire not_new_n5484_;
  wire not_new_n7763_;
  wire not_new_n9312_;
  wire not_new_n10303_;
  wire not_new_n8004_;
  wire new_n1795_;
  wire not_new_n1601__6782230728490;
  wire new_n1360_;
  wire not_new_n591__113988951853731430;
  wire not_new_n10029_;
  wire not_new_n3333_;
  wire not_new_n1616__3430;
  wire new_n1324_;
  wire new_n3811_;
  wire new_n9939_;
  wire not_new_n604__2;
  wire not_new_n1600__24010;
  wire not_new_n1584__10;
  wire new_n7360_;
  wire new_n7987_;
  wire not_new_n1362_;
  wire not_new_n10342_;
  wire not_new_n8337_;
  wire not_pi056_0;
  wire new_n2765_;
  wire new_n7802_;
  wire not_new_n4579_;
  wire new_n10104_;
  wire not_new_n1589__1;
  wire not_pi039_2;
  wire not_new_n5221_;
  wire not_new_n1009__7;
  wire new_n7677_;
  wire not_new_n8529_;
  wire not_new_n3281_;
  wire new_n10229_;
  wire not_new_n5776__0;
  wire new_n9598_;
  wire not_new_n9367_;
  wire not_new_n9285_;
  wire not_new_n7570_;
  wire new_n10175_;
  wire not_new_n9950__0;
  wire new_n6459_;
  wire not_new_n5791__0;
  wire not_new_n8149_;
  wire new_n4725_;
  wire and_new_n5097__new_n5098_;
  wire not_new_n7820_;
  wire po053;
  wire and_new_n1541__new_n2366_;
  wire not_new_n3338_;
  wire not_new_n2621_;
  wire not_new_n5871_;
  wire new_n1839_;
  wire or_not_new_n1279__not_new_n1277_;
  wire new_n8961_;
  wire not_new_n6822_;
  wire not_new_n608__7;
  wire new_n2644_;
  wire not_new_n6351_;
  wire not_new_n1375_;
  wire not_pi043_0;
  wire new_n5716_;
  wire new_n5263_;
  wire not_new_n9261_;
  wire not_new_n7521_;
  wire new_n1230_;
  wire not_new_n4700_;
  wire not_new_n6064_;
  wire not_new_n5678_;
  wire not_new_n9107_;
  wire new_n5061_;
  wire new_n1887_;
  wire not_new_n623__6;
  wire key_gate_29;
  wire not_new_n9464_;
  wire not_new_n3504_;
  wire not_new_n3545_;
  wire new_n7264_;
  wire not_pi043;
  wire not_new_n9437_;
  wire new_n3740_;
  wire not_new_n5800__0;
  wire new_n3533_;
  wire not_pi060_1;
  wire not_new_n9022_;
  wire new_n2689_;
  wire not_new_n4899__0;
  wire not_new_n5693_;
  wire not_new_n1017__0;
  wire new_n3608_;
  wire not_new_n8991_;
  wire not_new_n3532_;
  wire not_new_n618__8235430;
  wire not_new_n6492_;
  wire not_new_n3265_;
  wire not_new_n1027__5;
  wire new_n6836_;
  wire new_n1176_;
  wire new_n2240_;
  wire new_n8432_;
  wire not_new_n5893__0;
  wire not_new_n1651_;
  wire new_n3517_;
  wire not_new_n3038_;
  wire new_n1732_;
  wire new_n2038_;
  wire new_n7917_;
  wire not_new_n8868_;
  wire not_new_n1527_;
  wire new_n1849_;
  wire not_new_n6938_;
  wire key_gate_60;
  wire not_new_n1019__2;
  wire new_n1344_;
  wire not_new_n1204_;
  wire not_new_n618__5585458640832840070;
  wire not_new_n7285_;
  wire not_new_n676_;
  wire new_n5162_;
  wire new_n9772_;
  wire new_n5849_;
  wire new_n6585_;
  wire new_n7494_;
  wire not_new_n8118__1;
  wire new_n6692_;
  wire new_n10256_;
  wire not_new_n3479_;
  wire new_n9280_;
  wire not_new_n586__138412872010;
  wire new_n656_;
  wire not_new_n5905__0;
  wire not_new_n8147__0;
  wire not_new_n597__8235430;
  wire not_new_n608__2;
  wire new_n9934_;
  wire new_n10019_;
  wire new_n4457_;
  wire not_new_n645__57648010;
  wire not_new_n1601__968890104070;
  wire new_n3786_;
  wire not_new_n587__6;
  wire not_new_n6525__0;
  wire new_n5878_;
  wire and_and_new_n1839__new_n1842__new_n1840_;
  wire new_n7590_;
  wire not_new_n9249_;
  wire not_new_n6043_;
  wire not_new_n7709_;
  wire new_n8136_;
  wire not_new_n5351_;
  wire new_n1401_;
  wire new_n5541_;
  wire not_new_n10067_;
  wire not_new_n6510__0;
  wire not_new_n609__168070;
  wire not_new_n2656_;
  wire not_new_n6600_;
  wire not_new_n3302_;
  wire new_n3371_;
  wire not_new_n5900__1;
  wire not_new_n8211_;
  wire new_n4154_;
  wire new_n9152_;
  wire new_n1792_;
  wire not_new_n4687_;
  wire new_n5239_;
  wire not_new_n8973__0;
  wire not_new_n10114_;
  wire not_new_n1580__168070;
  wire new_n1972_;
  wire new_n8040_;
  wire not_new_n5780_;
  wire not_new_n970_;
  wire not_new_n4461_;
  wire not_pi154_0;
  wire not_pi034_0;
  wire new_n6997_;
  wire new_n7569_;
  wire not_new_n607__490;
  wire not_new_n8496_;
  wire not_new_n1925_;
  wire new_n8500_;
  wire new_n3163_;
  wire new_n6315_;
  wire new_n7818_;
  wire new_n5236_;
  wire new_n7729_;
  wire not_new_n1061__3430;
  wire new_n7284_;
  wire not_new_n621__16284135979104490;
  wire new_n8398_;
  wire not_new_n625__39098210485829880490;
  wire not_new_n8743_;
  wire new_n1528_;
  wire new_n7432_;
  wire not_new_n2527_;
  wire not_new_n3026_;
  wire new_n9822_;
  wire new_n9542_;
  wire new_n6418_;
  wire new_n4961_;
  wire not_new_n928__168070;
  wire or_or_not_new_n1782__not_new_n1783__not_new_n1785_;
  wire not_new_n1596__403536070;
  wire new_n7094_;
  wire new_n9776_;
  wire not_new_n1599__7;
  wire not_new_n5767_;
  wire not_new_n665_;
  wire not_new_n3000_;
  wire not_new_n6103_;
  wire not_new_n7361_;
  wire new_n2642_;
  wire new_n4950_;
  wire new_n5319_;
  wire not_new_n2322_;
  wire not_new_n1598__9;
  wire not_new_n5385_;
  wire not_new_n647__8;
  wire new_n6964_;
  wire not_new_n9372__0;
  wire and_new_n1266__new_n1970_;
  wire not_new_n7627__1;
  wire not_new_n2571_;
  wire not_new_n5099_;
  wire new_n5078_;
  wire not_new_n644__5585458640832840070;
  wire not_new_n6077_;
  wire not_new_n5092__0;
  wire new_n3308_;
  wire new_n8696_;
  wire and_new_n4403__new_n4407_;
  wire not_new_n601__490;
  wire not_new_n8165__0;
  wire new_n9856_;
  wire new_n2762_;
  wire not_new_n6321_;
  wire not_new_n1012__3;
  wire new_n1978_;
  wire not_new_n4417_;
  wire new_n3299_;
  wire not_new_n4724__0;
  wire new_n617_;
  wire new_n5490_;
  wire new_n8838_;
  wire not_new_n9787_;
  wire not_new_n714_;
  wire po031;
  wire not_new_n1534__24010;
  wire not_new_n5373_;
  wire not_new_n5554_;
  wire not_new_n648__8235430;
  wire new_n9144_;
  wire new_n9091_;
  wire not_new_n8523_;
  wire new_n3879_;
  wire new_n4255_;
  wire not_new_n8425_;
  wire not_new_n8893_;
  wire not_new_n9357__0;
  wire not_new_n7428_;
  wire not_new_n6527__0;
  wire new_n7488_;
  wire not_new_n5738_;
  wire not_new_n1761_;
  wire not_new_n1016_;
  wire not_new_n1063__138412872010;
  wire key_gate_45;
  wire not_new_n583__0;
  wire not_new_n8870__0;
  wire new_n6120_;
  wire new_n8780_;
  wire new_n7454_;
  wire new_n9019_;
  wire not_new_n3900_;
  wire not_new_n3754_;
  wire new_n6241_;
  wire new_n5343_;
  wire new_n1967_;
  wire new_n2751_;
  wire new_n9649_;
  wire or_not_new_n9523__1_not_new_n9327__1;
  wire not_new_n9746_;
  wire new_n6265_;
  wire not_new_n8252_;
  wire not_new_n5165_;
  wire po181;
  wire key_gate_65;
  wire new_n1669_;
  wire not_new_n8105__1;
  wire not_new_n1585__968890104070;
  wire not_new_n1617__0;
  wire not_new_n626__1577753820348458066150427430;
  wire new_n4050_;
  wire not_new_n3933_;
  wire not_new_n589__3430;
  wire not_new_n4767_;
  wire not_new_n4782__0;
  wire or_or_not_pi269_2_not_pi248_2_not_pi257_2;
  wire new_n8703_;
  wire new_n5306_;
  wire not_new_n1606__2;
  wire new_n7883_;
  wire not_new_n1584__168070;
  wire new_n4952_;
  wire new_n9788_;
  wire not_pi117_0;
  wire new_n3075_;
  wire new_n9761_;
  wire not_new_n4798__0;
  wire not_new_n719__1;
  wire not_new_n1728__6782230728490;
  wire new_n2934_;
  wire new_n3144_;
  wire not_new_n928__9;
  wire new_n1855_;
  wire not_new_n2210_;
  wire new_n2977_;
  wire not_new_n1006__0;
  wire not_new_n6912_;
  wire new_n5957_;
  wire not_new_n5741_;
  wire not_new_n6517__0;
  wire new_n9043_;
  wire not_new_n3858_;
  wire new_n8441_;
  wire new_n7990_;
  wire not_new_n1055__403536070;
  wire not_new_n1807_;
  wire new_n1335_;
  wire not_new_n6520_;
  wire new_n7466_;
  wire new_n2510_;
  wire not_new_n613_;
  wire not_new_n9109_;
  wire new_n2941_;
  wire new_n9607_;
  wire not_pi174;
  wire new_n5666_;
  wire not_new_n9933__0;
  wire not_new_n1069__70;
  wire not_new_n2349_;
  wire new_n9204_;
  wire new_n6969_;
  wire not_new_n2774_;
  wire not_new_n8874__1;
  wire not_new_n2509__3430;
  wire not_new_n597_;
  wire new_n1647_;
  wire new_n3038_;
  wire new_n5231_;
  wire new_n6222_;
  wire new_n7908_;
  wire new_n10239_;
  wire not_new_n1612__3430;
  wire not_new_n642__16284135979104490;
  wire new_n955_;
  wire not_new_n9668_;
  wire new_n1689_;
  wire new_n2684_;
  wire not_new_n752_;
  wire and_new_n6673__new_n6668_;
  wire not_new_n1996_;
  wire not_new_n4114__0;
  wire not_new_n3459_;
  wire not_new_n581__6;
  wire not_new_n596__3430;
  wire new_n7661_;
  wire not_new_n591__403536070;
  wire new_n7433_;
  wire not_pi063_0;
  wire not_new_n2299__0;
  wire not_new_n1045__70;
  wire not_new_n7677_;
  wire key_gate_13;
  wire new_n7009_;
  wire not_new_n9429_;
  wire new_n2343_;
  wire not_new_n1583__113988951853731430;
  wire new_n6970_;
  wire not_new_n6317_;
  wire new_n8665_;
  wire not_new_n4761_;
  wire not_new_n587__8235430;
  wire not_new_n1601__1;
  wire not_new_n8911_;
  wire not_new_n2116_;
  wire new_n4236_;
  wire not_new_n1320_;
  wire new_n6917_;
  wire new_n8281_;
  wire not_new_n1606__5;
  wire not_new_n4033_;
  wire new_n719_;
  wire not_new_n7790_;
  wire not_new_n4741_;
  wire not_new_n1596__39098210485829880490;
  wire new_n5808_;
  wire new_n8831_;
  wire new_n4462_;
  wire new_n6084_;
  wire not_new_n9026_;
  wire new_n8613_;
  wire not_new_n9625__0;
  wire new_n6656_;
  wire new_n9985_;
  wire not_new_n1938__0;
  wire po165;
  wire not_new_n8576_;
  wire not_new_n7439__1;
  wire not_new_n7640__0;
  wire not_new_n4839__1;
  wire new_n9734_;
  wire new_n2101_;
  wire new_n6134_;
  wire new_n2357_;
  wire not_new_n2822_;
  wire new_n10210_;
  wire not_new_n4351__0;
  wire not_new_n1603__10;
  wire not_new_n8136_;
  wire not_new_n600__9;
  wire not_new_n7307_;
  wire new_n7813_;
  wire new_n8396_;
  wire not_new_n626__19773267430;
  wire new_n9277_;
  wire not_new_n4524_;
  wire new_n5038_;
  wire new_n7666_;
  wire new_n8250_;
  wire new_n5180_;
  wire new_n8173_;
  wire not_new_n4277_;
  wire not_new_n2968_;
  wire new_n3074_;
  wire not_new_n3350_;
  wire not_new_n928__968890104070;
  wire not_new_n5432__0;
  wire not_new_n6208_;
  wire not_new_n9512__1;
  wire po259;
  wire new_n8979_;
  wire not_new_n1037__8;
  wire new_n7804_;
  wire new_n8555_;
  wire new_n8546_;
  wire not_new_n4931_;
  wire new_n4714_;
  wire new_n7764_;
  wire not_pi032;
  wire new_n8326_;
  wire new_n9654_;
  wire not_new_n1031__19773267430;
  wire not_new_n6074_;
  wire not_new_n928__8235430;
  wire new_n8266_;
  wire not_new_n1053__19773267430;
  wire not_new_n5630_;
  wire not_new_n8133__0;
  wire new_n5653_;
  wire not_new_n6622_;
  wire new_n9858_;
  wire new_n3121_;
  wire not_new_n2856_;
  wire new_n8820_;
  wire not_new_n8945_;
  wire not_new_n9326_;
  wire not_new_n4466__0;
  wire not_new_n621__70;
  wire new_n1676_;
  wire not_new_n722_;
  wire new_n8797_;
  wire new_n6412_;
  wire not_new_n1584__19773267430;
  wire not_po296_273687473400809163430;
  wire not_new_n5298_;
  wire new_n4733_;
  wire not_new_n7033__0;
  wire or_not_new_n5463__not_new_n5680__1;
  wire new_n2225_;
  wire new_n686_;
  wire new_n4102_;
  wire new_n2537_;
  wire not_new_n8947_;
  wire not_new_n5248_;
  wire new_n4576_;
  wire not_new_n4171_;
  wire not_new_n581__93874803376477543056490;
  wire not_new_n8135__0;
  wire new_n4276_;
  wire new_n6952_;
  wire not_new_n3467_;
  wire new_n6357_;
  wire not_new_n3752_;
  wire not_new_n7934__0;
  wire not_new_n7863__0;
  wire new_n9467_;
  wire not_new_n7750_;
  wire not_new_n1728__168070;
  wire new_n6744_;
  wire new_n6812_;
  wire not_new_n6002_;
  wire or_not_new_n9361__not_new_n9358__0;
  wire new_n1919_;
  wire new_n5022_;
  wire new_n7628_;
  wire not_new_n5891__0;
  wire not_new_n10104_;
  wire new_n6486_;
  wire not_new_n629__1;
  wire or_not_new_n5291__not_new_n5290_;
  wire not_new_n3147_;
  wire new_n6679_;
  wire not_new_n9646_;
  wire not_new_n1604__16284135979104490;
  wire and_new_n8723__new_n1174_;
  wire not_new_n1631__4;
  wire not_new_n3184__332329305696010;
  wire not_new_n9503_;
  wire new_n1520_;
  wire not_new_n1353_;
  wire not_new_n10001_;
  wire new_n6364_;
  wire not_new_n7313_;
  wire new_n8522_;
  wire not_new_n9809_;
  wire not_new_n5728_;
  wire not_new_n1576__1176490;
  wire not_new_n5028_;
  wire not_new_n4128__0;
  wire new_n6399_;
  wire not_new_n8818_;
  wire not_new_n741__0;
  wire not_pi149_0;
  wire new_n7857_;
  wire and_new_n2048__new_n2051_;
  wire not_new_n944_;
  wire new_n10057_;
  wire not_new_n9523__0;
  wire new_n4193_;
  wire not_new_n1071__10;
  wire new_n6583_;
  wire not_new_n7599__1;
  wire not_new_n6953_;
  wire new_n2542_;
  wire not_new_n2209_;
  wire new_n6340_;
  wire not_new_n5186_;
  wire new_n2302_;
  wire not_new_n8443__0;
  wire new_n3815_;
  wire new_n4331_;
  wire new_n5670_;
  wire not_new_n7606__0;
  wire new_n4897_;
  wire po194;
  wire not_new_n601__9;
  wire and_new_n1451__new_n2679_;
  wire new_n6935_;
  wire not_new_n8431_;
  wire new_n7816_;
  wire new_n5091_;
  wire new_n6328_;
  wire new_n2033_;
  wire new_n10078_;
  wire new_n6044_;
  wire not_new_n6998_;
  wire new_n9980_;
  wire not_new_n9628_;
  wire not_new_n5770_;
  wire not_new_n8949_;
  wire not_new_n10113_;
  wire not_new_n4080_;
  wire not_new_n4222_;
  wire not_new_n9613_;
  wire not_new_n9402_;
  wire new_n2502_;
  wire not_new_n630__70;
  wire new_n8103_;
  wire not_new_n4194_;
  wire new_n7419_;
  wire not_new_n7643__1;
  wire new_n3923_;
  wire not_new_n2836_;
  wire not_pi038_1;
  wire new_n9002_;
  wire not_new_n602__6;
  wire not_new_n635__1176490;
  wire not_new_n635_;
  wire and_and_and_not_pi056_1_not_pi055_1_not_pi054_1_not_pi053_1;
  wire not_new_n1581__113988951853731430;
  wire new_n8377_;
  wire not_new_n2840_;
  wire new_n2622_;
  wire key_gate_108;
  wire not_new_n640__8235430;
  wire not_new_n3998__0;
  wire new_n4026_;
  wire not_new_n4516_;
  wire new_n4666_;
  wire not_new_n631__47475615099430;
  wire new_n9942_;
  wire not_new_n603__490;
  wire not_new_n621__403536070;
  wire not_new_n4185_;
  wire key_gate_27;
  wire new_n1703_;
  wire new_n9279_;
  wire not_new_n3184__8235430;
  wire not_new_n1784_;
  wire new_n4636_;
  wire new_n9421_;
  wire not_new_n1055__5;
  wire not_new_n6137_;
  wire or_or_not_new_n1806__not_new_n1807__not_new_n1809_;
  wire not_new_n8128_;
  wire not_pi187;
  wire not_new_n618__168070;
  wire new_n4972_;
  wire not_new_n1600__6;
  wire not_pi141_0;
  wire not_new_n5996_;
  wire not_new_n1019__1;
  wire new_n1546_;
  wire new_n1436_;
  wire new_n8484_;
  wire not_new_n6024_;
  wire not_pi064_16284135979104490;
  wire new_n7672_;
  wire not_new_n640__19773267430;
  wire new_n5934_;
  wire new_n6081_;
  wire not_new_n8847_;
  wire not_new_n8678_;
  wire new_n6310_;
  wire new_n4126_;
  wire not_new_n6308_;
  wire not_new_n6966_;
  wire new_n6024_;
  wire new_n3946_;
  wire not_new_n9647__0;
  wire new_n7837_;
  wire new_n7015_;
  wire new_n3846_;
  wire not_new_n1043__47475615099430;
  wire not_pi110;
  wire not_new_n6974__47475615099430;
  wire not_new_n5617__0;
  wire new_n5221_;
  wire not_new_n8779_;
  wire not_pi129;
  wire new_n9157_;
  wire not_new_n626__2824752490;
  wire not_new_n7666__1;
  wire not_new_n9756_;
  wire new_n6708_;
  wire not_new_n2725_;
  wire not_new_n8581_;
  wire not_new_n1552_;
  wire not_new_n1051__57648010;
  wire new_n587_;
  wire new_n929_;
  wire not_new_n5772__0;
  wire new_n6137_;
  wire not_pi266_1;
  wire not_new_n7893_;
  wire not_new_n1059__490;
  wire not_new_n2675_;
  wire not_new_n1534__138412872010;
  wire not_new_n7173_;
  wire new_n9308_;
  wire not_new_n617__8235430;
  wire not_new_n5900__2;
  wire not_new_n2779_;
  wire not_new_n6757_;
  wire not_new_n3315__797922662976120010;
  wire not_new_n1067__5;
  wire po290;
  wire or_or_not_new_n8696__not_new_n8690__not_new_n8689_;
  wire not_new_n5697_;
  wire new_n9640_;
  wire not_new_n7962_;
  wire new_n2952_;
  wire not_new_n6531_;
  wire new_n2252_;
  wire new_n1294_;
  wire not_new_n5888_;
  wire not_new_n4599_;
  wire not_new_n1613__8;
  wire new_n6503_;
  wire not_new_n634__47475615099430;
  wire new_n7056_;
  wire not_new_n10231_;
  wire new_n6802_;
  wire not_new_n4979_;
  wire new_n9619_;
  wire not_new_n578_;
  wire not_new_n647__4;
  wire not_new_n3402_;
  wire new_n1451_;
  wire new_n7835_;
  wire new_n3174_;
  wire new_n9182_;
  wire not_new_n1047_;
  wire not_new_n8810_;
  wire not_new_n608__3;
  wire not_new_n8146__0;
  wire not_new_n928__4;
  wire not_new_n1583__10;
  wire not_new_n1639_;
  wire new_n8655_;
  wire not_new_n629__8;
  wire not_new_n7905_;
  wire new_n8695_;
  wire new_n1968_;
  wire not_new_n1039__1176490;
  wire and_not_pi037_2_not_pi036_2;
  wire not_new_n9348_;
  wire not_new_n2721_;
  wire new_n694_;
  wire not_new_n643__2;
  wire new_n1926_;
  wire not_new_n634__273687473400809163430;
  wire new_n588_;
  wire not_new_n3568_;
  wire not_new_n1536__16284135979104490;
  wire not_new_n6352_;
  wire new_n3744_;
  wire not_new_n9479_;
  wire not_new_n633__9;
  wire not_new_n9069_;
  wire new_n1303_;
  wire not_new_n635__0;
  wire new_n9225_;
  wire new_n6362_;
  wire not_new_n5049_;
  wire not_new_n8898__1;
  wire not_new_n994__70;
  wire new_n4633_;
  wire not_new_n631__113988951853731430;
  wire new_n8730_;
  wire new_n3580_;
  wire new_n1295_;
  wire new_n6139_;
  wire not_po296_138412872010;
  wire not_pi101;
  wire new_n8845_;
  wire new_n9812_;
  wire new_n9428_;
  wire new_n3779_;
  wire new_n2500_;
  wire not_new_n630__968890104070;
  wire not_new_n626__168070;
  wire not_new_n9909_;
  wire new_n968_;
  wire not_new_n7511_;
  wire not_new_n4645_;
  wire not_new_n6445_;
  wire not_new_n6982__1;
  wire new_n9670_;
  wire not_new_n9357_;
  wire not_new_n9668__0;
  wire not_new_n617__4;
  wire not_new_n8995__0;
  wire not_new_n644__403536070;
  wire not_new_n632__168070;
  wire not_new_n9506__1;
  wire not_new_n5732_;
  wire not_new_n7655__0;
  wire new_n2016_;
  wire new_n4530_;
  wire not_new_n926__0;
  wire not_new_n6481__0;
  wire new_n7887_;
  wire not_new_n2583_;
  wire not_new_n5822_;
  wire new_n6940_;
  wire not_new_n7392_;
  wire not_new_n4937__1;
  wire new_n8330_;
  wire not_new_n9397__0;
  wire not_new_n1576__4;
  wire not_new_n9095_;
  wire not_new_n3292_;
  wire not_new_n6456_;
  wire not_new_n2754_;
  wire new_n5785_;
  wire not_new_n593_;
  wire not_new_n9191_;
  wire not_new_n9423_;
  wire not_new_n4447_;
  wire not_new_n4711_;
  wire not_new_n585__168070;
  wire key_gate_47;
  wire not_new_n1959_;
  wire not_new_n8610_;
  wire new_n4742_;
  wire not_new_n1600__19773267430;
  wire new_n6444_;
  wire new_n6302_;
  wire not_new_n5953_;
  wire not_new_n4337__0;
  wire not_new_n617__168070;
  wire not_new_n8068_;
  wire new_n4801_;
  wire not_new_n1534__16284135979104490;
  wire not_new_n1015__4;
  wire not_new_n5814_;
  wire new_n4008_;
  wire new_n6738_;
  wire not_new_n7301_;
  wire new_n2849_;
  wire not_new_n2934_;
  wire new_n7368_;
  wire new_n7546_;
  wire new_n10305_;
  wire not_new_n4145_;
  wire or_not_new_n5276__not_new_n5277_;
  wire not_new_n1480_;
  wire not_new_n9719_;
  wire not_pi241;
  wire new_n6028_;
  wire not_new_n659_;
  wire new_n2236_;
  wire not_new_n7655_;
  wire not_new_n5778__0;
  wire not_new_n4254_;
  wire po025;
  wire not_new_n4147_;
  wire not_new_n9962_;
  wire new_n2750_;
  wire not_new_n4514_;
  wire new_n2662_;
  wire not_pi146_2;
  wire not_new_n2948_;
  wire not_new_n736__1;
  wire new_n8767_;
  wire not_new_n9506__0;
  wire new_n4006_;
  wire new_n6881_;
  wire new_n7496_;
  wire not_new_n635__138412872010;
  wire not_pi139;
  wire new_n2578_;
  wire new_n5360_;
  wire new_n3449_;
  wire new_n3158_;
  wire or_not_new_n2555__not_new_n2554_;
  wire new_n3723_;
  wire not_new_n1057__9;
  wire not_new_n631__168070;
  wire new_n2425_;
  wire not_new_n8121_;
  wire new_n8875_;
  wire new_n3126_;
  wire not_pi178_1;
  wire not_new_n1597__70;
  wire not_new_n5279_;
  wire not_new_n8827_;
  wire new_n2585_;
  wire not_new_n1156_;
  wire new_n6342_;
  wire not_new_n5674_;
  wire not_new_n5762_;
  wire new_n1198_;
  wire not_new_n3284_;
  wire not_new_n3708_;
  wire not_new_n775_;
  wire not_new_n643__168070;
  wire key_gate_125;
  wire not_new_n3484_;
  wire po192;
  wire not_new_n1601__490;
  wire new_n10163_;
  wire not_new_n7744_;
  wire new_n2122_;
  wire not_new_n1583__16284135979104490;
  wire new_n10301_;
  wire new_n6006_;
  wire new_n3146_;
  wire new_n8826_;
  wire new_n4588_;
  wire new_n3870_;
  wire not_new_n1037__9;
  wire not_new_n8596__0;
  wire new_n2742_;
  wire new_n5592_;
  wire not_new_n7460_;
  wire not_new_n1171_;
  wire not_new_n9501__0;
  wire new_n5684_;
  wire new_n7584_;
  wire not_new_n1942_;
  wire new_n9202_;
  wire new_n6131_;
  wire new_n1367_;
  wire not_new_n682_;
  wire not_new_n1581__57648010;
  wire new_n991_;
  wire new_n5844_;
  wire new_n2987_;
  wire new_n3764_;
  wire not_new_n8260_;
  wire not_new_n4142_;
  wire new_n2120_;
  wire new_n5202_;
  wire not_new_n3703_;
  wire not_new_n4621_;
  wire new_n612_;
  wire not_new_n4141_;
  wire new_n7262_;
  wire not_new_n9767_;
  wire new_n6693_;
  wire not_new_n7434_;
  wire not_new_n4494__0;
  wire not_new_n1538__19773267430;
  wire not_new_n1043__0;
  wire and_new_n5289__new_n5287_;
  wire not_new_n6921_;
  wire not_new_n1067__138412872010;
  wire not_new_n4541_;
  wire not_new_n1597__8235430;
  wire new_n1155_;
  wire not_new_n6562_;
  wire new_n8975_;
  wire not_new_n3315__47475615099430;
  wire new_n7933_;
  wire not_new_n3175_;
  wire new_n9718_;
  wire new_n4997_;
  wire not_new_n1301_;
  wire not_new_n1538__9;
  wire not_new_n1585_;
  wire new_n9630_;
  wire new_n1190_;
  wire not_new_n639__2;
  wire not_new_n738_;
  wire new_n6557_;
  wire new_n2766_;
  wire not_new_n9228_;
  wire not_new_n4732_;
  wire new_n9510_;
  wire not_new_n8212_;
  wire not_new_n5319_;
  wire not_new_n626_;
  wire and_and_new_n1991__new_n1994__new_n1992_;
  wire not_new_n5796_;
  wire not_new_n601__138412872010;
  wire not_new_n1616__1;
  wire new_n9508_;
  wire not_new_n984__968890104070;
  wire new_n7924_;
  wire new_n6260_;
  wire new_n1018_;
  wire new_n1586_;
  wire not_new_n9515__0;
  wire not_pi131_1;
  wire not_new_n4940_;
  wire not_pi024_0;
  wire not_new_n1594_;
  wire not_new_n6544__0;
  wire new_n6639_;
  wire not_new_n2750_;
  wire not_new_n597__797922662976120010;
  wire new_n8031_;
  wire new_n6118_;
  wire new_n9162_;
  wire new_n6883_;
  wire new_n6783_;
  wire new_n1398_;
  wire new_n7492_;
  wire not_new_n10077_;
  wire new_n1841_;
  wire new_n2481_;
  wire not_new_n3995__0;
  wire not_new_n4811__0;
  wire not_new_n6204_;
  wire not_new_n4032__1;
  wire not_new_n4440_;
  wire not_new_n633_;
  wire not_new_n7098_;
  wire not_pi012;
  wire not_new_n10060_;
  wire not_new_n4999__2;
  wire not_new_n1055__7;
  wire not_new_n4945_;
  wire not_new_n3386_;
  wire not_new_n991_;
  wire not_new_n591__16284135979104490;
  wire not_new_n6914_;
  wire not_new_n7263_;
  wire not_new_n3473_;
  wire not_new_n599__3;
  wire not_po298_3430;
  wire not_new_n6972_;
  wire not_new_n729__0;
  wire not_new_n1003__5;
  wire not_new_n8880__0;
  wire not_new_n4970__0;
  wire new_n7283_;
  wire not_new_n649_;
  wire new_n3825_;
  wire not_pi201;
  wire not_po296_2824752490;
  wire new_n4367_;
  wire new_n9895_;
  wire not_new_n7605__1;
  wire not_new_n1597__2326305139872070;
  wire not_new_n1589__24010;
  wire new_n9288_;
  wire new_n3791_;
  wire not_new_n3128_;
  wire not_new_n8858__0;
  wire new_n1585_;
  wire not_pi021_0;
  wire and_new_n3001__new_n998_;
  wire not_new_n5516_;
  wire not_new_n4772_;
  wire new_n6309_;
  wire not_new_n602__9;
  wire not_new_n2323_;
  wire not_new_n7761_;
  wire or_not_new_n2151__not_new_n2148_;
  wire not_new_n618__2326305139872070;
  wire new_n6703_;
  wire not_new_n10337_;
  wire not_new_n4118__1;
  wire not_new_n1983_;
  wire not_new_n4087_;
  wire not_new_n5265_;
  wire new_n9183_;
  wire not_new_n4168__0;
  wire new_n6147_;
  wire not_pi275;
  wire not_new_n9233_;
  wire key_gate_103;
  wire new_n3732_;
  wire new_n1276_;
  wire not_new_n1019__6;
  wire not_new_n631__6782230728490;
  wire not_new_n8926_;
  wire new_n6463_;
  wire or_not_new_n4414__0_not_new_n1010__3;
  wire not_new_n1061_;
  wire not_po298_8;
  wire not_new_n773_;
  wire not_new_n3238_;
  wire not_new_n7531_;
  wire new_n3226_;
  wire not_new_n9795_;
  wire new_n684_;
  wire not_new_n6644_;
  wire new_n4334_;
  wire new_n6393_;
  wire not_new_n1576__5;
  wire new_n5257_;
  wire new_n7065_;
  wire new_n2701_;
  wire new_n5607_;
  wire not_new_n6501__0;
  wire not_new_n1061__168070;
  wire new_n9042_;
  wire new_n579_;
  wire or_not_new_n6334__not_new_n6232__0;
  wire new_n8411_;
  wire not_new_n1576__6;
  wire not_new_n2509__70;
  wire new_n6445_;
  wire not_new_n7409_;
  wire not_new_n8645_;
  wire not_new_n1039__19773267430;
  wire not_new_n618__39098210485829880490;
  wire new_n3345_;
  wire new_n8969_;
  wire new_n8353_;
  wire new_n2719_;
  wire new_n2037_;
  wire not_new_n10030_;
  wire not_new_n587__113988951853731430;
  wire new_n4437_;
  wire not_new_n5784__0;
  wire not_new_n7752__1;
  wire not_new_n9872__0;
  wire not_new_n4753__0;
  wire new_n4464_;
  wire new_n10208_;
  wire not_new_n2886_;
  wire new_n5441_;
  wire not_new_n1035__4;
  wire new_n9633_;
  wire new_n9447_;
  wire new_n6794_;
  wire new_n4879_;
  wire new_n7440_;
  wire not_new_n647__2824752490;
  wire new_n8990_;
  wire not_new_n3184_;
  wire not_new_n9407_;
  wire not_new_n4159_;
  wire new_n5854_;
  wire not_new_n605__2;
  wire not_new_n625__1;
  wire not_new_n10085_;
  wire not_new_n4998_;
  wire not_new_n5063_;
  wire new_n9557_;
  wire not_new_n3143_;
  wire new_n9851_;
  wire not_new_n6910_;
  wire new_n9725_;
  wire not_new_n7360__1;
  wire not_new_n7541_;
  wire not_new_n923_;
  wire or_not_new_n2854__not_new_n2853_;
  wire new_n7095_;
  wire new_n5572_;
  wire new_n8086_;
  wire not_new_n9947__0;
  wire not_new_n7623_;
  wire not_new_n722__0;
  wire not_new_n2002_;
  wire not_new_n6189_;
  wire not_new_n581__3;
  wire new_n1825_;
  wire new_n1800_;
  wire not_new_n2104_;
  wire not_new_n6618_;
  wire new_n5036_;
  wire and_new_n6993__new_n7526_;
  wire not_new_n7350_;
  wire not_new_n1603_;
  wire not_new_n7863_;
  wire not_new_n1031__490;
  wire and_new_n1746__new_n1747_;
  wire new_n3937_;
  wire not_po296_1915812313805664144010;
  wire not_new_n9378__0;
  wire new_n4204_;
  wire or_not_new_n1291__not_new_n1289_;
  wire not_new_n586__19773267430;
  wire not_new_n3184__1;
  wire new_n2798_;
  wire new_n6560_;
  wire not_new_n7605__0;
  wire not_new_n4375_;
  wire not_new_n4421__0;
  wire not_new_n6467_;
  wire new_n2158_;
  wire not_new_n8412_;
  wire po057;
  wire not_new_n698_;
  wire not_new_n9293_;
  wire not_new_n1536__490;
  wire not_new_n9148_;
  wire not_new_n3111_;
  wire not_new_n624__113988951853731430;
  wire not_new_n1961_;
  wire new_n7767_;
  wire new_n7325_;
  wire not_new_n5899__1;
  wire new_n4862_;
  wire not_new_n989__168070;
  wire not_new_n5501_;
  wire not_new_n2867_;
  wire not_new_n3006_;
  wire or_or_not_new_n1561__not_new_n2464__not_new_n1391_;
  wire not_pi145_1;
  wire or_not_new_n1544__not_new_n1358_;
  wire new_n1869_;
  wire new_n8660_;
  wire new_n4564_;
  wire new_n2911_;
  wire new_n5595_;
  wire not_new_n7482_;
  wire new_n8545_;
  wire new_n946_;
  wire not_new_n2205_;
  wire not_new_n1069__1;
  wire not_new_n5834_;
  wire not_new_n601__6782230728490;
  wire new_n4486_;
  wire new_n3572_;
  wire not_new_n647__6782230728490;
  wire new_n8066_;
  wire not_new_n1303_;
  wire not_new_n9250_;
  wire new_n6895_;
  wire not_new_n4020_;
  wire not_new_n7591_;
  wire new_n5385_;
  wire new_n2828_;
  wire new_n10112_;
  wire not_new_n9499_;
  wire not_new_n7696_;
  wire not_new_n2952_;
  wire not_new_n6194_;
  wire not_new_n585__57648010;
  wire not_new_n3384__4;
  wire not_new_n4665_;
  wire new_n6308_;
  wire new_n10319_;
  wire po276;
  wire new_n7953_;
  wire not_pi077;
  wire not_new_n1857_;
  wire not_new_n611__0;
  wire new_n9860_;
  wire not_new_n1065__113988951853731430;
  wire new_n2930_;
  wire or_not_new_n3145__not_new_n3146_;
  wire new_n1639_;
  wire not_new_n9732_;
  wire not_new_n6503__1;
  wire new_n6370_;
  wire not_new_n6482__0;
  wire not_new_n599__70;
  wire not_new_n989__2326305139872070;
  wire not_new_n618__2;
  wire new_n10324_;
  wire not_pi268_2;
  wire not_pi167_3;
  wire new_n8885_;
  wire new_n8999_;
  wire new_n627_;
  wire not_new_n3543_;
  wire new_n6341_;
  wire new_n2057_;
  wire not_new_n1047__3;
  wire and_new_n1033__new_n3404_;
  wire new_n697_;
  wire not_new_n1063__8235430;
  wire not_pi127;
  wire po235;
  wire not_new_n4280_;
  wire not_new_n8834_;
  wire not_new_n3110_;
  wire not_pi022_0;
  wire new_n7351_;
  wire not_new_n1631__968890104070;
  wire not_new_n2152_;
  wire or_not_new_n1473__not_new_n2722_;
  wire new_n963_;
  wire new_n7646_;
  wire not_new_n5578_;
  wire new_n4556_;
  wire new_n1894_;
  wire new_n9390_;
  wire new_n3029_;
  wire not_new_n6534__0;
  wire not_new_n5977_;
  wire not_new_n5486__0;
  wire po160;
  wire new_n9481_;
  wire not_new_n1061__6;
  wire not_new_n4928__1;
  wire not_new_n6060_;
  wire new_n2756_;
  wire not_new_n7034__0;
  wire not_new_n2809_;
  wire new_n1275_;
  wire not_new_n6288_;
  wire new_n4974_;
  wire not_new_n6049_;
  wire not_pi156_0;
  wire not_new_n1209_;
  wire new_n5011_;
  wire new_n8485_;
  wire new_n10138_;
  wire not_new_n1288_;
  wire not_new_n7078_;
  wire new_n9665_;
  wire or_not_new_n3375__2_not_new_n3387__1;
  wire not_new_n755_;
  wire not_new_n5984_;
  wire new_n654_;
  wire new_n1709_;
  wire not_new_n3307_;
  wire new_n8370_;
  wire not_new_n9807_;
  wire not_new_n8676_;
  wire new_n7540_;
  wire not_new_n9927_;
  wire new_n4819_;
  wire not_new_n9935__0;
  wire and_and_new_n1858__new_n1861__new_n1859_;
  wire new_n9835_;
  wire not_new_n626__273687473400809163430;
  wire not_new_n6672_;
  wire new_n6916_;
  wire new_n2740_;
  wire new_n8189_;
  wire new_n9495_;
  wire not_new_n1051__403536070;
  wire not_new_n1069__3;
  wire key_gate_31;
  wire new_n10158_;
  wire not_new_n645__5;
  wire new_n7642_;
  wire not_new_n5333_;
  wire or_not_new_n5766__1_not_new_n6140_;
  wire new_n9852_;
  wire not_new_n5575_;
  wire new_n6851_;
  wire not_new_n9402__1;
  wire new_n4542_;
  wire not_new_n6929_;
  wire new_n7117_;
  wire not_new_n1189_;
  wire new_n4303_;
  wire new_n9353_;
  wire and_and_new_n1217__new_n1218__new_n1220_;
  wire new_n1879_;
  wire new_n3366_;
  wire new_n9588_;
  wire not_new_n1536__2824752490;
  wire new_n6747_;
  wire not_new_n7022_;
  wire not_new_n5592_;
  wire new_n6030_;
  wire not_new_n7545_;
  wire not_new_n1585__168070;
  wire new_n3091_;
  wire new_n6886_;
  wire new_n6214_;
  wire not_new_n1065__19773267430;
  wire not_new_n4129__2;
  wire not_new_n8915_;
  wire new_n7746_;
  wire new_n670_;
  wire not_new_n3187_;
  wire new_n2597_;
  wire not_new_n642__47475615099430;
  wire new_n10147_;
  wire not_new_n610__490;
  wire not_pi237;
  wire new_n2518_;
  wire not_new_n1843__0;
  wire not_new_n1434_;
  wire not_new_n8013_;
  wire not_new_n6455_;
  wire not_new_n9646__0;
  wire new_n2170_;
  wire new_n9517_;
  wire not_new_n602__8;
  wire new_n3173_;
  wire new_n5391_;
  wire new_n10303_;
  wire not_new_n9299_;
  wire not_new_n9951__2;
  wire not_new_n6776_;
  wire new_n2523_;
  wire new_n3287_;
  wire not_new_n5576_;
  wire not_new_n642_;
  wire new_n7811_;
  wire not_new_n8059_;
  wire new_n7921_;
  wire not_new_n596__19773267430;
  wire not_new_n9162_;
  wire not_new_n8349_;
  wire new_n1237_;
  wire new_n9368_;
  wire not_pi147_3;
  wire not_new_n614_;
  wire not_new_n10305_;
  wire not_new_n6061_;
  wire new_n4341_;
  wire not_pi170_0;
  wire or_not_new_n3914__not_new_n3969_;
  wire not_new_n2596_;
  wire not_new_n3137_;
  wire not_new_n7660__0;
  wire not_new_n1004__0;
  wire not_new_n5541_;
  wire not_new_n1603__7;
  wire and_new_n1739__new_n1740_;
  wire new_n7160_;
  wire new_n3708_;
  wire not_new_n9359_;
  wire new_n1370_;
  wire new_n2419_;
  wire not_new_n600__24010;
  wire not_new_n9236_;
  wire new_n5991_;
  wire new_n9773_;
  wire not_new_n3412_;
  wire new_n5855_;
  wire new_n1988_;
  wire not_new_n5121_;
  wire not_new_n3371_;
  wire new_n5333_;
  wire not_new_n6003_;
  wire not_new_n9220_;
  wire new_n5630_;
  wire not_new_n7766_;
  wire not_new_n3324__0;
  wire or_not_new_n2801__not_new_n2800_;
  wire not_new_n8149__0;
  wire not_new_n1549_;
  wire new_n7128_;
  wire new_n4147_;
  wire po071;
  wire new_n973_;
  wire not_new_n1537__4;
  wire new_n775_;
  wire not_new_n8143__0;
  wire not_new_n647__2;
  wire new_n8482_;
  wire new_n5338_;
  wire not_new_n2557_;
  wire new_n5056_;
  wire new_n6804_;
  wire not_new_n2525_;
  wire new_n7774_;
  wire or_or_not_new_n1323__not_new_n1321__not_new_n2230_;
  wire not_new_n2686_;
  wire not_new_n4225_;
  wire not_new_n4268_;
  wire new_n2846_;
  wire new_n3392_;
  wire not_new_n1631__24010;
  wire new_n3426_;
  wire not_new_n4693_;
  wire new_n7981_;
  wire not_new_n1584__2;
  wire not_new_n3229_;
  wire new_n1273_;
  wire new_n4293_;
  wire not_new_n621__2326305139872070;
  wire not_new_n6653_;
  wire not_new_n606__2;
  wire new_n9470_;
  wire new_n3658_;
  wire not_new_n3311__24010;
  wire new_n3860_;
  wire new_n4137_;
  wire not_new_n10227_;
  wire not_new_n1061__8235430;
  wire not_new_n1964_;
  wire not_new_n632__6782230728490;
  wire and_new_n1215__new_n1780_;
  wire new_n9979_;
  wire new_n6574_;
  wire key_gate_26;
  wire not_new_n1045__797922662976120010;
  wire new_n7787_;
  wire new_n9422_;
  wire not_new_n3873_;
  wire not_pi173;
  wire not_new_n9384__0;
  wire not_new_n4320_;
  wire not_new_n1037__2326305139872070;
  wire not_new_n735__0;
  wire new_n5739_;
  wire not_new_n618__6;
  wire new_n9226_;
  wire or_or_not_new_n2537__not_new_n2541__not_new_n1423_;
  wire new_n6949_;
  wire new_n7309_;
  wire not_new_n4136__1;
  wire not_new_n5579__0;
  wire new_n2891_;
  wire new_n4007_;
  wire not_new_n9277_;
  wire not_new_n1924_;
  wire or_not_new_n1311__not_new_n1309_;
  wire new_n2338_;
  wire not_new_n606__3430;
  wire new_n2077_;
  wire not_pi139_2;
  wire new_n9803_;
  wire new_n8988_;
  wire new_n9135_;
  wire not_new_n617__16284135979104490;
  wire not_new_n1882_;
  wire new_n6930_;
  wire not_new_n8892_;
  wire not_new_n603__138412872010;
  wire not_new_n621__57648010;
  wire not_new_n3387__5;
  wire not_new_n8714_;
  wire not_new_n8885__0;
  wire new_n6591_;
  wire new_n2455_;
  wire new_n3898_;
  wire not_new_n7606__2;
  wire not_new_n4036_;
  wire not_pi261_2;
  wire new_n9951_;
  wire not_new_n1594__9;
  wire new_n1579_;
  wire not_new_n4976_;
  wire not_new_n3211_;
  wire not_new_n8264_;
  wire and_and_new_n3750__new_n3753__new_n3759_;
  wire not_new_n2131_;
  wire not_new_n1583__332329305696010;
  wire new_n2182_;
  wire new_n9378_;
  wire new_n7840_;
  wire new_n6817_;
  wire not_new_n1623__0;
  wire not_new_n5138_;
  wire not_new_n1016__3;
  wire not_new_n5161_;
  wire and_new_n4937__new_n5303_;
  wire not_new_n5296_;
  wire not_new_n4910_;
  wire not_new_n3315__113988951853731430;
  wire new_n3996_;
  wire new_n4584_;
  wire new_n6868_;
  wire not_new_n5472__0;
  wire not_pi175;
  wire not_new_n9278_;
  wire not_new_n9890_;
  wire not_new_n7934_;
  wire not_new_n8245_;
  wire new_n7823_;
  wire not_new_n2180_;
  wire not_new_n1536__1;
  wire not_new_n1002__3;
  wire not_new_n9806_;
  wire not_new_n5948_;
  wire new_n9560_;
  wire not_new_n617__24010;
  wire not_new_n7989_;
  wire new_n2971_;
  wire new_n8217_;
  wire new_n6973_;
  wire not_new_n8780_;
  wire not_new_n618__4;
  wire new_n1306_;
  wire not_new_n4480_;
  wire not_new_n2906_;
  wire not_new_n7672__0;
  wire not_new_n3852_;
  wire not_new_n7042__0;
  wire not_new_n3913__1;
  wire not_new_n644__5;
  wire not_new_n624__16284135979104490;
  wire not_new_n10316_;
  wire new_n5884_;
  wire new_n2539_;
  wire not_new_n2537_;
  wire new_n1291_;
  wire not_new_n8595__0;
  wire new_n979_;
  wire new_n7944_;
  wire not_new_n9586_;
  wire new_n1738_;
  wire new_n1623_;
  wire not_new_n3899_;
  wire not_new_n1069__403536070;
  wire new_n9635_;
  wire not_new_n1623_;
  wire new_n1591_;
  wire new_n2324_;
  wire not_new_n3498_;
  wire new_n6806_;
  wire new_n2388_;
  wire not_new_n10057_;
  wire not_new_n611__10;
  wire new_n9264_;
  wire new_n8595_;
  wire not_new_n3057_;
  wire not_new_n9126_;
  wire not_new_n8241_;
  wire not_new_n6149_;
  wire new_n4116_;
  wire not_new_n6234__1;
  wire not_new_n6602_;
  wire new_n646_;
  wire not_pi064_47475615099430;
  wire not_new_n1597__6;
  wire not_pi062_1;
  wire not_new_n1019__0;
  wire and_new_n1877__new_n1880_;
  wire not_new_n3377_;
  wire new_n9862_;
  wire not_new_n5263_;
  wire not_new_n1268_;
  wire new_n6096_;
  wire not_new_n9527_;
  wire not_new_n4841__0;
  wire key_gate_40;
  wire new_n4494_;
  wire new_n8863_;
  wire new_n5824_;
  wire not_new_n1041__403536070;
  wire not_new_n1069__47475615099430;
  wire po227;
  wire po008;
  wire not_new_n4498__0;
  wire new_n637_;
  wire new_n3028_;
  wire new_n9977_;
  wire new_n5128_;
  wire not_new_n8984__1;
  wire not_new_n8820_;
  wire not_new_n5633_;
  wire new_n9138_;
  wire or_not_new_n1566__not_new_n2489_;
  wire new_n4247_;
  wire not_pi046_2;
  wire not_new_n994__5;
  wire not_new_n2338__0;
  wire not_new_n625__2824752490;
  wire new_n1845_;
  wire po264;
  wire not_new_n1600__10;
  wire not_new_n1598__5;
  wire not_new_n9465_;
  wire not_new_n5102__0;
  wire not_new_n591__490;
  wire not_new_n629__7;
  wire not_new_n631__32199057558131797268376070;
  wire new_n6773_;
  wire not_new_n5985_;
  wire not_new_n3905_;
  wire not_new_n1059__2;
  wire or_not_new_n3100__not_new_n3099_;
  wire not_new_n6443__0;
  wire not_new_n10037_;
  wire not_new_n5798__1;
  wire or_not_new_n8696__not_new_n8690_;
  wire new_n9878_;
  wire new_n7565_;
  wire not_new_n1053__332329305696010;
  wire not_new_n1631__10;
  wire not_new_n1607__57648010;
  wire or_not_new_n2756__not_new_n2755_;
  wire new_n4414_;
  wire new_n7572_;
  wire new_n9207_;
  wire not_new_n4321_;
  wire new_n3069_;
  wire not_new_n4019_;
  wire new_n10277_;
  wire not_pi141_2;
  wire new_n4630_;
  wire new_n10197_;
  wire not_new_n3496_;
  wire new_n7107_;
  wire not_new_n5419_;
  wire new_n1567_;
  wire new_n4182_;
  wire not_new_n10013_;
  wire new_n7481_;
  wire not_new_n9013_;
  wire new_n9211_;
  wire not_new_n1588__2;
  wire new_n7120_;
  wire new_n5880_;
  wire new_n3142_;
  wire not_new_n2826_;
  wire not_new_n4129__0;
  wire new_n6329_;
  wire new_n2075_;
  wire not_new_n1728__5;
  wire not_new_n5018_;
  wire not_new_n5905_;
  wire new_n8542_;
  wire not_new_n1588__332329305696010;
  wire new_n3778_;
  wire new_n733_;
  wire new_n5606_;
  wire not_new_n598__16284135979104490;
  wire not_new_n3146_;
  wire not_new_n1589__47475615099430;
  wire new_n4224_;
  wire new_n2317_;
  wire new_n1875_;
  wire new_n6070_;
  wire not_new_n8170_;
  wire new_n3824_;
  wire not_new_n8008_;
  wire not_new_n3090_;
  wire not_new_n585__1176490;
  wire not_new_n7665__1;
  wire not_new_n3285_;
  wire not_new_n6974__6782230728490;
  wire po171;
  wire not_new_n3989_;
  wire not_new_n5858_;
  wire new_n1837_;
  wire not_new_n9460_;
  wire not_new_n3930__0;
  wire not_new_n3202_;
  wire or_or_or_not_new_n2740__not_new_n2743__not_new_n2742__not_new_n2744_;
  wire new_n6323_;
  wire not_new_n643__19773267430;
  wire new_n6631_;
  wire not_new_n605__10;
  wire new_n5518_;
  wire not_pi168_0;
  wire new_n1923_;
  wire not_new_n2347_;
  wire not_new_n6004_;
  wire new_n8224_;
  wire new_n10264_;
  wire new_n4361_;
  wire new_n6511_;
  wire new_n6996_;
  wire not_new_n8604_;
  wire new_n2123_;
  wire new_n7366_;
  wire new_n6361_;
  wire po260;
  wire not_new_n1603__968890104070;
  wire new_n9017_;
  wire not_new_n2262_;
  wire new_n2809_;
  wire not_new_n6524__0;
  wire not_new_n581__24010;
  wire new_n4815_;
  wire not_new_n589__57648010;
  wire new_n7653_;
  wire not_new_n6443__10;
  wire not_new_n1867_;
  wire key_gate_99;
  wire new_n745_;
  wire new_n7081_;
  wire not_new_n9014_;
  wire new_n1743_;
  wire new_n1994_;
  wire not_new_n7441_;
  wire not_new_n1580__2;
  wire not_new_n598__968890104070;
  wire not_new_n1067__0;
  wire not_new_n644__6;
  wire not_new_n8647_;
  wire new_n5220_;
  wire not_pi164_0;
  wire new_n8935_;
  wire not_new_n10228_;
  wire new_n10309_;
  wire not_new_n1538__7;
  wire not_new_n9956_;
  wire not_new_n5118_;
  wire or_not_new_n3103__not_new_n3102_;
  wire not_new_n5448_;
  wire new_n5275_;
  wire not_new_n10055_;
  wire not_new_n989__4;
  wire new_n3204_;
  wire not_new_n6280_;
  wire key_gate_80;
  wire not_new_n606__0;
  wire not_new_n4777__0;
  wire not_new_n5910_;
  wire not_new_n3914__0;
  wire not_new_n5490__0;
  wire not_new_n8495_;
  wire new_n5744_;
  wire not_new_n6699_;
  wire new_n8704_;
  wire not_new_n733__0;
  wire new_n9848_;
  wire not_new_n631__1176490;
  wire not_new_n6976__0;
  wire new_n5589_;
  wire not_new_n8256_;
  wire new_n4141_;
  wire not_new_n1055__5585458640832840070;
  wire not_new_n1284_;
  wire not_new_n10009__0;
  wire not_new_n1027__70;
  wire new_n4954_;
  wire new_n2889_;
  wire new_n4863_;
  wire not_new_n994__8235430;
  wire new_n4384_;
  wire not_new_n2964_;
  wire new_n9545_;
  wire not_new_n10042_;
  wire not_new_n627__5;
  wire new_n2437_;
  wire not_new_n1534__3430;
  wire new_n7451_;
  wire new_n7919_;
  wire not_new_n8354_;
  wire new_n3759_;
  wire new_n1716_;
  wire new_n1989_;
  wire not_new_n4122__0;
  wire not_new_n3915_;
  wire not_pi240;
  wire not_new_n3972_;
  wire not_new_n7933_;
  wire new_n9789_;
  wire not_new_n3246_;
  wire not_new_n3920__0;
  wire not_new_n3372__5585458640832840070;
  wire not_new_n1023__3;
  wire not_new_n7345__0;
  wire not_new_n647__168070;
  wire not_new_n5299_;
  wire new_n3752_;
  wire new_n8739_;
  wire new_n5313_;
  wire not_new_n4016__0;
  wire new_n7644_;
  wire not_new_n1584__7;
  wire new_n2152_;
  wire not_new_n1483_;
  wire not_new_n6118_;
  wire not_new_n646__3;
  wire not_new_n8026_;
  wire not_new_n6025_;
  wire new_n2560_;
  wire not_new_n629__1176490;
  wire new_n2125_;
  wire not_new_n3261_;
  wire not_new_n8690_;
  wire new_n9149_;
  wire new_n5317_;
  wire not_pi097;
  wire not_new_n1037__24010;
  wire not_new_n4130__2;
  wire new_n4127_;
  wire new_n6239_;
  wire new_n7374_;
  wire new_n3868_;
  wire not_new_n7268_;
  wire not_new_n7575_;
  wire and_and_new_n6373__new_n6254__new_n6402_;
  wire new_n2855_;
  wire new_n3490_;
  wire not_new_n1616_;
  wire new_n5115_;
  wire not_new_n4518_;
  wire new_n3881_;
  wire new_n5138_;
  wire new_n4177_;
  wire new_n1057_;
  wire po173;
  wire not_new_n1015_;
  wire not_new_n626__32199057558131797268376070;
  wire not_new_n4961_;
  wire not_new_n5613_;
  wire not_new_n9877_;
  wire not_new_n5088_;
  wire not_new_n6232__0;
  wire new_n7396_;
  wire new_n1429_;
  wire not_new_n635__3430;
  wire and_not_pi034_2_not_pi033_4;
  wire not_new_n5471_;
  wire not_new_n6627_;
  wire key_gate_119;
  wire not_new_n8313_;
  wire new_n1177_;
  wire new_n8823_;
  wire not_new_n7655__2;
  wire not_new_n593__2;
  wire not_new_n9946_;
  wire new_n5839_;
  wire new_n2081_;
  wire not_new_n6443__113988951853731430;
  wire not_pi037;
  wire not_new_n7739_;
  wire not_new_n5327_;
  wire not_new_n4157__1;
  wire new_n1386_;
  wire not_new_n4208_;
  wire new_n3865_;
  wire not_new_n10287_;
  wire new_n5254_;
  wire not_new_n7055_;
  wire not_new_n1584__1176490;
  wire new_n8118_;
  wire not_new_n976_;
  wire not_new_n7700_;
  wire not_new_n1069__1176490;
  wire not_new_n3452_;
  wire new_n8249_;
  wire not_new_n5827_;
  wire not_new_n1786_;
  wire not_new_n7354__1;
  wire new_n1345_;
  wire not_new_n1037__3430;
  wire new_n8429_;
  wire not_new_n3830_;
  wire new_n9831_;
  wire not_new_n5288_;
  wire not_new_n597__5;
  wire new_n7092_;
  wire not_new_n2929_;
  wire not_new_n4410_;
  wire new_n1993_;
  wire not_new_n10092_;
  wire not_new_n7018__2;
  wire not_new_n1611__2326305139872070;
  wire not_new_n1611__57648010;
  wire new_n4474_;
  wire not_new_n4760__0;
  wire not_new_n8715__0;
  wire new_n641_;
  wire not_new_n9393_;
  wire not_new_n9928_;
  wire new_n2155_;
  wire not_new_n7003_;
  wire new_n1865_;
  wire not_new_n639__8;
  wire not_new_n4026_;
  wire not_new_n6495__0;
  wire not_new_n589__797922662976120010;
  wire new_n2808_;
  wire new_n1411_;
  wire new_n5270_;
  wire not_new_n1581__6;
  wire new_n9375_;
  wire new_n1685_;
  wire new_n1613_;
  wire not_new_n10325_;
  wire new_n6026_;
  wire new_n8027_;
  wire new_n9573_;
  wire not_new_n1299_;
  wire not_new_n9853_;
  wire not_new_n4650_;
  wire new_n1239_;
  wire new_n1278_;
  wire not_new_n1041__2824752490;
  wire not_new_n632__9;
  wire not_pi188;
  wire new_n6480_;
  wire not_po298_5585458640832840070;
  wire new_n9224_;
  wire not_new_n4111_;
  wire not_new_n10131_;
  wire not_new_n5605_;
  wire new_n6060_;
  wire not_new_n9397_;
  wire po229;
  wire not_new_n629__968890104070;
  wire not_new_n8993_;
  wire new_n3487_;
  wire new_n4811_;
  wire not_new_n4053_;
  wire not_new_n9426__0;
  wire not_new_n4173__0;
  wire or_or_not_new_n1958__not_new_n1959__not_new_n1961_;
  wire or_or_not_new_n1243__not_new_n1241__not_new_n1850_;
  wire new_n1258_;
  wire new_n7712_;
  wire not_new_n600__138412872010;
  wire new_n3207_;
  wire new_n6101_;
  wire not_new_n1580__3430;
  wire new_n1881_;
  wire new_n7704_;
  wire not_new_n7740_;
  wire new_n5136_;
  wire new_n8531_;
  wire not_new_n5477_;
  wire not_new_n8437_;
  wire new_n5089_;
  wire new_n3698_;
  wire not_new_n1607__3;
  wire new_n4442_;
  wire not_new_n1357_;
  wire not_new_n7009__0;
  wire not_new_n4491_;
  wire new_n6848_;
  wire not_new_n1607__70;
  wire not_pi136_1;
  wire not_new_n2261_;
  wire not_new_n1373_;
  wire new_n10251_;
  wire not_new_n4077_;
  wire not_new_n7342__1;
  wire not_new_n1604__138412872010;
  wire new_n6211_;
  wire not_new_n9764_;
  wire and_and_new_n1463__new_n1465__new_n1464_;
  wire new_n6596_;
  wire new_n653_;
  wire new_n4848_;
  wire new_n9854_;
  wire new_n4330_;
  wire new_n8498_;
  wire new_n6957_;
  wire not_new_n8141_;
  wire not_new_n7113_;
  wire not_new_n5967_;
  wire not_new_n3715_;
  wire not_new_n6289_;
  wire new_n3451_;
  wire not_new_n5814__0;
  wire new_n4468_;
  wire not_new_n1612__968890104070;
  wire or_or_not_new_n1055__168070_not_new_n6325__not_new_n6373__1;
  wire new_n7219_;
  wire new_n9298_;
  wire not_new_n621__6;
  wire not_new_n4806__0;
  wire new_n5208_;
  wire new_n5720_;
  wire not_new_n7615_;
  wire new_n2191_;
  wire not_new_n634__3;
  wire new_n4332_;
  wire new_n1236_;
  wire not_new_n2790_;
  wire not_new_n9794_;
  wire not_new_n3886_;
  wire not_new_n989__5;
  wire not_new_n7795__0;
  wire not_new_n6719_;
  wire not_pi058_2;
  wire new_n6629_;
  wire or_not_new_n2774__not_new_n2773_;
  wire not_new_n10263_;
  wire not_new_n5757_;
  wire not_new_n6640__0;
  wire not_new_n1603__2326305139872070;
  wire new_n8327_;
  wire new_n2950_;
  wire not_new_n2849_;
  wire new_n2704_;
  wire not_pi265_0;
  wire not_new_n942_;
  wire not_new_n634__6;
  wire new_n8937_;
  wire not_new_n8193_;
  wire new_n4157_;
  wire not_new_n4958__0;
  wire not_new_n9906_;
  wire new_n2354_;
  wire new_n8256_;
  wire not_pi064_10;
  wire new_n1469_;
  wire or_not_new_n8713__not_new_n8715_;
  wire not_new_n3264_;
  wire new_n9139_;
  wire not_pi013_0;
  wire not_new_n1053__968890104070;
  wire new_n1455_;
  wire not_pi064_968890104070;
  wire new_n4704_;
  wire new_n6095_;
  wire not_new_n4783_;
  wire not_new_n8150__0;
  wire not_new_n6536__0;
  wire new_n5436_;
  wire new_n9898_;
  wire not_new_n642__6;
  wire not_new_n597__968890104070;
  wire not_new_n4762_;
  wire not_new_n7294_;
  wire new_n1217_;
  wire not_new_n1952_;
  wire not_new_n4030_;
  wire not_new_n3236_;
  wire not_new_n3839_;
  wire not_new_n6486__1;
  wire not_new_n642__4;
  wire new_n1816_;
  wire not_new_n9506_;
  wire not_new_n608__9;
  wire not_new_n3226_;
  wire new_n2117_;
  wire new_n3773_;
  wire not_new_n648__70;
  wire not_new_n8452_;
  wire new_n2307_;
  wire not_new_n4094_;
  wire not_new_n4034_;
  wire not_new_n636__4;
  wire not_new_n602__10;
  wire new_n2590_;
  wire not_new_n644__1;
  wire not_new_n7682_;
  wire new_n2100_;
  wire not_new_n7494_;
  wire not_new_n1572__0;
  wire not_new_n4088_;
  wire not_new_n4551_;
  wire not_new_n8859__0;
  wire and_not_pi056_1_not_pi055_1;
  wire new_n4876_;
  wire not_new_n984__10;
  wire not_new_n6594_;
  wire new_n4399_;
  wire not_new_n8903_;
  wire new_n4568_;
  wire not_new_n989__57648010;
  wire not_new_n775__3;
  wire not_new_n1047__138412872010;
  wire not_new_n3212_;
  wire not_new_n9697_;
  wire not_new_n1573_;
  wire new_n10077_;
  wire po076;
  wire not_new_n603__1;
  wire not_new_n7430__1;
  wire not_new_n8028_;
  wire not_new_n10168_;
  wire new_n965_;
  wire new_n1588_;
  wire not_new_n1611__16284135979104490;
  wire not_new_n7688_;
  wire new_n5649_;
  wire not_new_n1536__1176490;
  wire not_new_n9789_;
  wire new_n8876_;
  wire new_n4131_;
  wire not_new_n9246_;
  wire not_new_n5312_;
  wire new_n4287_;
  wire or_not_new_n3167__not_new_n3166_;
  wire new_n8422_;
  wire new_n6538_;
  wire not_new_n1010__3;
  wire not_new_n8514_;
  wire not_new_n1045__3;
  wire not_new_n725_;
  wire new_n3719_;
  wire not_new_n9669_;
  wire not_new_n8884__0;
  wire new_n1665_;
  wire not_new_n2781_;
  wire not_new_n7660_;
  wire not_new_n6280__0;
  wire not_new_n2113_;
  wire not_new_n2997_;
  wire not_new_n640__16284135979104490;
  wire not_po296_1070069044235980333563563003849377848070;
  wire new_n5736_;
  wire new_n9916_;
  wire new_n4003_;
  wire not_new_n9960__0;
  wire not_new_n5145_;
  wire new_n3137_;
  wire or_not_new_n2989__not_new_n3826_;
  wire new_n6063_;
  wire not_new_n5305_;
  wire new_n4903_;
  wire and_new_n2219__new_n2222_;
  wire not_pi015_0;
  wire not_new_n3185__5;
  wire not_new_n3948_;
  wire new_n8925_;
  wire not_new_n1005__4;
  wire new_n5842_;
  wire not_new_n5058_;
  wire new_n7373_;
  wire new_n6283_;
  wire new_n2505_;
  wire not_new_n1599__4;
  wire not_new_n8881_;
  wire or_or_not_new_n6348__not_new_n6232__2_not_new_n6234__1;
  wire new_n3737_;
  wire not_new_n8798_;
  wire not_new_n9932__0;
  wire new_n2601_;
  wire new_n4432_;
  wire new_n7448_;
  wire not_new_n8161_;
  wire not_new_n623__1;
  wire not_new_n5735_;
  wire not_new_n2095_;
  wire new_n2725_;
  wire and_new_n2354__new_n2353_;
  wire new_n922_;
  wire new_n2764_;
  wire not_new_n8281__0;
  wire not_new_n9551_;
  wire or_or_not_new_n2910__not_new_n2913__not_new_n2912_;
  wire new_n1705_;
  wire not_new_n8037_;
  wire not_new_n1589__5;
  wire not_new_n9739_;
  wire new_n6523_;
  wire not_new_n2561_;
  wire new_n2611_;
  wire new_n10121_;
  wire new_n1183_;
  wire new_n8454_;
  wire or_not_new_n2863__not_new_n2862_;
  wire new_n5213_;
  wire new_n7370_;
  wire not_new_n5128_;
  wire not_new_n7844_;
  wire not_new_n1537__3;
  wire new_n6530_;
  wire not_new_n1016__0;
  wire not_new_n619__1176490;
  wire not_new_n1031__403536070;
  wire new_n9155_;
  wire new_n9456_;
  wire new_n8915_;
  wire not_new_n3185__4;
  wire new_n5159_;
  wire new_n3082_;
  wire not_new_n9912_;
  wire not_new_n2114_;
  wire not_new_n5087__0;
  wire not_new_n4641_;
  wire new_n2113_;
  wire new_n10151_;
  wire not_new_n640__8;
  wire not_new_n587__2;
  wire new_n5131_;
  wire not_new_n606__9;
  wire new_n8139_;
  wire not_new_n4796_;
  wire new_n7736_;
  wire not_new_n8794__0;
  wire not_new_n7149_;
  wire not_new_n10243_;
  wire new_n3234_;
  wire not_pi179_3;
  wire not_new_n9279_;
  wire new_n7357_;
  wire not_new_n4974__1;
  wire new_n3557_;
  wire not_new_n3934_;
  wire new_n6171_;
  wire new_n8628_;
  wire new_n10069_;
  wire new_n9461_;
  wire not_new_n9486__0;
  wire not_new_n1597__138412872010;
  wire not_pi010;
  wire new_n7114_;
  wire not_new_n7746_;
  wire not_new_n3828_;
  wire not_new_n3932__0;
  wire po274;
  wire not_new_n5452__1;
  wire not_new_n5398_;
  wire not_new_n605__6;
  wire not_new_n10266_;
  wire not_new_n5887__0;
  wire new_n5297_;
  wire new_n9579_;
  wire not_new_n6742_;
  wire new_n3893_;
  wire not_new_n3698_;
  wire or_or_not_new_n6354__not_new_n6373__8_not_new_n6355_;
  wire new_n5105_;
  wire new_n4030_;
  wire not_new_n963_;
  wire new_n2507_;
  wire not_new_n1259_;
  wire new_n8760_;
  wire not_new_n1631__6;
  wire not_new_n4839__0;
  wire new_n7938_;
  wire new_n8050_;
  wire new_n3373_;
  wire new_n4309_;
  wire new_n7918_;
  wire new_n3432_;
  wire not_pi257_4;
  wire not_new_n9810_;
  wire new_n9355_;
  wire po088;
  wire not_new_n4553_;
  wire new_n7821_;
  wire not_new_n10201_;
  wire not_new_n6528__0;
  wire not_new_n4326_;
  wire not_new_n3315__7;
  wire po212;
  wire new_n2028_;
  wire new_n4543_;
  wire not_new_n5163_;
  wire not_new_n1004__7;
  wire new_n5118_;
  wire not_new_n648__10;
  wire not_new_n2986_;
  wire not_new_n3505_;
  wire not_new_n8815_;
  wire new_n8963_;
  wire new_n5805_;
  wire new_n2011_;
  wire not_pi177_3;
  wire not_new_n6322_;
  wire not_new_n601__8;
  wire or_or_or_not_new_n2982__not_new_n2985__not_new_n2984__not_new_n2986_;
  wire not_new_n2910_;
  wire not_new_n1519_;
  wire not_new_n632__113988951853731430;
  wire new_n621_;
  wire new_n7717_;
  wire not_new_n1207_;
  wire not_new_n636__16284135979104490;
  wire new_n9775_;
  wire not_new_n9930_;
  wire new_n6617_;
  wire not_new_n9890__1;
  wire new_n7861_;
  wire new_n1600_;
  wire not_new_n2866_;
  wire not_pi040_2;
  wire not_new_n609__1176490;
  wire new_n7179_;
  wire not_new_n1536__47475615099430;
  wire new_n6601_;
  wire and_new_n3375__new_n3387_;
  wire new_n2279_;
  wire not_new_n5556_;
  wire not_new_n4450_;
  wire new_n5634_;
  wire not_pi064_57648010;
  wire and_new_n3076__new_n998_;
  wire new_n8942_;
  wire not_new_n1604__5;
  wire new_n10181_;
  wire new_n1606_;
  wire not_new_n9961_;
  wire new_n10196_;
  wire new_n10194_;
  wire new_n5571_;
  wire not_new_n632__7;
  wire new_n6749_;
  wire not_new_n1045__4;
  wire not_new_n4617_;
  wire not_new_n626__2326305139872070;
  wire not_new_n9623__0;
  wire not_new_n928__138412872010;
  wire not_new_n9432_;
  wire new_n3724_;
  wire not_new_n4337_;
  wire new_n7253_;
  wire new_n4380_;
  wire not_new_n8262__0;
  wire new_n7208_;
  wire new_n8229_;
  wire not_new_n1407_;
  wire or_not_new_n2665__not_new_n2664_;
  wire new_n2777_;
  wire not_new_n618__138412872010;
  wire new_n704_;
  wire not_new_n4306_;
  wire new_n7877_;
  wire new_n2139_;
  wire not_new_n1004__5;
  wire not_new_n8516_;
  wire not_new_n7652__0;
  wire not_pi196;
  wire not_new_n5786_;
  wire not_new_n7195_;
  wire not_new_n591__3;
  wire not_new_n7031__0;
  wire not_new_n1591__332329305696010;
  wire new_n4046_;
  wire not_new_n7759__2;
  wire or_not_new_n1547__not_new_n1364_;
  wire not_new_n5987_;
  wire new_n3380_;
  wire or_not_new_n1773__not_new_n1213_;
  wire not_new_n1580__2824752490;
  wire new_n2621_;
  wire or_not_new_n1469__not_new_n3820_;
  wire not_new_n3713_;
  wire new_n9488_;
  wire not_new_n7248_;
  wire not_new_n2853_;
  wire new_n7515_;
  wire new_n9374_;
  wire new_n8219_;
  wire not_new_n9494_;
  wire po265;
  wire new_n1465_;
  wire not_new_n5618_;
  wire not_new_n6569_;
  wire not_new_n6467__0;
  wire not_new_n4666_;
  wire not_new_n1612__797922662976120010;
  wire not_new_n600__6;
  wire not_new_n2846_;
  wire new_n9486_;
  wire not_new_n4966__0;
  wire not_new_n6891_;
  wire not_new_n1711_;
  wire not_new_n4760__1;
  wire not_new_n5865_;
  wire not_new_n4256_;
  wire new_n7781_;
  wire new_n2065_;
  wire new_n7292_;
  wire not_new_n3542_;
  wire new_n7782_;
  wire not_new_n8884__1;
  wire not_new_n9874__0;
  wire not_new_n5435__0;
  wire new_n4277_;
  wire new_n5748_;
  wire new_n4533_;
  wire new_n6441_;
  wire not_new_n9893_;
  wire not_new_n596__8235430;
  wire not_new_n9575_;
  wire not_new_n1047__7;
  wire not_new_n1049__19773267430;
  wire not_new_n4997__0;
  wire new_n9221_;
  wire not_new_n1275_;
  wire new_n5713_;
  wire not_new_n9092__0;
  wire new_n2079_;
  wire not_pi159_0;
  wire not_new_n3267_;
  wire not_new_n638__93874803376477543056490;
  wire new_n1882_;
  wire not_new_n3563_;
  wire not_new_n6992__0;
  wire or_or_or_not_new_n2892__not_new_n2895__not_new_n2894__not_new_n2896_;
  wire new_n8516_;
  wire key_gate_55;
  wire not_new_n632__490;
  wire or_or_not_new_n6343__not_new_n6344__not_new_n6345_;
  wire new_n3196_;
  wire not_new_n8264__0;
  wire new_n5419_;
  wire new_n7533_;
  wire not_new_n8057_;
  wire po092;
  wire not_new_n1057__168070;
  wire new_n3678_;
  wire new_n8538_;
  wire not_new_n5880_;
  wire not_pi135;
  wire not_new_n1031__24010;
  wire new_n4808_;
  wire not_new_n9103__0;
  wire new_n771_;
  wire not_new_n775__24010;
  wire new_n5243_;
  wire new_n2319_;
  wire not_new_n3581_;
  wire not_new_n1598__6782230728490;
  wire new_n5076_;
  wire new_n5985_;
  wire not_new_n7137__0;
  wire new_n982_;
  wire new_n1918_;
  wire not_new_n7453_;
  wire not_new_n1681_;
  wire not_new_n4578_;
  wire not_new_n7459_;
  wire new_n4178_;
  wire not_new_n9560_;
  wire not_new_n1071__6782230728490;
  wire not_po296_113988951853731430;
  wire new_n3362_;
  wire not_new_n4137__2;
  wire not_new_n1150__0;
  wire new_n2493_;
  wire or_not_new_n5095__1_not_new_n4899__1;
  wire not_new_n9097__0;
  wire not_new_n4900_;
  wire new_n9960_;
  wire and_new_n6357__new_n6356_;
  wire new_n3518_;
  wire not_new_n1584__16284135979104490;
  wire not_new_n3369_;
  wire new_n6644_;
  wire new_n3150_;
  wire not_new_n637__3;
  wire not_new_n632__8;
  wire not_new_n5950_;
  wire new_n6273_;
  wire new_n6752_;
  wire not_new_n8828__1;
  wire new_n3882_;
  wire not_new_n5580_;
  wire new_n1069_;
  wire new_n3032_;
  wire new_n9676_;
  wire not_new_n7102_;
  wire not_new_n6329_;
  wire not_new_n633__2824752490;
  wire not_new_n8941_;
  wire not_new_n8594_;
  wire not_new_n717_;
  wire not_new_n3980_;
  wire po153;
  wire new_n7982_;
  wire not_new_n4765__1;
  wire not_new_n1271_;
  wire new_n9700_;
  wire new_n624_;
  wire new_n2216_;
  wire new_n10189_;
  wire not_new_n7655__1;
  wire new_n9246_;
  wire new_n6532_;
  wire not_new_n5913_;
  wire new_n774_;
  wire new_n7074_;
  wire not_new_n3712_;
  wire not_new_n2953_;
  wire not_new_n1599__70;
  wire not_new_n5807_;
  wire new_n8980_;
  wire key_gate_70;
  wire new_n1534_;
  wire not_new_n8862_;
  wire not_new_n1348_;
  wire not_new_n8899__1;
  wire new_n10145_;
  wire not_new_n635__403536070;
  wire not_new_n642__2824752490;
  wire not_new_n6990_;
  wire not_new_n594__5;
  wire not_new_n984__1176490;
  wire not_new_n5048_;
  wire new_n4762_;
  wire not_new_n3456_;
  wire not_new_n8007_;
  wire new_n5298_;
  wire new_n3241_;
  wire not_new_n1597__1176490;
  wire not_pi188_0;
  wire not_new_n9358__1;
  wire new_n6963_;
  wire not_new_n994__168070;
  wire new_n8240_;
  wire not_new_n7417_;
  wire new_n6423_;
  wire not_new_n4953_;
  wire new_n8199_;
  wire new_n8639_;
  wire not_pi161_2;
  wire not_pi039;
  wire new_n7157_;
  wire not_new_n5787__0;
  wire new_n6662_;
  wire new_n6025_;
  wire new_n4580_;
  wire new_n2220_;
  wire not_pi100;
  wire not_new_n5409_;
  wire and_and_new_n1222__new_n1223__new_n1225_;
  wire new_n7016_;
  wire not_new_n8563_;
  wire not_new_n8215_;
  wire not_new_n604__70;
  wire and_new_n2325__new_n2332_;
  wire new_n9459_;
  wire new_n6325_;
  wire not_new_n3845_;
  wire new_n717_;
  wire new_n10044_;
  wire new_n8920_;
  wire new_n586_;
  wire not_new_n6066_;
  wire and_new_n2369__new_n2368_;
  wire new_n1193_;
  wire new_n4023_;
  wire not_new_n6052_;
  wire not_new_n7308_;
  wire new_n3096_;
  wire new_n2555_;
  wire not_new_n4776_;
  wire new_n8479_;
  wire not_new_n7621__0;
  wire not_new_n8077_;
  wire not_new_n6506__0;
  wire not_new_n1598__403536070;
  wire not_new_n4706_;
  wire new_n3797_;
  wire not_new_n1411_;
  wire not_new_n1616__5;
  wire not_new_n9254_;
  wire not_new_n641__2824752490;
  wire new_n7856_;
  wire new_n5487_;
  wire not_new_n1576__0;
  wire not_pi248_3;
  wire not_new_n633__0;
  wire new_n2256_;
  wire new_n4285_;
  wire new_n8181_;
  wire not_new_n9398_;
  wire po211;

  not g_0 (not_new_n606__10, new_n606_);
  not g_1 (not_new_n5274_, new_n5274_);
  or g_2 (or_not_new_n8595__not_new_n8593_, not_new_n8595_, not_new_n8593_);
  and g_3 (new_n1462_, new_n3738_, and_and_new_n3732__new_n3735__new_n3741_);
  not g_4 (not_new_n1604__8235430, new_n1604_);
  not g_5 (not_new_n7527_, new_n7527_);
  not g_6 (not_new_n7662__1, new_n7662_);
  not g_7 (not_new_n1536__6, new_n1536_);
  or g_8 (new_n6543_, not_new_n6739_, not_new_n6793_);
  or g_9 (new_n9836_, not_new_n9505_, not_new_n9504_);
  not g_10 (not_new_n1053__6782230728490, new_n1053_);
  not g_11 (not_new_n626__1176490, new_n626_);
  not g_12 (not_new_n597__10, new_n597_);
  not g_13 (not_new_n1057__3, new_n1057_);
  not g_14 (not_new_n3375__3, new_n3375_);
  or g_15 (new_n9101_, not_new_n9186_, not_new_n8943_);
  not g_16 (not_new_n587__168070, new_n587_);
  not g_17 (not_new_n7988_, new_n7988_);
  not g_18 (new_n5783_, new_n633_);
  not g_19 (not_new_n4169_, new_n4169_);
  not g_20 (new_n4782_, new_n1604_);
  not g_21 (not_new_n4764__0, new_n4764_);
  not g_22 (not_new_n4420__0, new_n4420_);
  not g_23 (not_new_n6810_, new_n6810_);
  not g_24 (not_new_n606_, new_n606_);
  not g_25 (not_new_n647__8235430, new_n647_);
  or g_26 (new_n7680_, not_new_n8042_, not_new_n8041_);
  not g_27 (not_new_n7687_, new_n7687_);
  or g_28 (new_n6471_, not_new_n6779_, not_new_n6634_);
  or g_29 (new_n8437_, not_new_n8091_, not_new_n8266__2);
  not g_30 (not_new_n4817_, new_n4817_);
  not g_31 (not_new_n965_, new_n965_);
  not g_32 (not_new_n962_, new_n962_);
  or g_33 (new_n2638_, not_new_n610__490, not_new_n4456__0);
  not g_34 (not_new_n1597__168070, new_n1597_);
  not g_35 (new_n1838_, new_n946_);
  or g_36 (new_n5737_, not_new_n6041_, not_new_n5899_);
  not g_37 (not_new_n8197_, new_n8197_);
  not g_38 (not_new_n1596__113988951853731430, new_n1596_);
  not g_39 (not_new_n6722_, new_n6722_);
  or g_40 (new_n5308_, not_new_n5102__0, not_new_n5306_);
  and g_41 (new_n5030_, new_n5125_, new_n5127_);
  and g_42 (new_n1355_, new_n2372_, and_new_n2374__new_n2373_);
  not g_43 (not_new_n5806__0, new_n5806_);
  or g_44 (new_n3171_, not_new_n928__16284135979104490, not_new_n1053__4);
  not g_45 (not_new_n8720_, new_n8720_);
  and g_46 (new_n1504_, new_n1505_, new_n3031_);
  or g_47 (new_n6559_, not_new_n6831_, not_new_n6830_);
  not g_48 (not_new_n7012_, new_n7012_);
  not g_49 (not_new_n4907_, new_n4907_);
  not g_50 (not_new_n9608_, new_n9608_);
  not g_51 (not_new_n1067__70, new_n1067_);
  not g_52 (not_new_n9565_, new_n9565_);
  or g_53 (new_n10067_, not_new_n10046_, not_new_n10042_);
  not g_54 (not_new_n3099_, new_n3099_);
  not g_55 (not_new_n7038_, new_n7038_);
  and g_56 (and_new_n6362__new_n6430_, new_n6430_, new_n6362_);
  not g_57 (not_new_n1018__4, new_n1018_);
  or g_58 (new_n10300_, not_new_n9934_, not_new_n630__5585458640832840070);
  not g_59 (not_new_n597__47475615099430, new_n597_);
  not g_60 (not_new_n594__24010, new_n594_);
  or g_61 (new_n1996_, not_pi174, not_new_n586__490);
  not g_62 (not_new_n8837_, new_n8837_);
  or g_63 (new_n8300_, not_new_n635__138412872010, not_new_n8107_);
  or g_64 (new_n6168_, not_new_n6021_, not_new_n5896_);
  not g_65 (not_new_n4012_, new_n4012_);
  or g_66 (new_n773_, not_new_n3240_, not_new_n3241_);
  not g_67 (not_new_n1233_, new_n1233_);
  not g_68 (not_new_n4929__0, new_n4929_);
  or g_69 (new_n9412_, not_new_n637__332329305696010, not_new_n1065__113988951853731430);
  not g_70 (not_new_n7395_, new_n7395_);
  or g_71 (new_n3853_, not_new_n6443__490, not_new_n622__70);
  not g_72 (new_n9050_, new_n8978_);
  or g_73 (new_n7429_, not_new_n6974__8235430, not_new_n758_);
  or g_74 (new_n8566_, not_new_n1063__57648010, not_new_n8163__0);
  or g_75 (new_n4401_, not_new_n650_, not_new_n4285_);
  not g_76 (not_new_n9205_, new_n9205_);
  not g_77 (new_n8867_, new_n1059_);
  not g_78 (not_new_n2852_, new_n2852_);
  not g_79 (not_new_n1728__1176490, new_n1728_);
  not g_80 (not_new_n4714_, new_n4714_);
  not g_81 (not_po296_29286449308136415160327158440136953416342323212091034008010, po296);
  not g_82 (not_new_n1269_, new_n1269_);
  not g_83 (not_new_n593__3, new_n593_);
  not g_84 (not_new_n4559_, new_n4559_);
  not g_85 (new_n7206_, new_n7000_);
  or g_86 (new_n2722_, not_new_n2721_, not_new_n3372__3);
  not g_87 (new_n8132_, new_n629_);
  or g_88 (new_n1158_, not_new_n3846_, not_new_n3845_);
  and g_89 (new_n7576_, new_n7852_, new_n7851_);
  and g_90 (and_new_n9879__new_n10247_, new_n9879_, new_n10247_);
  not g_91 (not_new_n6503_, new_n6503_);
  not g_92 (not_new_n1602__332329305696010, new_n1602_);
  not g_93 (not_new_n5085_, new_n5085_);
  not g_94 (not_new_n6266_, new_n6266_);
  not g_95 (not_new_n632__3, new_n632_);
  or g_96 (new_n5414_, not_new_n5412_, not_new_n5413_);
  not g_97 (not_new_n6484_, new_n6484_);
  or g_98 (new_n6750_, not_new_n1596__168070, not_new_n6541_);
  not g_99 (not_new_n7215_, new_n7215_);
  or g_100 (or_not_new_n6240__not_new_n6330_, not_new_n6240_, not_new_n6330_);
  and g_101 (new_n6326_, new_n6395_, and_new_n6375__new_n6382_);
  not g_102 (not_new_n9868__0, new_n9868_);
  not g_103 (not_new_n5879_, new_n5879_);
  and g_104 (and_and_new_n3804__new_n3807__new_n3813_, and_new_n3804__new_n3807_, new_n3813_);
  not g_105 (not_new_n638__968890104070, new_n638_);
  and g_106 (new_n5846_, and_new_n5748__new_n6116_, new_n6115_);
  buf g_107 (po005, pi198);
  or g_108 (new_n693_, not_new_n3051_, not_new_n1517_);
  or g_109 (new_n2450_, not_new_n1071__0, not_new_n598__57648010);
  not g_110 (not_new_n3008_, new_n3008_);
  not g_111 (not_new_n5857_, new_n5857_);
  not g_112 (not_new_n627__10, new_n627_);
  not g_113 (not_new_n8122_, new_n8122_);
  or g_114 (new_n765_, not_new_n3187_, not_new_n3186_);
  not g_115 (not_new_n606__8235430, new_n606_);
  not g_116 (not_new_n9241_, new_n9241_);
  not g_117 (not_new_n615__0, new_n615_);
  and g_118 (new_n6234_, and_and_new_n6326__new_n6241__new_n6227_, new_n6396_);
  not g_119 (not_new_n1017__5, new_n1017_);
  not g_120 (not_new_n1422_, new_n1422_);
  or g_121 (or_not_new_n2928__not_new_n2931_, not_new_n2928_, not_new_n2931_);
  not g_122 (not_new_n7641__0, new_n7641_);
  not g_123 (not_new_n633__19773267430, new_n633_);
  not g_124 (not_new_n4930__0, new_n4930_);
  and g_125 (new_n8926_, and_new_n8997__new_n8998_, new_n9000_);
  or g_126 (new_n3030_, not_new_n1599__2, not_new_n581__3430);
  not g_127 (new_n7634_, new_n640_);
  and g_128 (new_n1540_, new_n3593_, new_n3592_);
  and g_129 (new_n7082_, new_n6964_, new_n7240_);
  not g_130 (not_new_n7233_, new_n7233_);
  or g_131 (new_n7282_, not_new_n724__0, not_new_n7038__0);
  not g_132 (not_pi016_0, pi016);
  and g_133 (new_n5510_, new_n5659_, new_n5660_);
  not g_134 (not_new_n7651__1, new_n7651_);
  or g_135 (new_n689_, not_new_n1508_, not_new_n3035_);
  or g_136 (new_n7034_, not_new_n7420_, not_new_n7419_);
  not g_137 (not_new_n5956_, new_n5956_);
  not g_138 (not_new_n8244__0, new_n8244_);
  not g_139 (not_pi192_0, pi192);
  or g_140 (new_n9197_, not_new_n648__113988951853731430, not_new_n8840_);
  or g_141 (new_n9850_, not_new_n626__32199057558131797268376070, not_new_n9388_);
  or g_142 (new_n8349_, not_new_n8080_, not_new_n8348_);
  or g_143 (po078, not_new_n1205_, key_gate_110);
  or g_144 (new_n1790_, not_new_n585__1, not_pi255);
  not g_145 (not_new_n9911_, new_n9911_);
  not g_146 (not_new_n636__2, new_n636_);
  and g_147 (new_n5493_, and_new_n5582__new_n5648_, new_n5647_);
  or g_148 (new_n2712_, not_new_n2710_, not_new_n2711_);
  not g_149 (not_new_n6789_, new_n6789_);
  not g_150 (not_new_n10144_, new_n10144_);
  not g_151 (not_pi168_1, pi168);
  not g_152 (new_n9010_, new_n8956_);
  or g_153 (new_n6414_, or_not_new_n6250__not_new_n6371_, not_new_n1607__9);
  and g_154 (new_n4917_, new_n5212_, new_n5215_);
  not g_155 (not_new_n6635__5, new_n6635_);
  not g_156 (not_new_n5046_, new_n5046_);
  not g_157 (not_po298_0, po298);
  not g_158 (not_new_n7086_, new_n7086_);
  not g_159 (not_new_n3832_, new_n3832_);
  or g_160 (new_n6933_, not_new_n6518__0, not_new_n637__403536070);
  not g_161 (new_n6526_, new_n1055_);
  or g_162 (new_n8480_, not_new_n624__968890104070, not_new_n8108__0);
  not g_163 (not_new_n6532__0, new_n6532_);
  not g_164 (not_new_n4611_, new_n4611_);
  and g_165 (and_new_n3729__new_n3726_, new_n3726_, new_n3729_);
  not g_166 (not_new_n637__47475615099430, new_n637_);
  not g_167 (not_new_n634__70, new_n634_);
  or g_168 (new_n3165_, not_new_n928__332329305696010, not_new_n1057__3);
  not g_169 (new_n9933_, new_n625_);
  or g_170 (new_n4661_, not_pi178_2, not_new_n4448_);
  not g_171 (not_new_n1061__10, new_n1061_);
  or g_172 (new_n6635_, not_new_n6781_, not_new_n6824_);
  or g_173 (new_n4469_, not_new_n4715_, not_new_n4714_);
  or g_174 (new_n9056_, new_n627_, new_n1055_);
  or g_175 (new_n10065_, not_new_n10222_, not_new_n9981_);
  not g_176 (not_pi128_0, pi128);
  not g_177 (not_new_n607__70, new_n607_);
  not g_178 (not_new_n630__47475615099430, new_n630_);
  or g_179 (new_n5300_, not_new_n5056__0, not_new_n5255_);
  not g_180 (not_new_n10016__0, new_n10016_);
  not g_181 (not_new_n9627_, new_n9627_);
  not g_182 (new_n4424_, new_n1006_);
  or g_183 (new_n6826_, not_new_n6451__0, not_new_n6597_);
  not g_184 (not_new_n629__4, new_n629_);
  not g_185 (not_new_n3958_, new_n3958_);
  not g_186 (not_new_n3184__968890104070, new_n3184_);
  not g_187 (not_new_n1065__7, new_n1065_);
  not g_188 (not_new_n8011_, new_n8011_);
  not g_189 (not_new_n8104_, new_n8104_);
  not g_190 (not_new_n7421__1, new_n7421_);
  not g_191 (not_new_n1607_, new_n1607_);
  not g_192 (not_new_n591__19773267430, new_n591_);
  and g_193 (new_n8947_, new_n9082_, new_n8970_);
  or g_194 (new_n9025_, not_new_n8995_, not_new_n8799_);
  not g_195 (not_new_n5515__0, new_n5515_);
  not g_196 (not_new_n596__3, key_gate_88);
  not g_197 (not_new_n6002__0, new_n6002_);
  not g_198 (not_new_n6515_, new_n6515_);
  or g_199 (new_n7139_, not_new_n7251_, not_new_n7250_);
  not g_200 (not_new_n5878__2, new_n5878_);
  not g_201 (not_new_n9675_, new_n9675_);
  or g_202 (po133, not_new_n3480_, not_new_n3481_);
  not g_203 (not_new_n9398__0, new_n9398_);
  not g_204 (not_new_n5150_, new_n5150_);
  not g_205 (new_n4838_, new_n4773_);
  not g_206 (not_new_n1387_, new_n1387_);
  not g_207 (not_new_n3228_, new_n3228_);
  not g_208 (new_n7334_, new_n7018_);
  or g_209 (new_n1646_, not_pi037, not_new_n1631__3);
  or g_210 (new_n6209_, not_new_n6208_, not_new_n6072_);
  not g_211 (new_n4084_, pi253);
  not g_212 (not_new_n8325_, new_n8325_);
  not g_213 (not_new_n1601__1176490, new_n1601_);
  not g_214 (new_n4799_, new_n1061_);
  not g_215 (new_n5909_, new_n5809_);
  not g_216 (not_new_n632__138412872010, new_n632_);
  not g_217 (not_new_n7697_, new_n7697_);
  and g_218 (new_n9981_, new_n10064_, new_n9856_);
  not g_219 (not_new_n10213_, new_n10213_);
  not g_220 (not_new_n1536__39098210485829880490, new_n1536_);
  not g_221 (not_new_n994__8, new_n994_);
  not g_222 (not_new_n5597_, new_n5597_);
  not g_223 (not_new_n7040_, new_n7040_);
  or g_224 (new_n8503_, not_new_n8253__0, not_new_n8222_);
  not g_225 (new_n5468_, pi145);
  not g_226 (not_new_n8022_, new_n8022_);
  not g_227 (not_new_n1176_, new_n1176_);
  not g_228 (new_n7412_, new_n7031_);
  not g_229 (not_new_n633__5585458640832840070, new_n633_);
  not g_230 (new_n9709_, new_n9419_);
  and g_231 (new_n8664_, new_n8594_, new_n8770_);
  not g_232 (not_new_n7265_, new_n7265_);
  or g_233 (new_n5577_, not_new_n5576_, not_new_n5511_);
  not g_234 (not_new_n646__168070, new_n646_);
  not g_235 (not_new_n4127__0, new_n4127_);
  not g_236 (new_n4234_, new_n707_);
  not g_237 (not_po296_302268019717750559482470516839540966128657419430, po296);
  or g_238 (new_n9090_, new_n625_, new_n1602_);
  not g_239 (not_new_n598__168070, new_n598_);
  not g_240 (not_new_n8951_, new_n8951_);
  not g_241 (not_new_n9491__1, new_n9491_);
  or g_242 (new_n5366_, not_new_n1602__10, not_new_n4956__0);
  not g_243 (new_n7657_, new_n643_);
  not g_244 (not_pi145_0, pi145);
  not g_245 (not_pi113_0, pi113);
  not g_246 (not_new_n6048_, new_n6048_);
  or g_247 (new_n956_, or_or_not_new_n1279__not_new_n1277__not_new_n2021_, not_new_n2020_);
  not g_248 (not_new_n5266_, new_n5266_);
  not g_249 (new_n7230_, new_n7148_);
  or g_250 (or_not_new_n1806__not_new_n1807_, not_new_n1807_, not_new_n1806_);
  or g_251 (new_n1684_, key_gate_30, not_new_n596__1176490);
  not g_252 (not_new_n5446__0, new_n5446_);
  not g_253 (not_new_n5898__1, new_n5898_);
  or g_254 (new_n5832_, not_new_n6164_, not_new_n6165_);
  not g_255 (new_n8869_, new_n1061_);
  or g_256 (new_n3632_, not_pi182_0, not_new_n984__2824752490);
  or g_257 (new_n7805_, not_new_n7774_, not_new_n7618_);
  not g_258 (not_new_n5563_, new_n5563_);
  or g_259 (new_n959_, or_or_not_new_n1291__not_new_n1289__not_new_n2078_, not_new_n2077_);
  and g_260 (new_n1222_, and_and_new_n1746__new_n1747__new_n1749_, new_n1748_);
  or g_261 (or_or_not_new_n2964__not_new_n2967__not_new_n2966_, not_new_n2966_, or_not_new_n2964__not_new_n2967_);
  not g_262 (not_new_n9420_, new_n9420_);
  not g_263 (not_new_n6944_, new_n6944_);
  or g_264 (new_n2021_, not_new_n7682_, not_new_n1583__490);
  not g_265 (not_new_n1017__7, new_n1017_);
  not g_266 (not_new_n8501_, new_n8501_);
  not g_267 (not_new_n1003__4, new_n1003_);
  not g_268 (not_new_n5157_, new_n5157_);
  not g_269 (new_n8602_, new_n1047_);
  or g_270 (new_n9506_, not_new_n9699_, not_new_n9464_);
  and g_271 (new_n6333_, new_n6236_, and_and_and_new_n1043__new_n6232__new_n6229__new_n6317_);
  and g_272 (and_new_n2521__new_n2520_, new_n2520_, new_n2521_);
  or g_273 (new_n8734_, not_new_n8629_, not_new_n1037__2824752490);
  or g_274 (po066, not_new_n1193_, key_gate_62);
  not g_275 (not_new_n6242__2, new_n6242_);
  not g_276 (not_new_n1591__3430, new_n1591_);
  not g_277 (not_new_n3149_, new_n3149_);
  not g_278 (not_new_n1003__1, new_n1003_);
  or g_279 (new_n7833_, not_new_n637__2824752490, not_new_n7642_);
  xor g_280 (key_gate_22, key_22, new_n1657_);
  not g_281 (not_new_n4725__0, new_n4725_);
  not g_282 (not_new_n1028__70, new_n1028_);
  not g_283 (not_new_n1071__490, new_n1071_);
  or g_284 (po225, or_or_not_new_n2617__not_new_n2621__not_new_n1439_, not_new_n1438_);
  not g_285 (not_new_n9358__0, new_n9358_);
  or g_286 (new_n9146_, not_new_n9144_, not_new_n8953_);
  not g_287 (not_new_n7379_, new_n7379_);
  or g_288 (new_n4622_, not_new_n4421_, not_new_n1007__3);
  or g_289 (new_n3385_, not_pi053_0, not_new_n1534__16284135979104490);
  and g_290 (new_n1549_, new_n3611_, new_n3610_);
  not g_291 (not_new_n8118__2, new_n8118_);
  not g_292 (not_new_n1612__3, new_n1612_);
  not g_293 (not_po296_597682638941559493067901192655856192170251494124306816490, po296);
  not g_294 (not_new_n775__8, new_n775_);
  or g_295 (new_n2838_, not_new_n613__2, not_new_n1600__1);
  not g_296 (not_new_n6928_, new_n6928_);
  not g_297 (not_new_n639__24010, new_n639_);
  or g_298 (or_not_pi269_1_not_pi260_1, not_pi260_1, not_pi269_1);
  not g_299 (not_new_n3996_, new_n3996_);
  and g_300 (new_n8207_, new_n8467_, new_n8287_);
  not g_301 (not_new_n634__138412872010, new_n634_);
  not g_302 (not_new_n3454_, new_n3454_);
  not g_303 (new_n8603_, new_n1049_);
  and g_304 (new_n3998_, new_n4069_, new_n4070_);
  not g_305 (not_pi110_0, pi110);
  or g_306 (new_n10243_, not_new_n10241_, not_new_n10242_);
  not g_307 (not_new_n4549_, new_n4549_);
  not g_308 (not_new_n589__1, new_n589_);
  not g_309 (not_new_n646__19773267430, new_n646_);
  not g_310 (new_n6924_, new_n6604_);
  or g_311 (new_n9209_, not_new_n8829__0, not_new_n631__1915812313805664144010);
  not g_312 (not_new_n5991_, new_n5991_);
  not g_313 (not_new_n9121_, new_n9121_);
  not g_314 (not_new_n1583__1, new_n1583_);
  not g_315 (not_new_n1537__113988951853731430, new_n1537_);
  not g_316 (not_new_n10103__0, new_n10103_);
  or g_317 (new_n8331_, not_new_n8121__0, not_new_n8304__0);
  not g_318 (not_new_n8162__0, new_n8162_);
  or g_319 (new_n1740_, not_pi084, not_new_n1728__8);
  not g_320 (not_new_n2913_, new_n2913_);
  not g_321 (not_new_n1235_, new_n1235_);
  not g_322 (not_new_n587__10, new_n587_);
  or g_323 (new_n2506_, or_not_new_n4410__not_new_n609_, not_new_n611_);
  not g_324 (not_pi046_1, pi046);
  not g_325 (not_new_n2655_, new_n2655_);
  not g_326 (new_n6249_, new_n623_);
  or g_327 (or_not_new_n3088__not_new_n3087_, not_new_n3088_, not_new_n3087_);
  or g_328 (new_n1731_, not_new_n1728_, not_pi075);
  not g_329 (not_new_n6152_, new_n6152_);
  not g_330 (not_new_n1037__403536070, new_n1037_);
  not g_331 (not_pi028, pi028);
  not g_332 (not_new_n5890__1, new_n5890_);
  or g_333 (or_not_pi064_5585458640832840070_not_new_n4019__0, not_new_n4019__0, not_pi064_5585458640832840070);
  or g_334 (new_n7201_, not_new_n7077_, not_new_n7199_);
  not g_335 (not_new_n1560_, new_n1560_);
  or g_336 (or_or_not_new_n1255__not_new_n1253__not_new_n1907_, not_new_n1907_, or_not_new_n1255__not_new_n1253_);
  not g_337 (not_new_n10214_, new_n10214_);
  or g_338 (new_n10018_, not_new_n10132_, not_new_n10133_);
  or g_339 (new_n2064_, not_new_n1591__24010, not_new_n8918_);
  or g_340 (new_n9151_, not_new_n8982_, not_new_n9013_);
  not g_341 (not_pi120_0, pi120);
  not g_342 (not_new_n6818_, new_n6818_);
  not g_343 (not_new_n10321_, new_n10321_);
  not g_344 (not_new_n5413_, new_n5413_);
  not g_345 (not_new_n7219_, new_n7219_);
  and g_346 (and_and_new_n3768__new_n3771__new_n3777_, new_n3777_, and_new_n3768__new_n3771_);
  or g_347 (new_n9210_, not_new_n1043__138412872010, not_new_n8827_);
  or g_348 (or_or_not_new_n1554__not_new_n2429__not_new_n1377_, or_not_new_n1554__not_new_n2429_, not_new_n1377_);
  or g_349 (new_n5693_, not_new_n1017__7, not_new_n5457__0);
  not g_350 (not_new_n6686_, new_n6686_);
  or g_351 (new_n2801_, not_new_n4127__1, not_new_n994__9);
  not g_352 (not_new_n5517__0, new_n5517_);
  or g_353 (new_n7346_, not_new_n775__3, not_new_n7102_);
  not g_354 (not_pi115, pi115);
  or g_355 (new_n3886_, not_new_n626__490, not_new_n1576__16284135979104490);
  or g_356 (new_n6558_, not_new_n6952_, not_new_n6951_);
  or g_357 (new_n3225_, not_new_n633__7, not_new_n589__57648010);
  not g_358 (not_new_n6890_, new_n6890_);
  not g_359 (not_new_n7903_, new_n7903_);
  not g_360 (new_n6281_, new_n1035_);
  not g_361 (not_new_n1045__39098210485829880490, new_n1045_);
  not g_362 (not_new_n9512_, new_n9512_);
  or g_363 (new_n2208_, not_new_n4123_, not_new_n585__968890104070);
  not g_364 (not_new_n7258_, new_n7258_);
  not g_365 (not_new_n7755__0, new_n7755_);
  and g_366 (new_n8269_, new_n8567_, new_n8566_);
  or g_367 (new_n5009_, not_new_n5335_, not_new_n5336_);
  not g_368 (not_new_n6568_, new_n6568_);
  not g_369 (not_new_n8886__0, new_n8886_);
  not g_370 (not_new_n611__138412872010, new_n611_);
  or g_371 (new_n9185_, not_new_n9097__0, not_new_n1598__138412872010);
  and g_372 (new_n7701_, new_n7774_, new_n7956_);
  not g_373 (not_new_n3435_, new_n3435_);
  not g_374 (not_new_n605__0, new_n605_);
  not g_375 (not_new_n3227_, new_n3227_);
  or g_376 (new_n3233_, not_new_n644__7, not_new_n589__138412872010);
  not g_377 (not_new_n5878_, new_n5878_);
  not g_378 (not_new_n1372_, new_n1372_);
  not g_379 (not_new_n4014__3, new_n4014_);
  or g_380 (new_n6429_, or_or_not_new_n6343__not_new_n6344__not_new_n6345_, not_new_n6242__4);
  not g_381 (not_new_n9497_, new_n9497_);
  not g_382 (not_new_n7924_, new_n7924_);
  not g_383 (not_new_n1361_, new_n1361_);
  not g_384 (not_new_n7921_, new_n7921_);
  not g_385 (not_new_n581__17984650426474121466202803405696493492512490, new_n581_);
  not g_386 (not_new_n5812__0, new_n5812_);
  or g_387 (or_not_new_n4831__not_new_n4789_, not_new_n4789_, not_new_n4831_);
  or g_388 (po073, not_new_n1200_, key_gate_51);
  not g_389 (not_new_n8812_, new_n8812_);
  or g_390 (or_not_new_n2831__not_new_n1481_, not_new_n1481_, not_new_n2831_);
  not g_391 (not_new_n6443__8235430, new_n6443_);
  or g_392 (new_n7561_, not_new_n6999__1, not_new_n7033__1);
  or g_393 (new_n7519_, not_new_n7003__0, not_new_n7036__0);
  or g_394 (new_n6888_, not_new_n6626_, not_new_n6594_);
  not g_395 (not_new_n617__1915812313805664144010, new_n617_);
  or g_396 (new_n3035_, not_new_n1164_, not_new_n1027__57648010);
  and g_397 (new_n1533_, new_n3301_, new_n3303_);
  not g_398 (not_new_n5721_, new_n5721_);
  or g_399 (new_n6844_, not_new_n1043__24010, not_new_n6488__0);
  and g_400 (and_new_n3085__new_n998_, new_n998_, new_n3085_);
  not g_401 (not_new_n6617__1, new_n6617_);
  and g_402 (new_n4142_, pi261, pi259);
  not g_403 (not_po296_16284135979104490, po296);
  not g_404 (not_new_n1601__2326305139872070, new_n1601_);
  or g_405 (or_or_not_new_n1327__not_new_n1325__not_new_n2249_, or_not_new_n1327__not_new_n1325_, not_new_n2249_);
  or g_406 (new_n1028_, not_new_n3383_, not_new_n3382_);
  not g_407 (not_new_n1591__490, new_n1591_);
  not g_408 (not_new_n1574_, new_n1574_);
  or g_409 (new_n2392_, not_new_n603__7, not_new_n647__1);
  not g_410 (not_new_n4959_, new_n4959_);
  or g_411 (new_n5700_, not_new_n1018__7, not_new_n5455__0);
  not g_412 (not_new_n1829_, new_n1829_);
  not g_413 (not_new_n6233__2, new_n6233_);
  or g_414 (new_n7834_, not_new_n638__47475615099430, not_new_n7643_);
  not g_415 (not_new_n9425__0, new_n9425_);
  not g_416 (not_new_n4384_, new_n4384_);
  not g_417 (not_new_n1607__403536070, new_n1607_);
  or g_418 (new_n7395_, not_new_n7115__0, not_new_n7114_);
  or g_419 (new_n2699_, not_po296_63668057609090279857414351392240010, not_pi255_1);
  not g_420 (not_new_n2345_, new_n2345_);
  not g_421 (not_new_n1631__9, key_gate_76);
  and g_422 (new_n611_, new_n590_, new_n988_);
  not g_423 (not_new_n10038_, new_n10038_);
  not g_424 (not_new_n7562_, new_n7562_);
  not g_425 (not_new_n5439__0, new_n5439_);
  not g_426 (new_n5793_, new_n1055_);
  not g_427 (not_pi093, pi093);
  not g_428 (not_pi151_0, pi151);
  not g_429 (new_n4827_, new_n4739_);
  not g_430 (not_new_n6821_, new_n6821_);
  not g_431 (not_new_n3782_, new_n3782_);
  not g_432 (not_new_n7015_, new_n7015_);
  not g_433 (not_new_n9427__1, new_n9427_);
  not g_434 (not_new_n7605_, new_n7605_);
  or g_435 (new_n7213_, not_new_n7412__0, not_new_n6998__0);
  not g_436 (not_new_n8582_, new_n8582_);
  or g_437 (new_n9719_, not_new_n9512__2, not_new_n9378_);
  or g_438 (new_n3085_, not_new_n3372__13410686196639649008070, not_new_n641__2);
  not g_439 (not_new_n593__1, new_n593_);
  not g_440 (not_new_n1051__5, new_n1051_);
  not g_441 (not_new_n8772_, new_n8772_);
  or g_442 (new_n8287_, not_new_n8103_, not_new_n1047__8235430);
  not g_443 (not_new_n7643__0, new_n7643_);
  not g_444 (not_new_n1728__7, new_n1728_);
  not g_445 (not_new_n4752_, new_n4752_);
  not g_446 (not_pi064_6782230728490, pi064);
  or g_447 (new_n8717_, not_new_n1597__968890104070, not_new_n8656_);
  or g_448 (new_n3693_, not_po298_403536070, not_new_n645__9);
  not g_449 (not_new_n5440__1, new_n5440_);
  not g_450 (not_new_n4419_, new_n4419_);
  not g_451 (not_new_n7811_, new_n7811_);
  not g_452 (not_pi155, pi155);
  not g_453 (not_new_n4135__2, new_n4135_);
  not g_454 (not_new_n1606__7, new_n1606_);
  and g_455 (new_n606_, new_n3369_, new_n592_);
  or g_456 (new_n6731_, not_new_n640__57648010, not_new_n6512_);
  or g_457 (new_n3829_, not_new_n648__70, not_new_n6443__0);
  not g_458 (not_new_n6473__0, new_n6473_);
  or g_459 (new_n6705_, not_new_n6527_, not_new_n626__138412872010);
  not g_460 (not_new_n8272_, new_n8272_);
  not g_461 (not_new_n8227_, new_n8227_);
  or g_462 (or_not_new_n6343__not_new_n6344_, not_new_n6344_, not_new_n6343_);
  or g_463 (new_n4381_, not_new_n4310_, not_new_n4378_);
  or g_464 (new_n9830_, not_new_n9591_, not_new_n9828_);
  not g_465 (not_new_n4267_, new_n4267_);
  not g_466 (not_new_n3164_, new_n3164_);
  or g_467 (new_n8125_, not_new_n8306_, not_new_n8122_);
  not g_468 (not_new_n7812_, new_n7812_);
  not g_469 (not_new_n6990__0, new_n6990_);
  not g_470 (not_new_n9186_, new_n9186_);
  or g_471 (new_n8367_, not_new_n8082_, not_new_n8366_);
  not g_472 (not_new_n2017_, new_n2017_);
  or g_473 (new_n4613_, not_new_n4478_, not_new_n4479__0);
  or g_474 (new_n1636_, not_new_n596__0, key_gate_60);
  not g_475 (not_new_n607__168070, new_n607_);
  or g_476 (new_n3076_, not_new_n3372__39098210485829880490, not_new_n627__4);
  or g_477 (new_n5415_, not_new_n5000__0, not_new_n5264_);
  not g_478 (not_new_n1534__70, key_gate_5);
  or g_479 (new_n8299_, not_new_n8118_, not_new_n1045__968890104070);
  not g_480 (not_new_n1588__9, new_n1588_);
  or g_481 (new_n5735_, not_new_n5962_, not_new_n5959_);
  not g_482 (not_po296_47475615099430, po296);
  not g_483 (not_new_n4750_, new_n4750_);
  not g_484 (not_new_n9998_, new_n9998_);
  not g_485 (new_n7778_, new_n7652_);
  not g_486 (not_new_n643__0, new_n643_);
  or g_487 (new_n3218_, not_new_n1037__4, not_new_n3185__168070);
  or g_488 (new_n3125_, not_new_n629__5, not_new_n3315__3430);
  not g_489 (not_new_n1654_, key_gate_25);
  or g_490 (new_n7443_, not_new_n7129_, not_new_n775__968890104070);
  or g_491 (or_not_new_n6160__not_new_n6161_, not_new_n6161_, not_new_n6160_);
  or g_492 (new_n4110_, not_pi247_0, not_new_n4173_);
  or g_493 (new_n7035_, not_new_n7423_, not_new_n7422_);
  and g_494 (new_n8974_, new_n9297_, new_n9296_);
  and g_495 (new_n1243_, and_new_n1242__new_n1856_, new_n1855_);
  not g_496 (not_new_n589__63668057609090279857414351392240010, new_n589_);
  and g_497 (new_n6643_, new_n6956_, new_n6957_);
  not g_498 (not_new_n4234_, new_n4234_);
  or g_499 (or_not_new_n1287__not_new_n1285_, not_new_n1285_, not_new_n1287_);
  not g_500 (not_pi058_0, pi058);
  not g_501 (not_new_n6637_, new_n6637_);
  not g_502 (not_new_n625__6, new_n625_);
  or g_503 (new_n6368_, not_new_n6271_, not_new_n1045__24010);
  or g_504 (new_n2380_, not_new_n598__4, not_new_n1043__0);
  and g_505 (new_n7070_, new_n7027_, new_n7165_);
  not g_506 (not_new_n4954_, new_n4954_);
  or g_507 (new_n4065_, not_pi034_3, not_new_n3994_);
  or g_508 (new_n4676_, not_new_n4443__0, not_new_n1014__4);
  not g_509 (not_pi035_3, pi035);
  not g_510 (not_new_n7088_, new_n7088_);
  or g_511 (new_n690_, not_new_n1510_, not_new_n3038_);
  not g_512 (not_pi171, pi171);
  not g_513 (not_new_n595__10, new_n595_);
  or g_514 (new_n6866_, not_new_n6462_, or_not_new_n6541__0_not_new_n1596__1176490);
  or g_515 (new_n742_, not_new_n3258_, not_new_n3257_);
  not g_516 (not_new_n1371_, new_n1371_);
  or g_517 (new_n6608_, not_new_n6943_, not_new_n6944_);
  and g_518 (new_n8674_, new_n8730_, new_n8729_);
  not g_519 (not_new_n1049__16284135979104490, new_n1049_);
  not g_520 (not_new_n3219_, new_n3219_);
  not g_521 (not_new_n1596__9, new_n1596_);
  or g_522 (new_n7047_, not_new_n7568_, not_new_n7569_);
  or g_523 (new_n4853_, not_new_n4754_, not_new_n4845_);
  or g_524 (new_n8914_, not_new_n9269_, not_new_n9268_);
  not g_525 (new_n8004_, new_n7719_);
  or g_526 (new_n3563_, not_new_n1612__8235430, not_new_n2128__0);
  or g_527 (new_n4373_, not_new_n692_, not_new_n4264_);
  not g_528 (new_n5913_, new_n5748_);
  not g_529 (not_new_n5457__0, new_n5457_);
  or g_530 (new_n3850_, not_new_n617__490, not_new_n1576__10);
  and g_531 (new_n8671_, new_n8733_, new_n8670_);
  or g_532 (new_n9586_, not_new_n9335_, not_new_n9506_);
  and g_533 (new_n6610_, new_n6447_, new_n6775_);
  not g_534 (not_new_n635__2824752490, new_n635_);
  not g_535 (not_new_n3322_, new_n3322_);
  or g_536 (new_n3154_, not_new_n637__6, not_new_n581__1070069044235980333563563003849377848070);
  not g_537 (not_new_n4956__0, new_n4956_);
  or g_538 (or_or_or_not_new_n8528__not_new_n8429__not_new_n8457__not_new_n8458_, not_new_n8458_, or_or_not_new_n8528__not_new_n8429__not_new_n8457_);
  not g_539 (new_n5747_, new_n632_);
  not g_540 (not_new_n7859_, new_n7859_);
  or g_541 (new_n7045_, not_new_n7404_, not_new_n7405_);
  not g_542 (not_new_n7603__0, new_n7603_);
  and g_543 (new_n8930_, new_n9025_, new_n9027_);
  or g_544 (new_n4709_, not_new_n1019__3, not_new_n4433_);
  or g_545 (or_not_new_n2865__not_new_n2868_, not_new_n2868_, not_new_n2865_);
  not g_546 (not_new_n6250_, new_n6250_);
  not g_547 (not_new_n1576__2326305139872070, new_n1576_);
  or g_548 (po244, not_new_n3675_, not_new_n3674_);
  not g_549 (not_new_n9750_, new_n9750_);
  not g_550 (not_new_n5719_, new_n5719_);
  not g_551 (not_new_n638__168070, new_n638_);
  not g_552 (new_n6270_, new_n636_);
  or g_553 (new_n1030_, not_new_n3391_, not_new_n3392_);
  not g_554 (not_new_n1729_, new_n1729_);
  not g_555 (not_new_n989__490, new_n989_);
  not g_556 (not_new_n6345_, new_n6345_);
  not g_557 (not_new_n4139_, new_n4139_);
  not g_558 (not_new_n7643__2, new_n7643_);
  xnor g_559 (key_gate_34, key_34, new_n1675_);
  not g_560 (not_new_n9176_, new_n9176_);
  xnor g_561 (key_gate_53, not_new_n3922_, key_53);
  or g_562 (or_or_or_not_new_n2803__not_new_n2806__not_new_n2805__not_new_n2807_, not_new_n2807_, or_or_not_new_n2803__not_new_n2806__not_new_n2805_);
  not g_563 (not_new_n9915__0, new_n9915_);
  or g_564 (new_n8765_, not_new_n1603__2824752490, not_new_n8644_);
  not g_565 (not_new_n4269_, new_n4269_);
  or g_566 (new_n6561_, not_new_n6847_, not_new_n6846_);
  not g_567 (not_new_n604__968890104070, new_n604_);
  not g_568 (not_new_n8942_, new_n8942_);
  not g_569 (not_new_n6036_, new_n6036_);
  not g_570 (not_new_n587__5, new_n587_);
  not g_571 (not_new_n736__0, new_n736_);
  or g_572 (new_n3143_, not_new_n3315__403536070, not_new_n642__4);
  not g_573 (not_new_n1571_, new_n1571_);
  not g_574 (not_new_n4545_, new_n4545_);
  not g_575 (not_new_n7134_, new_n7134_);
  not g_576 (not_new_n3764_, new_n3764_);
  not g_577 (not_new_n6782_, new_n6782_);
  or g_578 (new_n2890_, not_new_n4126__1, not_new_n994__403536070);
  not g_579 (not_new_n581__1299348114471230201171721456984490, new_n581_);
  or g_580 (new_n5614_, not_new_n5500__0, not_new_n5499_);
  not g_581 (not_new_n2339_, new_n2339_);
  not g_582 (not_new_n4798_, new_n4798_);
  not g_583 (not_new_n7011__0, new_n7011_);
  not g_584 (not_new_n2434_, new_n2434_);
  not g_585 (not_new_n10178_, new_n10178_);
  or g_586 (new_n10215_, not_new_n9894_, not_new_n9863_);
  buf g_587 (po046, pi218);
  not g_588 (not_new_n1492_, new_n1492_);
  and g_589 (new_n4505_, new_n4703_, new_n4702_);
  or g_590 (new_n9792_, not_new_n9384_, not_new_n1602__332329305696010);
  not g_591 (not_new_n3257_, new_n3257_);
  or g_592 (new_n5304_, not_new_n4934_, not_new_n635__24010);
  or g_593 (or_not_new_n7664__0_not_new_n618__6782230728490, not_new_n618__6782230728490, not_new_n7664__0);
  not g_594 (not_new_n757_, new_n757_);
  not g_595 (not_new_n3208_, new_n3208_);
  not g_596 (new_n4260_, new_n662_);
  not g_597 (not_new_n8111__0, new_n8111_);
  not g_598 (not_new_n5560_, new_n5560_);
  or g_599 (new_n8965_, not_new_n8944_, not_new_n9101_);
  not g_600 (not_new_n5598_, new_n5598_);
  or g_601 (new_n9525_, not_new_n9450_, not_new_n9326_);
  not g_602 (not_new_n8982__0, new_n8982_);
  not g_603 (not_new_n5630__0, new_n5630_);
  not g_604 (not_new_n1601__39098210485829880490, new_n1601_);
  not g_605 (not_new_n6468_, new_n6468_);
  or g_606 (new_n7693_, not_new_n8058_, not_new_n8057_);
  or g_607 (new_n4185_, not_new_n4147_, not_pi260_4);
  or g_608 (new_n9127_, not_new_n640__6782230728490, not_new_n1604__138412872010);
  or g_609 (new_n2593_, not_new_n609__8, not_new_n4469_);
  not g_610 (not_new_n5528_, new_n5528_);
  not g_611 (not_pi005_0, pi005);
  and g_612 (new_n1218_, and_and_new_n1735__new_n1736__new_n1738_, new_n1737_);
  not g_613 (not_new_n5900__0, new_n5900_);
  or g_614 (new_n5148_, new_n626_, new_n1053_);
  or g_615 (new_n8754_, not_new_n8679_, not_new_n8595__4);
  not g_616 (not_pi274_1, pi274);
  or g_617 (new_n10280_, not_new_n10278_, not_new_n10152_);
  or g_618 (new_n2901_, not_new_n3311__490, not_new_n1035__1);
  or g_619 (new_n10275_, not_new_n1596__1915812313805664144010, not_new_n9945_);
  not g_620 (new_n4751_, new_n1049_);
  or g_621 (new_n2668_, not_new_n610__168070, not_new_n4459__0);
  not g_622 (not_new_n617__5585458640832840070, new_n617_);
  or g_623 (or_not_new_n9469__not_new_n9339_, not_new_n9469_, not_new_n9339_);
  not g_624 (new_n5770_, new_n630_);
  and g_625 (and_and_new_n1953__new_n1956__new_n1954_, new_n1954_, and_new_n1953__new_n1956_);
  not g_626 (not_new_n8547_, new_n8547_);
  not g_627 (not_new_n1041__168070, new_n1041_);
  not g_628 (not_new_n7711_, new_n7711_);
  not g_629 (not_new_n2533_, new_n2533_);
  and g_630 (new_n4138_, pi256, pi266);
  not g_631 (not_new_n7451__0, new_n7451_);
  or g_632 (new_n2385_, not_new_n1045__0, not_new_n598__5);
  and g_633 (new_n4781_, new_n4873_, new_n4872_);
  not g_634 (not_new_n5768_, new_n5768_);
  or g_635 (new_n2176_, not_new_n1581__2824752490, not_new_n8197_);
  or g_636 (new_n1644_, not_po296_3, not_pi028);
  or g_637 (new_n8743_, not_new_n8606_, not_new_n1154__0);
  or g_638 (new_n2670_, not_new_n1008__0, not_new_n608__168070);
  or g_639 (new_n3008_, not_new_n1155_, not_new_n1027__9);
  or g_640 (new_n5206_, not_new_n5063__0, not_new_n1596__8);
  and g_641 (new_n9984_, new_n9854_, new_n10078_);
  or g_642 (new_n2698_, not_new_n4452__0, not_new_n610__57648010);
  not g_643 (not_new_n9412__1, new_n9412_);
  not g_644 (not_new_n10035_, new_n10035_);
  or g_645 (new_n3627_, not_new_n961_, not_new_n1611__8235430);
  not g_646 (new_n9935_, new_n630_);
  not g_647 (new_n4785_, new_n1035_);
  or g_648 (new_n9814_, not_new_n9812_, not_new_n9813_);
  or g_649 (new_n4366_, not_new_n4305_, not_new_n4363_);
  or g_650 (new_n1713_, not_pi005_0, not_po296_332329305696010);
  not g_651 (not_pi142_3, pi142);
  or g_652 (new_n2375_, not_new_n1041__0, not_new_n598__3);
  not g_653 (not_new_n6927_, new_n6927_);
  not g_654 (not_new_n1631__138412872010, key_gate_76);
  not g_655 (not_new_n3916_, new_n3916_);
  not g_656 (not_new_n9291_, new_n9291_);
  not g_657 (not_new_n10045__0, new_n10045_);
  not g_658 (not_new_n624__19773267430, new_n624_);
  not g_659 (not_new_n3501_, new_n3501_);
  and g_660 (new_n1474_, new_n1592_, and_new_n3315__new_n923_);
  not g_661 (not_new_n8160_, new_n8160_);
  not g_662 (not_new_n3277_, new_n3277_);
  not g_663 (not_new_n2606_, new_n2606_);
  and g_664 (new_n1380_, new_n2436_, new_n2435_);
  not g_665 (not_new_n2229_, new_n2229_);
  not g_666 (not_new_n9541_, new_n9541_);
  or g_667 (new_n2571_, not_new_n606__5, not_new_n5489__0);
  not g_668 (not_new_n6991__0, new_n6991_);
  not g_669 (not_new_n4313_, new_n4313_);
  not g_670 (not_new_n9166_, new_n9166_);
  not g_671 (not_new_n8527_, new_n8527_);
  not g_672 (not_new_n7418_, new_n7418_);
  or g_673 (new_n1874_, not_new_n1591__4, not_new_n8819_);
  or g_674 (new_n4512_, not_new_n4511_, not_pi162_1);
  not g_675 (not_new_n1035__10, new_n1035_);
  not g_676 (not_new_n6546_, new_n6546_);
  and g_677 (new_n4791_, new_n4881_, new_n4880_);
  not g_678 (not_new_n2819_, new_n2819_);
  not g_679 (not_new_n601__8235430, new_n601_);
  not g_680 (not_new_n600__3, new_n600_);
  not g_681 (not_new_n9356_, new_n9356_);
  not g_682 (new_n5769_, new_n1600_);
  not g_683 (not_new_n2039_, new_n2039_);
  not g_684 (not_new_n5700_, new_n5700_);
  or g_685 (new_n7958_, not_new_n7602__0, not_new_n634__138412872010);
  or g_686 (new_n3741_, not_new_n3739_, not_new_n3740_);
  not g_687 (not_new_n9953__0, new_n9953_);
  not g_688 (not_new_n1043__490, new_n1043_);
  or g_689 (new_n3894_, not_new_n3896_, not_new_n3895_);
  not g_690 (not_new_n645__968890104070, new_n645_);
  or g_691 (or_not_new_n2946__not_new_n2949_, not_new_n2949_, not_new_n2946_);
  or g_692 (new_n7506_, not_new_n744__0, not_new_n7345__0);
  not g_693 (new_n8443_, new_n8178_);
  not g_694 (not_pi075, pi075);
  not g_695 (not_new_n1613__2824752490, new_n1613_);
  not g_696 (not_new_n641__3430, new_n641_);
  or g_697 (new_n3695_, not_new_n640__9, not_po298_2824752490);
  not g_698 (new_n4081_, pi251);
  not g_699 (not_new_n3961_, new_n3961_);
  not g_700 (not_new_n1366_, new_n1366_);
  not g_701 (not_pi064_113988951853731430, pi064);
  not g_702 (not_new_n2047_, new_n2047_);
  not g_703 (not_new_n1603__8, new_n1603_);
  or g_704 (new_n8325_, not_new_n8324_, not_new_n8209_);
  not g_705 (not_new_n1059__332329305696010, new_n1059_);
  or g_706 (new_n10169_, not_new_n10168_, not_new_n10318_);
  not g_707 (not_new_n594__10, new_n594_);
  not g_708 (not_new_n634__168070, new_n634_);
  and g_709 (and_new_n1053__new_n6232_, new_n6232_, new_n1053_);
  and g_710 (new_n6235_, new_n6317_, new_n6239_);
  not g_711 (not_new_n625__273687473400809163430, new_n625_);
  or g_712 (new_n644_, or_or_not_new_n1996__not_new_n1997__not_new_n1999_, not_new_n1998_);
  or g_713 (new_n5809_, not_new_n5918_, not_new_n6138_);
  or g_714 (new_n2160_, not_new_n4915_, not_new_n1589__403536070);
  or g_715 (new_n2811_, not_new_n602__8, not_new_n1478_);
  not g_716 (not_new_n6113_, new_n6113_);
  or g_717 (new_n2501_, not_new_n1606__0, not_new_n598__113988951853731430);
  or g_718 (new_n7271_, not_new_n7088_, not_new_n7270_);
  not g_719 (not_new_n6490__0, new_n6490_);
  or g_720 (new_n7423_, not_new_n759_, not_new_n6974__168070);
  not g_721 (not_new_n4728__0, new_n4728_);
  and g_722 (new_n6232_, new_n6370_, and_and_new_n6374__new_n6372__new_n6371_);
  not g_723 (not_new_n6941_, new_n6941_);
  or g_724 (new_n6779_, not_new_n6484_, not_new_n641__168070);
  or g_725 (new_n2979_, not_new_n602__2326305139872070, not_new_n648__3);
  or g_726 (new_n6112_, not_new_n624__1176490, not_new_n5744__0);
  not g_727 (not_new_n4993_, new_n4993_);
  and g_728 (new_n1409_, new_n987_, new_n1408_);
  not g_729 (not_new_n1049__2824752490, new_n1049_);
  not g_730 (not_new_n678_, new_n678_);
  or g_731 (new_n2864_, or_not_new_n2863__not_new_n2862_, not_new_n2861_);
  not g_732 (not_new_n8267__0, new_n8267_);
  not g_733 (not_new_n7927_, new_n7927_);
  not g_734 (not_new_n9272_, new_n9272_);
  or g_735 (po197, not_new_n1378_, or_or_not_new_n1554__not_new_n2429__not_new_n1377_);
  or g_736 (new_n4702_, not_new_n1018__3, not_new_n4435_);
  not g_737 (not_new_n3363_, new_n3363_);
  not g_738 (not_new_n8315_, new_n8315_);
  not g_739 (not_new_n1598__332329305696010, new_n1598_);
  not g_740 (not_new_n1589__1176490, new_n1589_);
  not g_741 (not_new_n598__6782230728490, new_n598_);
  not g_742 (not_new_n7461_, new_n7461_);
  or g_743 (new_n2074_, not_new_n588__1176490, not_pi114);
  not g_744 (not_new_n3310__8, new_n3310_);
  not g_745 (not_new_n5415_, new_n5415_);
  and g_746 (new_n9875_, new_n10065_, new_n10226_);
  not g_747 (not_new_n7393_, new_n7393_);
  or g_748 (new_n7315_, not_new_n7345_, not_new_n6985_);
  or g_749 (new_n9088_, not_new_n9085_, not_new_n9087_);
  and g_750 (new_n4317_, new_n4400_, new_n4401_);
  not g_751 (not_new_n8973_, new_n8973_);
  or g_752 (new_n989_, not_pi275_1, not_new_n1621_);
  or g_753 (new_n7375_, not_new_n7373_, not_new_n7323_);
  or g_754 (new_n5831_, not_new_n6145_, not_new_n6146_);
  not g_755 (not_new_n603__968890104070, new_n603_);
  not g_756 (not_new_n1061__1176490, new_n1061_);
  not g_757 (not_new_n3550_, new_n3550_);
  not g_758 (new_n3390_, new_n1029_);
  not g_759 (not_new_n2132_, new_n2132_);
  not g_760 (not_new_n9473_, new_n9473_);
  or g_761 (new_n2086_, not_new_n594__168070, not_new_n9969_);
  not g_762 (not_new_n4986_, new_n4986_);
  not g_763 (not_new_n10160_, new_n10160_);
  not g_764 (not_new_n7122_, new_n7122_);
  not g_765 (not_new_n1728__490, new_n1728_);
  not g_766 (not_new_n6234__0, new_n6234_);
  not g_767 (not_new_n628__3, new_n628_);
  not g_768 (not_new_n4730_, new_n4730_);
  not g_769 (not_new_n640__403536070, new_n640_);
  not g_770 (not_new_n1055__797922662976120010, new_n1055_);
  not g_771 (not_new_n5292_, new_n5292_);
  or g_772 (new_n7228_, not_new_n7225_, not_new_n728_);
  or g_773 (new_n3209_, not_new_n589__10, not_new_n629__7);
  and g_774 (and_new_n7791__new_n7786_, new_n7786_, new_n7791_);
  not g_775 (not_new_n4387_, new_n4387_);
  not g_776 (not_new_n8809_, new_n8809_);
  not g_777 (not_new_n10153_, new_n10153_);
  not g_778 (not_new_n648__6, new_n648_);
  or g_779 (or_not_new_n2944__not_new_n2943_, not_new_n2944_, not_new_n2943_);
  not g_780 (not_new_n5481_, new_n5481_);
  not g_781 (not_new_n7014__2, new_n7014_);
  not g_782 (not_new_n1602__7, new_n1602_);
  not g_783 (not_new_n4248_, new_n4248_);
  not g_784 (not_new_n8265_, new_n8265_);
  not g_785 (not_new_n1051__6782230728490, new_n1051_);
  or g_786 (new_n4966_, not_new_n1055__9, not_new_n627__24010);
  not g_787 (not_new_n8526_, new_n8526_);
  and g_788 (and_and_new_n1896__new_n1899__new_n1897_, new_n1897_, and_new_n1896__new_n1899_);
  or g_789 (new_n7441_, not_new_n755_, not_new_n6974__19773267430);
  or g_790 (new_n619_, not_new_n2302_, or_or_not_new_n2300__not_new_n2301__not_new_n2303_);
  or g_791 (new_n9260_, not_new_n9259_, not_new_n9258_);
  not g_792 (not_new_n1057__4, new_n1057_);
  and g_793 (and_new_n1539__new_n2356_, new_n2356_, new_n1539_);
  and g_794 (and_new_n8837__new_n9203_, new_n8837_, new_n9203_);
  not g_795 (new_n6518_, new_n1065_);
  not g_796 (not_new_n3811_, new_n3811_);
  not g_797 (not_new_n1601__2824752490, new_n1601_);
  or g_798 (po273, or_or_or_not_new_n2785__not_new_n2788__not_new_n2787__not_new_n2789_, not_new_n2786_);
  not g_799 (not_new_n5740_, new_n5740_);
  not g_800 (not_new_n9376__0, new_n9376_);
  not g_801 (not_pi275_1, pi275);
  not g_802 (not_new_n7477_, new_n7477_);
  or g_803 (new_n6181_, not_new_n5781__0, not_new_n645__1176490);
  not g_804 (not_new_n605__4, new_n605_);
  not g_805 (not_new_n6558_, new_n6558_);
  not g_806 (new_n5454_, pi139);
  or g_807 (new_n5326_, not_new_n1607__6, not_new_n5058__0);
  or g_808 (new_n1051_, not_new_n3447_, not_new_n3448_);
  not g_809 (not_new_n3205_, new_n3205_);
  not g_810 (not_new_n1596__24010, new_n1596_);
  not g_811 (new_n4321_, new_n711_);
  not g_812 (not_new_n612_, new_n612_);
  and g_813 (new_n8924_, new_n628_, new_n1039_);
  or g_814 (new_n8764_, not_new_n8596__2, not_new_n8685_);
  or g_815 (new_n10334_, not_new_n1067__2326305139872070, not_new_n9914_);
  and g_816 (new_n1496_, new_n3019_, new_n1497_);
  not g_817 (not_new_n734_, new_n734_);
  or g_818 (new_n9254_, not_new_n9160_, not_new_n8966__0);
  or g_819 (new_n2485_, not_new_n598__47475615099430, not_new_n1598__0);
  or g_820 (new_n2797_, not_new_n6968_, not_new_n595__6);
  not g_821 (not_new_n639__5, new_n639_);
  or g_822 (new_n7556_, not_new_n7153__0, not_new_n7309_);
  not g_823 (not_new_n4756__0, new_n4756_);
  not g_824 (not_new_n10058_, new_n10058_);
  not g_825 (not_new_n1018__1, new_n1018_);
  not g_826 (not_new_n5082__0, new_n5082_);
  or g_827 (new_n4713_, not_new_n4712_, not_new_n4711_);
  or g_828 (po067, key_gate_118, not_new_n1194_);
  not g_829 (not_new_n4304_, new_n4304_);
  not g_830 (not_new_n4115__2, new_n4115_);
  or g_831 (new_n10295_, not_new_n629__113988951853731430, not_new_n9938_);
  not g_832 (not_new_n3311__3430, new_n3311_);
  not g_833 (not_pi255_1, pi255);
  not g_834 (not_new_n9057_, new_n9057_);
  not g_835 (not_new_n6023_, new_n6023_);
  not g_836 (not_new_n1061__24010, new_n1061_);
  or g_837 (new_n2695_, not_new_n605__57648010, not_new_n5475_);
  not g_838 (not_new_n937_, new_n937_);
  or g_839 (new_n8361_, not_new_n1604__57648010, not_new_n8141_);
  not g_840 (not_new_n931_, new_n931_);
  not g_841 (new_n7225_, new_n6993_);
  or g_842 (new_n7340_, not_new_n775__1, not_new_n7100_);
  not g_843 (not_new_n1603__3430, new_n1603_);
  not g_844 (not_new_n7127_, new_n7127_);
  or g_845 (new_n6793_, not_new_n6456_, not_new_n6544_);
  or g_846 (new_n3822_, not_new_n1590_, not_new_n8598_);
  or g_847 (new_n2568_, not_new_n4466__0, not_new_n610__5);
  not g_848 (not_new_n5870_, new_n5870_);
  not g_849 (not_new_n1014__5, new_n1014_);
  or g_850 (new_n6735_, not_new_n6658_, not_new_n6450_);
  not g_851 (not_new_n1605__3, new_n1605_);
  or g_852 (new_n9124_, not_new_n9123_, not_new_n8898__0);
  not g_853 (not_new_n3221_, new_n3221_);
  or g_854 (new_n8514_, not_new_n8255_, not_new_n8441_);
  and g_855 (new_n7099_, new_n7336_, new_n7335_);
  not g_856 (not_new_n1534__968890104070, key_gate_5);
  xnor g_857 (key_gate_94, not_new_n1702_, key_94);
  not g_858 (not_new_n6516_, new_n6516_);
  or g_859 (new_n4188_, not_pi269_5, not_new_n4076_);
  and g_860 (new_n1379_, new_n2432_, new_n2433_);
  or g_861 (new_n3122_, not_new_n622__5, not_new_n3315__490);
  not g_862 (not_new_n2924_, new_n2924_);
  not g_863 (not_new_n2834_, new_n2834_);
  or g_864 (new_n7852_, not_new_n7631_, not_new_n625__968890104070);
  not g_865 (not_new_n7109__0, new_n7109_);
  or g_866 (or_or_not_new_n2973__not_new_n2976__not_new_n2975_, not_new_n2975_, or_not_new_n2973__not_new_n2976_);
  and g_867 (new_n1313_, new_n2194_, new_n2193_);
  or g_868 (new_n7814_, not_new_n1045__19773267430, not_new_n7611__1);
  not g_869 (not_new_n7582_, new_n7582_);
  not g_870 (not_new_n9921_, new_n9921_);
  not g_871 (not_new_n9035_, new_n9035_);
  not g_872 (not_new_n7731_, new_n7731_);
  not g_873 (not_new_n3258_, new_n3258_);
  and g_874 (new_n4759_, new_n4855_, new_n4854_);
  not g_875 (not_new_n7030_, new_n7030_);
  or g_876 (new_n2823_, not_new_n7048_, not_new_n595__9);
  not g_877 (not_new_n2882_, new_n2882_);
  not g_878 (not_new_n6136_, new_n6136_);
  not g_879 (not_new_n9354_, new_n9354_);
  not g_880 (not_new_n9879__0, new_n9879_);
  not g_881 (not_new_n1005__3, new_n1005_);
  and g_882 (and_new_n3016__new_n998_, new_n998_, new_n3016_);
  not g_883 (not_new_n770_, new_n770_);
  not g_884 (not_new_n4737__0, new_n4737_);
  not g_885 (not_new_n7501_, new_n7501_);
  not g_886 (not_new_n1154__0, new_n1154_);
  and g_887 (new_n8274_, new_n8587_, new_n8588_);
  not g_888 (not_new_n7155_, new_n7155_);
  not g_889 (not_new_n1013_, new_n1013_);
  or g_890 (new_n709_, not_new_n1495_, not_new_n3015_);
  or g_891 (new_n2907_, not_new_n647__2, not_new_n602__403536070);
  not g_892 (not_new_n4679_, new_n4679_);
  or g_893 (new_n6057_, not_new_n5993_, not_new_n5900_);
  not g_894 (not_new_n1588__6, new_n1588_);
  not g_895 (not_pi038_3, pi038);
  or g_896 (new_n2345_, or_not_new_n2343__not_new_n2344_, not_new_n1569_);
  not g_897 (not_new_n1184_, new_n1184_);
  not g_898 (not_new_n7278_, new_n7278_);
  not g_899 (not_new_n3447_, new_n3447_);
  not g_900 (not_new_n6520__0, new_n6520_);
  not g_901 (not_new_n1020__2, new_n1020_);
  not g_902 (not_new_n5847_, new_n5847_);
  or g_903 (po293, or_or_or_not_new_n2964__not_new_n2967__not_new_n2966__not_new_n2968_, not_new_n2965_);
  not g_904 (not_new_n3242_, new_n3242_);
  or g_905 (new_n3697_, not_new_n639__9, not_po298_19773267430);
  not g_906 (not_new_n1616__57648010, new_n1616_);
  or g_907 (new_n1173_, not_new_n3876_, not_new_n3875_);
  or g_908 (new_n7019_, not_new_n7355_, not_new_n7356_);
  not g_909 (not_new_n3142_, new_n3142_);
  not g_910 (not_new_n6281_, new_n6281_);
  or g_911 (new_n761_, not_new_n3232_, not_new_n3233_);
  not g_912 (not_new_n3693_, new_n3693_);
  not g_913 (not_new_n4422_, new_n4422_);
  and g_914 (new_n7580_, new_n7837_, new_n7573_);
  and g_915 (new_n8676_, new_n8591_, new_n8749_);
  not g_916 (not_new_n3223_, new_n3223_);
  not g_917 (not_new_n593__0, new_n593_);
  not g_918 (not_new_n5727_, new_n5727_);
  and g_919 (new_n8204_, new_n8311_, new_n8312_);
  or g_920 (new_n8719_, not_new_n8641_, not_new_n1065__332329305696010);
  not g_921 (not_new_n8539_, new_n8539_);
  not g_922 (not_new_n9530__0, new_n9530_);
  and g_923 (and_new_n1735__new_n1736_, new_n1735_, new_n1736_);
  not g_924 (not_new_n9208_, new_n9208_);
  or g_925 (new_n2508_, or_not_new_n5426__not_new_n605_, not_new_n611__1);
  not g_926 (not_new_n3330_, new_n3330_);
  not g_927 (not_new_n775__16284135979104490, new_n775_);
  not g_928 (not_new_n8679_, new_n8679_);
  or g_929 (new_n9427_, or_not_new_n9704__not_new_n9705_, not_new_n9593_);
  or g_930 (new_n9681_, not_new_n9679_, not_new_n9483_);
  not g_931 (not_new_n648__6782230728490, new_n648_);
  not g_932 (not_new_n9971_, new_n9971_);
  and g_933 (new_n1426_, new_n2558_, new_n2559_);
  not g_934 (not_new_n584_, new_n584_);
  not g_935 (not_pi272, pi272);
  not g_936 (not_new_n632__47475615099430, new_n632_);
  not g_937 (not_new_n2884_, new_n2884_);
  or g_938 (new_n3743_, not_new_n973_, not_new_n2228_);
  or g_939 (or_not_new_n618__2326305139872070_not_new_n8496_, not_new_n8496_, not_new_n618__2326305139872070);
  or g_940 (new_n7220_, not_new_n7219_, not_new_n7150_);
  or g_941 (new_n9692_, not_new_n9675_, not_new_n9511__0);
  or g_942 (new_n2614_, not_new_n1003_, not_new_n607__8);
  or g_943 (new_n10259_, not_new_n10257_, not_new_n10073__0);
  not g_944 (not_new_n3293_, new_n3293_);
  not g_945 (not_new_n2302_, new_n2302_);
  not g_946 (not_new_n5836_, new_n5836_);
  not g_947 (not_new_n4508__0, new_n4508_);
  not g_948 (not_new_n4187_, new_n4187_);
  not g_949 (not_new_n4119__2, new_n4119_);
  or g_950 (new_n3266_, not_new_n622__8, not_new_n3184__9);
  not g_951 (new_n4156_, new_n4144_);
  not g_952 (not_new_n1810_, new_n1810_);
  not g_953 (not_new_n581__39098210485829880490, new_n581_);
  not g_954 (not_new_n2151_, new_n2151_);
  and g_955 (new_n6349_, new_n6232_, new_n6252_);
  not g_956 (not_new_n7710_, new_n7710_);
  not g_957 (not_new_n2350_, new_n2350_);
  or g_958 (new_n2349_, not_new_n3387__4, not_new_n3384__5);
  not g_959 (not_new_n1588__10, new_n1588_);
  not g_960 (not_new_n3372__6, new_n3372_);
  or g_961 (new_n3664_, not_new_n989__4, not_pi218);
  not g_962 (not_new_n3127_, new_n3127_);
  and g_963 (new_n8079_, new_n8345_, new_n8282_);
  or g_964 (new_n5341_, not_new_n5339_, not_new_n5340_);
  not g_965 (not_new_n645__2326305139872070, new_n645_);
  not g_966 (new_n8827_, new_n631_);
  or g_967 (new_n942_, not_new_n1774_, or_or_or_not_new_n1773__not_new_n1213__not_new_n1214__not_new_n1775_);
  not g_968 (not_new_n1057__5, new_n1057_);
  not g_969 (not_new_n589__5, new_n589_);
  not g_970 (not_new_n2720_, new_n2720_);
  not g_971 (not_new_n8157__0, new_n8157_);
  not g_972 (not_new_n1599_, new_n1599_);
  not g_973 (not_new_n1594__1, new_n1594_);
  not g_974 (not_new_n3355_, new_n3355_);
  not g_975 (not_new_n4759_, new_n4759_);
  not g_976 (not_new_n4140_, new_n4140_);
  or g_977 (or_or_or_not_new_n2749__not_new_n2752__not_new_n2751__not_new_n2753_, not_new_n2753_, or_or_not_new_n2749__not_new_n2752__not_new_n2751_);
  not g_978 (not_new_n4746_, new_n4746_);
  not g_979 (not_new_n5761__0, new_n5761_);
  not g_980 (not_pi251_1, pi251);
  not g_981 (not_new_n3493_, new_n3493_);
  not g_982 (not_new_n4763_, new_n4763_);
  not g_983 (not_new_n4250_, new_n4250_);
  and g_984 (and_new_n9402__new_n9804_, new_n9804_, new_n9402_);
  not g_985 (not_new_n611__2, new_n611_);
  not g_986 (not_new_n1588__24010, new_n1588_);
  not g_987 (not_pi143_3, pi143);
  not g_988 (not_new_n7914_, new_n7914_);
  not g_989 (not_new_n9961__0, new_n9961_);
  xnor g_990 (key_gate_0, not_new_n1633_, key_0);
  or g_991 (new_n3355_, not_pi045_0, not_new_n1534__403536070);
  or g_992 (new_n7525_, not_new_n728__1, not_new_n7427__0);
  or g_993 (new_n8127_, or_not_new_n8411__not_new_n8293_, not_new_n8277_);
  not g_994 (not_new_n9317_, new_n9317_);
  not g_995 (not_new_n3224_, new_n3224_);
  not g_996 (not_pi168_3, pi168);
  not g_997 (not_new_n1981_, new_n1981_);
  and g_998 (and_new_n1896__new_n1899_, new_n1896_, new_n1899_);
  or g_999 (new_n3031_, not_new_n622__4, not_new_n3372__8235430);
  and g_1000 (new_n5494_, new_n5586_, new_n5651_);
  and g_1001 (new_n1204_, new_n1701_, new_n1703_);
  not g_1002 (not_new_n1588__5585458640832840070, new_n1588_);
  or g_1003 (new_n3616_, not_pi174_0, not_new_n984__490);
  or g_1004 (new_n698_, not_new_n3066_, not_new_n1522_);
  or g_1005 (new_n2461_, not_new_n4781__0, not_new_n597__2824752490);
  not g_1006 (not_new_n6987_, new_n6987_);
  not g_1007 (not_pi023_0, pi023);
  or g_1008 (new_n987_, not_new_n3384__3, not_new_n591_);
  or g_1009 (or_or_not_new_n2246__not_new_n2243__not_new_n2244_, or_not_new_n2246__not_new_n2243_, not_new_n2244_);
  or g_1010 (new_n6552_, not_new_n6911_, not_new_n6910_);
  not g_1011 (not_new_n1027__1915812313805664144010, new_n1027_);
  or g_1012 (new_n6203_, not_new_n5787__0, not_new_n643__403536070);
  not g_1013 (not_new_n7491_, new_n7491_);
  or g_1014 (new_n2327_, not_new_n7591_, not_new_n1583__16284135979104490);
  not g_1015 (not_new_n2266_, new_n2266_);
  or g_1016 (new_n9954_, not_new_n578_, not_new_n579_);
  not g_1017 (not_new_n7012__0, new_n7012_);
  not g_1018 (not_new_n4458_, new_n4458_);
  not g_1019 (not_new_n8831_, new_n8831_);
  not g_1020 (not_new_n588__1, new_n588_);
  or g_1021 (new_n7652_, not_new_n7616_, not_new_n647__2824752490);
  not g_1022 (not_new_n3707_, new_n3707_);
  not g_1023 (not_new_n630_, new_n630_);
  or g_1024 (or_not_new_n1405__not_new_n616_, not_new_n1405_, not_new_n616_);
  not g_1025 (not_new_n1591__6, new_n1591_);
  not g_1026 (not_new_n984__7, new_n984_);
  not g_1027 (not_new_n624__6, new_n624_);
  not g_1028 (not_new_n4173_, new_n4173_);
  not g_1029 (new_n4833_, new_n4742_);
  not g_1030 (not_new_n3996__0, new_n3996_);
  not g_1031 (not_new_n1536__19773267430, new_n1536_);
  not g_1032 (not_new_n643__10, new_n643_);
  or g_1033 (new_n6073_, not_new_n5848_, not_new_n5878__2);
  or g_1034 (new_n8340_, not_new_n8339_, not_new_n8338_);
  not g_1035 (not_new_n5465_, new_n5465_);
  not g_1036 (not_pi111, pi111);
  not g_1037 (not_new_n1611__968890104070, new_n1611_);
  or g_1038 (new_n2909_, not_new_n2906_, or_not_new_n2908__not_new_n2907_);
  buf g_1039 (po004, pi197);
  not g_1040 (not_new_n5942__0, new_n5942_);
  not g_1041 (not_new_n2509__4, new_n2509_);
  not g_1042 (not_new_n6072_, new_n6072_);
  not g_1043 (new_n8893_, new_n1596_);
  not g_1044 (not_po296_403536070, po296);
  not g_1045 (not_new_n9340_, new_n9340_);
  not g_1046 (not_new_n3139_, new_n3139_);
  not g_1047 (not_new_n639__3, new_n639_);
  or g_1048 (new_n4773_, not_new_n4775__0, not_new_n4837__0);
  not g_1049 (new_n7104_, new_n772_);
  or g_1050 (or_or_or_not_new_n2865__not_new_n2868__not_new_n2867__not_new_n2869_, not_new_n2869_, or_or_not_new_n2865__not_new_n2868__not_new_n2867_);
  not g_1051 (not_new_n681_, new_n681_);
  not g_1052 (not_new_n632__797922662976120010, new_n632_);
  not g_1053 (not_new_n6207_, new_n6207_);
  not g_1054 (not_new_n3716_, new_n3716_);
  not g_1055 (not_new_n10097_, new_n10097_);
  or g_1056 (new_n8552_, not_new_n8266__5, not_new_n8234_);
  not g_1057 (not_new_n5759__0, new_n5759_);
  or g_1058 (new_n8233_, not_new_n8543_, not_new_n8544_);
  not g_1059 (not_new_n9387_, new_n9387_);
  not g_1060 (new_n8841_, new_n648_);
  not g_1061 (not_new_n8294__0, new_n8294_);
  or g_1062 (po072, key_gate_91, not_new_n1199_);
  or g_1063 (new_n3382_, not_new_n1534__2326305139872070, not_pi052_0);
  not g_1064 (not_new_n4404_, new_n4404_);
  not g_1065 (not_new_n613__6, new_n613_);
  not g_1066 (not_new_n1601__332329305696010, new_n1601_);
  or g_1067 (new_n3022_, not_new_n3372__24010, not_new_n618__3);
  not g_1068 (not_new_n9389_, new_n9389_);
  not g_1069 (not_new_n3751_, new_n3751_);
  or g_1070 (new_n4665_, not_new_n4493_, not_new_n4494__0);
  not g_1071 (not_new_n8103_, new_n8103_);
  or g_1072 (new_n5014_, not_new_n5369_, not_new_n5368_);
  not g_1073 (not_new_n5190_, new_n5190_);
  not g_1074 (not_pi222, pi222);
  not g_1075 (not_new_n1169_, new_n1169_);
  or g_1076 (new_n9218_, not_new_n9216_, not_new_n9217_);
  or g_1077 (new_n3587_, not_new_n1612__113988951853731430, not_new_n2345__0);
  not g_1078 (not_new_n6291_, new_n6291_);
  or g_1079 (new_n1878_, not_new_n635_, not_new_n593__4);
  not g_1080 (not_new_n7354__0, new_n7354_);
  not g_1081 (not_new_n3372__8, new_n3372_);
  and g_1082 (new_n7573_, new_n7832_, new_n7769_);
  not g_1083 (not_new_n1065__5585458640832840070, new_n1065_);
  not g_1084 (not_pi177_1, pi177);
  not g_1085 (not_new_n7520_, new_n7520_);
  not g_1086 (not_new_n1580__797922662976120010, new_n1580_);
  not g_1087 (not_new_n3233_, new_n3233_);
  not g_1088 (not_new_n9704_, new_n9704_);
  or g_1089 (new_n4712_, not_new_n4434__0, not_pi171_3);
  or g_1090 (new_n5123_, not_new_n632__3430, not_new_n1037__8);
  not g_1091 (new_n8116_, new_n642_);
  not g_1092 (not_new_n4908_, new_n4908_);
  or g_1093 (new_n7731_, not_new_n8064_, not_new_n8065_);
  and g_1094 (new_n7085_, new_n7161_, new_n7256_);
  not g_1095 (not_new_n5938__0, new_n5938_);
  not g_1096 (not_po298_168070, po298);
  or g_1097 (new_n8182_, not_new_n8524_, not_new_n8523_);
  or g_1098 (new_n2645_, not_new_n5480_, not_new_n605__3430);
  or g_1099 (new_n4748_, not_new_n4877_, not_new_n4876_);
  not g_1100 (not_new_n7637_, new_n7637_);
  not g_1101 (not_new_n7739__0, new_n7739_);
  not g_1102 (not_new_n628__1, new_n628_);
  or g_1103 (new_n6634_, not_new_n1031__168070, not_new_n6548_);
  not g_1104 (not_new_n6539__0, new_n6539_);
  or g_1105 (new_n4663_, not_pi178_3, not_new_n4448__0);
  not g_1106 (not_new_n7889_, new_n7889_);
  not g_1107 (not_new_n4712_, new_n4712_);
  not g_1108 (new_n6723_, new_n6637_);
  or g_1109 (new_n3123_, not_new_n928__490, not_new_n1599__3);
  or g_1110 (new_n4393_, not_new_n4314_, not_new_n4390_);
  not g_1111 (not_new_n8683_, new_n8683_);
  not g_1112 (not_new_n9061_, new_n9061_);
  not g_1113 (not_new_n1523_, new_n1523_);
  or g_1114 (new_n10028_, not_new_n10102_, not_new_n10103_);
  not g_1115 (not_new_n8120__0, new_n8120_);
  not g_1116 (not_new_n1027__0, new_n1027_);
  or g_1117 (new_n2730_, not_new_n7065_, not_new_n595_);
  not g_1118 (not_new_n8888_, new_n8888_);
  not g_1119 (not_new_n7341_, new_n7341_);
  not g_1120 (not_new_n5255_, new_n5255_);
  not g_1121 (not_new_n9364_, new_n9364_);
  not g_1122 (not_new_n5675_, new_n5675_);
  not g_1123 (not_pi033_2, pi033);
  not g_1124 (not_new_n7891_, new_n7891_);
  not g_1125 (not_new_n10304_, new_n10304_);
  not g_1126 (not_new_n4731_, new_n4731_);
  or g_1127 (new_n3423_, not_new_n1594__3, not_new_n1007__1);
  not g_1128 (not_pi212, pi212);
  xnor g_1129 (key_gate_37, new_n3977_, key_37);
  or g_1130 (new_n4550_, new_n1018_, pi172);
  or g_1131 (new_n4624_, not_new_n4421__0, not_new_n1007__4);
  not g_1132 (not_new_n9869_, new_n9869_);
  not g_1133 (not_pi045_0, pi045);
  or g_1134 (new_n8314_, not_new_n8124_, not_new_n1051__8235430);
  not g_1135 (not_new_n8542_, new_n8542_);
  not g_1136 (not_new_n10238_, new_n10238_);
  not g_1137 (not_new_n1584__9, new_n1584_);
  not g_1138 (not_new_n7463_, new_n7463_);
  not g_1139 (not_new_n9522_, new_n9522_);
  not g_1140 (new_n6537_, new_n621_);
  and g_1141 (new_n1314_, new_n2196_, new_n2195_);
  not g_1142 (not_new_n4560_, new_n4560_);
  not g_1143 (not_new_n994__9, new_n994_);
  or g_1144 (new_n8715_, not_new_n1606__6, not_new_n8653_);
  not g_1145 (not_new_n4266_, new_n4266_);
  not g_1146 (not_new_n4876_, new_n4876_);
  not g_1147 (not_new_n605__7, new_n605_);
  not g_1148 (not_new_n9156_, new_n9156_);
  not g_1149 (not_new_n1613__47475615099430, new_n1613_);
  not g_1150 (new_n10177_, new_n10023_);
  not g_1151 (new_n4159_, new_n4083_);
  not g_1152 (not_new_n6656_, new_n6656_);
  not g_1153 (not_new_n4149_, new_n4149_);
  or g_1154 (or_not_new_n2785__not_new_n2788_, not_new_n2785_, not_new_n2788_);
  or g_1155 (new_n5697_, not_new_n5558_, not_new_n5695_);
  not g_1156 (not_new_n7054_, new_n7054_);
  not g_1157 (not_new_n5763__1, new_n5763_);
  or g_1158 (new_n9567_, not_new_n9749_, or_or_not_new_n9361__not_new_n9358__0_not_new_n9750_);
  not g_1159 (not_new_n7848_, new_n7848_);
  or g_1160 (new_n6391_, not_new_n6293_, not_new_n637__8235430);
  not g_1161 (new_n1624_, new_n997_);
  not g_1162 (new_n4017_, new_n3943_);
  or g_1163 (new_n3164_, not_new_n636__5, not_new_n3315__332329305696010);
  not g_1164 (not_new_n7324_, new_n7324_);
  or g_1165 (new_n2478_, not_new_n4122__0, not_new_n600__6782230728490);
  and g_1166 (new_n7706_, new_n7830_, new_n7582_);
  not g_1167 (not_new_n1845_, new_n1845_);
  and g_1168 (and_new_n2687__new_n2688_, new_n2688_, new_n2687_);
  not g_1169 (not_new_n6889_, new_n6889_);
  not g_1170 (not_new_n4830_, new_n4830_);
  or g_1171 (new_n4038_, not_new_n4031_, not_pi052_3);
  or g_1172 (new_n8551_, not_new_n8550_, not_new_n8456_);
  not g_1173 (not_new_n7791__0, new_n7791_);
  or g_1174 (new_n1712_, not_pi059, not_new_n1631__47475615099430);
  and g_1175 (and_new_n8731__new_n8730_, new_n8730_, new_n8731_);
  not g_1176 (not_new_n1292_, new_n1292_);
  not g_1177 (not_new_n596__138412872010, key_gate_88);
  or g_1178 (or_not_new_n1571__not_new_n2504_, not_new_n2504_, not_new_n1571_);
  not g_1179 (not_new_n3885_, new_n3885_);
  not g_1180 (not_new_n591__4, new_n591_);
  not g_1181 (not_new_n605__57648010, new_n605_);
  not g_1182 (not_pi039_1, pi039);
  or g_1183 (new_n1777_, not_new_n9954_, not_new_n594_);
  not g_1184 (not_new_n5867_, new_n5867_);
  not g_1185 (not_new_n627__3, new_n627_);
  not g_1186 (not_new_n10236_, new_n10236_);
  and g_1187 (new_n1480_, new_n2815_, new_n2814_);
  not g_1188 (not_new_n3673_, new_n3673_);
  not g_1189 (not_new_n7061_, new_n7061_);
  or g_1190 (or_or_not_new_n1844__not_new_n1845__not_new_n1847_, or_not_new_n1844__not_new_n1845_, not_new_n1847_);
  or g_1191 (new_n9841_, not_new_n1057__6782230728490, not_new_n9391_);
  or g_1192 (new_n2025_, not_new_n6557_, not_new_n1580__3430);
  not g_1193 (not_new_n6073_, new_n6073_);
  not g_1194 (not_po296_1176490, po296);
  or g_1195 (new_n6762_, not_new_n6519__0, not_new_n638__138412872010);
  or g_1196 (new_n2757_, not_new_n2754_, or_not_new_n2756__not_new_n2755_);
  or g_1197 (new_n7719_, not_new_n8003_, not_new_n8002_);
  and g_1198 (new_n7151_, new_n7539_, new_n7540_);
  not g_1199 (not_new_n3871_, new_n3871_);
  not g_1200 (not_new_n3987__0, key_gate_12);
  not g_1201 (not_new_n3719_, new_n3719_);
  not g_1202 (not_new_n590_, new_n590_);
  or g_1203 (new_n10327_, not_new_n10325_, not_new_n10165__0);
  not g_1204 (not_new_n605__8235430, new_n605_);
  not g_1205 (not_new_n1596__968890104070, new_n1596_);
  or g_1206 (new_n3352_, not_new_n3918__0, not_pi064_8235430);
  and g_1207 (and_new_n9356__new_n9738_, new_n9738_, new_n9356_);
  not g_1208 (not_new_n4903_, new_n4903_);
  or g_1209 (new_n5860_, not_new_n6147_, not_new_n6148_);
  and g_1210 (new_n7700_, and_new_n7597__new_n7953_, new_n7952_);
  not g_1211 (new_n7621_, new_n1598_);
  not g_1212 (not_new_n1035__2, new_n1035_);
  not g_1213 (not_new_n8844__0, new_n8844_);
  not g_1214 (not_new_n6974__2824752490, new_n6974_);
  or g_1215 (new_n6100_, not_new_n1047__490, not_new_n5739__0);
  not g_1216 (not_new_n1164_, new_n1164_);
  not g_1217 (not_new_n8785_, new_n8785_);
  not g_1218 (not_new_n582__0, new_n582_);
  not g_1219 (not_new_n1158__0, new_n1158_);
  not g_1220 (not_new_n645__3, new_n645_);
  not g_1221 (new_n6068_, new_n5814_);
  not g_1222 (not_new_n7628_, new_n7628_);
  and g_1223 (new_n8675_, new_n8747_, new_n8748_);
  not g_1224 (new_n9929_, new_n1061_);
  and g_1225 (new_n7140_, new_n7485_, new_n7486_);
  and g_1226 (new_n8677_, new_n8724_, new_n8726_);
  not g_1227 (not_new_n7431_, new_n7431_);
  not g_1228 (not_pi178, pi178);
  or g_1229 (new_n9494_, not_new_n9623_, not_new_n9622_);
  or g_1230 (new_n7036_, not_new_n7432_, not_new_n7431_);
  not g_1231 (not_new_n1059__16284135979104490, new_n1059_);
  not g_1232 (not_new_n6373__8, new_n6373_);
  or g_1233 (new_n3450_, not_new_n1537__8, not_pi106_0);
  not g_1234 (not_new_n7426_, new_n7426_);
  not g_1235 (not_new_n1602__2326305139872070, new_n1602_);
  not g_1236 (not_new_n5821_, new_n5821_);
  not g_1237 (not_new_n607__7, new_n607_);
  or g_1238 (new_n6672_, not_new_n6445_, not_new_n6671_);
  not g_1239 (not_new_n7985_, new_n7985_);
  or g_1240 (new_n5678_, not_new_n1014__6, not_new_n5676_);
  or g_1241 (new_n6217_, not_new_n627__8235430, not_new_n5793__0);
  or g_1242 (new_n2454_, not_new_n9870__0, not_new_n599__403536070);
  not g_1243 (not_new_n3184__0, new_n3184_);
  not g_1244 (new_n5800_, new_n643_);
  not g_1245 (not_pi179_0, pi179);
  not g_1246 (not_new_n1812_, new_n1812_);
  not g_1247 (not_pi162_2, pi162);
  or g_1248 (new_n4333_, or_not_new_n4291__not_new_n4326_, not_new_n4292_);
  or g_1249 (new_n9801_, not_new_n1603__332329305696010, not_new_n9408__0);
  not g_1250 (not_new_n9372_, new_n9372_);
  or g_1251 (new_n3720_, not_new_n3718_, not_new_n3719_);
  not g_1252 (not_new_n9426_, new_n9426_);
  or g_1253 (new_n6947_, not_new_n6641_, not_new_n6608_);
  or g_1254 (new_n9539_, new_n1049_, new_n648_);
  not g_1255 (not_new_n610__1, new_n610_);
  not g_1256 (not_new_n1555_, new_n1555_);
  or g_1257 (new_n10286_, not_new_n10015__0, not_new_n10014_);
  not g_1258 (not_new_n2444_, new_n2444_);
  not g_1259 (not_new_n1057__968890104070, new_n1057_);
  not g_1260 (not_new_n7579_, new_n7579_);
  not g_1261 (not_new_n8118__0, new_n8118_);
  not g_1262 (not_new_n7123_, new_n7123_);
  not g_1263 (not_new_n5170_, new_n5170_);
  not g_1264 (not_new_n1061__8, new_n1061_);
  or g_1265 (new_n732_, not_new_n3292_, not_new_n3291_);
  not g_1266 (not_new_n748_, new_n748_);
  or g_1267 (new_n1172_, not_new_n3873_, not_new_n3874_);
  not g_1268 (not_new_n596__797922662976120010, key_gate_88);
  not g_1269 (not_new_n7389_, new_n7389_);
  not g_1270 (not_new_n1604__2326305139872070, new_n1604_);
  not g_1271 (not_new_n9992_, new_n9992_);
  not g_1272 (not_new_n6227_, new_n6227_);
  not g_1273 (not_new_n637__16284135979104490, new_n637_);
  or g_1274 (or_not_new_n1567__not_new_n2494_, not_new_n2494_, not_new_n1567_);
  not g_1275 (not_new_n629__19773267430, new_n629_);
  or g_1276 (new_n6392_, not_new_n643__2824752490, not_new_n6294_);
  not g_1277 (not_pi053_0, pi053);
  or g_1278 (or_or_or_not_new_n1055__168070_not_new_n6325__not_new_n6373__1_not_new_n6317_, not_new_n6317_, or_or_not_new_n1055__168070_not_new_n6325__not_new_n6373__1);
  or g_1279 (new_n7997_, not_new_n7996_, not_new_n7995_);
  or g_1280 (new_n6727_, not_new_n1069__24010, not_new_n6515_);
  not g_1281 (new_n4074_, pi248);
  and g_1282 (new_n1369_, and_new_n2409__new_n2408_, new_n2407_);
  and g_1283 (new_n1494_, new_n3013_, new_n3012_);
  not g_1284 (not_new_n7279_, new_n7279_);
  not g_1285 (not_new_n9868_, new_n9868_);
  or g_1286 (new_n6534_, not_new_n6520_, not_new_n643__19773267430);
  not g_1287 (not_new_n6960_, new_n6960_);
  not g_1288 (not_new_n3122_, new_n3122_);
  not g_1289 (not_pi257_0, pi257);
  or g_1290 (new_n7238_, not_new_n7038_, not_new_n724_);
  or g_1291 (new_n9752_, not_new_n9486_, not_new_n1607__57648010);
  not g_1292 (not_new_n625__8235430, new_n625_);
  not g_1293 (not_new_n6461_, new_n6461_);
  not g_1294 (not_new_n8130__0, new_n8130_);
  or g_1295 (new_n9429_, not_new_n9806_, not_new_n9805_);
  not g_1296 (not_pi167_0, pi167);
  or g_1297 (new_n8466_, not_new_n648__2326305139872070, not_new_n8110__1);
  not g_1298 (not_new_n1887_, new_n1887_);
  not g_1299 (not_new_n1616__2, new_n1616_);
  not g_1300 (not_new_n640__4, new_n640_);
  not g_1301 (not_new_n5022_, new_n5022_);
  not g_1302 (not_new_n5360_, new_n5360_);
  or g_1303 (new_n10342_, not_new_n9917__0, not_new_n638__1577753820348458066150427430);
  not g_1304 (not_new_n2321_, new_n2321_);
  not g_1305 (not_new_n7430__0, new_n7430_);
  not g_1306 (not_new_n589__113988951853731430, new_n589_);
  or g_1307 (new_n4060_, not_new_n4017__2, not_new_n3986__0);
  not g_1308 (not_new_n597__9, new_n597_);
  not g_1309 (new_n5898_, new_n1035_);
  or g_1310 (new_n4360_, not_new_n4303_, not_new_n4357_);
  or g_1311 (new_n2004_, not_new_n9448_, not_new_n1584__70);
  not g_1312 (not_new_n618__113988951853731430, new_n618_);
  not g_1313 (not_new_n7714_, new_n7714_);
  or g_1314 (new_n5648_, not_pi148_1, not_new_n5507_);
  not g_1315 (not_new_n6232__1, new_n6232_);
  xnor g_1316 (key_gate_124, key_124, not_new_n3987_);
  not g_1317 (not_new_n1053__24010, new_n1053_);
  or g_1318 (new_n3611_, not_new_n953_, not_new_n1611__9);
  not g_1319 (not_new_n1065__4, new_n1065_);
  not g_1320 (not_new_n730__1, new_n730_);
  not g_1321 (new_n4275_, new_n655_);
  or g_1322 (new_n1916_, not_new_n648_, not_new_n593__6);
  or g_1323 (new_n8358_, not_new_n1069__57648010, not_new_n8146_);
  or g_1324 (new_n3455_, not_new_n1537__9, not_pi107_0);
  not g_1325 (not_new_n7984_, new_n7984_);
  not g_1326 (not_new_n5349_, new_n5349_);
  not g_1327 (not_new_n1604__2, new_n1604_);
  not g_1328 (not_new_n3341_, new_n3341_);
  not g_1329 (not_new_n9327_, new_n9327_);
  and g_1330 (new_n1228_, new_n3404_, new_n590_);
  not g_1331 (not_new_n2574_, new_n2574_);
  not g_1332 (not_new_n1014__2, new_n1014_);
  not g_1333 (not_new_n1028__8, new_n1028_);
  not g_1334 (not_new_n1061__490, new_n1061_);
  not g_1335 (not_new_n1589__6, new_n1589_);
  not g_1336 (not_new_n9881_, new_n9881_);
  and g_1337 (new_n5053_, new_n5245_, new_n4902_);
  or g_1338 (po149, not_new_n3524_, not_new_n3525_);
  not g_1339 (not_pi051_2, pi051);
  not g_1340 (not_new_n634__2326305139872070, new_n634_);
  not g_1341 (not_new_n1597__57648010, new_n1597_);
  not g_1342 (not_new_n1588__168070, new_n1588_);
  or g_1343 (po084, not_new_n1211_, key_gate_74);
  not g_1344 (not_new_n8950_, new_n8950_);
  not g_1345 (not_new_n635__2326305139872070, new_n635_);
  not g_1346 (not_new_n1049__8235430, new_n1049_);
  or g_1347 (new_n6885_, not_new_n6500__0, not_new_n622__403536070);
  or g_1348 (new_n9695_, not_new_n9326__1, or_not_new_n9327__0_not_new_n9524__0);
  not g_1349 (not_new_n4567_, new_n4567_);
  not g_1350 (not_new_n5755__0, new_n5755_);
  not g_1351 (not_new_n629__3, new_n629_);
  not g_1352 (not_new_n5758_, new_n5758_);
  or g_1353 (new_n7916_, not_new_n7848_, not_new_n7847_);
  not g_1354 (not_new_n7846_, new_n7846_);
  or g_1355 (new_n1986_, not_new_n8094_, not_new_n1581__10);
  not g_1356 (not_new_n3088_, new_n3088_);
  not g_1357 (not_new_n644__9, new_n644_);
  or g_1358 (new_n9839_, not_new_n9396_, not_new_n1059__2326305139872070);
  not g_1359 (not_new_n8935_, new_n8935_);
  not g_1360 (not_new_n3522_, new_n3522_);
  or g_1361 (new_n2111_, not_new_n587__57648010, not_pi148);
  or g_1362 (new_n2863_, not_new_n994__1176490, not_new_n4131__1);
  not g_1363 (not_new_n5549_, new_n5549_);
  not g_1364 (not_new_n1728__2, new_n1728_);
  and g_1365 (new_n8243_, new_n8459_, new_n8460_);
  not g_1366 (not_new_n8533_, new_n8533_);
  not g_1367 (not_new_n626__16284135979104490, new_n626_);
  not g_1368 (not_new_n610__9, new_n610_);
  and g_1369 (new_n8220_, new_n8379_, new_n8378_);
  or g_1370 (new_n2893_, not_new_n612__4, not_new_n4126__2);
  not g_1371 (not_pi179_1, pi179);
  not g_1372 (not_new_n8616_, new_n8616_);
  not g_1373 (not_new_n3773_, new_n3773_);
  or g_1374 (new_n6666_, not_new_n6665_, not_new_n6486_);
  not g_1375 (not_new_n6823_, new_n6823_);
  not g_1376 (new_n4794_, new_n1065_);
  not g_1377 (not_new_n6998__0, new_n6998_);
  not g_1378 (not_new_n616__0, new_n616_);
  not g_1379 (not_new_n6974_, new_n6974_);
  or g_1380 (new_n3550_, not_pi141_0, not_new_n1538__70);
  and g_1381 (and_new_n2652__new_n2651_, new_n2651_, new_n2652_);
  or g_1382 (new_n3734_, not_new_n626__10, not_new_n1053__7);
  not g_1383 (new_n9069_, new_n8884_);
  or g_1384 (new_n4667_, not_new_n4445_, not_new_n1013__3);
  not g_1385 (not_new_n3419_, new_n3419_);
  not g_1386 (not_new_n9922_, new_n9922_);
  not g_1387 (not_new_n621__168070, new_n621_);
  or g_1388 (new_n7769_, not_new_n1063__168070, not_new_n7656_);
  not g_1389 (not_new_n6334_, new_n6334_);
  not g_1390 (not_new_n3588_, new_n3588_);
  and g_1391 (new_n1235_, and_new_n1234__new_n1818_, new_n1817_);
  not g_1392 (not_new_n5201_, new_n5201_);
  not g_1393 (not_new_n3156_, new_n3156_);
  or g_1394 (new_n3006_, not_new_n1027__8, not_new_n1154_);
  not g_1395 (not_new_n5476__0, new_n5476_);
  not g_1396 (not_new_n7070_, new_n7070_);
  not g_1397 (not_new_n4968_, new_n4968_);
  not g_1398 (not_new_n3015_, new_n3015_);
  or g_1399 (new_n2159_, not_new_n1591__403536070, not_new_n8815_);
  not g_1400 (not_new_n8359_, new_n8359_);
  not g_1401 (not_new_n9180_, new_n9180_);
  not g_1402 (not_new_n633__1, new_n633_);
  and g_1403 (and_and_new_n1746__new_n1747__new_n1749_, and_new_n1746__new_n1747_, new_n1749_);
  not g_1404 (not_new_n6443__3, new_n6443_);
  not g_1405 (not_new_n1039__797922662976120010, new_n1039_);
  or g_1406 (new_n6811_, not_new_n6683__0, not_new_n6613_);
  or g_1407 (or_or_not_new_n1565__not_new_n2484__not_new_n1399_, or_not_new_n1565__not_new_n2484_, not_new_n1399_);
  or g_1408 (new_n3833_, not_new_n6443__2, not_new_n635__70);
  not g_1409 (not_new_n8968_, new_n8968_);
  not g_1410 (not_new_n8988_, new_n8988_);
  not g_1411 (not_new_n589__21838143759917965991093122527538323430, new_n589_);
  not g_1412 (not_new_n10106_, new_n10106_);
  or g_1413 (new_n10217_, not_new_n10106_, not_new_n10103__0);
  not g_1414 (new_n8877_, new_n646_);
  not g_1415 (not_new_n1180_, new_n1180_);
  not g_1416 (not_new_n6975__0, new_n6975_);
  not g_1417 (not_new_n3431_, new_n3431_);
  and g_1418 (new_n1502_, new_n3028_, new_n1503_);
  not g_1419 (not_new_n591__24010, new_n591_);
  or g_1420 (new_n6784_, not_new_n6572_, not_new_n6617__1);
  not g_1421 (not_new_n1594__3, new_n1594_);
  not g_1422 (not_new_n2033_, new_n2033_);
  and g_1423 (and_new_n1246__new_n1875_, new_n1875_, new_n1246_);
  not g_1424 (not_new_n3343_, new_n3343_);
  not g_1425 (not_new_n586__2, new_n586_);
  not g_1426 (not_new_n1041_, new_n1041_);
  not g_1427 (not_new_n9822_, new_n9822_);
  not g_1428 (not_new_n8244_, new_n8244_);
  not g_1429 (not_new_n8741_, new_n8741_);
  not g_1430 (not_new_n3513_, new_n3513_);
  not g_1431 (not_new_n8956_, new_n8956_);
  not g_1432 (not_new_n4421_, new_n4421_);
  or g_1433 (new_n8830_, not_new_n642__332329305696010, not_new_n1035__24010);
  not g_1434 (new_n8842_, new_n647_);
  not g_1435 (not_new_n5158_, new_n5158_);
  or g_1436 (new_n2612_, not_new_n2509__9, not_pi203);
  not g_1437 (new_n7795_, new_n7618_);
  not g_1438 (not_new_n9330_, new_n9330_);
  not g_1439 (not_new_n5187_, new_n5187_);
  not g_1440 (not_new_n1015__6, new_n1015_);
  not g_1441 (not_new_n3714_, new_n3714_);
  not g_1442 (not_new_n604__57648010, new_n604_);
  not g_1443 (not_new_n7753__2, new_n7753_);
  not g_1444 (not_new_n1489_, new_n1489_);
  not g_1445 (not_new_n683_, new_n683_);
  not g_1446 (not_new_n4833__1, new_n4833_);
  not g_1447 (not_pi041_3, pi041);
  not g_1448 (not_new_n4765_, new_n4765_);
  not g_1449 (not_new_n3842_, new_n3842_);
  not g_1450 (not_new_n6624_, new_n6624_);
  not g_1451 (not_new_n8849__0, new_n8849_);
  not g_1452 (not_new_n985_, new_n985_);
  not g_1453 (not_pi033_3, pi033);
  not g_1454 (not_new_n1609__0, new_n1609_);
  not g_1455 (not_new_n1047__0, new_n1047_);
  not g_1456 (not_new_n9376_, new_n9376_);
  or g_1457 (new_n9537_, not_new_n9373_, not_new_n9328_);
  or g_1458 (new_n8713_, not_new_n1155__0, not_new_n8654_);
  or g_1459 (new_n1846_, not_new_n588__4, not_pi102);
  not g_1460 (not_new_n6138__0, new_n6138_);
  not g_1461 (not_new_n8358_, new_n8358_);
  or g_1462 (new_n2549_, not_pi246, not_po296_13410686196639649008070);
  not g_1463 (not_new_n7084_, new_n7084_);
  and g_1464 (and_new_n9365__new_n9731_, new_n9365_, new_n9731_);
  not g_1465 (new_n2726_, new_n996_);
  not g_1466 (not_new_n713_, new_n713_);
  not g_1467 (not_new_n4958_, new_n4958_);
  not g_1468 (not_new_n1152__0, new_n1152_);
  not g_1469 (not_new_n1039__4, new_n1039_);
  not g_1470 (not_new_n645__16284135979104490, new_n645_);
  not g_1471 (new_n6482_, new_n628_);
  not g_1472 (new_n6023_, new_n5813_);
  not g_1473 (not_new_n3372__1176490, new_n3372_);
  or g_1474 (new_n9825_, not_new_n9386_, not_new_n1063__6782230728490);
  not g_1475 (not_new_n6373__5, new_n6373_);
  not g_1476 (not_new_n1027__8, new_n1027_);
  not g_1477 (not_new_n9891_, new_n9891_);
  or g_1478 (new_n3045_, not_new_n1604__2, not_new_n581__57648010);
  and g_1479 (new_n1195_, new_n1676_, new_n1674_);
  not g_1480 (not_new_n3185__57648010, new_n3185_);
  not g_1481 (not_new_n6985__1, new_n6985_);
  not g_1482 (not_new_n1175__1, new_n1175_);
  not g_1483 (not_pi163_1, pi163);
  not g_1484 (not_new_n3315__168070, new_n3315_);
  not g_1485 (not_new_n1660_, key_gate_42);
  or g_1486 (new_n9443_, not_new_n9811_, not_new_n9810_);
  or g_1487 (new_n3577_, not_new_n2261__0, not_new_n1612__6782230728490);
  not g_1488 (not_new_n5421_, new_n5421_);
  or g_1489 (new_n6037_, not_new_n1055__3430, not_new_n5791__1);
  or g_1490 (new_n7783_, not_new_n7606__0, not_new_n7605_);
  not g_1491 (not_pi260, pi260);
  and g_1492 (and_and_new_n6326__new_n6241__new_n6227_, and_new_n6326__new_n6241_, new_n6227_);
  not g_1493 (not_pi246_1, pi246);
  not g_1494 (not_new_n1598__0, new_n1598_);
  not g_1495 (not_new_n10256_, new_n10256_);
  or g_1496 (new_n3176_, not_new_n641__3, not_new_n3315__797922662976120010);
  not g_1497 (not_new_n7260__0, new_n7260_);
  or g_1498 (new_n9641_, not_new_n9637_, not_new_n9512_);
  and g_1499 (new_n1322_, new_n2234_, new_n2233_);
  or g_1500 (new_n7756_, not_new_n7659_, not_new_n7839_);
  not g_1501 (not_new_n5923_, new_n5923_);
  not g_1502 (not_new_n630__0, new_n630_);
  not g_1503 (not_new_n1071__403536070, new_n1071_);
  or g_1504 (new_n5241_, new_n1057_, new_n636_);
  not g_1505 (not_new_n4539_, new_n4539_);
  not g_1506 (not_new_n8155__0, new_n8155_);
  or g_1507 (new_n8750_, not_new_n8593__0, or_or_not_new_n8609__not_new_n8595__0_not_new_n1168__0);
  or g_1508 (new_n5583_, not_new_n5493_, not_new_n5581_);
  and g_1509 (new_n9504_, new_n9832_, new_n9831_);
  not g_1510 (not_new_n9288_, new_n9288_);
  not g_1511 (not_pi042_1, pi042);
  not g_1512 (not_new_n9409_, new_n9409_);
  not g_1513 (not_new_n1449_, new_n1449_);
  not g_1514 (not_new_n9762_, new_n9762_);
  not g_1515 (not_new_n1601__4, new_n1601_);
  not g_1516 (not_new_n601__57648010, new_n601_);
  not g_1517 (new_n8601_, new_n1051_);
  or g_1518 (new_n2268_, not_new_n1583__47475615099430, not_new_n7689_);
  or g_1519 (new_n6169_, not_new_n6060_, not_new_n5895_);
  or g_1520 (new_n2639_, not_po296_541169560379521116689596608490, not_pi248);
  not g_1521 (not_new_n5429_, new_n5429_);
  not g_1522 (not_new_n1337_, new_n1337_);
  not g_1523 (not_new_n3524_, new_n3524_);
  not g_1524 (not_new_n1611__403536070, new_n1611_);
  or g_1525 (new_n8453_, not_new_n8210_, not_new_n8452_);
  not g_1526 (not_new_n647__968890104070, new_n647_);
  not g_1527 (not_new_n7245_, new_n7245_);
  not g_1528 (not_new_n627__2326305139872070, new_n627_);
  not g_1529 (not_new_n7087_, new_n7087_);
  or g_1530 (new_n7226_, not_new_n6993_, not_new_n6994__0);
  not g_1531 (not_new_n633__138412872010, new_n633_);
  not g_1532 (not_new_n5488__0, new_n5488_);
  not g_1533 (not_new_n1613__797922662976120010, new_n1613_);
  or g_1534 (new_n3633_, not_new_n966_, not_new_n1611__2824752490);
  or g_1535 (new_n3907_, not_new_n1061__7, not_new_n9930_);
  not g_1536 (not_new_n7045__1, new_n7045_);
  or g_1537 (new_n2336_, not_new_n591__113988951853731430, not_new_n4761_);
  not g_1538 (not_new_n646__113988951853731430, new_n646_);
  or g_1539 (new_n1650_, not_pi026, not_po296_5);
  not g_1540 (not_new_n1613__2, new_n1613_);
  not g_1541 (not_new_n1188_, new_n1188_);
  not g_1542 (not_pi130_0, pi130);
  not g_1543 (not_new_n7309_, new_n7309_);
  not g_1544 (not_new_n8103__0, new_n8103_);
  not g_1545 (not_new_n7017__0, new_n7017_);
  or g_1546 (new_n6873_, not_new_n1597__168070, not_new_n6539__1);
  not g_1547 (new_n8872_, new_n1071_);
  or g_1548 (new_n5247_, new_n1057_, new_n636_);
  not g_1549 (not_po296_70, po296);
  or g_1550 (new_n2774_, not_new_n994__6, not_new_n4136__1);
  not g_1551 (not_new_n1059__2326305139872070, new_n1059_);
  not g_1552 (not_new_n3769_, new_n3769_);
  not g_1553 (not_new_n1588__968890104070, new_n1588_);
  not g_1554 (not_new_n994__2824752490, new_n994_);
  not g_1555 (not_new_n10335_, new_n10335_);
  not g_1556 (not_new_n1067__403536070, new_n1067_);
  or g_1557 (new_n8268_, not_new_n8166_, not_new_n8352_);
  not g_1558 (not_po298_6782230728490, po298);
  not g_1559 (not_new_n1602__6782230728490, new_n1602_);
  not g_1560 (not_new_n981_, new_n981_);
  not g_1561 (not_new_n9705_, new_n9705_);
  or g_1562 (new_n4098_, not_pi254_0, not_new_n4167_);
  or g_1563 (new_n5408_, not_new_n5077_, not_new_n5076_);
  not g_1564 (not_new_n8137_, new_n8137_);
  not g_1565 (not_new_n1607__490, new_n1607_);
  not g_1566 (not_new_n1576__6782230728490, new_n1576_);
  or g_1567 (new_n3565_, not_new_n2147__0, not_new_n1612__57648010);
  buf g_1568 (po026, pi238);
  and g_1569 (new_n9475_, new_n9498_, new_n9610_);
  not g_1570 (not_new_n595__8235430, new_n595_);
  not g_1571 (not_new_n9444_, new_n9444_);
  not g_1572 (new_n8123_, new_n1051_);
  and g_1573 (new_n8246_, new_n8475_, new_n8476_);
  or g_1574 (new_n2420_, not_new_n1059__0, not_new_n598__490);
  not g_1575 (not_new_n7357__1, new_n7357_);
  or g_1576 (new_n5829_, not_new_n6114_, not_new_n6113_);
  not g_1577 (not_new_n9728_, new_n9728_);
  or g_1578 (po119, not_new_n3410_, not_new_n3411_);
  not g_1579 (not_new_n5992_, new_n5992_);
  not g_1580 (not_new_n9466_, new_n9466_);
  not g_1581 (not_new_n642__6782230728490, new_n642_);
  not g_1582 (not_pi181_0, pi181);
  or g_1583 (new_n2885_, not_new_n1616__168070, not_new_n2882_);
  or g_1584 (or_or_not_new_n9361__not_new_n9358__0_not_new_n9750_, or_not_new_n9361__not_new_n9358__0, not_new_n9750_);
  not g_1585 (not_new_n6773_, new_n6773_);
  not g_1586 (new_n4262_, new_n693_);
  not g_1587 (not_new_n2267_, new_n2267_);
  or g_1588 (new_n5766_, not_new_n5806_, not_new_n621__1176490);
  not g_1589 (new_n4090_, pi259);
  not g_1590 (not_new_n7599__2, new_n7599_);
  not g_1591 (not_new_n6992__2, new_n6992_);
  not g_1592 (not_new_n1053__7, new_n1053_);
  not g_1593 (not_pi178_2, pi178);
  not g_1594 (not_new_n1358_, new_n1358_);
  or g_1595 (new_n4024_, not_pi061_2, not_new_n4023_);
  not g_1596 (not_new_n1611__797922662976120010, new_n1611_);
  and g_1597 (new_n1225_, and_new_n1760__new_n1759_, new_n1758_);
  not g_1598 (not_new_n1241_, new_n1241_);
  not g_1599 (not_new_n3933__0, new_n3933_);
  not g_1600 (new_n9913_, new_n637_);
  not g_1601 (not_new_n4801__0, new_n4801_);
  or g_1602 (new_n4407_, not_new_n4286_, not_new_n649_);
  or g_1603 (new_n2530_, not_new_n608__1, not_new_n1012__0);
  or g_1604 (new_n6756_, not_new_n1601__57648010, not_new_n6503__1);
  not g_1605 (not_new_n7608_, new_n7608_);
  or g_1606 (new_n3141_, not_new_n1037__3, not_new_n928__57648010);
  not g_1607 (not_new_n4109_, new_n4109_);
  or g_1608 (new_n7558_, not_new_n735__0, not_new_n7418__0);
  not g_1609 (not_new_n9615_, new_n9615_);
  not g_1610 (not_new_n4114_, new_n4114_);
  not g_1611 (not_new_n1588__57648010, new_n1588_);
  not g_1612 (not_new_n611__8235430, new_n611_);
  not g_1613 (not_new_n9654_, new_n9654_);
  not g_1614 (not_new_n1237_, new_n1237_);
  not g_1615 (not_new_n4289_, new_n4289_);
  not g_1616 (not_new_n1601__6, new_n1601_);
  or g_1617 (new_n8046_, not_new_n8045_, not_new_n7841_);
  or g_1618 (new_n9077_, new_n1603_, new_n639_);
  not g_1619 (not_new_n6557_, new_n6557_);
  not g_1620 (not_new_n1007__0, new_n1007_);
  not g_1621 (not_new_n3451_, new_n3451_);
  or g_1622 (new_n6993_, not_new_n729_, not_new_n7028_);
  and g_1623 (new_n1224_, and_and_new_n1754__new_n1755__new_n1757_, new_n1756_);
  or g_1624 (new_n9893_, not_new_n9977_, not_new_n10044_);
  not g_1625 (not_new_n6604_, new_n6604_);
  or g_1626 (new_n7052_, not_new_n7395_, not_new_n7396_);
  or g_1627 (new_n3722_, not_new_n2342_, not_new_n983_);
  or g_1628 (new_n3790_, not_new_n2057_, not_new_n3484_);
  not g_1629 (not_new_n1997_, new_n1997_);
  or g_1630 (new_n9283_, not_new_n9118__0, not_new_n9281_);
  not g_1631 (not_new_n630__4, new_n630_);
  or g_1632 (new_n3472_, not_new_n1536__2326305139872070, not_pi018_0);
  or g_1633 (new_n7526_, not_new_n7029__1, not_new_n6994__1);
  not g_1634 (not_new_n961_, new_n961_);
  not g_1635 (not_new_n5264_, new_n5264_);
  not g_1636 (not_new_n7008__0, new_n7008_);
  not g_1637 (not_new_n5766__0, new_n5766_);
  or g_1638 (new_n6157_, not_new_n5770__2, not_new_n1601__24010);
  not g_1639 (new_n4228_, new_n678_);
  not g_1640 (not_new_n8958_, new_n8958_);
  or g_1641 (po186, not_new_n1355_, not_new_n1356_);
  or g_1642 (new_n9833_, not_new_n643__39098210485829880490, not_new_n9397__0);
  or g_1643 (po177, not_new_n3580_, not_new_n3581_);
  not g_1644 (not_new_n4918_, new_n4918_);
  not g_1645 (new_n8879_, new_n1603_);
  or g_1646 (new_n6387_, not_new_n6266_, not_new_n1069__490);
  not g_1647 (not_new_n9933_, new_n9933_);
  not g_1648 (not_pi176_2, pi176);
  not g_1649 (not_new_n4784__0, new_n4784_);
  not g_1650 (not_new_n600__8, new_n600_);
  or g_1651 (new_n8459_, not_new_n1051__57648010, not_new_n8124__0);
  not g_1652 (not_new_n3877_, new_n3877_);
  or g_1653 (new_n3638_, not_new_n984__968890104070, not_pi185_0);
  not g_1654 (not_new_n9618_, new_n9618_);
  or g_1655 (new_n3480_, not_pi112_0, not_new_n1537__24010);
  or g_1656 (new_n5828_, not_new_n6110_, not_new_n6109_);
  not g_1657 (not_new_n1599__8235430, new_n1599_);
  or g_1658 (new_n8335_, not_new_n627__138412872010, not_new_n8157_);
  not g_1659 (not_new_n5764__1, new_n5764_);
  not g_1660 (not_new_n1600__6782230728490, new_n1600_);
  or g_1661 (new_n3025_, not_new_n617__4, not_new_n3372__168070);
  not g_1662 (not_new_n4319_, new_n4319_);
  not g_1663 (new_n8154_, new_n1057_);
  not g_1664 (not_new_n8899__2, new_n8899_);
  not g_1665 (not_new_n599__6, new_n599_);
  or g_1666 (new_n9671_, not_new_n9480_, not_new_n9670_);
  or g_1667 (new_n2154_, not_new_n1583__403536070, not_new_n7677_);
  not g_1668 (not_new_n1728_, new_n1728_);
  or g_1669 (new_n5528_, not_new_n5435_, not_pi132_1);
  and g_1670 (new_n1333_, new_n2288_, new_n2289_);
  not g_1671 (not_new_n8674_, new_n8674_);
  not g_1672 (not_new_n623__5, new_n623_);
  not g_1673 (not_new_n2869_, new_n2869_);
  or g_1674 (new_n4511_, not_new_n4415_, not_new_n4416_);
  not g_1675 (not_new_n632__1, new_n632_);
  or g_1676 (new_n5146_, not_new_n626__24010, not_new_n1053__9);
  not g_1677 (new_n10073_, new_n9901_);
  or g_1678 (new_n7529_, not_new_n7527_, not_new_n7528_);
  or g_1679 (new_n3147_, not_new_n928__2824752490, not_new_n1069__3);
  not g_1680 (not_new_n626__70, new_n626_);
  or g_1681 (new_n9071_, not_new_n633__6782230728490, not_new_n9070_);
  not g_1682 (not_new_n8158__1, new_n8158_);
  not g_1683 (new_n8850_, new_n621_);
  or g_1684 (new_n8992_, new_n1037_, new_n632_);
  not g_1685 (not_pi144, pi144);
  or g_1686 (new_n750_, not_new_n3209_, not_new_n3208_);
  not g_1687 (not_new_n1631__1176490, key_gate_76);
  or g_1688 (new_n7885_, not_new_n7855__0, not_new_n7632__0);
  not g_1689 (not_new_n9902_, new_n9902_);
  and g_1690 (new_n3964_, and_and_and_not_pi056_1_not_pi055_1_not_pi054_1_not_pi053_1, not_pi052_1);
  or g_1691 (new_n2494_, not_new_n599__2326305139872070, not_new_n9961__0);
  not g_1692 (not_new_n4742_, new_n4742_);
  not g_1693 (not_new_n1027__168070, new_n1027_);
  not g_1694 (not_new_n9837_, new_n9837_);
  not g_1695 (not_pi216, pi216);
  not g_1696 (not_new_n10244_, new_n10244_);
  not g_1697 (not_new_n742__0, new_n742_);
  or g_1698 (new_n8419_, not_new_n8418_, not_new_n8343_);
  not g_1699 (not_new_n1399_, new_n1399_);
  not g_1700 (not_new_n9184_, new_n9184_);
  not g_1701 (not_new_n3310__0, new_n3310_);
  not g_1702 (not_new_n638__2, new_n638_);
  not g_1703 (not_new_n7011_, new_n7011_);
  not g_1704 (not_new_n9490_, new_n9490_);
  not g_1705 (not_pi003_0, pi003);
  not g_1706 (not_new_n1536__8235430, new_n1536_);
  or g_1707 (new_n5812_, not_new_n5996_, not_new_n6051_);
  not g_1708 (not_new_n1601_, new_n1601_);
  or g_1709 (new_n3859_, not_new_n6443__168070, not_new_n625__70);
  or g_1710 (new_n8415_, not_new_n8203_, not_new_n8248__1);
  not g_1711 (not_new_n9958_, new_n9958_);
  not g_1712 (not_new_n2509__7, new_n2509_);
  or g_1713 (new_n6401_, not_new_n6297_, not_new_n624__8235430);
  not g_1714 (not_new_n6778_, new_n6778_);
  and g_1715 (and_new_n4580__new_n4649_, new_n4649_, new_n4580_);
  not g_1716 (not_new_n8909_, new_n8909_);
  not g_1717 (not_new_n6567_, new_n6567_);
  not g_1718 (not_new_n7741__0, new_n7741_);
  or g_1719 (new_n1012_, not_new_n3345_, not_new_n3346_);
  not g_1720 (not_new_n637__5, new_n637_);
  not g_1721 (not_new_n8240_, new_n8240_);
  or g_1722 (new_n2045_, not_new_n1591__3430, not_new_n8919_);
  not g_1723 (not_new_n6472__0, new_n6472_);
  not g_1724 (not_new_n7742__0, new_n7742_);
  or g_1725 (new_n7224_, not_new_n7430_, not_new_n6992_);
  not g_1726 (not_new_n1333_, new_n1333_);
  not g_1727 (not_new_n1053__57648010, new_n1053_);
  not g_1728 (not_new_n5359_, new_n5359_);
  not g_1729 (not_new_n1581__0, new_n1581_);
  or g_1730 (new_n9672_, not_new_n9668_, not_new_n9511_);
  or g_1731 (new_n7760_, not_new_n7654_, not_new_n7937_);
  not g_1732 (not_new_n2683_, new_n2683_);
  not g_1733 (not_new_n7092_, new_n7092_);
  not g_1734 (not_new_n6324_, new_n6324_);
  or g_1735 (po167, not_new_n3561_, not_new_n3560_);
  not g_1736 (not_new_n720_, new_n720_);
  not g_1737 (not_new_n736__2, new_n736_);
  not g_1738 (not_new_n4308_, new_n4308_);
  not g_1739 (not_new_n4488_, new_n4488_);
  not g_1740 (not_new_n6974__6, new_n6974_);
  or g_1741 (new_n930_, not_new_n1023__0, or_not_new_n1027__not_new_n1028__0);
  not g_1742 (not_new_n639__332329305696010, new_n639_);
  not g_1743 (new_n1768_, new_n928_);
  and g_1744 (new_n594_, new_n1577_, new_n3387_);
  and g_1745 (new_n9463_, new_n9334_, new_n9328_);
  and g_1746 (new_n8799_, new_n8992_, new_n8991_);
  not g_1747 (not_new_n599__57648010, new_n599_);
  not g_1748 (not_new_n5459__0, new_n5459_);
  or g_1749 (new_n5968_, not_new_n5791_, not_new_n1055__70);
  not g_1750 (not_new_n1581__968890104070, new_n1581_);
  or g_1751 (new_n7988_, not_new_n7665__1, not_new_n1596__2824752490);
  not g_1752 (not_new_n625__70, new_n625_);
  not g_1753 (not_new_n2573_, new_n2573_);
  not g_1754 (not_new_n9204_, new_n9204_);
  not g_1755 (new_n2114_, new_n645_);
  or g_1756 (new_n2290_, not_new_n8097_, not_new_n1581__332329305696010);
  or g_1757 (new_n1820_, not_new_n594__1, not_new_n9873_);
  not g_1758 (not_new_n7490_, new_n7490_);
  and g_1759 (new_n9473_, and_new_n9512__new_n9773_, new_n9772_);
  not g_1760 (not_new_n604__3430, new_n604_);
  not g_1761 (not_new_n585__70, new_n585_);
  or g_1762 (new_n2230_, not_new_n7676_, not_new_n1583__968890104070);
  not g_1763 (not_new_n7535_, new_n7535_);
  or g_1764 (new_n10322_, not_new_n10022_, not_new_n10177_);
  not g_1765 (not_new_n4297_, new_n4297_);
  or g_1766 (new_n2458_, not_new_n4126__0, not_new_n600__2824752490);
  not g_1767 (new_n7004_, new_n725_);
  or g_1768 (new_n6604_, not_new_n6922_, not_new_n6923_);
  or g_1769 (new_n9682_, not_new_n9510__0, not_new_n9542_);
  or g_1770 (new_n7991_, not_new_n7990_, not_new_n7867_);
  not g_1771 (not_new_n8033_, new_n8033_);
  not g_1772 (not_new_n2318_, new_n2318_);
  or g_1773 (new_n10216_, not_new_n10029__2, not_new_n9866_);
  not g_1774 (not_new_n594__57648010, new_n594_);
  and g_1775 (new_n1290_, new_n2082_, new_n2081_);
  not g_1776 (not_new_n590__2, new_n590_);
  not g_1777 (not_new_n2499_, new_n2499_);
  and g_1778 (new_n1510_, new_n1511_, new_n3040_);
  not g_1779 (not_new_n2077_, new_n2077_);
  or g_1780 (new_n7553_, not_new_n734__0, not_new_n7409__0);
  or g_1781 (new_n8397_, not_new_n1065__6782230728490, not_new_n8162__1);
  not g_1782 (not_new_n10229_, new_n10229_);
  not g_1783 (not_new_n605__1, new_n605_);
  and g_1784 (and_new_n4348__new_n4301_, new_n4348_, new_n4301_);
  or g_1785 (new_n9252_, not_new_n8853_, not_new_n1600__138412872010);
  not g_1786 (not_new_n4354_, new_n4354_);
  not g_1787 (not_new_n625__6782230728490, new_n625_);
  not g_1788 (not_new_n7753__1, new_n7753_);
  or g_1789 (new_n3019_, not_new_n3372__3430, not_new_n619__2);
  not g_1790 (not_new_n8645__0, new_n8645_);
  or g_1791 (new_n6143_, not_new_n1598__490, not_new_n5765__0);
  and g_1792 (and_and_new_n3732__new_n3735__new_n3741_, and_new_n3732__new_n3735_, new_n3741_);
  not g_1793 (not_new_n2816_, new_n2816_);
  or g_1794 (new_n10099_, not_new_n9990_, not_new_n10097_);
  not g_1795 (not_new_n2804_, new_n2804_);
  or g_1796 (new_n3780_, not_new_n3779_, not_new_n3778_);
  not g_1797 (not_new_n625__10, new_n625_);
  not g_1798 (not_new_n2604_, new_n2604_);
  or g_1799 (new_n3105_, not_new_n581__4599865365447399609768010, not_new_n620__1);
  not g_1800 (new_n9388_, new_n1053_);
  or g_1801 (new_n6119_, not_new_n6118_, not_new_n6117_);
  or g_1802 (new_n9733_, not_new_n1045__5585458640832840070, not_new_n9363_);
  not g_1803 (not_new_n8250__0, new_n8250_);
  not g_1804 (not_pi141_3, pi141);
  not g_1805 (new_n4828_, new_n4800_);
  or g_1806 (new_n9790_, not_new_n9620__0, not_new_n9788_);
  not g_1807 (not_pi105_0, pi105);
  not g_1808 (not_new_n2019_, new_n2019_);
  not g_1809 (not_new_n4912_, new_n4912_);
  or g_1810 (new_n998_, not_new_n3314_, not_new_n3313_);
  or g_1811 (new_n8446_, not_new_n8088_, not_new_n8244__1);
  not g_1812 (not_new_n9170_, new_n9170_);
  not g_1813 (not_new_n585__24010, new_n585_);
  not g_1814 (not_new_n8132__0, new_n8132_);
  or g_1815 (new_n8737_, not_new_n1176__0, not_new_n8614_);
  not g_1816 (not_new_n1283_, new_n1283_);
  not g_1817 (not_new_n587_, new_n587_);
  not g_1818 (not_new_n1051_, new_n1051_);
  or g_1819 (new_n7828_, not_new_n7653_, not_new_n1057__8235430);
  not g_1820 (not_new_n1059__5, new_n1059_);
  not g_1821 (not_new_n6796_, new_n6796_);
  not g_1822 (not_new_n9262_, new_n9262_);
  not g_1823 (not_new_n8148__0, new_n8148_);
  not g_1824 (not_pi118_0, pi118);
  not g_1825 (not_new_n1589__0, new_n1589_);
  or g_1826 (new_n5358_, not_new_n630__168070, not_new_n4986__0);
  or g_1827 (new_n7825_, not_new_n7572_, not_new_n7824_);
  or g_1828 (new_n9212_, not_new_n1041__19773267430, not_new_n8826_);
  or g_1829 (new_n4881_, not_new_n4832_, not_new_n4789__0);
  not g_1830 (new_n4953_, new_n629_);
  not g_1831 (not_new_n8798__1, new_n8798_);
  or g_1832 (new_n4752_, not_new_n4733__0, not_new_n4816__0);
  or g_1833 (new_n7156_, not_new_n7266_, not_new_n7137_);
  or g_1834 (new_n2397_, not_new_n603__8, not_new_n626__1);
  not g_1835 (not_new_n994__47475615099430, new_n994_);
  not g_1836 (not_new_n6005_, new_n6005_);
  not g_1837 (not_new_n2897_, new_n2897_);
  not g_1838 (not_new_n5334_, new_n5334_);
  not g_1839 (not_new_n3311__5, new_n3311_);
  not g_1840 (not_new_n7036_, new_n7036_);
  not g_1841 (not_new_n3336_, new_n3336_);
  not g_1842 (not_new_n1547_, new_n1547_);
  or g_1843 (new_n2724_, or_or_not_new_n1473__not_new_n2722__not_new_n2723_, not_new_n936_);
  or g_1844 (new_n4052_, not_new_n4000__0, not_new_n3978__0);
  not g_1845 (new_n5442_, pi134);
  not g_1846 (not_new_n6310_, new_n6310_);
  or g_1847 (new_n1014_, not_new_n3349_, not_new_n3350_);
  not g_1848 (new_n4253_, new_n698_);
  and g_1849 (new_n1257_, new_n1927_, new_n1928_);
  not g_1850 (not_pi268_1, pi268);
  not g_1851 (not_pi041_2, pi041);
  not g_1852 (not_new_n4452__0, new_n4452_);
  not g_1853 (not_pi112, pi112);
  not g_1854 (not_new_n6632_, new_n6632_);
  not g_1855 (not_new_n1051__8, new_n1051_);
  not g_1856 (not_new_n8403_, new_n8403_);
  and g_1857 (and_new_n4984__new_n5390_, new_n5390_, new_n4984_);
  or g_1858 (new_n9728_, not_new_n9683_, not_new_n9484__0);
  not g_1859 (not_new_n928__490, new_n928_);
  not g_1860 (new_n6657_, new_n6534_);
  and g_1861 (new_n5848_, new_n5977_, new_n5726_);
  or g_1862 (new_n2583_, not_new_n609__7, not_new_n4468_);
  not g_1863 (not_new_n6156_, new_n6156_);
  not g_1864 (new_n6527_, new_n1053_);
  not g_1865 (not_new_n756_, new_n756_);
  not g_1866 (not_new_n1536__113988951853731430, new_n1536_);
  not g_1867 (not_new_n6355_, new_n6355_);
  or g_1868 (new_n3562_, not_new_n1538__8235430, not_pi147_0);
  not g_1869 (not_new_n5094_, new_n5094_);
  not g_1870 (not_pi070, pi070);
  not g_1871 (not_pi220, pi220);
  not g_1872 (not_new_n6599_, new_n6599_);
  not g_1873 (not_new_n581__3430, new_n581_);
  not g_1874 (not_new_n1245_, new_n1245_);
  or g_1875 (new_n9053_, not_new_n8985_, not_new_n8802_);
  not g_1876 (not_new_n1587_, new_n1587_);
  or g_1877 (new_n9136_, not_new_n633__47475615099430, not_new_n1067__2824752490);
  not g_1878 (not_new_n3324_, new_n3324_);
  not g_1879 (not_new_n9194_, new_n9194_);
  or g_1880 (new_n6188_, not_new_n5991_, not_new_n6187_);
  not g_1881 (not_new_n4826_, new_n4826_);
  not g_1882 (not_new_n3761_, new_n3761_);
  not g_1883 (not_new_n5994_, new_n5994_);
  and g_1884 (new_n6967_, new_n7179_, new_n6961_);
  or g_1885 (new_n3566_, not_new_n1538__403536070, not_pi149_0);
  not g_1886 (not_new_n10100__0, new_n10100_);
  or g_1887 (new_n5003_, not_new_n5295_, not_new_n5296_);
  or g_1888 (or_or_not_new_n2847__not_new_n2850__not_new_n2849_, or_not_new_n2847__not_new_n2850_, not_new_n2849_);
  not g_1889 (not_new_n601__6, new_n601_);
  not g_1890 (not_new_n6537__0, new_n6537_);
  not g_1891 (not_new_n5020_, new_n5020_);
  not g_1892 (not_new_n1011__1, new_n1011_);
  not g_1893 (not_new_n3389_, new_n3389_);
  not g_1894 (not_new_n1051__4, new_n1051_);
  not g_1895 (not_new_n7736_, new_n7736_);
  not g_1896 (not_new_n7495_, new_n7495_);
  and g_1897 (new_n598_, new_n1611_, new_n1588_);
  not g_1898 (not_new_n1003__2, new_n1003_);
  not g_1899 (not_new_n1580__1176490, new_n1580_);
  or g_1900 (or_not_new_n8528__not_new_n8429_, not_new_n8528_, not_new_n8429_);
  not g_1901 (new_n6487_, new_n635_);
  or g_1902 (new_n10247_, not_new_n1047__16284135979104490, not_new_n9878_);
  not g_1903 (not_new_n2802_, new_n2802_);
  not g_1904 (not_new_n5520_, new_n5520_);
  not g_1905 (not_new_n9018_, new_n9018_);
  and g_1906 (new_n1511_, new_n3039_, new_n998_);
  not g_1907 (not_new_n1596__4, new_n1596_);
  not g_1908 (not_new_n626__1915812313805664144010, new_n626_);
  or g_1909 (new_n5167_, new_n1067_, new_n633_);
  and g_1910 (po111, key_gate_101, pi090);
  not g_1911 (not_new_n3323_, new_n3323_);
  or g_1912 (or_not_new_n2838__not_new_n2841_, not_new_n2838_, not_new_n2841_);
  or g_1913 (or_or_not_new_n2527__not_new_n2531__not_new_n1421_, or_not_new_n2527__not_new_n2531_, not_new_n1421_);
  not g_1914 (not_new_n640__47475615099430, new_n640_);
  not g_1915 (not_new_n632__70, new_n632_);
  or g_1916 (or_not_new_n3113__not_new_n3112_, not_new_n3113_, not_new_n3112_);
  or g_1917 (or_not_new_n1299__not_new_n1297_, not_new_n1297_, not_new_n1299_);
  not g_1918 (not_new_n1229_, new_n1229_);
  not g_1919 (not_new_n5890__0, new_n5890_);
  not g_1920 (new_n9514_, new_n9406_);
  not g_1921 (not_new_n8979_, new_n8979_);
  or g_1922 (new_n4741_, not_new_n4797_, or_not_new_n4829__not_new_n4794_);
  or g_1923 (new_n2323_, not_new_n3366__0, not_new_n926_);
  not g_1924 (not_new_n5890__3, new_n5890_);
  or g_1925 (new_n9272_, not_new_n8879__0, not_new_n639__2326305139872070);
  or g_1926 (new_n4347_, not_new_n4340_, not_new_n4297_);
  not g_1927 (not_new_n5102_, new_n5102_);
  or g_1928 (new_n4778_, not_new_n4835__0, not_new_n4780__0);
  or g_1929 (new_n7305_, not_new_n7284_, not_new_n7160__0);
  or g_1930 (new_n2653_, not_new_n609__24010, not_new_n4458_);
  not g_1931 (not_new_n3278_, new_n3278_);
  not g_1932 (not_new_n2773_, new_n2773_);
  not g_1933 (not_new_n7014__1, new_n7014_);
  not g_1934 (not_new_n8117_, new_n8117_);
  not g_1935 (not_new_n6283_, new_n6283_);
  not g_1936 (not_new_n589__32199057558131797268376070, new_n589_);
  not g_1937 (not_new_n658_, new_n658_);
  not g_1938 (not_new_n10149_, new_n10149_);
  buf g_1939 (po016, pi209);
  not g_1940 (not_new_n6340_, new_n6340_);
  not g_1941 (not_new_n994__490, new_n994_);
  not g_1942 (not_new_n8221_, new_n8221_);
  not g_1943 (not_new_n5770__0, new_n5770_);
  or g_1944 (new_n2565_, not_new_n5489_, not_new_n605__5);
  or g_1945 (new_n7632_, not_new_n639__19773267430, not_new_n7633_);
  not g_1946 (not_new_n1049__10, new_n1049_);
  and g_1947 (and_new_n3750__new_n3753_, new_n3753_, new_n3750_);
  or g_1948 (new_n1027_, not_new_n3386_, not_new_n3385_);
  or g_1949 (new_n9156_, not_new_n8837__1, not_new_n9021_);
  not g_1950 (new_n4973_, new_n645_);
  or g_1951 (new_n1779_, not_new_n591__0, not_new_n1031__0);
  not g_1952 (not_new_n593__10, new_n593_);
  and g_1953 (new_n6616_, new_n6848_, new_n6849_);
  not g_1954 (not_new_n4079_, new_n4079_);
  or g_1955 (new_n3617_, not_new_n1611__490, not_new_n956_);
  not g_1956 (not_new_n9434_, new_n9434_);
  not g_1957 (not_new_n9071_, new_n9071_);
  not g_1958 (new_n8648_, new_n1600_);
  not g_1959 (not_new_n4481__0, new_n4481_);
  not g_1960 (not_new_n622__16284135979104490, new_n622_);
  or g_1961 (new_n7503_, not_new_n7502_, not_new_n7501_);
  not g_1962 (not_pi102_0, pi102);
  not g_1963 (not_new_n7401_, new_n7401_);
  not g_1964 (not_new_n1067__10, new_n1067_);
  or g_1965 (new_n2251_, not_new_n1584__6782230728490, not_new_n9439_);
  not g_1966 (not_new_n6995__0, new_n6995_);
  not g_1967 (not_new_n604__8235430, new_n604_);
  or g_1968 (or_not_new_n2883__not_new_n2886_, not_new_n2883_, not_new_n2886_);
  not g_1969 (not_new_n644__273687473400809163430, new_n644_);
  not g_1970 (new_n4956_, new_n625_);
  not g_1971 (not_new_n1616__168070, new_n1616_);
  and g_1972 (new_n9343_, new_n9656_, new_n9653_);
  xnor g_1973 (key_gate_67, new_n1645_, key_67);
  or g_1974 (new_n9723_, not_new_n9682_, not_new_n9372__0);
  not g_1975 (not_new_n5440_, new_n5440_);
  not g_1976 (not_new_n656_, new_n656_);
  not g_1977 (not_new_n6610_, new_n6610_);
  and g_1978 (and_new_n1274__new_n2008_, new_n2008_, new_n1274_);
  not g_1979 (not_new_n8306_, new_n8306_);
  or g_1980 (new_n8317_, not_new_n8316_, not_new_n8207_);
  or g_1981 (new_n6745_, not_new_n6625__0, not_new_n6586_);
  not g_1982 (not_new_n1516_, new_n1516_);
  or g_1983 (new_n8021_, not_new_n7885_, not_new_n7750__0);
  and g_1984 (new_n7089_, new_n7012_, new_n7161_);
  or g_1985 (or_or_not_new_n1482__not_new_n2858__not_new_n2857_, not_new_n2857_, or_not_new_n1482__not_new_n2858_);
  not g_1986 (not_new_n1524_, new_n1524_);
  and g_1987 (and_new_n3073__new_n998_, new_n998_, new_n3073_);
  or g_1988 (new_n4654_, not_pi179_3, not_new_n4450_);
  not g_1989 (not_new_n1012_, new_n1012_);
  and g_1990 (new_n9996_, new_n10161_, new_n9862_);
  not g_1991 (not_new_n3418_, new_n3418_);
  or g_1992 (new_n7294_, not_new_n7415__0, not_new_n6995__0);
  not g_1993 (not_new_n718_, new_n718_);
  not g_1994 (not_new_n728__0, new_n728_);
  not g_1995 (not_new_n1423_, new_n1423_);
  or g_1996 (new_n8362_, not_new_n640__138412872010, not_new_n8143_);
  not g_1997 (not_new_n7034_, new_n7034_);
  not g_1998 (new_n7158_, new_n6983_);
  not g_1999 (not_new_n610__8, new_n610_);
  not g_2000 (not_new_n7113__0, new_n7113_);
  not g_2001 (not_new_n6210_, new_n6210_);
  not g_2002 (not_pi173_0, pi173);
  not g_2003 (new_n8642_, new_n1171_);
  not g_2004 (not_new_n6598_, new_n6598_);
  not g_2005 (not_new_n2111_, new_n2111_);
  not g_2006 (not_new_n769_, new_n769_);
  and g_2007 (and_new_n6403__new_n6402_, new_n6402_, new_n6403_);
  not g_2008 (not_new_n7620_, new_n7620_);
  or g_2009 (new_n3080_, not_new_n1035__2, not_new_n581__797922662976120010);
  or g_2010 (new_n10142_, not_new_n1598__2326305139872070, not_new_n621__5585458640832840070);
  or g_2011 (or_not_new_n2935__not_new_n2934_, not_new_n2935_, not_new_n2934_);
  not g_2012 (not_new_n4078_, new_n4078_);
  not g_2013 (not_new_n3372__0, new_n3372_);
  not g_2014 (not_new_n650_, new_n650_);
  or g_2015 (new_n9663_, not_new_n9412__0, not_new_n9594_);
  not g_2016 (not_new_n5793_, new_n5793_);
  not g_2017 (not_new_n5852_, new_n5852_);
  or g_2018 (new_n6071_, not_new_n5878__1, not_new_n5726_);
  not g_2019 (not_new_n600__4, new_n600_);
  or g_2020 (new_n9174_, not_new_n9062_, not_new_n9059__0);
  not g_2021 (new_n4073_, pi274);
  not g_2022 (not_new_n5790__0, new_n5790_);
  not g_2023 (not_new_n7826_, new_n7826_);
  or g_2024 (or_or_not_new_n1287__not_new_n1285__not_new_n2059_, not_new_n2059_, or_not_new_n1287__not_new_n1285_);
  not g_2025 (not_new_n2766_, new_n2766_);
  and g_2026 (new_n1452_, and_new_n1451__new_n2679_, new_n2678_);
  not g_2027 (not_new_n5024_, new_n5024_);
  not g_2028 (not_new_n5878__3, new_n5878_);
  or g_2029 (new_n6828_, not_new_n6493__0, not_new_n1051__24010);
  not g_2030 (not_new_n4793_, new_n4793_);
  or g_2031 (new_n4340_, not_new_n4294_, not_new_n4333_);
  not g_2032 (not_new_n3796_, new_n3796_);
  or g_2033 (new_n6720_, not_new_n1065__168070, not_new_n6531__0);
  not g_2034 (not_new_n1004_, new_n1004_);
  or g_2035 (or_not_new_n8609__not_new_n8595__0, not_new_n8595__0, not_new_n8609_);
  not g_2036 (not_new_n6995__2, new_n6995_);
  not g_2037 (not_new_n3914__1, new_n3914_);
  not g_2038 (not_new_n4944__0, new_n4944_);
  not g_2039 (not_new_n7266_, new_n7266_);
  not g_2040 (not_new_n5672_, new_n5672_);
  not g_2041 (not_new_n7375_, new_n7375_);
  not g_2042 (not_new_n5907_, new_n5907_);
  not g_2043 (not_new_n631__70, new_n631_);
  not g_2044 (not_new_n6148_, new_n6148_);
  not g_2045 (not_new_n1583__3430, new_n1583_);
  or g_2046 (new_n5322_, not_new_n4922_, not_new_n1037__10);
  not g_2047 (not_new_n1321_, new_n1321_);
  not g_2048 (not_new_n2813_, new_n2813_);
  or g_2049 (new_n9577_, not_new_n9575_, not_new_n9576_);
  not g_2050 (not_new_n4690_, new_n4690_);
  not g_2051 (not_new_n5920_, new_n5920_);
  not g_2052 (not_new_n9588_, new_n9588_);
  not g_2053 (not_new_n1998_, new_n1998_);
  not g_2054 (not_new_n1010__5, new_n1010_);
  not g_2055 (not_new_n2744_, new_n2744_);
  or g_2056 (new_n4183_, not_pi248_3, not_new_n4146_);
  not g_2057 (not_new_n7032__0, new_n7032_);
  not g_2058 (not_new_n5941_, new_n5941_);
  xor g_2059 (key_gate_81, key_81, not_pi033_0);
  not g_2060 (not_new_n3485_, new_n3485_);
  not g_2061 (not_new_n6226__0, new_n6226_);
  not g_2062 (not_new_n7771__0, new_n7771_);
  not g_2063 (not_new_n1305_, new_n1305_);
  or g_2064 (new_n7499_, not_new_n7436__1, not_new_n724__1);
  not g_2065 (not_new_n3809_, new_n3809_);
  or g_2066 (new_n7688_, not_new_n7979_, not_new_n7980_);
  not g_2067 (not_new_n4416_, new_n4416_);
  and g_2068 (new_n9482_, and_new_n9510__new_n9851_, new_n9850_);
  not g_2069 (new_n4160_, new_n4151_);
  not g_2070 (not_new_n7445__0, new_n7445_);
  not g_2071 (not_pi145_3, pi145);
  not g_2072 (not_pi131_0, pi131);
  not g_2073 (not_new_n641__70, new_n641_);
  not g_2074 (not_new_n2584_, new_n2584_);
  not g_2075 (not_new_n3029_, new_n3029_);
  not g_2076 (not_pi115_0, pi115);
  and g_2077 (and_and_new_n3780__new_n3783__new_n3789_, new_n3789_, and_new_n3780__new_n3783_);
  not g_2078 (not_new_n585__1, new_n585_);
  or g_2079 (new_n9780_, not_new_n9381_, not_new_n1600__6782230728490);
  not g_2080 (not_new_n593__7, new_n593_);
  not g_2081 (not_new_n4589_, new_n4589_);
  or g_2082 (po198, or_or_not_new_n1555__not_new_n2434__not_new_n1379_, not_new_n1380_);
  or g_2083 (new_n5252_, not_new_n626__168070, not_new_n1053__10);
  not g_2084 (not_new_n3907_, new_n3907_);
  not g_2085 (not_new_n1053_, new_n1053_);
  not g_2086 (not_new_n3184__138412872010, new_n3184_);
  not g_2087 (new_n5743_, new_n1045_);
  or g_2088 (new_n6080_, not_new_n5890_, not_new_n5859_);
  or g_2089 (new_n4070_, not_new_n3997__0, not_new_n4013__0);
  not g_2090 (not_new_n2635_, new_n2635_);
  not g_2091 (not_new_n8828__0, new_n8828_);
  not g_2092 (not_new_n3106_, new_n3106_);
  not g_2093 (not_new_n589__657123623635342801395430, new_n589_);
  not g_2094 (not_new_n597__6, new_n597_);
  not g_2095 (not_new_n641__3, new_n641_);
  or g_2096 (new_n633_, not_new_n2074_, or_or_not_new_n2072__not_new_n2073__not_new_n2075_);
  or g_2097 (new_n9666_, new_n637_, new_n1065_);
  not g_2098 (new_n8168_, new_n621_);
  not g_2099 (not_new_n10286_, new_n10286_);
  not g_2100 (not_new_n6466_, new_n6466_);
  not g_2101 (not_new_n2972_, new_n2972_);
  or g_2102 (new_n978_, not_new_n2286_, or_or_not_new_n1335__not_new_n1333__not_new_n2287_);
  not g_2103 (not_new_n631__16284135979104490, new_n631_);
  not g_2104 (not_new_n1597__3, new_n1597_);
  not g_2105 (not_new_n617__7, new_n617_);
  not g_2106 (not_new_n2703_, new_n2703_);
  not g_2107 (not_new_n2943_, new_n2943_);
  not g_2108 (not_new_n3158_, new_n3158_);
  not g_2109 (not_new_n9869__0, new_n9869_);
  or g_2110 (new_n7210_, not_new_n7031_, not_new_n732_);
  not g_2111 (new_n4155_, new_n4077_);
  and g_2112 (new_n6311_, new_n627_, new_n6284_);
  or g_2113 (new_n2559_, not_pi272, not_po296_93874803376477543056490);
  not g_2114 (not_new_n3201_, new_n3201_);
  and g_2115 (new_n6581_, new_n6457_, new_n6712_);
  not g_2116 (not_new_n7673_, new_n7673_);
  not g_2117 (not_new_n9369_, new_n9369_);
  or g_2118 (new_n8184_, not_new_n8547_, not_new_n8546_);
  not g_2119 (not_new_n4453_, new_n4453_);
  or g_2120 (new_n6854_, not_new_n1039__8235430, not_new_n6482__2);
  not g_2121 (not_new_n599__24010, new_n599_);
  not g_2122 (not_new_n651_, new_n651_);
  not g_2123 (not_new_n1587__0, new_n1587_);
  not g_2124 (not_new_n1008__0, new_n1008_);
  and g_2125 (new_n5879_, new_n6100_, new_n6101_);
  not g_2126 (not_new_n2228_, new_n2228_);
  not g_2127 (not_new_n588__3, new_n588_);
  or g_2128 (or_or_not_new_n1259__not_new_n1257__not_new_n1926_, or_not_new_n1259__not_new_n1257_, not_new_n1926_);
  not g_2129 (new_n9013_, new_n8844_);
  not g_2130 (not_new_n4336_, new_n4336_);
  and g_2131 (and_new_n2327__new_n2328_, new_n2327_, new_n2328_);
  not g_2132 (not_po298_8235430, po298);
  not g_2133 (not_new_n626__93874803376477543056490, new_n626_);
  or g_2134 (new_n1725_, not_po296_797922662976120010, not_pi001_0);
  or g_2135 (new_n5271_, not_new_n4945__1, not_new_n5035_);
  not g_2136 (not_pi064_6, pi064);
  or g_2137 (new_n8504_, not_new_n8170__1, not_new_n1597__19773267430);
  not g_2138 (not_pi050_3, pi050);
  or g_2139 (new_n5368_, not_new_n5069_, not_new_n5068_);
  not g_2140 (not_new_n3863_, new_n3863_);
  not g_2141 (not_new_n603__403536070, new_n603_);
  not g_2142 (not_new_n5804__0, new_n5804_);
  or g_2143 (new_n4615_, not_new_n4423_, not_new_n1006__3);
  or g_2144 (new_n7274_, not_new_n7090_, not_new_n7272_);
  or g_2145 (or_not_new_n4818__not_new_n4749_, not_new_n4749_, not_new_n4818_);
  or g_2146 (new_n6145_, not_new_n6017_, not_new_n5890__3);
  and g_2147 (new_n9338_, new_n9331_, new_n9336_);
  not g_2148 (not_pi269_5, pi269);
  or g_2149 (new_n7446_, not_new_n775__6782230728490, not_new_n7130_);
  not g_2150 (new_n6677_, new_n6494_);
  or g_2151 (or_not_new_n1844__not_new_n1845_, not_new_n1844_, not_new_n1845_);
  not g_2152 (not_new_n3091_, new_n3091_);
  not g_2153 (not_new_n8270_, new_n8270_);
  or g_2154 (new_n2606_, not_new_n2603_, or_not_new_n2605__not_new_n2604_);
  or g_2155 (new_n4459_, not_new_n4635_, not_new_n4634_);
  or g_2156 (or_or_or_not_new_n2910__not_new_n2913__not_new_n2912__not_new_n2914_, not_new_n2914_, or_or_not_new_n2910__not_new_n2913__not_new_n2912_);
  not g_2157 (not_new_n4787__1, new_n4787_);
  not g_2158 (not_new_n10029__1, new_n10029_);
  not g_2159 (not_new_n7152_, new_n7152_);
  or g_2160 (new_n7302_, not_new_n7202_, not_new_n6983__1);
  not g_2161 (not_pi082, pi082);
  not g_2162 (not_new_n4126__2, new_n4126_);
  not g_2163 (not_new_n2685_, new_n2685_);
  not g_2164 (not_new_n7232_, new_n7232_);
  or g_2165 (new_n8793_, not_new_n1159__1, not_new_n8597_);
  not g_2166 (not_new_n984__8235430, new_n984_);
  or g_2167 (new_n9529_, not_new_n1043__968890104070, not_new_n9509_);
  not g_2168 (not_new_n5837_, new_n5837_);
  not g_2169 (not_new_n8807_, new_n8807_);
  or g_2170 (new_n4944_, not_new_n5112_, not_new_n4959_);
  or g_2171 (new_n2361_, not_new_n4748__0, not_new_n597__0);
  not g_2172 (new_n9366_, new_n1047_);
  and g_2173 (new_n3925_, new_n4029_, new_n3945_);
  not g_2174 (not_new_n5417_, new_n5417_);
  not g_2175 (not_new_n603__8235430, new_n603_);
  or g_2176 (new_n2362_, not_new_n628__1, not_new_n603__1);
  not g_2177 (not_new_n5768__0, new_n5768_);
  not g_2178 (not_new_n1010__6, new_n1010_);
  not g_2179 (not_new_n618__93874803376477543056490, new_n618_);
  not g_2180 (not_new_n989__1, new_n989_);
  not g_2181 (not_new_n645__0, new_n645_);
  or g_2182 (new_n9093_, new_n630_, new_n1601_);
  not g_2183 (new_n4025_, new_n3945_);
  and g_2184 (new_n7714_, new_n7866_, new_n7865_);
  not g_2185 (not_new_n593__138412872010, new_n593_);
  and g_2186 (new_n6321_, new_n6373_, new_n6409_);
  not g_2187 (not_pi243, pi243);
  not g_2188 (not_new_n8266_, new_n8266_);
  not g_2189 (not_new_n7300_, new_n7300_);
  and g_2190 (new_n1439_, new_n2620_, new_n2622_);
  or g_2191 (new_n7853_, not_new_n7776_, not_new_n7575_);
  or g_2192 (or_not_new_n2962__not_new_n2961_, not_new_n2962_, not_new_n2961_);
  or g_2193 (new_n6215_, not_new_n5907_, not_new_n5874_);
  not g_2194 (not_new_n10103_, new_n10103_);
  or g_2195 (new_n3507_, not_new_n1613__19773267430, not_new_n2204_);
  not g_2196 (not_new_n3746_, new_n3746_);
  not g_2197 (not_new_n8578_, new_n8578_);
  or g_2198 (new_n1920_, not_pi170, not_new_n586__8);
  not g_2199 (not_new_n638__70, new_n638_);
  and g_2200 (new_n8951_, new_n9136_, new_n8803_);
  not g_2201 (not_new_n4435_, new_n4435_);
  not g_2202 (not_new_n6779_, new_n6779_);
  or g_2203 (new_n3114_, not_new_n928__9, not_new_n1596__3);
  not g_2204 (not_new_n600__2326305139872070, new_n600_);
  or g_2205 (or_not_new_n2792__not_new_n2791_, not_new_n2791_, not_new_n2792_);
  not g_2206 (not_new_n4658_, new_n4658_);
  not g_2207 (not_new_n589__2326305139872070, new_n589_);
  not g_2208 (not_new_n5504_, new_n5504_);
  not g_2209 (not_new_n6902_, new_n6902_);
  not g_2210 (not_pi185, pi185);
  or g_2211 (new_n3098_, not_new_n928__3, not_new_n1043__3);
  not g_2212 (new_n5745_, new_n1047_);
  not g_2213 (not_new_n8637_, new_n8637_);
  not g_2214 (not_new_n8920_, new_n8920_);
  or g_2215 (new_n7350_, not_new_n771_, not_new_n6974__3);
  or g_2216 (new_n3303_, not_new_n1626__1, not_new_n1020__1);
  not g_2217 (not_new_n2135_, new_n2135_);
  not g_2218 (not_new_n1598__47475615099430, new_n1598_);
  not g_2219 (not_new_n3359_, new_n3359_);
  not g_2220 (not_new_n1435_, new_n1435_);
  or g_2221 (new_n6777_, not_new_n626__6782230728490, not_new_n6527__1);
  not g_2222 (not_new_n6926_, new_n6926_);
  or g_2223 (new_n632_, or_or_not_new_n1782__not_new_n1783__not_new_n1785_, not_new_n1784_);
  not g_2224 (not_new_n7647_, new_n7647_);
  not g_2225 (not_new_n984__9, new_n984_);
  not g_2226 (not_new_n8846__0, new_n8846_);
  not g_2227 (not_pi136, pi136);
  not g_2228 (new_n4735_, new_n1043_);
  not g_2229 (not_new_n6481__1, new_n6481_);
  not g_2230 (new_n7003_, new_n727_);
  not g_2231 (not_new_n730__0, new_n730_);
  or g_2232 (new_n9547_, not_new_n634__113988951853731430, not_new_n1047__6782230728490);
  or g_2233 (or_not_new_n1235__not_new_n1233_, not_new_n1233_, not_new_n1235_);
  or g_2234 (new_n9166_, not_new_n1596__47475615099430, not_new_n618__797922662976120010);
  or g_2235 (new_n3896_, not_new_n9924_, not_new_n627__3430);
  or g_2236 (new_n8520_, not_new_n8132__0, not_new_n1600__403536070);
  not g_2237 (not_pi186, pi186);
  not g_2238 (not_new_n679_, new_n679_);
  or g_2239 (new_n8026_, not_new_n7924_, not_new_n8025_);
  or g_2240 (new_n8385_, not_new_n8262_, not_new_n8368_);
  not g_2241 (not_new_n3978_, new_n3978_);
  or g_2242 (new_n5932_, not_new_n628__1176490, not_new_n5913_);
  not g_2243 (not_new_n3906_, new_n3906_);
  or g_2244 (po240, not_new_n3667_, not_new_n3666_);
  not g_2245 (not_new_n8794_, new_n8794_);
  not g_2246 (new_n6250_, new_n619_);
  not g_2247 (not_new_n1031__6, new_n1031_);
  not g_2248 (not_new_n2469_, new_n2469_);
  not g_2249 (not_new_n2738_, new_n2738_);
  or g_2250 (new_n1796_, not_new_n1581__0, not_new_n8184_);
  not g_2251 (not_new_n8900__0, new_n8900_);
  not g_2252 (not_new_n4558_, new_n4558_);
  not g_2253 (new_n9541_, new_n9372_);
  not g_2254 (not_new_n7032_, new_n7032_);
  or g_2255 (new_n10195_, not_new_n10061_, not_new_n10032_);
  not g_2256 (not_new_n1597_, new_n1597_);
  not g_2257 (new_n4101_, pi252);
  not g_2258 (not_new_n8250_, new_n8250_);
  not g_2259 (not_new_n984__5, new_n984_);
  not g_2260 (not_new_n1005__2, new_n1005_);
  or g_2261 (new_n8431_, not_new_n8359_, not_new_n8266_);
  not g_2262 (not_new_n8927_, new_n8927_);
  or g_2263 (new_n3251_, not_new_n589__5585458640832840070, not_new_n1045__5);
  or g_2264 (new_n5929_, not_new_n5749_, not_new_n1039__70);
  not g_2265 (not_new_n648__9, new_n648_);
  not g_2266 (not_new_n989__797922662976120010, new_n989_);
  not g_2267 (not_new_n6460_, new_n6460_);
  and g_2268 (and_new_n1270__new_n1989_, new_n1989_, new_n1270_);
  not g_2269 (not_new_n2000_, new_n2000_);
  not g_2270 (not_new_n1589__8235430, new_n1589_);
  or g_2271 (new_n8991_, new_n628_, new_n1039_);
  not g_2272 (not_new_n636__2824752490, new_n636_);
  not g_2273 (not_new_n9863_, new_n9863_);
  or g_2274 (new_n4555_, not_new_n4504_, not_new_n4554_);
  or g_2275 (new_n5705_, not_new_n5452__0, not_pi139_2);
  not g_2276 (not_new_n1596__332329305696010, new_n1596_);
  not g_2277 (not_new_n640__0, new_n640_);
  or g_2278 (new_n4859_, not_new_n4842_, not_new_n4762__0);
  not g_2279 (not_new_n1588__1, new_n1588_);
  not g_2280 (not_new_n8543_, new_n8543_);
  or g_2281 (new_n9958_, not_new_n10259_, not_new_n10258_);
  not g_2282 (not_new_n628__168070, new_n628_);
  or g_2283 (new_n2008_, not_new_n5020_, not_new_n1589__70);
  not g_2284 (not_new_n645__24010, new_n645_);
  not g_2285 (new_n7624_, new_n1599_);
  or g_2286 (new_n2922_, not_new_n7054_, not_new_n595__2824752490);
  not g_2287 (not_new_n7226_, new_n7226_);
  not g_2288 (not_new_n4651_, new_n4651_);
  not g_2289 (not_new_n589__4599865365447399609768010, new_n589_);
  not g_2290 (not_pi228, pi228);
  not g_2291 (not_new_n1041__47475615099430, new_n1041_);
  not g_2292 (not_pi163_0, pi163);
  or g_2293 (new_n4548_, not_pi171_1, not_new_n1019__2);
  not g_2294 (not_new_n8266__3, new_n8266_);
  not g_2295 (new_n6275_, new_n634_);
  or g_2296 (new_n5567_, not_pi143_1, not_new_n5462_);
  or g_2297 (new_n9303_, not_new_n8869_, not_new_n643__16284135979104490);
  or g_2298 (or_or_not_new_n1562__not_new_n2469__not_new_n1393_, not_new_n1393_, or_not_new_n1562__not_new_n2469_);
  not g_2299 (new_n6647_, new_n6538_);
  not g_2300 (not_new_n7016__0, new_n7016_);
  not g_2301 (not_new_n3116_, new_n3116_);
  not g_2302 (new_n4965_, new_n627_);
  or g_2303 (po054, key_gate_0, key_gate_68);
  or g_2304 (new_n6683_, not_new_n6493_, not_new_n1051__3430);
  not g_2305 (new_n6818_, new_n6640_);
  not g_2306 (not_new_n1059__10, new_n1059_);
  not g_2307 (not_new_n648__273687473400809163430, new_n648_);
  and g_2308 (new_n3974_, not_pi048_3, not_pi047_3);
  or g_2309 (new_n7892_, not_new_n1065__2824752490, not_new_n7655__1);
  and g_2310 (new_n6576_, new_n6836_, new_n6656_);
  not g_2311 (not_new_n5205_, new_n5205_);
  and g_2312 (and_and_and_new_n6422__new_n6426__new_n6360__new_n6359_, and_and_new_n6422__new_n6426__new_n6360_, new_n6359_);
  not g_2313 (not_pi132_3, pi132);
  not g_2314 (not_new_n2224_, new_n2224_);
  not g_2315 (not_pi050_2, pi050);
  or g_2316 (new_n2671_, not_new_n606__168070, not_new_n5482__0);
  not g_2317 (not_new_n1602__8235430, new_n1602_);
  not g_2318 (not_new_n5067_, new_n5067_);
  not g_2319 (new_n10038_, new_n9919_);
  or g_2320 (new_n8070_, not_new_n7650__0, not_new_n627__19773267430);
  not g_2321 (not_new_n597__1176490, new_n597_);
  not g_2322 (not_new_n738__1, new_n738_);
  not g_2323 (not_new_n8053_, new_n8053_);
  or g_2324 (new_n2149_, not_new_n587__2824752490, not_pi150);
  or g_2325 (new_n6813_, not_new_n6613__0, not_new_n6454_);
  not g_2326 (not_new_n1978_, new_n1978_);
  or g_2327 (new_n8000_, not_new_n7666__1, not_new_n7874_);
  not g_2328 (not_new_n7871_, new_n7871_);
  not g_2329 (not_new_n1675_, key_gate_34);
  or g_2330 (new_n9223_, not_new_n619__403536070, not_new_n8959_);
  not g_2331 (not_new_n1027__273687473400809163430, new_n1027_);
  or g_2332 (new_n6373_, not_new_n618__403536070, not_new_n6303_);
  and g_2333 (new_n1252_, and_and_new_n1896__new_n1899__new_n1897_, new_n1898_);
  not g_2334 (not_new_n1591__168070, new_n1591_);
  or g_2335 (new_n2358_, not_pi265_0, not_new_n600__0);
  not g_2336 (not_new_n6285_, new_n6285_);
  not g_2337 (not_new_n3141_, new_n3141_);
  not g_2338 (not_new_n775__1176490, new_n775_);
  not g_2339 (not_new_n1581__332329305696010, new_n1581_);
  not g_2340 (not_new_n3559_, new_n3559_);
  not g_2341 (not_pi140_3, pi140);
  not g_2342 (not_new_n1536__968890104070, new_n1536_);
  not g_2343 (not_new_n611__3430, new_n611_);
  or g_2344 (new_n9689_, not_new_n9659_, not_new_n9402__1);
  not g_2345 (not_pi057_3, pi057);
  or g_2346 (new_n10187_, not_new_n10002_, not_new_n10186_);
  or g_2347 (new_n2960_, not_new_n604__6782230728490, not_new_n644__3);
  and g_2348 (new_n8245_, new_n8468_, new_n8469_);
  or g_2349 (new_n1997_, not_new_n587__490, not_pi142);
  or g_2350 (new_n7531_, not_new_n7222__0, not_new_n7529_);
  not g_2351 (not_new_n1534_, key_gate_5);
  not g_2352 (not_new_n5808_, new_n5808_);
  not g_2353 (not_new_n7983_, new_n7983_);
  not g_2354 (not_new_n6243_, new_n6243_);
  not g_2355 (new_n4981_, new_n1065_);
  or g_2356 (new_n7542_, not_new_n7001__1, not_new_n7034__1);
  or g_2357 (new_n7518_, not_new_n7433__0, not_new_n727__0);
  not g_2358 (not_new_n7327_, new_n7327_);
  not g_2359 (not_new_n5725_, new_n5725_);
  not g_2360 (not_new_n604__4, new_n604_);
  not g_2361 (not_new_n6801_, new_n6801_);
  not g_2362 (not_new_n5546_, new_n5546_);
  not g_2363 (not_new_n7281_, new_n7281_);
  or g_2364 (new_n9310_, not_new_n8867_, not_new_n644__16284135979104490);
  not g_2365 (not_new_n631__797922662976120010, new_n631_);
  not g_2366 (not_new_n4130__0, new_n4130_);
  not g_2367 (not_new_n8921_, new_n8921_);
  or g_2368 (new_n6653_, not_new_n1598__24010, not_new_n6537_);
  or g_2369 (new_n4055_, not_pi063_1, not_new_n3942_);
  or g_2370 (new_n3462_, not_pi020_0, not_new_n1536__47475615099430);
  not g_2371 (not_new_n1045__138412872010, new_n1045_);
  not g_2372 (not_new_n5025_, new_n5025_);
  not g_2373 (new_n4967_, new_n1059_);
  not g_2374 (not_new_n3392_, new_n3392_);
  not g_2375 (not_pi103_0, pi103);
  or g_2376 (new_n2352_, not_new_n642__1, not_new_n603_);
  or g_2377 (new_n5628_, not_new_n5529_, not_new_n5626_);
  not g_2378 (not_new_n8992__0, new_n8992_);
  or g_2379 (new_n6842_, not_new_n6476__0, not_new_n635__403536070);
  or g_2380 (new_n10041_, new_n628_, new_n1039_);
  not g_2381 (not_new_n4811_, new_n4811_);
  not g_2382 (not_new_n989__6782230728490, new_n989_);
  or g_2383 (new_n6403_, not_new_n6298_, not_new_n632__57648010);
  not g_2384 (not_new_n9925_, new_n9925_);
  not g_2385 (not_new_n585__8, new_n585_);
  not g_2386 (not_new_n8429_, new_n8429_);
  or g_2387 (new_n10340_, not_new_n638__225393402906922580878632490, not_new_n9917_);
  not g_2388 (not_new_n6480__0, new_n6480_);
  or g_2389 (new_n3595_, not_new_n1611__1, not_new_n945_);
  not g_2390 (not_new_n3169_, new_n3169_);
  and g_2391 (new_n10005_, new_n9857_, new_n10196_);
  not g_2392 (not_new_n3872_, new_n3872_);
  not g_2393 (not_new_n10290_, new_n10290_);
  not g_2394 (not_new_n2646_, new_n2646_);
  or g_2395 (new_n8587_, not_new_n8156__0, not_new_n1053__403536070);
  or g_2396 (new_n9679_, not_new_n9541_, not_new_n9510_);
  not g_2397 (not_new_n4252_, new_n4252_);
  not g_2398 (not_new_n2021_, new_n2021_);
  not g_2399 (not_pi170, pi170);
  not g_2400 (not_pi063_1, pi063);
  and g_2401 (new_n9451_, new_n1037_, new_n632_);
  or g_2402 (new_n10024_, not_new_n10214_, not_new_n10230_);
  and g_2403 (new_n9976_, new_n628_, new_n1039_);
  not g_2404 (not_new_n8169__0, new_n8169_);
  not g_2405 (not_new_n3731_, new_n3731_);
  not g_2406 (not_new_n7764_, new_n7764_);
  not g_2407 (not_new_n3870_, new_n3870_);
  or g_2408 (new_n8490_, not_new_n8127__1, not_new_n8333_);
  not g_2409 (not_new_n5637_, new_n5637_);
  not g_2410 (not_new_n588__1176490, new_n588_);
  not g_2411 (not_new_n5486_, new_n5486_);
  not g_2412 (not_new_n7354_, new_n7354_);
  not g_2413 (not_new_n7157_, new_n7157_);
  or g_2414 (new_n4408_, not_new_n681__0, or_not_new_n4319__0_not_new_n713_);
  or g_2415 (new_n4518_, new_n1008_, pi164);
  or g_2416 (new_n5998_, not_new_n630__1176490, not_new_n5773_);
  not g_2417 (not_new_n3283_, new_n3283_);
  and g_2418 (new_n585_, new_n1030_, new_n1029_);
  not g_2419 (not_new_n1601__403536070, new_n1601_);
  not g_2420 (not_new_n5257_, new_n5257_);
  and g_2421 (and_and_new_n2508__new_n2510__new_n2507_, and_new_n2508__new_n2510_, new_n2507_);
  not g_2422 (not_new_n6201_, new_n6201_);
  not g_2423 (not_new_n1008__5, new_n1008_);
  not g_2424 (not_new_n1345_, new_n1345_);
  xnor g_2425 (key_gate_92, key_92, not_new_n1678_);
  and g_2426 (new_n6230_, new_n6401_, and_new_n6403__new_n6402_);
  not g_2427 (not_new_n4571_, new_n4571_);
  or g_2428 (new_n5594_, not_new_n5495_, not_new_n5496__0);
  or g_2429 (new_n7388_, not_new_n7113__2, not_new_n7112_);
  not g_2430 (new_n7630_, new_n1601_);
  not g_2431 (not_new_n9158_, new_n9158_);
  or g_2432 (new_n3543_, not_new_n1612__7, not_new_n1938__0);
  not g_2433 (not_new_n6222_, new_n6222_);
  not g_2434 (not_new_n9431_, new_n9431_);
  not g_2435 (not_new_n618__490, new_n618_);
  not g_2436 (not_new_n4737_, new_n4737_);
  not g_2437 (not_new_n4749__1, new_n4749_);
  not g_2438 (not_new_n618__3430, new_n618_);
  not g_2439 (not_pi205, pi205);
  not g_2440 (not_new_n1598__24010, new_n1598_);
  and g_2441 (new_n9988_, new_n10215_, new_n10094_);
  not g_2442 (not_new_n4017__2, new_n4017_);
  not g_2443 (not_new_n9213_, new_n9213_);
  not g_2444 (not_new_n629__16284135979104490, new_n629_);
  not g_2445 (new_n9515_, new_n9382_);
  not g_2446 (not_new_n6278_, new_n6278_);
  not g_2447 (not_new_n618__3, new_n618_);
  or g_2448 (new_n2503_, not_new_n598__797922662976120010, not_new_n1605__0);
  not g_2449 (not_new_n597__19773267430, new_n597_);
  or g_2450 (new_n2258_, not_new_n621_, not_new_n593__6782230728490);
  not g_2451 (not_new_n586_, new_n586_);
  not g_2452 (not_pi147_4, pi147);
  or g_2453 (new_n639_, not_new_n2150_, or_or_not_new_n2151__not_new_n2148__not_new_n2149_);
  not g_2454 (not_pi100_0, pi100);
  not g_2455 (not_new_n3297_, new_n3297_);
  or g_2456 (new_n9171_, not_new_n8935_, not_new_n8845__1);
  not g_2457 (not_new_n3185__70, new_n3185_);
  or g_2458 (new_n10220_, not_new_n10108_, not_new_n10218_);
  not g_2459 (not_new_n6044_, new_n6044_);
  not g_2460 (not_new_n624__2326305139872070, new_n624_);
  not g_2461 (not_new_n7695_, new_n7695_);
  not g_2462 (not_new_n705_, new_n705_);
  not g_2463 (not_new_n4655_, new_n4655_);
  not g_2464 (not_new_n6578_, new_n6578_);
  or g_2465 (new_n2734_, not_new_n4121__1, not_new_n994__1);
  or g_2466 (new_n7450_, not_new_n748_, not_new_n6974__6782230728490);
  not g_2467 (not_new_n2797_, new_n2797_);
  xnor g_2468 (key_gate_21, not_new_n1639_, key_21);
  not g_2469 (not_new_n10252_, new_n10252_);
  or g_2470 (new_n7768_, not_new_n7649_, not_new_n1053__1176490);
  not g_2471 (not_new_n6646_, new_n6646_);
  not g_2472 (not_new_n1601__47475615099430, new_n1601_);
  not g_2473 (not_new_n4121_, new_n4121_);
  not g_2474 (not_new_n597__1, new_n597_);
  not g_2475 (not_new_n6807_, new_n6807_);
  not g_2476 (not_new_n3185__10, new_n3185_);
  not g_2477 (not_new_n3760_, new_n3760_);
  not g_2478 (not_new_n4429__0, new_n4429_);
  not g_2479 (not_new_n6571_, new_n6571_);
  not g_2480 (not_new_n638__8235430, new_n638_);
  and g_2481 (new_n1472_, new_n1033_, new_n1032_);
  not g_2482 (new_n8708_, new_n1596_);
  not g_2483 (not_new_n581__4599865365447399609768010, new_n581_);
  and g_2484 (new_n6606_, new_n6449_, new_n6766_);
  or g_2485 (new_n2534_, not_new_n1013_, not_new_n607__0);
  or g_2486 (new_n9137_, not_new_n9135_, not_new_n8951_);
  not g_2487 (not_new_n1522_, new_n1522_);
  or g_2488 (new_n2202_, not_new_n4779_, not_new_n591__138412872010);
  and g_2489 (new_n1347_, new_n2352_, and_new_n2354__new_n2353_);
  or g_2490 (new_n3653_, not_new_n1615__0, not_new_n1611__797922662976120010);
  or g_2491 (or_not_new_n3124__not_new_n3125_, not_new_n3125_, not_new_n3124_);
  not g_2492 (not_pi036_0, pi036);
  or g_2493 (new_n2844_, not_new_n602__490, not_new_n646__2);
  or g_2494 (po085, not_new_n1212_, key_gate_95);
  not g_2495 (not_new_n8350_, new_n8350_);
  or g_2496 (or_not_new_n2892__not_new_n2895_, not_new_n2895_, not_new_n2892_);
  not g_2497 (not_new_n5777__0, new_n5777_);
  not g_2498 (not_new_n10338_, new_n10338_);
  or g_2499 (new_n6922_, not_new_n1069__168070, not_new_n6515__0);
  not g_2500 (not_new_n635__10, new_n635_);
  not g_2501 (not_new_n3089_, new_n3089_);
  or g_2502 (new_n9564_, not_new_n9520__0, not_new_n9523__0);
  or g_2503 (or_or_not_new_n1560__not_new_n2459__not_new_n1389_, not_new_n1389_, or_not_new_n1560__not_new_n2459_);
  not g_2504 (not_new_n4957_, new_n4957_);
  not g_2505 (not_new_n619__2, new_n619_);
  not g_2506 (not_new_n5632_, new_n5632_);
  not g_2507 (not_new_n7730_, new_n7730_);
  not g_2508 (not_new_n633__1176490, new_n633_);
  not g_2509 (not_new_n1536__6782230728490, new_n1536_);
  or g_2510 (new_n6718_, not_new_n6717_, not_new_n6449_);
  and g_2511 (new_n10004_, new_n3891_, and_new_n10032__new_n580_);
  not g_2512 (not_new_n643__7, new_n643_);
  not g_2513 (not_new_n5966_, new_n5966_);
  or g_2514 (new_n5535_, not_new_n5440_, not_pi134_1);
  or g_2515 (new_n1778_, not_new_n593_, not_new_n642_);
  or g_2516 (new_n10193_, not_new_n10192_, not_new_n9899_);
  not g_2517 (not_new_n1684_, key_gate_58);
  or g_2518 (new_n5635_, not_new_n1009__6, not_new_n5433_);
  not g_2519 (new_n1914_, new_n950_);
  not g_2520 (not_new_n595__70, new_n595_);
  not g_2521 (not_new_n4479__0, new_n4479_);
  not g_2522 (new_n6663_, new_n6496_);
  or g_2523 (new_n4994_, not_new_n5208_, not_new_n4954_);
  or g_2524 (new_n6627_, not_new_n6804_, not_new_n6794_);
  not g_2525 (not_new_n8134__2, new_n8134_);
  not g_2526 (not_new_n9823_, new_n9823_);
  not g_2527 (not_new_n7258__0, new_n7258_);
  or g_2528 (new_n769_, not_new_n3194_, not_new_n3195_);
  or g_2529 (new_n1152_, not_new_n3834_, not_new_n3833_);
  not g_2530 (not_new_n8478_, new_n8478_);
  or g_2531 (new_n4337_, not_new_n705_, not_new_n4239_);
  or g_2532 (new_n9807_, not_new_n9400_, not_new_n645__2326305139872070);
  not g_2533 (not_new_n3888_, new_n3888_);
  not g_2534 (new_n8145_, new_n1071_);
  not g_2535 (not_new_n1596__273687473400809163430, new_n1596_);
  not g_2536 (not_new_n7186_, new_n7186_);
  not g_2537 (not_new_n4163__0, new_n4163_);
  not g_2538 (not_new_n3461_, new_n3461_);
  or g_2539 (po275, or_or_or_not_new_n2803__not_new_n2806__not_new_n2805__not_new_n2807_, not_new_n2804_);
  not g_2540 (not_new_n5561_, new_n5561_);
  not g_2541 (new_n1605_, new_n983_);
  not g_2542 (new_n7656_, new_n638_);
  not g_2543 (not_new_n5569_, new_n5569_);
  not g_2544 (not_new_n5032_, new_n5032_);
  or g_2545 (new_n999_, not_new_n3320_, not_new_n3319_);
  not g_2546 (not_new_n6482__2, new_n6482_);
  not g_2547 (not_new_n4672_, new_n4672_);
  not g_2548 (not_new_n598_, new_n598_);
  not g_2549 (new_n6691_, new_n6495_);
  or g_2550 (new_n5822_, not_new_n6189_, not_new_n6188_);
  or g_2551 (new_n8144_, not_new_n645__138412872010, not_new_n8145_);
  not g_2552 (new_n1597_, new_n977_);
  or g_2553 (new_n7311_, not_new_n736__0, not_new_n7018__0);
  not g_2554 (not_new_n9404_, new_n9404_);
  or g_2555 (new_n754_, not_new_n3217_, not_new_n3216_);
  not g_2556 (not_new_n1027__8235430, new_n1027_);
  or g_2557 (new_n10097_, not_new_n10035_, not_new_n9858_);
  not g_2558 (not_new_n586__7, new_n586_);
  not g_2559 (not_new_n7218_, new_n7218_);
  not g_2560 (not_new_n1630_, new_n1630_);
  not g_2561 (not_new_n4450__0, new_n4450_);
  or g_2562 (new_n6381_, not_new_n1600__3430, not_new_n6280__0);
  not g_2563 (not_new_n3315__968890104070, new_n3315_);
  not g_2564 (not_pi048_2, pi048);
  not g_2565 (not_new_n1838_, new_n1838_);
  or g_2566 (new_n3284_, not_new_n633__8, not_new_n3184__57648010);
  not g_2567 (not_new_n2828_, new_n2828_);
  or g_2568 (new_n8763_, not_new_n8684_, not_new_n8596__1);
  not g_2569 (not_new_n5776_, new_n5776_);
  or g_2570 (new_n3528_, not_pi130_0, not_new_n1538__0);
  not g_2571 (not_new_n6708_, new_n6708_);
  not g_2572 (not_new_n628__332329305696010, new_n628_);
  not g_2573 (not_new_n7939_, new_n7939_);
  or g_2574 (new_n2099_, not_new_n9342_, not_new_n1584__1176490);
  not g_2575 (not_new_n6062_, new_n6062_);
  not g_2576 (not_new_n986_, new_n986_);
  not g_2577 (not_new_n2919_, new_n2919_);
  not g_2578 (not_new_n5811_, new_n5811_);
  not g_2579 (new_n5926_, new_n5899_);
  and g_2580 (new_n1461_, and_and_new_n3804__new_n3807__new_n3813_, new_n3810_);
  or g_2581 (or_not_new_n2917__not_new_n2916_, not_new_n2916_, not_new_n2917_);
  not g_2582 (not_new_n581__138412872010, new_n581_);
  or g_2583 (new_n2486_, not_new_n597__47475615099430, not_new_n4769__0);
  and g_2584 (new_n4472_, new_n4587_, new_n4588_);
  not g_2585 (not_new_n5892_, new_n5892_);
  not g_2586 (not_new_n1827_, new_n1827_);
  or g_2587 (new_n4869_, not_new_n4837__1, not_new_n4775__1);
  or g_2588 (new_n6673_, not_new_n1041__3430, not_new_n6489_);
  not g_2589 (not_new_n9457_, new_n9457_);
  not g_2590 (not_new_n984__403536070, new_n984_);
  not g_2591 (new_n4968_, new_n644_);
  or g_2592 (new_n5616_, not_new_n5440__0, not_pi134_2);
  or g_2593 (po135, not_new_n3490_, not_new_n3491_);
  or g_2594 (new_n5323_, not_new_n5059_, not_new_n619__8);
  or g_2595 (new_n10205_, not_new_n10178_, not_new_n9905__1);
  not g_2596 (not_new_n6655__0, new_n6655_);
  or g_2597 (new_n1995_, not_new_n1272_, not_new_n1990_);
  not g_2598 (not_new_n5813_, new_n5813_);
  or g_2599 (new_n4086_, not_new_n4140_, not_new_n4159_);
  not g_2600 (not_new_n7967_, new_n7967_);
  or g_2601 (new_n948_, not_new_n1868_, or_or_not_new_n1247__not_new_n1245__not_new_n1869_);
  not g_2602 (not_new_n6764_, new_n6764_);
  or g_2603 (new_n5646_, not_new_n1010__6, not_new_n5518_);
  not g_2604 (not_new_n653_, new_n653_);
  or g_2605 (new_n9241_, not_new_n9239_, not_new_n9240_);
  and g_2606 (new_n9478_, new_n9817_, and_new_n9412__new_n9818_);
  not g_2607 (not_new_n6249_, new_n6249_);
  not g_2608 (not_new_n645__403536070, new_n645_);
  or g_2609 (new_n2381_, not_new_n597__4, not_new_n4726__0);
  not g_2610 (not_new_n3315__1176490, new_n3315_);
  and g_2611 (po096, pi075, key_gate_101);
  or g_2612 (new_n3064_, not_new_n638__4, not_new_n3372__16284135979104490);
  not g_2613 (new_n4170_, new_n4102_);
  not g_2614 (not_new_n4951_, new_n4951_);
  or g_2615 (or_not_new_n4814__not_new_n4734_, not_new_n4734_, not_new_n4814_);
  or g_2616 (new_n8094_, not_new_n8407_, not_new_n8404_);
  not g_2617 (not_new_n1613__6, new_n1613_);
  not g_2618 (not_new_n1618_, new_n1618_);
  not g_2619 (new_n8634_, new_n1151_);
  not g_2620 (not_new_n7806_, new_n7806_);
  not g_2621 (not_new_n3173_, new_n3173_);
  not g_2622 (not_new_n5877_, new_n5877_);
  not g_2623 (not_new_n604__7, new_n604_);
  not g_2624 (not_new_n634__10, new_n634_);
  or g_2625 (po184, not_new_n1351_, not_new_n1352_);
  and g_2626 (new_n7722_, new_n8014_, new_n7770_);
  not g_2627 (not_new_n1007__1, new_n1007_);
  not g_2628 (not_new_n7804_, new_n7804_);
  and g_2629 (new_n6360_, new_n6425_, new_n6424_);
  or g_2630 (new_n10252_, not_new_n10250_, not_new_n10052__0);
  not g_2631 (not_new_n998_, new_n998_);
  not g_2632 (not_new_n5019_, new_n5019_);
  or g_2633 (new_n3902_, not_new_n9928_, not_new_n1059__7);
  or g_2634 (new_n4191_, not_pi273_1, not_new_n4110_);
  or g_2635 (new_n3157_, not_new_n638__6, not_new_n581__7490483309651862334944941026945644936490);
  or g_2636 (new_n5689_, not_new_n5685_, or_not_new_n5460__not_new_n5686__1);
  not g_2637 (not_new_n10302_, new_n10302_);
  or g_2638 (new_n3482_, not_new_n1536__113988951853731430, not_pi016_0);
  not g_2639 (not_new_n5657_, new_n5657_);
  not g_2640 (not_new_n4777_, new_n4777_);
  not g_2641 (new_n8609_, new_n1037_);
  not g_2642 (not_new_n586__10, new_n586_);
  not g_2643 (not_new_n3502_, new_n3502_);
  not g_2644 (not_new_n2038_, new_n2038_);
  or g_2645 (po258, not_new_n3703_, not_new_n3702_);
  or g_2646 (new_n3103_, not_new_n3315__7, not_new_n628__5);
  not g_2647 (not_pi066_0, pi066);
  not g_2648 (not_new_n1585__57648010, new_n1585_);
  not g_2649 (not_new_n3838_, new_n3838_);
  or g_2650 (new_n8899_, or_not_new_n9176__not_new_n9177_, not_new_n9065_);
  not g_2651 (not_new_n1534__9, key_gate_5);
  not g_2652 (not_new_n589__93874803376477543056490, new_n589_);
  or g_2653 (new_n1003_, not_new_n3327_, not_new_n3328_);
  not g_2654 (not_new_n9487_, new_n9487_);
  and g_2655 (new_n7571_, new_n7768_, new_n7821_);
  or g_2656 (new_n6216_, not_new_n5791__2, not_new_n1055__24010);
  not g_2657 (not_new_n588__57648010, new_n588_);
  and g_2658 (new_n1269_, new_n1984_, new_n1985_);
  not g_2659 (not_new_n633__490, new_n633_);
  not g_2660 (not_new_n3775_, new_n3775_);
  not g_2661 (not_new_n8116_, new_n8116_);
  not g_2662 (not_new_n1562_, new_n1562_);
  not g_2663 (not_new_n7340_, new_n7340_);
  not g_2664 (not_new_n9867_, new_n9867_);
  not g_2665 (not_new_n1588__16284135979104490, new_n1588_);
  not g_2666 (not_new_n625__2326305139872070, new_n625_);
  not g_2667 (not_new_n7837__0, new_n7837_);
  not g_2668 (not_new_n1450_, new_n1450_);
  or g_2669 (new_n10192_, new_n1051_, new_n647_);
  not g_2670 (not_new_n9573_, new_n9573_);
  not g_2671 (not_new_n9260_, new_n9260_);
  not g_2672 (not_new_n7980_, new_n7980_);
  or g_2673 (new_n9312_, not_new_n8862_, not_new_n636__332329305696010);
  not g_2674 (not_new_n8457_, new_n8457_);
  or g_2675 (new_n3151_, not_new_n633__6, not_new_n581__152867006319425761937651857692768264010);
  not g_2676 (new_n7162_, new_n6997_);
  or g_2677 (new_n10240_, not_new_n10061__0, not_new_n10238_);
  not g_2678 (not_new_n9400_, new_n9400_);
  not g_2679 (not_new_n4547_, new_n4547_);
  or g_2680 (new_n7057_, not_new_n7484_, not_new_n7483_);
  or g_2681 (new_n10297_, not_new_n10296_, not_new_n10295_);
  or g_2682 (new_n2005_, not_new_n1581__70, not_new_n8189_);
  not g_2683 (not_new_n7717_, new_n7717_);
  or g_2684 (new_n9424_, not_new_n9599_, not_new_n9600_);
  not g_2685 (not_new_n2843_, new_n2843_);
  not g_2686 (not_new_n641__168070, new_n641_);
  not g_2687 (new_n7329_, new_n7153_);
  not g_2688 (new_n6277_, new_n647_);
  not g_2689 (not_new_n8418_, new_n8418_);
  not g_2690 (not_new_n8458_, new_n8458_);
  and g_2691 (new_n6318_, new_n6232_, new_n6282_);
  not g_2692 (not_new_n5882__0, new_n5882_);
  not g_2693 (not_pi036_3, pi036);
  not g_2694 (not_new_n7941_, new_n7941_);
  not g_2695 (not_new_n8187_, new_n8187_);
  not g_2696 (not_new_n1538__8, new_n1538_);
  and g_2697 (new_n6589_, new_n6748_, new_n6747_);
  not g_2698 (not_new_n630__2, new_n630_);
  or g_2699 (new_n5834_, not_new_n6201_, not_new_n6200_);
  not g_2700 (not_new_n632__57648010, new_n632_);
  and g_2701 (new_n5049_, new_n5227_, new_n4904_);
  not g_2702 (not_new_n591__3430, new_n591_);
  not g_2703 (new_n4163_, new_n4089_);
  not g_2704 (not_new_n6613__0, new_n6613_);
  not g_2705 (not_new_n8304_, new_n8304_);
  and g_2706 (new_n8802_, new_n9052_, new_n9051_);
  or g_2707 (new_n5539_, not_pi135_1, not_new_n1005__5);
  not g_2708 (not_new_n1568_, new_n1568_);
  and g_2709 (and_and_new_n6422__new_n6426__new_n6360_, new_n6360_, and_new_n6422__new_n6426_);
  not g_2710 (not_new_n617__39098210485829880490, new_n617_);
  not g_2711 (not_new_n631__6, new_n631_);
  and g_2712 (new_n9454_, new_n9528_, and_new_n9525__new_n9526_);
  not g_2713 (not_new_n6550_, new_n6550_);
  not g_2714 (not_new_n2474_, new_n2474_);
  or g_2715 (new_n7898_, not_new_n7934_, not_new_n7897_);
  not g_2716 (not_new_n9459_, new_n9459_);
  not g_2717 (not_new_n5921_, new_n5921_);
  or g_2718 (po288, or_or_or_not_new_n2919__not_new_n2922__not_new_n2921__not_new_n2923_, not_new_n2920_);
  not g_2719 (not_new_n1031__1176490, new_n1031_);
  or g_2720 (new_n5212_, not_new_n5045_, not_new_n5211_);
  not g_2721 (not_new_n8143_, new_n8143_);
  not g_2722 (not_pi268_0, pi268);
  or g_2723 (new_n2582_, not_new_n2509__6, not_pi200);
  not g_2724 (not_new_n1028__5, new_n1028_);
  not g_2725 (not_new_n1047__1, new_n1047_);
  or g_2726 (new_n940_, not_new_n1024__1, not_new_n1023__2);
  not g_2727 (not_new_n1155__0, new_n1155_);
  and g_2728 (and_and_not_pi040_1_not_pi039_1_not_pi042_1, and_not_pi040_1_not_pi039_1, not_pi042_1);
  not g_2729 (not_new_n7363__0, new_n7363_);
  not g_2730 (not_new_n587__2326305139872070, new_n587_);
  or g_2731 (new_n4716_, not_new_n4412_, not_new_n1020__5);
  not g_2732 (not_new_n617_, new_n617_);
  not g_2733 (not_new_n5741__1, new_n5741_);
  not g_2734 (not_new_n5346_, new_n5346_);
  not g_2735 (not_new_n7035__1, new_n7035_);
  not g_2736 (not_pi217, pi217);
  not g_2737 (not_new_n2921_, new_n2921_);
  not g_2738 (not_new_n5434_, new_n5434_);
  not g_2739 (not_new_n1316_, new_n1316_);
  or g_2740 (new_n2497_, not_new_n600__16284135979104490, not_new_n4072__0);
  not g_2741 (not_new_n641__4, new_n641_);
  or g_2742 (new_n3899_, not_new_n3900_, not_new_n3901_);
  and g_2743 (new_n9859_, new_n10112_, new_n10111_);
  not g_2744 (not_new_n6767_, new_n6767_);
  not g_2745 (not_new_n5911_, new_n5911_);
  not g_2746 (not_new_n5874_, new_n5874_);
  not g_2747 (not_new_n3185__8, new_n3185_);
  or g_2748 (or_not_new_n8799__0_not_new_n8996__0, not_new_n8799__0, not_new_n8996__0);
  and g_2749 (new_n4750_, new_n4849_, new_n4848_);
  not g_2750 (not_new_n1063__4, new_n1063_);
  not g_2751 (not_new_n7657_, new_n7657_);
  not g_2752 (not_pi144_1, pi144);
  not g_2753 (not_new_n1598__3430, new_n1598_);
  not g_2754 (not_new_n1601__5585458640832840070, new_n1601_);
  not g_2755 (not_new_n1007__3, new_n1007_);
  not g_2756 (not_new_n606__6, new_n606_);
  not g_2757 (not_new_n6969_, new_n6969_);
  not g_2758 (not_new_n595__168070, new_n595_);
  not g_2759 (not_new_n1055__39098210485829880490, new_n1055_);
  not g_2760 (not_new_n1960_, new_n1960_);
  or g_2761 (new_n8098_, or_not_new_n8413__not_new_n8252_, not_new_n8276_);
  or g_2762 (new_n2609_, not_po296_1577753820348458066150427430, not_pi256);
  not g_2763 (not_new_n7059_, new_n7059_);
  or g_2764 (new_n5116_, not_new_n4945__0, not_new_n5115_);
  not g_2765 (not_new_n8560_, new_n8560_);
  not g_2766 (not_new_n7140_, new_n7140_);
  not g_2767 (not_new_n637__968890104070, new_n637_);
  not g_2768 (new_n3940_, pi036);
  not g_2769 (not_new_n8618__0, new_n8618_);
  not g_2770 (not_new_n1061__19773267430, new_n1061_);
  and g_2771 (and_and_new_n2181__new_n2184__new_n2182_, and_new_n2181__new_n2184_, new_n2182_);
  not g_2772 (not_new_n5715_, new_n5715_);
  or g_2773 (new_n8774_, not_new_n8621_, not_new_n1165__0);
  not g_2774 (not_new_n1594__8, new_n1594_);
  not g_2775 (not_new_n1065__24010, new_n1065_);
  not g_2776 (new_n5150_, new_n5078_);
  not g_2777 (not_new_n1591__0, new_n1591_);
  or g_2778 (new_n1814_, not_new_n1584__1, not_new_n9346_);
  not g_2779 (not_new_n3743_, new_n3743_);
  and g_2780 (po102, pi081, key_gate_101);
  not g_2781 (not_new_n6371_, new_n6371_);
  and g_2782 (new_n5843_, new_n5921_, new_n6099_);
  or g_2783 (new_n4106_, not_pi258_0, not_new_n4171_);
  not g_2784 (not_new_n5798__2, new_n5798_);
  or g_2785 (new_n4184_, not_new_n4176_, not_new_n4074_);
  not g_2786 (new_n2171_, new_n625_);
  and g_2787 (new_n9476_, and_new_n9402__new_n9804_, new_n9803_);
  or g_2788 (new_n8971_, not_new_n641__57648010, not_new_n1031__57648010);
  not g_2789 (not_new_n4184_, new_n4184_);
  or g_2790 (new_n5224_, not_new_n5223_, not_new_n4998__0);
  or g_2791 (new_n8285_, not_new_n1037__57648010, not_new_n8111_);
  or g_2792 (or_or_not_new_n3914__not_new_n3969__not_new_n4014_, not_new_n4014_, or_not_new_n3914__not_new_n3969_);
  not g_2793 (new_n6515_, new_n646_);
  xnor g_2794 (key_gate_61, new_n1663_, key_61);
  not g_2795 (not_new_n3469_, new_n3469_);
  or g_2796 (new_n1987_, not_new_n1580__70, not_new_n6463_);
  not g_2797 (not_new_n9676_, new_n9676_);
  or g_2798 (new_n3941_, or_or_not_new_n3965__not_new_n3966__not_new_n3968_, not_new_n3967_);
  not g_2799 (not_new_n9386__0, new_n9386_);
  and g_2800 (new_n5052_, and_new_n5083__new_n5411_, new_n5410_);
  not g_2801 (not_new_n5256_, new_n5256_);
  or g_2802 (new_n3666_, not_pi219, not_new_n989__5);
  not g_2803 (not_new_n7105_, new_n7105_);
  not g_2804 (not_new_n1004__1, new_n1004_);
  not g_2805 (not_pi120, pi120);
  not g_2806 (not_new_n8259_, new_n8259_);
  not g_2807 (not_new_n5842_, new_n5842_);
  not g_2808 (not_new_n2950_, new_n2950_);
  not g_2809 (not_new_n581__4, new_n581_);
  not g_2810 (not_new_n3376_, new_n3376_);
  not g_2811 (not_new_n9634_, new_n9634_);
  not g_2812 (not_new_n994__2326305139872070, new_n994_);
  not g_2813 (not_new_n7255_, new_n7255_);
  or g_2814 (new_n6938_, not_new_n6638_, not_new_n6761__0);
  not g_2815 (not_new_n10330_, new_n10330_);
  or g_2816 (new_n9612_, not_new_n1603__6782230728490, not_new_n639__16284135979104490);
  or g_2817 (new_n7618_, not_new_n7793_, not_new_n7615_);
  or g_2818 (new_n5869_, not_new_n6186_, not_new_n6185_);
  not g_2819 (not_new_n7522_, new_n7522_);
  not g_2820 (new_n6649_, new_n6473_);
  and g_2821 (new_n4484_, new_n4629_, new_n4630_);
  not g_2822 (not_new_n6147_, new_n6147_);
  or g_2823 (po075, not_new_n1202_, key_gate_127);
  not g_2824 (new_n1886_, new_n634_);
  and g_2825 (new_n1485_, new_n2937_, new_n1486_);
  not g_2826 (not_new_n4073_, new_n4073_);
  not g_2827 (not_new_n4163_, new_n4163_);
  not g_2828 (not_new_n1600_, new_n1600_);
  not g_2829 (not_pi036_1, pi036);
  not g_2830 (not_new_n8243_, new_n8243_);
  not g_2831 (new_n4922_, new_n632_);
  and g_2832 (and_new_n3058__new_n998_, new_n998_, new_n3058_);
  not g_2833 (not_new_n627__2, new_n627_);
  not g_2834 (not_new_n1581__70, new_n1581_);
  not g_2835 (new_n2228_, new_n622_);
  not g_2836 (not_new_n5240__0, new_n5240_);
  or g_2837 (new_n7061_, not_new_n7511_, not_new_n7512_);
  not g_2838 (new_n7129_, new_n752_);
  not g_2839 (not_new_n6628_, new_n6628_);
  not g_2840 (not_new_n7611__0, new_n7611_);
  and g_2841 (new_n1365_, and_new_n2399__new_n2398_, new_n2397_);
  not g_2842 (not_new_n629__138412872010, new_n629_);
  not g_2843 (not_new_n2243_, new_n2243_);
  or g_2844 (new_n1797_, not_new_n6553_, not_new_n1580__1);
  not g_2845 (not_new_n1806_, new_n1806_);
  not g_2846 (new_n6474_, new_n648_);
  or g_2847 (new_n4350_, not_new_n4250_, not_new_n700_);
  not g_2848 (not_new_n631__9, new_n631_);
  not g_2849 (not_pi275_0, pi275);
  not g_2850 (not_new_n8740_, new_n8740_);
  not g_2851 (not_new_n1594__6, new_n1594_);
  not g_2852 (not_new_n6713_, new_n6713_);
  not g_2853 (not_new_n4479_, new_n4479_);
  not g_2854 (not_new_n636__6, new_n636_);
  or g_2855 (new_n8185_, not_new_n8552_, not_new_n8551_);
  not g_2856 (not_new_n2674_, new_n2674_);
  or g_2857 (new_n4021_, not_new_n4020_, not_pi035_3);
  not g_2858 (not_new_n4550_, new_n4550_);
  or g_2859 (or_not_new_n1327__not_new_n1325_, not_new_n1327_, not_new_n1325_);
  or g_2860 (new_n4194_, not_new_n4173__0, not_new_n4109_);
  not g_2861 (not_new_n5949_, new_n5949_);
  or g_2862 (new_n4858_, not_new_n4763_, not_new_n1596__7);
  not g_2863 (not_new_n1053__6, new_n1053_);
  or g_2864 (new_n6185_, not_new_n1069__70, not_new_n5782__0);
  or g_2865 (po151, not_new_n3529_, not_new_n3528_);
  not g_2866 (not_new_n6451_, new_n6451_);
  and g_2867 (and_new_n3732__new_n3735_, new_n3735_, new_n3732_);
  or g_2868 (new_n5680_, not_new_n5464_, not_new_n5565_);
  or g_2869 (new_n5242_, not_new_n5000_, not_new_n5241_);
  not g_2870 (not_pi022, pi022);
  or g_2871 (new_n3545_, not_new_n1612__8, not_new_n1957__0);
  or g_2872 (new_n1699_, key_gate_20, not_new_n596__19773267430);
  or g_2873 (new_n4822_, not_new_n1041__7, not_new_n4813_);
  not g_2874 (not_new_n4157_, new_n4157_);
  not g_2875 (not_new_n3326_, new_n3326_);
  not g_2876 (new_n9708_, new_n9423_);
  not g_2877 (not_new_n1598__8235430, new_n1598_);
  or g_2878 (new_n5352_, not_new_n1600__9, not_new_n4953_);
  and g_2879 (new_n5872_, new_n6197_, new_n5916_);
  and g_2880 (new_n4779_, new_n4871_, new_n4870_);
  or g_2881 (new_n5140_, not_new_n4930__1, not_new_n4933__0);
  not g_2882 (not_pi045, pi045);
  not g_2883 (not_new_n1415_, new_n1415_);
  not g_2884 (not_pi174_0, pi174);
  not g_2885 (not_new_n607__2, new_n607_);
  not g_2886 (not_new_n5794__1, new_n5794_);
  or g_2887 (new_n3645_, not_new_n1611__332329305696010, not_new_n978_);
  or g_2888 (new_n3747_, not_new_n3746_, not_new_n3745_);
  not g_2889 (not_new_n647__113988951853731430, new_n647_);
  or g_2890 (new_n2842_, not_pi258, not_po296_6168735096280623662907561568153897267931784070);
  not g_2891 (not_new_n9755_, new_n9755_);
  xor g_2892 (key_gate_104, key_104, not_new_n3990_);
  not g_2893 (not_new_n9446_, new_n9446_);
  not g_2894 (not_new_n8236_, new_n8236_);
  or g_2895 (or_or_not_new_n3397__not_new_n3398__not_new_n1761_, or_not_new_n3397__not_new_n3398_, not_new_n1761_);
  not g_2896 (not_new_n6663__0, new_n6663_);
  or g_2897 (new_n10294_, not_new_n10156__0, not_new_n10292_);
  or g_2898 (new_n7199_, not_new_n7170_, not_new_n6983__0);
  or g_2899 (new_n7796_, not_new_n1049__8235430, not_new_n7598_);
  not g_2900 (not_new_n3017_, new_n3017_);
  not g_2901 (not_new_n2820_, new_n2820_);
  or g_2902 (new_n9511_, not_new_n1057__968890104070, not_new_n636__2326305139872070);
  not g_2903 (not_new_n7776_, new_n7776_);
  not g_2904 (not_new_n6412_, new_n6412_);
  not g_2905 (new_n6047_, new_n5797_);
  not g_2906 (not_new_n1067__1176490, new_n1067_);
  not g_2907 (new_n8849_, new_n617_);
  not g_2908 (not_new_n641__10, new_n641_);
  not g_2909 (not_new_n8266__2, new_n8266_);
  and g_2910 (new_n1301_, new_n2136_, new_n2137_);
  or g_2911 (new_n10212_, not_new_n9854__2, or_not_new_n10045__1_not_new_n9855__1);
  not g_2912 (not_new_n1031_, new_n1031_);
  or g_2913 (new_n3346_, not_new_n3920__0, not_pi064_24010);
  or g_2914 (new_n5633_, or_not_new_n5436__not_new_n5630__1, not_new_n5629_);
  not g_2915 (not_new_n2142_, new_n2142_);
  not g_2916 (not_new_n5042_, new_n5042_);
  not g_2917 (not_new_n10209_, new_n10209_);
  not g_2918 (not_new_n9149_, new_n9149_);
  not g_2919 (not_new_n620__3, new_n620_);
  or g_2920 (new_n9902_, not_new_n10068_, not_new_n10067_);
  not g_2921 (not_new_n9905_, new_n9905_);
  or g_2922 (new_n5345_, not_new_n1598__10, not_new_n4950__0);
  or g_2923 (new_n3088_, not_new_n648__5, not_new_n3315__2);
  not g_2924 (not_new_n8983__0, new_n8983_);
  not g_2925 (not_new_n710_, new_n710_);
  not g_2926 (not_new_n1895_, new_n1895_);
  not g_2927 (not_new_n6962_, new_n6962_);
  or g_2928 (new_n5858_, not_new_n6132_, not_new_n6131_);
  or g_2929 (new_n660_, not_new_n3138_, or_not_new_n3140__not_new_n3139_);
  not g_2930 (not_new_n619__19773267430, new_n619_);
  not g_2931 (not_new_n9135_, new_n9135_);
  or g_2932 (new_n2761_, not_new_n7063_, not_new_n595__2);
  or g_2933 (new_n5287_, or_not_new_n5203__not_new_n5087__0, not_new_n5079__0);
  not g_2934 (not_new_n2727_, new_n2727_);
  not g_2935 (not_new_n1566_, new_n1566_);
  not g_2936 (new_n7841_, new_n7756_);
  or g_2937 (new_n6439_, or_or_not_new_n6354__not_new_n6373__8_not_new_n6355_, not_new_n6233__2);
  not g_2938 (not_pi052_3, pi052);
  not g_2939 (not_new_n3204_, new_n3204_);
  or g_2940 (new_n3467_, not_pi019_0, not_new_n1536__332329305696010);
  not g_2941 (not_new_n6860_, new_n6860_);
  buf g_2942 (po011, pi204);
  not g_2943 (not_new_n8131_, new_n8131_);
  and g_2944 (new_n4297_, and_and_new_n4298__new_n4341__new_n4345_, new_n4342_);
  or g_2945 (new_n2424_, not_new_n9971__0, not_new_n599__3430);
  or g_2946 (new_n7153_, not_new_n7328_, not_new_n7000_);
  not g_2947 (not_new_n1594__168070, new_n1594_);
  not g_2948 (not_new_n4434__0, new_n4434_);
  or g_2949 (new_n4640_, not_new_n4639_, not_new_n4638_);
  not g_2950 (not_new_n1538__332329305696010, new_n1538_);
  or g_2951 (new_n966_, not_new_n2172_, or_or_not_new_n1311__not_new_n1309__not_new_n2173_);
  and g_2952 (new_n9332_, new_n9604_, new_n9603_);
  not g_2953 (not_new_n3520_, new_n3520_);
  or g_2954 (po087, not_new_n3381_, not_new_n3380_);
  not g_2955 (not_new_n1611__113988951853731430, new_n1611_);
  or g_2956 (new_n6193_, not_new_n5988_, not_new_n6192_);
  not g_2957 (not_pi267_0, pi267);
  not g_2958 (not_new_n625__332329305696010, new_n625_);
  not g_2959 (not_new_n3184__47475615099430, new_n3184_);
  not g_2960 (not_pi170_2, pi170);
  or g_2961 (new_n7200_, not_new_n7025__0, not_new_n742__0);
  or g_2962 (new_n3670_, not_new_n989__7, not_pi221);
  or g_2963 (new_n6156_, not_new_n5861_, not_new_n5892_);
  not g_2964 (not_new_n8817_, new_n8817_);
  not g_2965 (new_n4976_, new_n1069_);
  not g_2966 (not_new_n1603__3, new_n1603_);
  not g_2967 (not_new_n4816_, new_n4816_);
  or g_2968 (new_n7290_, not_new_n7288_, not_new_n7094_);
  or g_2969 (new_n9512_, not_new_n1599__138412872010, not_new_n622__332329305696010);
  or g_2970 (new_n6127_, not_new_n1607__8, not_new_n5885__0);
  or g_2971 (new_n751_, not_new_n3211_, not_new_n3210_);
  and g_2972 (new_n1220_, new_n1743_, and_new_n1745__new_n1744_);
  not g_2973 (not_new_n8194_, new_n8194_);
  not g_2974 (not_new_n1648_, key_gate_49);
  not g_2975 (not_new_n1538__797922662976120010, new_n1538_);
  not g_2976 (not_new_n9905__0, new_n9905_);
  not g_2977 (not_new_n5766_, new_n5766_);
  not g_2978 (not_new_n1608_, new_n1608_);
  not g_2979 (not_new_n8435_, new_n8435_);
  and g_2980 (and_new_n1222__new_n1223_, new_n1223_, new_n1222_);
  not g_2981 (not_new_n1612__113988951853731430, new_n1612_);
  not g_2982 (not_new_n591__47475615099430, new_n591_);
  not g_2983 (not_new_n5474_, new_n5474_);
  or g_2984 (new_n2082_, not_new_n6464_, not_new_n1580__1176490);
  not g_2985 (not_new_n4775__1, new_n4775_);
  or g_2986 (new_n2687_, not_new_n2686_, not_new_n611__19773267430);
  or g_2987 (new_n8056_, not_new_n7644__0, not_new_n643__6782230728490);
  or g_2988 (new_n8518_, not_new_n8517_, not_new_n8438_);
  not g_2989 (not_new_n601__1176490, new_n601_);
  and g_2990 (and_new_n9512__new_n9773_, new_n9773_, new_n9512_);
  not g_2991 (not_pi137, pi137);
  not g_2992 (not_new_n624__968890104070, new_n624_);
  not g_2993 (not_new_n1613__968890104070, new_n1613_);
  not g_2994 (not_new_n6812__0, new_n6812_);
  not g_2995 (not_new_n6463_, new_n6463_);
  not g_2996 (not_new_n1447_, new_n1447_);
  or g_2997 (new_n5548_, pi138, new_n1002_);
  and g_2998 (new_n9347_, new_n9559_, new_n9562_);
  not g_2999 (not_new_n5169_, new_n5169_);
  not g_3000 (not_pi264, pi264);
  not g_3001 (not_pi132, pi132);
  not g_3002 (not_new_n4840_, new_n4840_);
  or g_3003 (new_n2850_, not_new_n6969_, not_new_n595__490);
  or g_3004 (new_n1900_, not_new_n1252_, not_new_n1895_);
  not g_3005 (new_n6755_, new_n6629_);
  or g_3006 (new_n6416_, not_new_n620__6, not_new_n6248_);
  not g_3007 (not_new_n5824_, new_n5824_);
  not g_3008 (not_pi045_2, pi045);
  not g_3009 (not_new_n618__24010, new_n618_);
  or g_3010 (or_not_new_n1545__not_new_n1360_, not_new_n1545_, not_new_n1360_);
  or g_3011 (new_n1726_, key_gate_65, not_new_n596__797922662976120010);
  not g_3012 (not_new_n2956_, new_n2956_);
  not g_3013 (not_new_n8899_, new_n8899_);
  not g_3014 (not_new_n7073_, new_n7073_);
  and g_3015 (and_and_new_n2124__new_n2127__new_n2125_, and_new_n2124__new_n2127_, new_n2125_);
  or g_3016 (new_n2619_, not_po296_11044276742439206463052992010, not_pi266);
  not g_3017 (not_new_n4443_, new_n4443_);
  not g_3018 (not_new_n621__47475615099430, new_n621_);
  not g_3019 (not_new_n1792_, new_n1792_);
  not g_3020 (not_new_n2793_, new_n2793_);
  not g_3021 (not_new_n2073_, new_n2073_);
  not g_3022 (not_new_n647__490, new_n647_);
  or g_3023 (po168, not_new_n3563_, not_new_n3562_);
  not g_3024 (not_new_n1063__3430, new_n1063_);
  not g_3025 (not_new_n3970_, new_n3970_);
  not g_3026 (not_po296_5080218607396233653221881976522165017724345248360010, po296);
  not g_3027 (not_new_n4032__0, new_n4032_);
  or g_3028 (new_n3876_, not_new_n1576__968890104070, not_new_n638__490);
  not g_3029 (not_new_n7597__0, new_n7597_);
  or g_3030 (new_n4687_, not_new_n4685_, not_new_n4561_);
  not g_3031 (new_n7125_, new_n756_);
  or g_3032 (new_n2700_, not_new_n1020__0, not_new_n608__57648010);
  or g_3033 (new_n1783_, not_pi131, not_new_n587__0);
  not g_3034 (not_new_n3455_, new_n3455_);
  not g_3035 (not_new_n647__3430, new_n647_);
  not g_3036 (not_new_n621__9, new_n621_);
  not g_3037 (new_n2142_, new_n962_);
  or g_3038 (new_n4745_, or_not_new_n4837__not_new_n4772_, not_new_n4775_);
  or g_3039 (new_n3252_, not_new_n635__8, not_new_n3184__2);
  buf g_3040 (po009, pi202);
  not g_3041 (not_new_n1607__0, new_n1607_);
  not g_3042 (not_new_n1581_, new_n1581_);
  not g_3043 (not_new_n4114__2, new_n4114_);
  not g_3044 (not_new_n588__7, new_n588_);
  not g_3045 (not_new_n7412__1, new_n7412_);
  not g_3046 (not_new_n8124__0, new_n8124_);
  or g_3047 (new_n5013_, not_new_n5361_, not_new_n5362_);
  or g_3048 (new_n580_, not_new_n9921_, not_new_n1053_);
  not g_3049 (new_n7607_, new_n1037_);
  or g_3050 (new_n3556_, not_new_n1538__24010, not_pi144_0);
  not g_3051 (not_new_n618__1, new_n618_);
  or g_3052 (new_n6382_, not_new_n6223_, not_new_n6310_);
  not g_3053 (not_new_n1585__24010, new_n1585_);
  not g_3054 (not_new_n621__8, new_n621_);
  not g_3055 (not_new_n591__1, new_n591_);
  and g_3056 (and_new_n8724__new_n8726_, new_n8724_, new_n8726_);
  not g_3057 (not_new_n2926_, new_n2926_);
  and g_3058 (new_n1209_, new_n1718_, new_n1716_);
  not g_3059 (not_new_n581__32199057558131797268376070, new_n581_);
  not g_3060 (not_new_n3315__9, new_n3315_);
  or g_3061 (new_n6164_, not_new_n6020_, not_new_n5811__0);
  or g_3062 (po226, not_new_n1441_, not_new_n1440_);
  not g_3063 (not_new_n5483__0, new_n5483_);
  not g_3064 (not_new_n1596__2326305139872070, new_n1596_);
  not g_3065 (not_new_n2731_, new_n2731_);
  not g_3066 (not_new_n3203_, new_n3203_);
  not g_3067 (not_new_n1160_, new_n1160_);
  and g_3068 (and_and_new_n2327__new_n2328__new_n2331_, new_n2331_, and_new_n2327__new_n2328_);
  or g_3069 (or_not_new_n4829__not_new_n4794_, not_new_n4829_, not_new_n4794_);
  not g_3070 (not_new_n4899_, new_n4899_);
  not g_3071 (not_new_n1055__113988951853731430, new_n1055_);
  or g_3072 (new_n6841_, not_new_n6487__2, not_new_n1045__57648010);
  not g_3073 (not_new_n6635__3, new_n6635_);
  not g_3074 (not_new_n9955_, new_n9955_);
  not g_3075 (new_n8560_, new_n8236_);
  or g_3076 (new_n1901_, not_pi169, not_new_n586__7);
  not g_3077 (new_n4737_, new_n1039_);
  not g_3078 (not_new_n5219_, new_n5219_);
  not g_3079 (not_new_n727__1, new_n727_);
  and g_3080 (new_n8252_, new_n8498_, new_n8497_);
  or g_3081 (new_n2860_, not_po296_302268019717750559482470516839540966128657419430, not_pi260_0);
  not g_3082 (not_new_n3981__1, new_n3981_);
  not g_3083 (not_new_n9886_, new_n9886_);
  not g_3084 (not_new_n7454__2, new_n7454_);
  not g_3085 (not_new_n5055_, new_n5055_);
  not g_3086 (not_new_n607__3430, new_n607_);
  not g_3087 (not_new_n6753_, new_n6753_);
  or g_3088 (new_n3042_, not_new_n581__8235430, not_new_n1603__2);
  or g_3089 (or_not_new_n2565__not_new_n2564_, not_new_n2565_, not_new_n2564_);
  or g_3090 (new_n3313_, not_pi056_0, not_new_n1534__0);
  or g_3091 (new_n9520_, new_n1037_, new_n632_);
  or g_3092 (or_not_new_n1263__not_new_n1261_, not_new_n1261_, not_new_n1263_);
  not g_3093 (not_new_n6830_, new_n6830_);
  not g_3094 (not_new_n624__3, new_n624_);
  not g_3095 (not_new_n1443_, new_n1443_);
  not g_3096 (not_pi170_3, pi170);
  not g_3097 (new_n6999_, new_n735_);
  not g_3098 (not_new_n623_, new_n623_);
  or g_3099 (new_n9489_, or_not_new_n9694__not_new_n9634_, not_new_n9508_);
  or g_3100 (new_n9774_, not_new_n622__2326305139872070, not_new_n9417_);
  not g_3101 (not_new_n4788_, new_n4788_);
  not g_3102 (not_new_n5059__0, new_n5059_);
  not g_3103 (not_new_n1059__138412872010, new_n1059_);
  not g_3104 (new_n8167_, new_n1069_);
  or g_3105 (new_n3594_, not_pi163_0, not_new_n984__1);
  not g_3106 (not_new_n6221_, new_n6221_);
  or g_3107 (new_n8350_, not_new_n8164_, not_new_n1061__403536070);
  and g_3108 (new_n1489_, and_new_n2998__new_n998_, new_n2996_);
  or g_3109 (new_n2779_, not_new_n595__4, not_new_n7068_);
  or g_3110 (new_n3763_, not_new_n618__9, not_new_n1596__6);
  or g_3111 (new_n6099_, not_new_n6097_, not_new_n6098_);
  or g_3112 (new_n7165_, new_n775_, new_n745_);
  or g_3113 (new_n9919_, not_new_n648__39098210485829880490, not_new_n1049__16284135979104490);
  or g_3114 (new_n3839_, not_new_n6443__5, not_new_n4720_);
  not g_3115 (not_new_n613__2, new_n613_);
  not g_3116 (not_new_n1006_, new_n1006_);
  or g_3117 (new_n1674_, not_pi018, not_po296_3430);
  not g_3118 (not_new_n1045__8, new_n1045_);
  and g_3119 (and_new_n8692__new_n8691_, new_n8692_, new_n8691_);
  not g_3120 (not_new_n8640_, new_n8640_);
  or g_3121 (new_n8034_, not_new_n7638__0, not_new_n645__19773267430);
  not g_3122 (new_n6501_, new_n629_);
  not g_3123 (not_new_n10250_, new_n10250_);
  not g_3124 (not_new_n9452_, new_n9452_);
  buf g_3125 (po017, pi210);
  or g_3126 (new_n691_, not_new_n1512_, not_new_n3041_);
  or g_3127 (new_n3847_, not_new_n618__10, not_new_n6443__9);
  not g_3128 (not_new_n9905__1, new_n9905_);
  not g_3129 (not_new_n3109_, new_n3109_);
  not g_3130 (not_new_n1071__19773267430, new_n1071_);
  and g_3131 (po097, key_gate_101, pi076);
  or g_3132 (new_n3806_, not_new_n1037__6, not_new_n632__10);
  not g_3133 (not_new_n3546_, new_n3546_);
  not g_3134 (not_new_n5900__4, new_n5900_);
  not g_3135 (not_new_n4927_, new_n4927_);
  and g_3136 (new_n5040_, new_n5191_, new_n5283_);
  and g_3137 (new_n9465_, new_n9337_, new_n9592_);
  not g_3138 (not_new_n8113__0, new_n8113_);
  not g_3139 (new_n8645_, new_n1165_);
  not g_3140 (not_pi059, pi059);
  or g_3141 (new_n1753_, not_pi096, not_new_n1728__19773267430);
  not g_3142 (not_new_n6846_, new_n6846_);
  not g_3143 (not_new_n3299_, new_n3299_);
  or g_3144 (new_n4599_, not_new_n4475__0, not_new_n4474_);
  not g_3145 (not_new_n631__8235430, new_n631_);
  and g_3146 (new_n8955_, new_n8801_, new_n9152_);
  not g_3147 (not_new_n5963_, new_n5963_);
  not g_3148 (not_new_n1728__24010, new_n1728_);
  and g_3149 (and_new_n10047__new_n10048_, new_n10047_, new_n10048_);
  or g_3150 (new_n6109_, not_new_n5762__0, not_new_n5964_);
  not g_3151 (not_new_n10090_, new_n10090_);
  not g_3152 (not_new_n1201_, new_n1201_);
  and g_3153 (new_n5027_, and_new_n5268__new_n5267_, new_n5101_);
  not g_3154 (not_new_n4631_, new_n4631_);
  not g_3155 (not_new_n639__1, new_n639_);
  not g_3156 (not_new_n5829_, new_n5829_);
  not g_3157 (not_new_n598__8, new_n598_);
  not g_3158 (not_pi138_0, pi138);
  or g_3159 (new_n2325_, not_new_n1341_, not_new_n623_);
  not g_3160 (not_pi114_0, pi114);
  not g_3161 (not_new_n640_, new_n640_);
  not g_3162 (not_new_n5213_, new_n5213_);
  not g_3163 (not_new_n3048_, new_n3048_);
  and g_3164 (new_n7582_, new_n7828_, new_n7579_);
  not g_3165 (not_new_n9631_, new_n9631_);
  not g_3166 (not_new_n6634__2, new_n6634_);
  or g_3167 (new_n2084_, not_new_n1589__168070, not_new_n5017_);
  not g_3168 (not_new_n9888_, new_n9888_);
  not g_3169 (not_new_n642__1, new_n642_);
  not g_3170 (not_new_n7439_, new_n7439_);
  not g_3171 (new_n7742_, new_n619_);
  or g_3172 (or_not_new_n5184__not_new_n5183_, not_new_n5183_, not_new_n5184_);
  not g_3173 (not_new_n4048_, new_n4048_);
  not g_3174 (not_new_n4717_, new_n4717_);
  or g_3175 (new_n4028_, not_new_n4017__1, not_new_n3986_);
  or g_3176 (new_n3717_, not_new_n620__2, not_po298_5585458640832840070);
  not g_3177 (new_n8146_, new_n646_);
  not g_3178 (not_new_n4762__0, new_n4762_);
  not g_3179 (not_new_n5777_, new_n5777_);
  not g_3180 (not_new_n5383_, new_n5383_);
  or g_3181 (new_n2126_, not_new_n591__57648010, not_new_n4791_);
  not g_3182 (new_n9932_, new_n1602_);
  not g_3183 (not_new_n5878__0, new_n5878_);
  not g_3184 (not_new_n5271_, new_n5271_);
  and g_3185 (new_n8962_, new_n9231_, new_n9230_);
  or g_3186 (new_n5249_, not_new_n4944_, not_new_n5248_);
  not g_3187 (not_new_n8106__2, new_n8106_);
  not g_3188 (not_new_n3366_, new_n3366_);
  or g_3189 (new_n8058_, not_new_n7940_, not_new_n7758_);
  not g_3190 (not_new_n3288_, new_n3288_);
  not g_3191 (not_new_n679__0, new_n679_);
  or g_3192 (new_n9052_, new_n1057_, new_n636_);
  not g_3193 (not_new_n5789__0, new_n5789_);
  not g_3194 (not_new_n9805_, new_n9805_);
  or g_3195 (new_n10060_, not_new_n10059_, not_new_n10006_);
  or g_3196 (new_n720_, not_new_n3266_, not_new_n3265_);
  not g_3197 (not_new_n9352_, new_n9352_);
  not g_3198 (not_new_n5450__0, new_n5450_);
  not g_3199 (not_new_n6997_, new_n6997_);
  not g_3200 (not_new_n1601__7, new_n1601_);
  not g_3201 (not_new_n700_, new_n700_);
  not g_3202 (new_n10228_, new_n10029_);
  not g_3203 (not_new_n5027_, new_n5027_);
  not g_3204 (not_new_n9119__0, new_n9119_);
  not g_3205 (not_new_n1545_, new_n1545_);
  not g_3206 (not_new_n5887_, new_n5887_);
  or g_3207 (new_n7482_, not_new_n7480_, not_new_n7481_);
  not g_3208 (not_new_n603__3, new_n603_);
  not g_3209 (not_new_n7041__1, new_n7041_);
  not g_3210 (not_new_n1849_, new_n1849_);
  not g_3211 (not_new_n5786__0, new_n5786_);
  not g_3212 (not_new_n638__13410686196639649008070, new_n638_);
  not g_3213 (not_new_n6169_, new_n6169_);
  not g_3214 (not_new_n601__10, new_n601_);
  not g_3215 (new_n2019_, new_n643_);
  not g_3216 (new_n6484_, new_n1031_);
  or g_3217 (new_n7297_, not_new_n7293_, not_new_n7159_);
  not g_3218 (not_new_n7418__1, new_n7418_);
  not g_3219 (not_new_n618__6782230728490, new_n618_);
  not g_3220 (not_new_n8324_, new_n8324_);
  not g_3221 (not_new_n3917__0, key_gate_70);
  not g_3222 (not_po298_797922662976120010, po298);
  not g_3223 (new_n10214_, new_n9948_);
  not g_3224 (not_new_n3396_, new_n3396_);
  or g_3225 (new_n9693_, not_new_n9394__0, not_new_n9584__0);
  not g_3226 (not_new_n5014_, new_n5014_);
  not g_3227 (not_new_n1900_, new_n1900_);
  not g_3228 (not_new_n629__168070, new_n629_);
  not g_3229 (new_n8278_, new_n8169_);
  not g_3230 (not_po298_70, po298);
  not g_3231 (new_n9943_, new_n1597_);
  not g_3232 (not_new_n3315__24010, new_n3315_);
  or g_3233 (or_not_new_n4291__not_new_n4326_, not_new_n4291_, not_new_n4326_);
  and g_3234 (new_n4410_, new_n4585_, new_n4581_);
  or g_3235 (new_n6014_, not_new_n617__1176490, not_new_n5912_);
  not g_3236 (not_new_n3140_, new_n3140_);
  or g_3237 (new_n5654_, not_new_n1011__8, not_new_n5472__0);
  or g_3238 (new_n9110_, new_n1599_, new_n622_);
  not g_3239 (not_new_n3727_, new_n3727_);
  or g_3240 (new_n5576_, new_n1012_, pi146);
  and g_3241 (and_and_and_new_n1043__new_n6232__new_n6229__new_n6317_, and_and_new_n1043__new_n6232__new_n6229_, new_n6317_);
  not g_3242 (not_new_n6974__1176490, new_n6974_);
  or g_3243 (new_n4740_, not_new_n4802_, or_not_new_n4827__not_new_n4799_);
  not g_3244 (not_new_n7430__2, new_n7430_);
  or g_3245 (new_n6900_, not_new_n625__138412872010, not_new_n6507__1);
  or g_3246 (new_n3377_, or_not_pi245_0_not_new_n1625_, not_new_n3318__1);
  or g_3247 (new_n1798_, not_new_n8901_, not_new_n1591__0);
  or g_3248 (new_n4181_, not_new_n4145_, not_pi274_2);
  not g_3249 (not_new_n9546_, new_n9546_);
  not g_3250 (not_new_n1028__7, new_n1028_);
  not g_3251 (not_new_n9978_, new_n9978_);
  not g_3252 (not_new_n1616__490, new_n1616_);
  or g_3253 (new_n2284_, not_new_n585__2326305139872070, not_new_n4119_);
  not g_3254 (not_new_n7007__1, new_n7007_);
  or g_3255 (new_n8771_, not_new_n8594_, not_new_n8686_);
  not g_3256 (not_new_n1178_, new_n1178_);
  not g_3257 (not_new_n1581__10, new_n1581_);
  or g_3258 (new_n1951_, not_new_n1589__8, not_new_n5003_);
  or g_3259 (new_n6908_, not_new_n6512__0, not_new_n640__403536070);
  not g_3260 (not_new_n5895_, new_n5895_);
  not g_3261 (not_new_n6361_, new_n6361_);
  not g_3262 (not_new_n6871_, new_n6871_);
  and g_3263 (new_n9333_, new_n9332_, new_n9605_);
  and g_3264 (and_and_new_n6244__new_n6372__new_n1596_, new_n1596_, and_new_n6244__new_n6372_);
  not g_3265 (not_new_n624__24010, new_n624_);
  not g_3266 (not_new_n3874_, new_n3874_);
  not g_3267 (not_new_n3213_, new_n3213_);
  not g_3268 (not_new_n641__19773267430, new_n641_);
  not g_3269 (not_new_n10019_, new_n10019_);
  not g_3270 (not_pi125_0, pi125);
  not g_3271 (not_new_n4091_, new_n4091_);
  or g_3272 (new_n7806_, not_new_n7700_, not_new_n7805_);
  or g_3273 (new_n3021_, not_new_n581__10, not_new_n1596__2);
  not g_3274 (not_new_n8445_, new_n8445_);
  and g_3275 (new_n3932_, new_n4002_, new_n4008_);
  or g_3276 (new_n10071_, not_new_n9902_, not_new_n10041_);
  not g_3277 (not_new_n4155__1, new_n4155_);
  not g_3278 (not_new_n8852_, new_n8852_);
  or g_3279 (new_n2830_, not_new_n4118__2, not_new_n3310__6);
  or g_3280 (new_n4371_, not_new_n4265_, not_new_n660_);
  not g_3281 (not_new_n1591__24010, new_n1591_);
  or g_3282 (new_n4650_, not_new_n1028__10, not_new_n4491__0);
  not g_3283 (not_new_n7018_, new_n7018_);
  xnor g_3284 (key_gate_74, key_74, not_new_n1723_);
  and g_3285 (and_new_n3061__new_n998_, new_n998_, new_n3061_);
  not g_3286 (not_pi134_3, pi134);
  or g_3287 (new_n7278_, not_new_n7439__0, not_new_n7004__0);
  not g_3288 (new_n4249_, new_n669_);
  or g_3289 (new_n6490_, not_new_n6477_, not_new_n624__57648010);
  not g_3290 (not_new_n9510__0, new_n9510_);
  not g_3291 (not_new_n7813_, new_n7813_);
  or g_3292 (new_n4359_, not_new_n664_, not_new_n4257_);
  or g_3293 (new_n9219_, not_new_n9158_, not_new_n8957_);
  not g_3294 (not_new_n1850_, new_n1850_);
  not g_3295 (not_new_n624_, new_n624_);
  or g_3296 (new_n7265_, not_new_n7045__0, not_new_n718__0);
  not g_3297 (new_n7170_, new_n6991_);
  not g_3298 (new_n4257_, new_n696_);
  not g_3299 (not_new_n8280_, new_n8280_);
  or g_3300 (new_n3307_, not_new_n5733__0, not_new_n1585__113988951853731430);
  or g_3301 (new_n3659_, not_new_n632__9, not_po298_2);
  not g_3302 (not_new_n627__490, new_n627_);
  not g_3303 (not_new_n7735__3, new_n7735_);
  or g_3304 (new_n8399_, not_new_n638__5585458640832840070, not_new_n8150__1);
  or g_3305 (new_n8390_, not_new_n8139__0, not_new_n8368__0);
  not g_3306 (not_new_n5414_, new_n5414_);
  or g_3307 (new_n760_, not_new_n3231_, not_new_n3230_);
  not g_3308 (not_new_n1163__0, new_n1163_);
  or g_3309 (new_n4063_, not_new_n3948_, not_pi053_3);
  not g_3310 (not_new_n631__968890104070, new_n631_);
  not g_3311 (new_n7932_, new_n7666_);
  not g_3312 (not_new_n9743_, new_n9743_);
  not g_3313 (not_new_n10132_, new_n10132_);
  not g_3314 (not_new_n6538_, new_n6538_);
  not g_3315 (not_new_n6475__0, new_n6475_);
  not g_3316 (not_new_n9471_, new_n9471_);
  not g_3317 (not_new_n1315_, new_n1315_);
  or g_3318 (new_n5691_, not_new_n1017__6, not_new_n5457_);
  not g_3319 (not_new_n8166_, new_n8166_);
  not g_3320 (not_pi133, pi133);
  not g_3321 (not_new_n10066_, new_n10066_);
  or g_3322 (new_n2574_, not_new_n1017_, not_new_n607__4);
  not g_3323 (not_new_n3968_, new_n3968_);
  or g_3324 (new_n2377_, not_new_n603__4, not_new_n635__1);
  or g_3325 (new_n5404_, not_new_n1061__70, not_new_n4970_);
  or g_3326 (or_or_not_new_n2208__not_new_n2205__not_new_n2206_, or_not_new_n2208__not_new_n2205_, not_new_n2206_);
  not g_3327 (not_new_n3508_, new_n3508_);
  not g_3328 (not_new_n1049__490, new_n1049_);
  not g_3329 (not_new_n645__490, new_n645_);
  or g_3330 (new_n1652_, not_new_n1631__5, not_pi039);
  not g_3331 (not_new_n6271_, new_n6271_);
  not g_3332 (not_pi269, pi269);
  not g_3333 (not_new_n1457_, new_n1457_);
  not g_3334 (not_new_n1008__2, new_n1008_);
  or g_3335 (new_n3422_, not_new_n1536__8235430, not_pi028_0);
  not g_3336 (new_n7601_, new_n1041_);
  not g_3337 (not_new_n1063__10, new_n1063_);
  not g_3338 (not_pi270_1, pi270);
  not g_3339 (not_new_n5749__1, new_n5749_);
  not g_3340 (not_new_n1047__968890104070, new_n1047_);
  not g_3341 (not_new_n6886_, new_n6886_);
  not g_3342 (not_new_n1768_, new_n1768_);
  and g_3343 (new_n8700_, new_n8597_, new_n8782_);
  not g_3344 (not_new_n5297_, new_n5297_);
  not g_3345 (not_pi064, pi064);
  not g_3346 (not_new_n3387__1, new_n3387_);
  not g_3347 (not_new_n3836_, new_n3836_);
  not g_3348 (not_pi257, pi257);
  not g_3349 (not_new_n603__332329305696010, new_n603_);
  or g_3350 (new_n7050_, not_new_n7381_, not_new_n7382_);
  or g_3351 (new_n1764_, not_pi130, not_new_n587_);
  or g_3352 (new_n9199_, not_new_n9198_, not_new_n9197_);
  not g_3353 (not_pi109_0, pi109);
  not g_3354 (not_new_n8179_, new_n8179_);
  not g_3355 (not_new_n2509__8235430, new_n2509_);
  not g_3356 (not_new_n3924__0, new_n3924_);
  not g_3357 (not_new_n6306_, new_n6306_);
  not g_3358 (not_new_n5096__0, new_n5096_);
  or g_3359 (new_n1730_, not_new_n925__0, not_new_n3324__0);
  not g_3360 (new_n6660_, new_n6528_);
  or g_3361 (new_n6428_, not_new_n6233__0, or_or_not_new_n6340__not_new_n6341__not_new_n6342_);
  not g_3362 (not_new_n7314_, new_n7314_);
  not g_3363 (not_new_n9763_, new_n9763_);
  and g_3364 (and_new_n2662__new_n2661_, new_n2661_, new_n2662_);
  and g_3365 (new_n5029_, new_n5119_, new_n4900_);
  not g_3366 (not_new_n589__5585458640832840070, new_n589_);
  not g_3367 (not_new_n8286__1, new_n8286_);
  or g_3368 (new_n7022_, not_new_n7359_, not_new_n7358_);
  not g_3369 (new_n7409_, new_n7032_);
  not g_3370 (not_new_n628__0, new_n628_);
  and g_3371 (new_n3929_, new_n3938_, new_n4021_);
  not g_3372 (not_new_n4825__1, new_n4825_);
  and g_3373 (new_n1545_, new_n3603_, new_n3602_);
  not g_3374 (not_pi138_2, pi138);
  or g_3375 (new_n4579_, not_new_n4451_, not_new_n4578_);
  or g_3376 (new_n2213_, not_new_n9441_, not_new_n1584__138412872010);
  not g_3377 (not_new_n4954__0, new_n4954_);
  not g_3378 (not_new_n1059__24010, new_n1059_);
  and g_3379 (new_n8800_, new_n9004_, new_n9003_);
  or g_3380 (new_n4626_, not_new_n4625_, not_new_n4624_);
  not g_3381 (not_new_n3578_, new_n3578_);
  not g_3382 (not_new_n7177_, new_n7177_);
  or g_3383 (new_n7176_, not_new_n6960_, not_new_n6991_);
  or g_3384 (new_n4368_, not_new_n4263_, not_new_n693_);
  not g_3385 (not_new_n9177_, new_n9177_);
  not g_3386 (not_new_n5893_, new_n5893_);
  not g_3387 (not_new_n8996_, new_n8996_);
  not g_3388 (not_new_n3356_, new_n3356_);
  not g_3389 (not_new_n7058_, new_n7058_);
  or g_3390 (new_n3099_, not_new_n581__93874803376477543056490, not_new_n631__6);
  not g_3391 (not_new_n8118_, new_n8118_);
  not g_3392 (not_new_n10312_, new_n10312_);
  not g_3393 (not_new_n8866_, new_n8866_);
  not g_3394 (not_pi187_0, pi187);
  not g_3395 (not_new_n989__2, new_n989_);
  not g_3396 (not_new_n581__7, new_n581_);
  or g_3397 (new_n1821_, not_new_n628_, not_new_n593__1);
  not g_3398 (not_new_n1010_, new_n1010_);
  and g_3399 (new_n9477_, new_n9332_, new_n9655_);
  not g_3400 (not_new_n6584_, new_n6584_);
  not g_3401 (not_new_n9516_, new_n9516_);
  not g_3402 (not_new_n5109_, new_n5109_);
  or g_3403 (new_n1757_, not_new_n1728__47475615099430, not_pi071);
  not g_3404 (not_new_n627__8235430, new_n627_);
  not g_3405 (not_new_n6443__5, new_n6443_);
  not g_3406 (not_new_n8126_, new_n8126_);
  or g_3407 (new_n3079_, not_new_n3372__273687473400809163430, not_new_n626__4);
  not g_3408 (not_new_n1605__5, new_n1605_);
  not g_3409 (not_new_n595__332329305696010, new_n595_);
  and g_3410 (new_n7071_, new_n7174_, new_n7175_);
  not g_3411 (not_new_n2265_, new_n2265_);
  not g_3412 (not_new_n646__5, new_n646_);
  not g_3413 (not_new_n1600__3430, new_n1600_);
  not g_3414 (not_new_n7082_, new_n7082_);
  and g_3415 (new_n8960_, new_n9224_, new_n9223_);
  not g_3416 (not_new_n7487_, new_n7487_);
  not g_3417 (not_new_n8266__1, new_n8266_);
  not g_3418 (not_new_n8000_, new_n8000_);
  not g_3419 (not_new_n1045__2326305139872070, new_n1045_);
  or g_3420 (new_n4648_, not_new_n1028__9, not_new_n4491_);
  not g_3421 (new_n1574_, new_n8598_);
  not g_3422 (not_new_n9597_, new_n9597_);
  not g_3423 (not_new_n2857_, new_n2857_);
  not g_3424 (not_new_n5567_, new_n5567_);
  not g_3425 (not_new_n622__10, new_n622_);
  or g_3426 (new_n3597_, not_new_n1611__2, not_new_n946_);
  or g_3427 (new_n6669_, not_new_n635__57648010, not_new_n6476_);
  or g_3428 (new_n2561_, not_new_n5488__0, not_new_n606__4);
  not g_3429 (not_new_n8857_, new_n8857_);
  not g_3430 (not_new_n989__113988951853731430, new_n989_);
  not g_3431 (not_new_n8978__0, new_n8978_);
  or g_3432 (new_n3168_, not_new_n1055__3, not_new_n928__2326305139872070);
  not g_3433 (not_new_n8140_, new_n8140_);
  or g_3434 (new_n9419_, or_not_new_n9719__not_new_n9718_, not_new_n9628_);
  and g_3435 (and_and_new_n2276__new_n2279__new_n2277_, and_new_n2276__new_n2279_, new_n2277_);
  not g_3436 (not_new_n8878__0, new_n8878_);
  or g_3437 (new_n1711_, not_new_n596__47475615099430, key_gate_7);
  not g_3438 (new_n8892_, new_n618_);
  or g_3439 (new_n8388_, not_new_n625__16284135979104490, not_new_n8138__0);
  not g_3440 (not_new_n8451_, new_n8451_);
  not g_3441 (not_new_n9182_, new_n9182_);
  and g_3442 (and_new_n6374__new_n6372_, new_n6372_, new_n6374_);
  and g_3443 (new_n1433_, new_n2590_, new_n2592_);
  not g_3444 (not_new_n1071__5, new_n1071_);
  or g_3445 (new_n6852_, not_new_n1039__1176490, not_new_n6482__1);
  not g_3446 (not_new_n1039__47475615099430, new_n1039_);
  not g_3447 (new_n8643_, new_n1167_);
  and g_3448 (and_new_n9915__new_n10334_, new_n9915_, new_n10334_);
  or g_3449 (new_n7186_, not_new_n738_, not_new_n7183_);
  not g_3450 (not_new_n4415__0, new_n4415_);
  or g_3451 (new_n6039_, not_new_n626__403536070, not_new_n5794__1);
  not g_3452 (not_new_n1669_, key_gate_13);
  not g_3453 (not_new_n4967_, new_n4967_);
  not g_3454 (not_new_n933__0, new_n933_);
  not g_3455 (new_n6521_, new_n644_);
  or g_3456 (or_not_new_n4228__not_new_n4329_, not_new_n4228_, not_new_n4329_);
  not g_3457 (not_new_n7664_, new_n7664_);
  not g_3458 (not_new_n1023__1, new_n1023_);
  and g_3459 (new_n9987_, new_n9863_, new_n9856_);
  not g_3460 (not_new_n606__7, new_n606_);
  not g_3461 (not_new_n10195_, new_n10195_);
  not g_3462 (new_n8105_, new_n648_);
  or g_3463 (new_n7960_, not_new_n7795__0, not_new_n7736_);
  not g_3464 (new_n5788_, new_n644_);
  or g_3465 (new_n9819_, not_new_n9409_, not_new_n637__2326305139872070);
  not g_3466 (not_new_n7836_, new_n7836_);
  not g_3467 (not_new_n6482_, new_n6482_);
  not g_3468 (not_new_n1049__6, new_n1049_);
  not g_3469 (new_n4166_, new_n4094_);
  or g_3470 (new_n4608_, not_new_n4425_, not_new_n1005__3);
  not g_3471 (not_new_n627__47475615099430, new_n627_);
  not g_3472 (not_new_n1596__8, new_n1596_);
  not g_3473 (not_new_n8608_, new_n8608_);
  xor g_3474 (key_gate_32, not_new_n3982_, key_32);
  not g_3475 (not_new_n3151_, new_n3151_);
  not g_3476 (not_new_n8035_, new_n8035_);
  not g_3477 (not_new_n1020__6, new_n1020_);
  not g_3478 (not_new_n581__52433383167563036344614587188619514555430, new_n581_);
  or g_3479 (new_n5958_, not_new_n5957_, not_new_n5956_);
  not g_3480 (not_new_n2981_, new_n2981_);
  not g_3481 (not_new_n9506__3, new_n9506_);
  not g_3482 (not_new_n6847_, new_n6847_);
  not g_3483 (not_new_n8139_, new_n8139_);
  or g_3484 (new_n986_, or_not_new_n1024__2_not_new_n1028__3, not_new_n3387__2);
  or g_3485 (new_n7996_, not_new_n7622__1, not_new_n617__47475615099430);
  not g_3486 (new_n9944_, new_n617_);
  or g_3487 (new_n7557_, not_new_n7329_, not_new_n7555_);
  or g_3488 (new_n9628_, new_n621_, new_n1598_);
  or g_3489 (or_or_not_new_n8609__not_new_n8595__0_not_new_n1168__0, or_not_new_n8609__not_new_n8595__0, not_new_n1168__0);
  not g_3490 (not_pi039_3, pi039);
  not g_3491 (new_n4268_, new_n658_);
  not g_3492 (not_new_n3660_, new_n3660_);
  not g_3493 (not_new_n1597__113988951853731430, new_n1597_);
  not g_3494 (not_new_n7571_, new_n7571_);
  not g_3495 (not_new_n8739_, new_n8739_);
  or g_3496 (new_n10135_, new_n630_, new_n1601_);
  or g_3497 (new_n4463_, not_new_n4673_, not_new_n4672_);
  not g_3498 (not_new_n4032_, new_n4032_);
  or g_3499 (new_n2390_, not_new_n598__6, not_new_n1047__0);
  not g_3500 (not_new_n4013__0, new_n4013_);
  or g_3501 (new_n7023_, not_new_n7341_, not_new_n7340_);
  not g_3502 (not_new_n618_, new_n618_);
  or g_3503 (po220, or_or_not_new_n2567__not_new_n2571__not_new_n1429_, not_new_n1428_);
  or g_3504 (or_not_new_n1565__not_new_n2484_, not_new_n2484_, not_new_n1565_);
  or g_3505 (or_not_new_n4246__not_new_n4350_, not_new_n4350_, not_new_n4246_);
  and g_3506 (new_n4753_, new_n4850_, new_n4851_);
  xnor g_3507 (key_gate_64, not_new_n1666_, key_64);
  or g_3508 (new_n4015_, not_new_n3953_, not_new_n4014__3);
  or g_3509 (new_n6018_, not_new_n5770__1, not_new_n1601__3430);
  not g_3510 (not_new_n3310__9, new_n3310_);
  or g_3511 (new_n2746_, not_new_n634__2, not_new_n602__1);
  not g_3512 (not_new_n6505__0, new_n6505_);
  not g_3513 (not_new_n1979_, new_n1979_);
  not g_3514 (not_new_n6443__19773267430, new_n6443_);
  not g_3515 (new_n5885_, new_n619_);
  not g_3516 (not_new_n8392__0, new_n8392_);
  or g_3517 (new_n7537_, not_new_n7149_, not_new_n7150__0);
  or g_3518 (or_not_new_n2346__not_new_n2347_, not_new_n2347_, not_new_n2346_);
  or g_3519 (new_n2692_, not_new_n2509__8235430, not_pi211);
  not g_3520 (not_new_n4998__0, new_n4998_);
  or g_3521 (new_n7435_, not_new_n6974__403536070, not_new_n753_);
  not g_3522 (not_new_n3184__2, new_n3184_);
  not g_3523 (not_new_n1043__3430, new_n1043_);
  or g_3524 (new_n4522_, new_n1007_, pi165);
  or g_3525 (or_not_new_n1882__not_new_n1883_, not_new_n1882_, not_new_n1883_);
  or g_3526 (new_n2106_, not_new_n593__1176490, not_new_n646_);
  or g_3527 (new_n9073_, not_new_n8803_, not_new_n8899_);
  and g_3528 (new_n1444_, and_new_n2647__new_n2648_, new_n2649_);
  and g_3529 (new_n9346_, new_n9567_, new_n9570_);
  not g_3530 (not_new_n10045_, new_n10045_);
  or g_3531 (new_n1984_, not_new_n1585__10, not_new_n5730_);
  not g_3532 (not_new_n7877_, new_n7877_);
  not g_3533 (new_n7014_, new_n718_);
  or g_3534 (new_n9667_, not_new_n9506__0, not_new_n9584_);
  not g_3535 (not_new_n4172_, new_n4172_);
  not g_3536 (not_new_n1065__0, new_n1065_);
  not g_3537 (not_new_n9356__0, new_n9356_);
  not g_3538 (not_new_n7057_, new_n7057_);
  not g_3539 (not_new_n4704_, new_n4704_);
  or g_3540 (new_n5542_, not_new_n5498_, not_new_n5541_);
  not g_3541 (not_new_n6791_, new_n6791_);
  not g_3542 (not_new_n6617_, new_n6617_);
  or g_3543 (new_n7109_, not_new_n7073_, not_new_n7324_);
  not g_3544 (not_new_n581__168070, new_n581_);
  not g_3545 (new_n9907_, new_n1069_);
  not g_3546 (not_new_n1596__5, new_n1596_);
  or g_3547 (new_n5134_, not_new_n5132_, not_new_n5032_);
  not g_3548 (not_new_n4999__3, new_n4999_);
  not g_3549 (not_new_n6942_, new_n6942_);
  not g_3550 (not_new_n5124_, new_n5124_);
  not g_3551 (not_new_n5901__0, new_n5901_);
  not g_3552 (not_new_n4274_, new_n4274_);
  or g_3553 (new_n934_, not_new_n1623__0, not_new_n3384__0);
  not g_3554 (not_pi064_3, pi064);
  or g_3555 (new_n2709_, or_not_new_n1469__not_new_n3820_, not_new_n3819_);
  and g_3556 (new_n1430_, new_n2578_, new_n2579_);
  or g_3557 (new_n5655_, not_pi147_4, not_new_n5473__0);
  not g_3558 (not_new_n1243_, new_n1243_);
  not g_3559 (not_new_n624__7, new_n624_);
  not g_3560 (new_n8722_, new_n8625_);
  not g_3561 (not_new_n5573_, new_n5573_);
  not g_3562 (not_new_n4833_, new_n4833_);
  or g_3563 (new_n5373_, not_new_n4980__0, not_new_n1603__10);
  not g_3564 (not_new_n633__8235430, new_n633_);
  or g_3565 (new_n2107_, not_new_n591__8235430, not_new_n4793_);
  not g_3566 (not_new_n8133_, new_n8133_);
  or g_3567 (new_n1660_, not_new_n596__8, key_gate_93);
  or g_3568 (new_n4376_, not_new_n659_, not_new_n4266_);
  not g_3569 (not_new_n3495_, new_n3495_);
  not g_3570 (not_new_n5332_, new_n5332_);
  or g_3571 (or_not_new_n3134__not_new_n3133_, not_new_n3133_, not_new_n3134_);
  not g_3572 (not_new_n1580__6782230728490, new_n1580_);
  and g_3573 (new_n6611_, new_n6955_, new_n6650_);
  not g_3574 (new_n4284_, new_n650_);
  not g_3575 (not_new_n5071_, new_n5071_);
  not g_3576 (not_new_n1604__6, new_n1604_);
  not g_3577 (not_po296_2115876138024253916377293617876786762900601936010, po296);
  or g_3578 (new_n9086_, new_n1069_, new_n646_);
  not g_3579 (not_new_n2962_, new_n2962_);
  or g_3580 (new_n2877_, not_new_n7056_, not_new_n595__168070);
  and g_3581 (new_n595_, new_n1595_, new_n1475_);
  or g_3582 (new_n2802_, or_not_new_n2801__not_new_n2800_, not_new_n2799_);
  not g_3583 (not_new_n626__5585458640832840070, new_n626_);
  not g_3584 (not_new_n4923_, new_n4923_);
  or g_3585 (new_n5133_, not_new_n631__24010, not_new_n1043__9);
  not g_3586 (not_new_n7276_, new_n7276_);
  not g_3587 (not_new_n9081_, new_n9081_);
  not g_3588 (not_new_n612__5, new_n612_);
  not g_3589 (not_new_n934_, new_n934_);
  not g_3590 (not_new_n637__403536070, new_n637_);
  not g_3591 (not_new_n6876_, new_n6876_);
  or g_3592 (new_n8440_, not_new_n8215_, not_new_n8266__4);
  not g_3593 (not_new_n597__113988951853731430, new_n597_);
  not g_3594 (not_new_n3185__2, new_n3185_);
  or g_3595 (new_n5658_, not_new_n5579__0, not_new_n5656_);
  or g_3596 (new_n2832_, not_new_n595__10, not_new_n7052_);
  not g_3597 (not_new_n7633__0, new_n7633_);
  not g_3598 (not_new_n4439__0, new_n4439_);
  not g_3599 (not_new_n622__332329305696010, new_n622_);
  not g_3600 (not_new_n5896_, new_n5896_);
  or g_3601 (new_n2665_, not_new_n5482_, not_new_n605__168070);
  not g_3602 (not_new_n625__13410686196639649008070, new_n625_);
  not g_3603 (not_new_n999__0, new_n999_);
  or g_3604 (new_n5711_, not_new_n5428_, not_new_n1020__7);
  not g_3605 (not_new_n7560_, new_n7560_);
  or g_3606 (new_n3878_, not_new_n1576__6782230728490, not_new_n643__490);
  or g_3607 (new_n9813_, not_new_n1069__968890104070, not_new_n9405_);
  or g_3608 (new_n9035_, new_n624_, new_n1041_);
  not g_3609 (not_new_n1059__8235430, new_n1059_);
  not g_3610 (not_pi049_0, pi049);
  not g_3611 (not_new_n599_, new_n599_);
  not g_3612 (not_pi064_403536070, pi064);
  not g_3613 (not_new_n9775_, new_n9775_);
  not g_3614 (not_new_n8168__0, new_n8168_);
  not g_3615 (not_new_n9953_, new_n9953_);
  not g_3616 (not_po296_2569235775210588780886114772242356213216070, po296);
  not g_3617 (not_new_n5455_, new_n5455_);
  or g_3618 (new_n9083_, not_new_n8986_, not_new_n8805_);
  not g_3619 (not_new_n6614_, new_n6614_);
  or g_3620 (new_n8616_, not_new_n8738_, not_new_n8737_);
  or g_3621 (new_n8956_, not_new_n9009_, not_new_n9169_);
  not g_3622 (not_new_n928__2, new_n928_);
  not g_3623 (not_pi214, pi214);
  and g_3624 (new_n7698_, new_n7799_, new_n7798_);
  or g_3625 (new_n6859_, not_new_n6702_, not_new_n6496__1);
  not g_3626 (not_new_n1280_, new_n1280_);
  not g_3627 (not_new_n9749_, new_n9749_);
  not g_3628 (not_new_n602__24010, new_n602_);
  not g_3629 (not_new_n7316_, new_n7316_);
  not g_3630 (new_n8857_, new_n1063_);
  not g_3631 (not_new_n671_, new_n671_);
  not g_3632 (new_n4263_, new_n661_);
  not g_3633 (not_new_n9969_, new_n9969_);
  not g_3634 (not_new_n1594__24010, new_n1594_);
  not g_3635 (not_new_n2577_, new_n2577_);
  not g_3636 (not_new_n3790_, new_n3790_);
  not g_3637 (not_new_n1603__4, new_n1603_);
  not g_3638 (not_new_n4125__2, new_n4125_);
  or g_3639 (new_n8524_, not_new_n8226_, not_new_n8258_);
  or g_3640 (new_n5256_, not_new_n4937__1, not_new_n5121_);
  not g_3641 (not_pi013, pi013);
  or g_3642 (new_n7391_, not_new_n7023__0, not_new_n6981__0);
  not g_3643 (not_new_n9392_, new_n9392_);
  or g_3644 (new_n2430_, not_new_n598__24010, not_new_n1063__0);
  not g_3645 (new_n8158_, new_n1053_);
  or g_3646 (new_n3201_, not_new_n618__6, not_new_n589__6);
  and g_3647 (new_n6577_, new_n6696_, new_n6445_);
  not g_3648 (not_new_n581__9095436801298611408202050198891430, new_n581_);
  or g_3649 (or_not_new_n2818__not_new_n2817_, not_new_n2817_, not_new_n2818_);
  not g_3650 (not_new_n6242__5, new_n6242_);
  not g_3651 (not_new_n4017_, new_n4017_);
  not g_3652 (not_new_n3320_, new_n3320_);
  not g_3653 (new_n7103_, new_n771_);
  not g_3654 (not_new_n6974__7, new_n6974_);
  not g_3655 (not_new_n6974__0, new_n6974_);
  or g_3656 (new_n5795_, not_new_n647__168070, not_new_n5759_);
  or g_3657 (new_n9645_, not_new_n9614_, not_new_n9501_);
  not g_3658 (not_new_n8603_, new_n8603_);
  not g_3659 (not_new_n3372__2326305139872070, new_n3372_);
  not g_3660 (not_new_n4414_, new_n4414_);
  not g_3661 (not_new_n6022_, new_n6022_);
  not g_3662 (not_new_n640__332329305696010, new_n640_);
  not g_3663 (new_n9060_, new_n8977_);
  not g_3664 (not_pi148_1, pi148);
  not g_3665 (not_new_n1588__1176490, new_n1588_);
  or g_3666 (new_n2837_, not_new_n2834_, or_not_new_n2836__not_new_n2835_);
  not g_3667 (not_pi256, pi256);
  not g_3668 (not_new_n4789__0, new_n4789_);
  not g_3669 (not_new_n6894_, new_n6894_);
  or g_3670 (new_n7689_, not_new_n8001_, not_new_n8000_);
  not g_3671 (not_new_n9578_, new_n9578_);
  not g_3672 (not_pi037_0, pi037);
  or g_3673 (new_n9193_, not_new_n8842_, not_new_n1051__19773267430);
  and g_3674 (new_n8206_, and_new_n8104__new_n8464_, new_n8463_);
  not g_3675 (not_new_n605__9, new_n605_);
  or g_3676 (new_n2013_, not_new_n1588__490, not_new_n1057_);
  not g_3677 (not_new_n1588__47475615099430, new_n1588_);
  or g_3678 (new_n5002_, not_new_n5424_, not_new_n5425_);
  and g_3679 (and_new_n2295__new_n2298_, new_n2298_, new_n2295_);
  or g_3680 (new_n2007_, not_new_n8920_, not_new_n1591__70);
  not g_3681 (not_new_n1024_, new_n1024_);
  not g_3682 (not_new_n602__2, new_n602_);
  or g_3683 (new_n3851_, not_new_n621__70, not_new_n6443__70);
  not g_3684 (not_new_n7773__1, new_n7773_);
  or g_3685 (new_n3272_, not_new_n625__8, not_new_n3184__490);
  not g_3686 (not_new_n9090_, new_n9090_);
  and g_3687 (new_n5850_, new_n5990_, new_n6050_);
  not g_3688 (not_new_n9911__0, new_n9911_);
  not g_3689 (not_new_n9836_, new_n9836_);
  not g_3690 (not_new_n8589_, new_n8589_);
  or g_3691 (or_not_new_n2595__not_new_n2594_, not_new_n2594_, not_new_n2595_);
  not g_3692 (not_new_n4466_, new_n4466_);
  or g_3693 (new_n6379_, not_new_n629__8235430, not_new_n6258_);
  not g_3694 (not_new_n5003_, new_n5003_);
  not g_3695 (not_pi146, pi146);
  not g_3696 (not_new_n681__0, new_n681_);
  or g_3697 (new_n4882_, not_new_n4741_, not_new_n1067__7);
  not g_3698 (not_new_n5899_, new_n5899_);
  not g_3699 (new_n4824_, new_n4810_);
  or g_3700 (po070, not_new_n1197_, key_gate_11);
  not g_3701 (not_new_n1175__0, new_n1175_);
  not g_3702 (not_new_n6302_, new_n6302_);
  or g_3703 (new_n9055_, not_new_n8938_, not_new_n9053_);
  and g_3704 (new_n8945_, and_new_n8984__new_n9245_, new_n9244_);
  not g_3705 (not_new_n9689_, new_n9689_);
  or g_3706 (new_n3488_, not_new_n1594__1176490, not_new_n1012__1);
  not g_3707 (not_new_n1469_, new_n1469_);
  not g_3708 (new_n5240_, new_n5000_);
  not g_3709 (not_new_n1598__2, new_n1598_);
  not g_3710 (not_pi140_2, pi140);
  not g_3711 (not_new_n600__490, new_n600_);
  or g_3712 (new_n2280_, not_new_n1332_, not_new_n2275_);
  or g_3713 (new_n6861_, not_new_n1607__10, not_new_n6620_);
  or g_3714 (new_n10136_, not_new_n10018_, not_new_n10135_);
  or g_3715 (or_new_n1031__new_n1037_, new_n1031_, new_n1037_);
  not g_3716 (not_new_n5203__0, new_n5203_);
  not g_3717 (not_new_n9002_, new_n9002_);
  not g_3718 (not_new_n4290_, new_n4290_);
  not g_3719 (new_n5189_, new_n5069_);
  and g_3720 (new_n3959_, and_not_pi034_1_not_pi033_3, not_pi035_1);
  or g_3721 (new_n2274_, not_new_n1589__47475615099430, not_new_n4917_);
  or g_3722 (new_n6111_, not_new_n5756__0, not_new_n1041__70);
  not g_3723 (not_new_n6411_, new_n6411_);
  not g_3724 (not_pi245_0, pi245);
  not g_3725 (not_new_n600__2824752490, new_n600_);
  not g_3726 (not_new_n5883_, new_n5883_);
  not g_3727 (not_new_n9583_, new_n9583_);
  or g_3728 (new_n7550_, not_new_n7549_, not_new_n7548_);
  not g_3729 (not_new_n8562_, new_n8562_);
  not g_3730 (not_new_n9790_, new_n9790_);
  or g_3731 (new_n7862_, not_new_n1597__8235430, not_new_n7663_);
  xor g_3732 (key_gate_75, new_n3921_, key_75);
  not g_3733 (not_new_n600__16284135979104490, new_n600_);
  not g_3734 (not_new_n4506__0, new_n4506_);
  not g_3735 (not_new_n8214_, new_n8214_);
  not g_3736 (not_new_n6032_, new_n6032_);
  or g_3737 (new_n1163_, not_new_n3855_, not_new_n3856_);
  or g_3738 (new_n1799_, not_new_n1589__0, not_new_n5001_);
  not g_3739 (new_n8886_, new_n1601_);
  or g_3740 (new_n9926_, not_new_n1055__39098210485829880490, not_new_n627__16284135979104490);
  not g_3741 (not_new_n4562_, new_n4562_);
  not g_3742 (not_new_n2736_, new_n2736_);
  and g_3743 (new_n8938_, new_n9054_, new_n8983_);
  not g_3744 (not_new_n5740__1, new_n5740_);
  not g_3745 (not_new_n6192_, new_n6192_);
  not g_3746 (not_new_n3078_, new_n3078_);
  or g_3747 (new_n2787_, not_new_n2784_, not_new_n1616__5);
  not g_3748 (not_new_n5447_, new_n5447_);
  not g_3749 (not_new_n3184__1176490, new_n3184_);
  or g_3750 (new_n8781_, not_new_n8709__0, not_new_n8779__0);
  not g_3751 (not_new_n6495_, new_n6495_);
  or g_3752 (new_n5873_, not_new_n6206_, not_new_n6207_);
  not g_3753 (not_new_n637__9, new_n637_);
  not g_3754 (not_new_n4448__0, new_n4448_);
  not g_3755 (not_new_n1053__8235430, new_n1053_);
  and g_3756 (new_n3985_, new_n4057_, new_n4058_);
  not g_3757 (new_n6995_, new_n733_);
  not g_3758 (not_new_n2818_, new_n2818_);
  not g_3759 (not_new_n6078_, new_n6078_);
  and g_3760 (and_new_n9888__new_n10254_, new_n9888_, new_n10254_);
  not g_3761 (not_new_n5789_, new_n5789_);
  or g_3762 (new_n5949_, not_new_n5948_, not_new_n5795__0);
  or g_3763 (new_n8275_, not_new_n8256_, not_new_n8223_);
  or g_3764 (new_n6702_, not_new_n6481__0, not_new_n6654_);
  and g_3765 (new_n1311_, new_n2178_, and_new_n1310__new_n2179_);
  not g_3766 (not_new_n5224_, new_n5224_);
  not g_3767 (not_new_n1071__4, new_n1071_);
  not g_3768 (not_new_n602__3, new_n602_);
  not g_3769 (not_new_n2429_, new_n2429_);
  not g_3770 (not_new_n617__490, new_n617_);
  or g_3771 (new_n5367_, not_new_n5365_, not_new_n5366_);
  or g_3772 (new_n3663_, not_new_n624__9, not_po298_4);
  not g_3773 (not_new_n1041__490, new_n1041_);
  or g_3774 (po080, not_new_n1207_, key_gate_113);
  not g_3775 (not_new_n9859_, new_n9859_);
  not g_3776 (not_new_n7509_, new_n7509_);
  not g_3777 (not_new_n7552_, new_n7552_);
  not g_3778 (not_new_n7229_, new_n7229_);
  and g_3779 (and_new_n1310__new_n2179_, new_n1310_, new_n2179_);
  xnor g_3780 (key_gate_36, new_n3929_, key_36);
  not g_3781 (not_new_n633__70, new_n633_);
  not g_3782 (not_pi051_1, pi051);
  or g_3783 (new_n5153_, not_new_n5085_, not_new_n4902_);
  or g_3784 (new_n5901_, not_new_n5850_, not_new_n6049_);
  not g_3785 (new_n4265_, new_n692_);
  or g_3786 (new_n2403_, not_new_n4137__0, not_new_n600__9);
  not g_3787 (not_new_n1581__2, new_n1581_);
  or g_3788 (new_n5108_, not_new_n1047__8, not_new_n5105_);
  buf g_3789 (po010, pi203);
  or g_3790 (new_n5679_, not_new_n5462__0, not_pi143_2);
  not g_3791 (not_new_n10008__0, new_n10008_);
  not g_3792 (not_new_n636__6782230728490, new_n636_);
  or g_3793 (new_n2102_, not_new_n1591__1176490, not_new_n8814_);
  or g_3794 (new_n10180_, not_new_n633__5585458640832840070, not_new_n1067__332329305696010);
  or g_3795 (new_n2679_, not_po296_1299348114471230201171721456984490, not_pi250_1);
  not g_3796 (not_new_n1591__2, new_n1591_);
  or g_3797 (new_n6887_, not_new_n6886_, not_new_n6807_);
  not g_3798 (not_new_n1047__16284135979104490, new_n1047_);
  not g_3799 (not_new_n2524_, new_n2524_);
  not g_3800 (not_new_n2665_, new_n2665_);
  not g_3801 (not_new_n597__7, new_n597_);
  not g_3802 (not_new_n4743_, new_n4743_);
  not g_3803 (not_new_n10279_, new_n10279_);
  not g_3804 (not_new_n5964_, new_n5964_);
  not g_3805 (not_new_n633__3, new_n633_);
  or g_3806 (new_n1942_, not_new_n4137_, not_new_n585__9);
  or g_3807 (new_n5142_, not_new_n5033_, not_new_n5140_);
  or g_3808 (new_n4496_, not_new_n4567_, not_new_n4568_);
  not g_3809 (not_new_n1494_, new_n1494_);
  not g_3810 (not_new_n8203_, new_n8203_);
  and g_3811 (and_new_n9525__new_n9526_, new_n9525_, new_n9526_);
  or g_3812 (or_not_new_n6226__not_new_n6323_, not_new_n6226_, not_new_n6323_);
  or g_3813 (new_n747_, not_new_n3202_, not_new_n3203_);
  or g_3814 (new_n9177_, not_new_n9064_, not_new_n9175_);
  xor g_3815 (key_gate_3, key_3, new_n1633_);
  not g_3816 (not_new_n3696_, new_n3696_);
  not g_3817 (not_new_n8127__0, new_n8127_);
  not g_3818 (not_new_n1028__0, new_n1028_);
  or g_3819 (new_n2231_, not_new_n5818_, not_new_n1585__968890104070);
  or g_3820 (new_n6856_, not_new_n6854_, not_new_n6855_);
  not g_3821 (not_pi059_0, pi059);
  not g_3822 (not_new_n8904_, new_n8904_);
  not g_3823 (not_new_n975_, new_n975_);
  or g_3824 (new_n5073_, not_new_n5270_, not_new_n5173_);
  not g_3825 (not_new_n595__403536070, new_n595_);
  not g_3826 (not_new_n4727_, new_n4727_);
  and g_3827 (and_new_n1463__new_n1465_, new_n1465_, new_n1463_);
  not g_3828 (not_new_n3503_, new_n3503_);
  not g_3829 (not_new_n5348_, new_n5348_);
  not g_3830 (not_new_n581__273687473400809163430, new_n581_);
  or g_3831 (new_n6889_, not_new_n1600__168070, not_new_n6501__0);
  not g_3832 (not_new_n1379_, new_n1379_);
  not g_3833 (not_new_n1589__16284135979104490, new_n1589_);
  or g_3834 (new_n6932_, not_new_n6531__2, not_new_n1065__8235430);
  not g_3835 (not_new_n8449_, new_n8449_);
  or g_3836 (new_n9057_, new_n644_, new_n1059_);
  not g_3837 (not_new_n7045_, new_n7045_);
  or g_3838 (new_n3235_, not_new_n589__968890104070, not_new_n636__7);
  not g_3839 (not_new_n6293_, new_n6293_);
  not g_3840 (not_new_n9533_, new_n9533_);
  or g_3841 (new_n3655_, not_new_n641__7, not_po298_0);
  or g_3842 (new_n3197_, not_new_n589__4, not_new_n624__7);
  not g_3843 (not_new_n7810_, new_n7810_);
  not g_3844 (not_new_n4151_, new_n4151_);
  not g_3845 (not_new_n9929_, new_n9929_);
  or g_3846 (new_n2914_, not_pi266_0, not_po296_35561530251773635572553173835655155124070416738520070);
  or g_3847 (new_n9605_, new_n1603_, new_n639_);
  not g_3848 (not_new_n608__168070, new_n608_);
  and g_3849 (new_n4482_, new_n4623_, new_n4622_);
  or g_3850 (new_n7169_, not_new_n744_, not_new_n7026_);
  or g_3851 (new_n7983_, not_new_n7742__0, not_new_n1607__3430);
  or g_3852 (new_n4349_, not_new_n4299_, not_new_n4351__0);
  or g_3853 (new_n3750_, not_new_n3748_, not_new_n3749_);
  or g_3854 (new_n4456_, not_new_n4613_, not_new_n4614_);
  or g_3855 (new_n8735_, not_new_n1035__3430, not_new_n8608_);
  or g_3856 (new_n1000_, not_new_n3323_, not_new_n3322_);
  not g_3857 (not_new_n2170_, new_n2170_);
  not g_3858 (not_new_n9212_, new_n9212_);
  not g_3859 (new_n6994_, new_n728_);
  or g_3860 (new_n1873_, not_new_n6561_, not_new_n1580__5);
  not g_3861 (new_n3474_, new_n1061_);
  not g_3862 (not_new_n1612__9, new_n1612_);
  not g_3863 (not_new_n3849_, new_n3849_);
  not g_3864 (not_new_n4818__0, new_n4818_);
  not g_3865 (not_new_n2728_, new_n2728_);
  or g_3866 (po170, not_new_n3567_, not_new_n3566_);
  not g_3867 (not_new_n609__57648010, new_n609_);
  not g_3868 (not_new_n8776_, new_n8776_);
  or g_3869 (new_n5959_, not_new_n5958_, not_new_n5845_);
  not g_3870 (not_new_n989__138412872010, new_n989_);
  not g_3871 (not_new_n643__2824752490, new_n643_);
  not g_3872 (not_new_n5072_, new_n5072_);
  or g_3873 (new_n3561_, not_new_n1612__1176490, not_new_n2109__0);
  not g_3874 (not_new_n4644_, new_n4644_);
  not g_3875 (new_n4229_, new_n677_);
  or g_3876 (new_n10299_, not_new_n10297_, not_new_n10138_);
  not g_3877 (not_new_n4180_, new_n4180_);
  or g_3878 (new_n725_, not_new_n3275_, not_new_n3276_);
  not g_3879 (not_new_n1598__57648010, new_n1598_);
  or g_3880 (or_not_new_n2955__not_new_n2958_, not_new_n2955_, not_new_n2958_);
  and g_3881 (and_new_n3049__new_n998_, new_n3049_, new_n998_);
  or g_3882 (new_n8407_, not_new_n8241_, not_new_n8405_);
  or g_3883 (new_n6005_, not_new_n5768_, not_new_n1600__10);
  not g_3884 (not_new_n10222_, new_n10222_);
  not g_3885 (not_new_n1433_, new_n1433_);
  not g_3886 (not_new_n8568_, new_n8568_);
  or g_3887 (new_n2898_, not_new_n632__2, not_new_n602__57648010);
  or g_3888 (new_n4213_, not_new_n4089_, not_pi261_2);
  not g_3889 (not_new_n1031__2, new_n1031_);
  and g_3890 (new_n9997_, new_n10124_, new_n10021_);
  not g_3891 (new_n7606_, new_n628_);
  not g_3892 (new_n8644_, new_n1166_);
  or g_3893 (po209, not_new_n1402_, or_or_not_new_n1566__not_new_n2489__not_new_n1401_);
  or g_3894 (po243, not_new_n3673_, not_new_n3672_);
  not g_3895 (not_new_n8178__0, new_n8178_);
  not g_3896 (not_new_n952_, new_n952_);
  not g_3897 (not_new_n6619_, new_n6619_);
  or g_3898 (new_n2022_, not_new_n5824_, not_new_n1585__490);
  not g_3899 (not_new_n5938_, new_n5938_);
  or g_3900 (new_n7562_, not_new_n7560_, not_new_n7561_);
  not g_3901 (not_new_n602__70, new_n602_);
  or g_3902 (new_n4707_, not_new_n4506__0, not_new_n4505_);
  or g_3903 (new_n1635_, not_po296_0, not_pi031);
  not g_3904 (not_pi129_1, pi129);
  or g_3905 (new_n5316_, not_new_n4923_, not_new_n628__168070);
  or g_3906 (new_n4327_, not_new_n4330_, or_or_not_new_n4228__not_new_n4329__not_new_n710_);
  not g_3907 (not_new_n1534__168070, key_gate_5);
  or g_3908 (new_n5910_, not_new_n5854_, not_new_n5887_);
  not g_3909 (new_n5174_, new_n5073_);
  or g_3910 (new_n671_, not_new_n3086_, or_not_new_n3088__not_new_n3087_);
  not g_3911 (new_n6506_, new_n1601_);
  not g_3912 (not_new_n1596__7, new_n1596_);
  not g_3913 (not_new_n9514_, new_n9514_);
  not g_3914 (not_new_n585__0, new_n585_);
  or g_3915 (new_n3503_, not_new_n1613__403536070, not_new_n2166_);
  not g_3916 (not_new_n1049__6782230728490, new_n1049_);
  not g_3917 (not_new_n644__138412872010, new_n644_);
  not g_3918 (not_new_n6474__1, new_n6474_);
  not g_3919 (not_new_n1580__70, new_n1580_);
  not g_3920 (not_new_n4071__2, new_n4071_);
  not g_3921 (not_new_n6683_, new_n6683_);
  or g_3922 (new_n3046_, not_new_n3372__138412872010, not_new_n640__4);
  not g_3923 (not_new_n9976_, new_n9976_);
  or g_3924 (new_n9963_, not_new_n10294_, not_new_n10293_);
  and g_3925 (new_n8670_, new_n8735_, new_n8734_);
  not g_3926 (not_new_n9363_, new_n9363_);
  not g_3927 (not_new_n3315__5585458640832840070, new_n3315_);
  not g_3928 (not_new_n1049__70, new_n1049_);
  not g_3929 (not_new_n7625__0, new_n7625_);
  or g_3930 (new_n4546_, new_n1019_, pi171);
  not g_3931 (not_new_n3844_, new_n3844_);
  and g_3932 (new_n5426_, new_n5583_, new_n5587_);
  not g_3933 (not_new_n4123__2, new_n4123_);
  not g_3934 (not_new_n9614__0, new_n9614_);
  not g_3935 (not_new_n4975_, new_n4975_);
  not g_3936 (new_n6271_, new_n635_);
  xor g_3937 (key_gate_56, new_n3992_, key_56);
  or g_3938 (new_n6195_, not_new_n5798__2, not_new_n1065__3430);
  or g_3939 (new_n7068_, not_new_n7556_, not_new_n7557_);
  not g_3940 (not_new_n5772_, new_n5772_);
  not g_3941 (not_new_n7351_, new_n7351_);
  not g_3942 (new_n9658_, new_n9500_);
  not g_3943 (not_new_n9320_, new_n9320_);
  or g_3944 (new_n6894_, not_new_n6503__2, not_new_n1601__403536070);
  or g_3945 (new_n8913_, not_new_n9261_, not_new_n9262_);
  not g_3946 (not_new_n6948_, new_n6948_);
  not g_3947 (new_n9371_, new_n1051_);
  not g_3948 (not_new_n5801__0, new_n5801_);
  or g_3949 (new_n7969_, not_new_n624__19773267430, not_new_n7601__0);
  not g_3950 (new_n2085_, new_n959_);
  not g_3951 (not_pi256_0, pi256);
  not g_3952 (not_new_n1781__0, new_n1781_);
  not g_3953 (not_new_n3252_, new_n3252_);
  not g_3954 (not_pi211, pi211);
  not g_3955 (new_n1626_, new_n922_);
  not g_3956 (not_new_n6985_, new_n6985_);
  not g_3957 (not_new_n1277_, new_n1277_);
  not g_3958 (not_new_n7374_, new_n7374_);
  or g_3959 (new_n4048_, not_new_n4019_, not_new_n3981_);
  not g_3960 (not_new_n9032_, new_n9032_);
  and g_3961 (new_n1557_, new_n3627_, new_n3626_);
  or g_3962 (new_n2293_, not_new_n5010_, not_new_n1589__332329305696010);
  not g_3963 (not_new_n6809_, new_n6809_);
  and g_3964 (new_n1530_, new_n932_, new_n997_);
  or g_3965 (new_n7907_, not_new_n646__2824752490, not_new_n7660_);
  not g_3966 (not_new_n7636_, new_n7636_);
  not g_3967 (not_new_n3259_, new_n3259_);
  or g_3968 (new_n3274_, not_new_n639__8, not_new_n3184__3430);
  not g_3969 (not_new_n639__797922662976120010, new_n639_);
  or g_3970 (or_or_not_new_n2300__not_new_n2301__not_new_n2303_, not_new_n2303_, or_not_new_n2300__not_new_n2301_);
  not g_3971 (new_n1857_, new_n947_);
  or g_3972 (new_n707_, not_new_n3003_, not_new_n1491_);
  or g_3973 (new_n7605_, not_new_n7607_, not_new_n632__19773267430);
  not g_3974 (new_n6633_, new_n1035_);
  or g_3975 (new_n8792_, not_new_n8595__6, not_new_n8616_);
  not g_3976 (not_new_n2009_, new_n2009_);
  and g_3977 (new_n1219_, new_n1741_, and_and_new_n1739__new_n1740__new_n1742_);
  not g_3978 (not_new_n8465_, new_n8465_);
  or g_3979 (new_n9062_, not_new_n1061__138412872010, not_new_n643__2326305139872070);
  or g_3980 (new_n5570_, not_new_n5465_, not_pi144_1);
  or g_3981 (new_n2026_, not_new_n8813_, not_new_n1591__490);
  not g_3982 (not_pi133_1, pi133);
  not g_3983 (not_new_n1165__0, new_n1165_);
  or g_3984 (new_n4708_, not_new_n4706_, not_new_n4549_);
  or g_3985 (new_n3904_, not_new_n3906_, not_new_n10104_);
  not g_3986 (not_new_n9493_, new_n9493_);
  or g_3987 (new_n9832_, not_new_n1061__332329305696010, not_new_n9398_);
  not g_3988 (not_new_n1035__6, new_n1035_);
  not g_3989 (not_new_n611__1, new_n611_);
  not g_3990 (not_new_n1003__3, new_n1003_);
  not g_3991 (new_n8280_, new_n8104_);
  or g_3992 (new_n9402_, not_new_n645__332329305696010, not_new_n1071__138412872010);
  or g_3993 (new_n2536_, not_new_n2533_, or_not_new_n2535__not_new_n2534_);
  or g_3994 (new_n2379_, not_new_n9874__0, not_new_n599__4);
  and g_3995 (new_n9455_, and_new_n9696__new_n9695_, new_n9529_);
  not g_3996 (not_new_n4625_, new_n4625_);
  not g_3997 (new_n8996_, new_n8830_);
  not g_3998 (not_new_n3865_, new_n3865_);
  or g_3999 (new_n3609_, not_new_n1611__8, not_new_n952_);
  not g_4000 (new_n10107_, new_n10026_);
  not g_4001 (not_new_n5466_, new_n5466_);
  not g_4002 (not_new_n7606__1, new_n7606_);
  not g_4003 (not_new_n8257_, new_n8257_);
  not g_4004 (new_n9411_, new_n633_);
  not g_4005 (not_new_n1596__1, new_n1596_);
  or g_4006 (new_n6989_, or_not_new_n7316__not_new_n7186_, not_new_n7185_);
  or g_4007 (new_n7285_, not_new_n6992__0, not_new_n7430__0);
  or g_4008 (new_n4874_, not_new_n1604__7, not_new_n4783_);
  not g_4009 (not_new_n4207_, new_n4207_);
  not g_4010 (not_new_n2261__0, new_n2261_);
  not g_4011 (not_new_n1051__1176490, new_n1051_);
  or g_4012 (new_n8368_, not_new_n8136_, not_new_n1603__57648010);
  not g_4013 (not_new_n7654_, new_n7654_);
  not g_4014 (new_n9918_, new_n638_);
  not g_4015 (not_new_n1521_, new_n1521_);
  not g_4016 (not_new_n8112_, new_n8112_);
  not g_4017 (not_new_n3954_, new_n3954_);
  not g_4018 (not_new_n611__70, new_n611_);
  not g_4019 (not_new_n1584__332329305696010, new_n1584_);
  and g_4020 (and_and_new_n4295__new_n4334__new_n4338_, and_new_n4295__new_n4334_, new_n4338_);
  or g_4021 (or_not_new_n2319__not_new_n2320_, not_new_n2320_, not_new_n2319_);
  not g_4022 (not_new_n995_, new_n995_);
  not g_4023 (not_new_n1538__1176490, new_n1538_);
  or g_4024 (new_n7193_, not_new_n7021__0, not_new_n738__0);
  not g_4025 (not_new_n775__0, new_n775_);
  not g_4026 (not_new_n7349_, new_n7349_);
  not g_4027 (not_new_n3889_, new_n3889_);
  not g_4028 (not_new_n8878_, new_n8878_);
  not g_4029 (not_new_n4659_, new_n4659_);
  or g_4030 (new_n4227_, not_new_n4320_, not_new_n4404_);
  or g_4031 (new_n7291_, not_new_n7430__1, not_new_n6992__1);
  not g_4032 (not_new_n6693_, new_n6693_);
  or g_4033 (new_n1966_, not_new_n1584__9, not_new_n9340_);
  or g_4034 (new_n8424_, not_new_n8087_, not_new_n8175_);
  not g_4035 (not_new_n1572_, new_n1572_);
  not g_4036 (not_new_n1583__24010, new_n1583_);
  not g_4037 (not_new_n6342_, new_n6342_);
  and g_4038 (new_n7073_, new_n7318_, new_n7188_);
  and g_4039 (and_new_n6378__new_n6379_, new_n6379_, new_n6378_);
  not g_4040 (not_new_n645__3430, new_n645_);
  not g_4041 (not_new_n9760_, new_n9760_);
  not g_4042 (not_new_n1392_, new_n1392_);
  or g_4043 (new_n8303_, not_new_n8076_, not_new_n8302_);
  not g_4044 (not_new_n3372__332329305696010, new_n3372_);
  not g_4045 (not_new_n2283_, new_n2283_);
  not g_4046 (new_n6488_, new_n631_);
  or g_4047 (new_n3395_, not_new_n1020__2, not_new_n1594_);
  or g_4048 (new_n1715_, not_new_n1631__332329305696010, not_pi060);
  not g_4049 (not_new_n7622__1, new_n7622_);
  or g_4050 (new_n7913_, not_new_n7912_, not_new_n7830_);
  or g_4051 (new_n2257_, not_new_n9963_, not_new_n594__6782230728490);
  or g_4052 (po077, not_new_n1204_, key_gate_94);
  not g_4053 (not_new_n9426__1, new_n9426_);
  not g_4054 (not_new_n1071__1, new_n1071_);
  not g_4055 (not_new_n7625_, new_n7625_);
  not g_4056 (not_new_n1002__2, new_n1002_);
  or g_4057 (new_n4551_, not_new_n4506_, not_new_n4550_);
  not g_4058 (not_new_n5794_, new_n5794_);
  not g_4059 (not_new_n3086_, new_n3086_);
  not g_4060 (not_new_n591__6782230728490, new_n591_);
  not g_4061 (not_new_n928__1176490, new_n928_);
  or g_4062 (new_n3379_, not_new_n1614_, not_new_n1729_);
  not g_4063 (not_new_n8540_, new_n8540_);
  not g_4064 (not_new_n1607__8, new_n1607_);
  not g_4065 (not_new_n2617_, new_n2617_);
  not g_4066 (not_new_n6029_, new_n6029_);
  or g_4067 (new_n5259_, not_new_n5084__0, not_new_n5216_);
  not g_4068 (not_new_n5747__0, new_n5747_);
  not g_4069 (not_po296_881247870897231951843937366879128181133112010, po296);
  not g_4070 (not_new_n1627_, new_n1627_);
  not g_4071 (not_pi160, pi160);
  not g_4072 (not_new_n7176_, new_n7176_);
  not g_4073 (not_new_n6485_, new_n6485_);
  not g_4074 (not_new_n9777_, new_n9777_);
  or g_4075 (new_n5563_, not_new_n5686_, not_new_n1016__5);
  not g_4076 (not_new_n5130_, new_n5130_);
  or g_4077 (or_not_new_n8781__not_new_n8701_, not_new_n8781_, not_new_n8701_);
  not g_4078 (not_pi265_2, pi265);
  not g_4079 (not_new_n1597__24010, new_n1597_);
  not g_4080 (not_new_n581__13410686196639649008070, new_n581_);
  not g_4081 (not_new_n6098_, new_n6098_);
  not g_4082 (not_new_n10016__1, new_n10016_);
  not g_4083 (not_new_n624__3430, new_n624_);
  or g_4084 (new_n1065_, not_new_n3482_, not_new_n3483_);
  not g_4085 (not_new_n3848_, new_n3848_);
  not g_4086 (not_new_n2172_, new_n2172_);
  or g_4087 (new_n6954_, not_new_n6526__0, not_new_n627__403536070);
  not g_4088 (new_n8852_, new_n1600_);
  or g_4089 (new_n3246_, not_new_n3184_, not_new_n647__8);
  not g_4090 (not_new_n3315__490, new_n3315_);
  not g_4091 (not_pi259_1, pi259);
  not g_4092 (not_new_n4500_, new_n4500_);
  not g_4093 (not_new_n4836_, new_n4836_);
  not g_4094 (not_new_n1603__332329305696010, new_n1603_);
  or g_4095 (new_n4128_, not_new_n4208_, not_new_n4207_);
  not g_4096 (not_new_n585__2824752490, new_n585_);
  and g_4097 (and_and_new_n1934__new_n1937__new_n1935_, and_new_n1934__new_n1937_, new_n1935_);
  not g_4098 (not_new_n4590_, new_n4590_);
  not g_4099 (not_new_n596__2824752490, key_gate_88);
  and g_4100 (new_n603_, new_n593_, new_n1611_);
  not g_4101 (not_new_n9373__2, new_n9373_);
  or g_4102 (new_n3359_, not_pi043_0, not_new_n1534__19773267430);
  and g_4103 (new_n5841_, new_n6045_, new_n5840_);
  not g_4104 (not_new_n8195_, new_n8195_);
  not g_4105 (not_new_n5500__0, new_n5500_);
  not g_4106 (not_new_n7712_, new_n7712_);
  or g_4107 (new_n730_, not_new_n3288_, not_new_n3287_);
  or g_4108 (new_n1911_, not_new_n1580__7, not_new_n6560_);
  not g_4109 (not_new_n626__7, new_n626_);
  not g_4110 (not_new_n5921__0, new_n5921_);
  or g_4111 (new_n1965_, not_new_n1585__9, not_new_n5836_);
  not g_4112 (not_new_n1053__138412872010, new_n1053_);
  not g_4113 (new_n4573_, new_n4494_);
  or g_4114 (new_n4475_, not_new_n4535_, not_new_n4536_);
  not g_4115 (not_new_n4467_, new_n4467_);
  not g_4116 (not_new_n1206_, new_n1206_);
  not g_4117 (not_new_n6473_, new_n6473_);
  not g_4118 (not_pi041_1, pi041);
  not g_4119 (not_new_n3191_, new_n3191_);
  or g_4120 (new_n713_, not_new_n1768_, not_new_n3315_);
  not g_4121 (not_new_n9405_, new_n9405_);
  and g_4122 (po098, key_gate_101, pi077);
  not g_4123 (not_new_n6172_, new_n6172_);
  not g_4124 (not_new_n633__2326305139872070, new_n633_);
  not g_4125 (not_new_n9723_, new_n9723_);
  not g_4126 (not_new_n9637__0, new_n9637_);
  or g_4127 (new_n5967_, not_new_n5748__0, not_new_n5919_);
  not g_4128 (not_new_n7050_, new_n7050_);
  not g_4129 (not_new_n3311__8, new_n3311_);
  not g_4130 (not_new_n4944_, new_n4944_);
  not g_4131 (not_pi173_1, pi173);
  or g_4132 (new_n7485_, not_new_n7448__0, not_new_n722__0);
  or g_4133 (new_n6918_, not_new_n645__403536070, not_new_n6514__0);
  not g_4134 (not_new_n971_, new_n971_);
  not g_4135 (not_new_n6489__0, new_n6489_);
  xnor g_4136 (key_gate_42, key_42, new_n1660_);
  not g_4137 (not_new_n3433_, new_n3433_);
  or g_4138 (new_n10328_, not_new_n9907_, not_new_n646__113988951853731430);
  or g_4139 (or_or_not_new_n8833__not_new_n8830__0_not_new_n9222_, or_not_new_n8833__not_new_n8830__0, not_new_n9222_);
  and g_4140 (new_n4899_, new_n5091_, new_n5092_);
  not g_4141 (not_pi122_0, pi122);
  not g_4142 (not_new_n8661_, new_n8661_);
  not g_4143 (new_n9409_, new_n1065_);
  or g_4144 (new_n5552_, not_new_n5706_, not_new_n1019__5);
  not g_4145 (new_n1776_, new_n942_);
  not g_4146 (not_new_n589__2824752490, new_n589_);
  and g_4147 (new_n7072_, new_n7187_, new_n6967_);
  not g_4148 (new_n6182_, new_n5868_);
  not g_4149 (not_new_n939_, new_n939_);
  not g_4150 (new_n6726_, new_n6636_);
  buf g_4151 (po052, pi276);
  or g_4152 (or_not_new_n10126__not_new_n10125_, not_new_n10125_, not_new_n10126_);
  not g_4153 (not_new_n4504_, new_n4504_);
  not g_4154 (not_new_n4947_, new_n4947_);
  not g_4155 (not_pi203, pi203);
  not g_4156 (not_new_n640__3, new_n640_);
  not g_4157 (not_new_n586__3, new_n586_);
  not g_4158 (not_new_n1809_, new_n1809_);
  or g_4159 (new_n3365_, not_new_n3927__0, not_pi064_968890104070);
  not g_4160 (not_new_n1585__4, new_n1585_);
  not g_4161 (not_new_n9316_, new_n9316_);
  not g_4162 (not_new_n638__57648010, new_n638_);
  not g_4163 (not_new_n7665_, new_n7665_);
  not g_4164 (not_new_n6138_, new_n6138_);
  not g_4165 (new_n8606_, new_n1041_);
  not g_4166 (not_new_n648__168070, new_n648_);
  not g_4167 (not_new_n609__3, new_n609_);
  not g_4168 (not_new_n1027__47475615099430, new_n1027_);
  not g_4169 (new_n6620_, new_n619_);
  not g_4170 (not_pi147_0, pi147);
  not g_4171 (not_new_n1607__9, new_n1607_);
  not g_4172 (new_n5205_, new_n5063_);
  not g_4173 (new_n10082_, new_n10007_);
  not g_4174 (not_new_n6974__57648010, new_n6974_);
  or g_4175 (new_n6890_, not_new_n6502__0, not_new_n629__403536070);
  not g_4176 (not_new_n1496_, new_n1496_);
  or g_4177 (new_n8389_, not_new_n8176_, not_new_n8388_);
  not g_4178 (not_new_n1255_, new_n1255_);
  not g_4179 (not_new_n10028_, new_n10028_);
  or g_4180 (new_n5611_, not_new_n5443__0, not_new_n1005__7);
  not g_4181 (not_new_n1584__138412872010, new_n1584_);
  not g_4182 (not_new_n5625_, new_n5625_);
  or g_4183 (new_n772_, not_new_n3219_, not_new_n3218_);
  not g_4184 (new_n9885_, new_n1041_);
  not g_4185 (not_new_n4131__2, new_n4131_);
  or g_4186 (new_n1762_, not_new_n941_, or_or_not_new_n3397__not_new_n3398__not_new_n1761_);
  not g_4187 (not_new_n8802_, new_n8802_);
  not g_4188 (not_new_n7593_, new_n7593_);
  or g_4189 (new_n8773_, not_new_n8687_, not_new_n8772_);
  not g_4190 (not_new_n7573_, new_n7573_);
  not g_4191 (not_new_n5751_, new_n5751_);
  or g_4192 (new_n9003_, new_n1047_, new_n634_);
  or g_4193 (new_n10125_, not_new_n9861_, not_new_n10036_);
  or g_4194 (or_not_new_n2910__not_new_n2913_, not_new_n2910_, not_new_n2913_);
  or g_4195 (new_n6815_, not_new_n6457_, not_new_n6613__1);
  not g_4196 (not_new_n994__403536070, new_n994_);
  not g_4197 (not_new_n1193_, new_n1193_);
  or g_4198 (new_n10236_, not_new_n647__113988951853731430, not_new_n9898_);
  or g_4199 (or_not_new_n3176__not_new_n3175_, not_new_n3176_, not_new_n3175_);
  or g_4200 (or_not_new_n2758__not_new_n2761_, not_new_n2761_, not_new_n2758_);
  or g_4201 (new_n4488_, not_new_n1010__2, not_new_n4510_);
  or g_4202 (or_or_not_new_n1901__not_new_n1902__not_new_n1904_, or_not_new_n1901__not_new_n1902_, not_new_n1904_);
  or g_4203 (new_n7495_, not_new_n7008__1, not_new_n7040__1);
  and g_4204 (new_n3969_, not_pi062_1, not_pi061_1);
  not g_4205 (not_new_n3424_, new_n3424_);
  not g_4206 (not_new_n2280__0, new_n2280_);
  not g_4207 (not_new_n4522_, new_n4522_);
  or g_4208 (new_n2138_, not_new_n8185_, not_new_n1581__57648010);
  and g_4209 (new_n7709_, new_n7860_, new_n7585_);
  or g_4210 (new_n5870_, not_new_n6190_, not_new_n6191_);
  not g_4211 (not_new_n7565_, new_n7565_);
  or g_4212 (new_n5019_, not_new_n5409_, not_new_n5408_);
  and g_4213 (and_and_new_n6365__new_n6439__new_n6438_, new_n6438_, and_new_n6365__new_n6439_);
  not g_4214 (not_pi271_1, pi271);
  or g_4215 (new_n1071_, not_new_n3497_, not_new_n3498_);
  not g_4216 (not_new_n4281_, new_n4281_);
  not g_4217 (not_new_n627__19773267430, new_n627_);
  and g_4218 (new_n4796_, new_n4884_, new_n4885_);
  not g_4219 (new_n7268_, new_n7138_);
  not g_4220 (not_new_n4999_, new_n4999_);
  or g_4221 (new_n2655_, not_new_n605__24010, not_new_n5481_);
  or g_4222 (new_n4114_, not_new_n4180_, not_new_n4179_);
  and g_4223 (new_n1373_, new_n2418_, new_n2417_);
  or g_4224 (new_n1657_, key_gate_41, not_new_n596__7);
  or g_4225 (new_n8577_, not_new_n8576_, not_new_n8447_);
  or g_4226 (po279, not_new_n2839_, or_or_or_not_new_n2838__not_new_n2841__not_new_n2840__not_new_n2842_);
  or g_4227 (new_n10040_, new_n624_, new_n1041_);
  or g_4228 (new_n9699_, not_new_n9373__1, not_new_n9463_);
  or g_4229 (new_n1169_, not_new_n3868_, not_new_n3867_);
  or g_4230 (new_n7469_, not_new_n7045__2, not_new_n7014__2);
  not g_4231 (new_n4835_, new_n4743_);
  not g_4232 (not_new_n6625__0, new_n6625_);
  not g_4233 (not_new_n972_, new_n972_);
  not g_4234 (not_new_n3159_, new_n3159_);
  not g_4235 (not_new_n1591__2326305139872070, new_n1591_);
  or g_4236 (or_or_not_new_n4228__not_new_n4329__not_new_n710_, or_not_new_n4228__not_new_n4329_, not_new_n710_);
  not g_4237 (not_new_n599__490, new_n599_);
  or g_4238 (or_not_new_n3158__not_new_n3157_, not_new_n3158_, not_new_n3157_);
  not g_4239 (not_new_n771_, new_n771_);
  not g_4240 (not_new_n1047__5, new_n1047_);
  not g_4241 (not_new_n9164_, new_n9164_);
  not g_4242 (not_new_n6710_, new_n6710_);
  not g_4243 (not_new_n7742_, new_n7742_);
  or g_4244 (new_n1861_, not_new_n1041_, not_new_n1588__4);
  not g_4245 (not_new_n5468__0, new_n5468_);
  or g_4246 (new_n4886_, not_new_n1063__7, not_new_n4740_);
  not g_4247 (new_n7116_, new_n747_);
  not g_4248 (not_new_n1602__797922662976120010, new_n1602_);
  or g_4249 (new_n3475_, not_pi111_0, not_new_n1537__3430);
  not g_4250 (not_new_n7048_, new_n7048_);
  and g_4251 (new_n5497_, new_n5603_, new_n5602_);
  not g_4252 (not_new_n1728__19773267430, new_n1728_);
  not g_4253 (new_n8045_, new_n7727_);
  or g_4254 (new_n7905_, not_new_n641__1176490, not_new_n7608_);
  or g_4255 (new_n3784_, not_new_n3396_, not_new_n1791_);
  or g_4256 (po179, not_new_n3585_, not_new_n3584_);
  or g_4257 (new_n9622_, not_new_n9416_, not_new_n9621_);
  and g_4258 (new_n4072_, new_n4174_, new_n4143_);
  not g_4259 (not_new_n10264_, new_n10264_);
  not g_4260 (not_new_n7652_, new_n7652_);
  and g_4261 (new_n8259_, new_n8530_, new_n8531_);
  not g_4262 (not_new_n1728__70, new_n1728_);
  and g_4263 (and_and_not_pi037_2_not_pi036_2_not_pi039_3, and_not_pi037_2_not_pi036_2, not_pi039_3);
  not g_4264 (not_new_n5480__0, new_n5480_);
  not g_4265 (not_new_n639__16284135979104490, new_n639_);
  or g_4266 (new_n9097_, new_n1599_, new_n622_);
  not g_4267 (not_po296_26517308458596534717790233816010, po296);
  or g_4268 (new_n6953_, not_new_n6524__2, not_new_n1055__403536070);
  or g_4269 (new_n5866_, not_new_n6170_, not_new_n6171_);
  not g_4270 (new_n2180_, new_n966_);
  or g_4271 (new_n8265_, not_new_n8179_, not_new_n1031__8235430);
  not g_4272 (not_new_n622__8, new_n622_);
  not g_4273 (not_new_n7935_, new_n7935_);
  not g_4274 (not_new_n8285_, new_n8285_);
  not g_4275 (not_new_n1053__168070, new_n1053_);
  or g_4276 (new_n4582_, not_pi179_2, not_new_n1011__2);
  or g_4277 (new_n5165_, not_new_n638__3430, not_new_n1063__8);
  or g_4278 (new_n3596_, not_new_n984__2, not_pi164_0);
  not g_4279 (not_new_n7373_, new_n7373_);
  not g_4280 (not_new_n4720_, new_n4720_);
  or g_4281 (new_n1593_, not_new_n922_, not_new_n1529_);
  or g_4282 (new_n6038_, not_new_n5875_, not_new_n6036_);
  not g_4283 (not_new_n3314_, new_n3314_);
  not g_4284 (not_new_n7037_, new_n7037_);
  or g_4285 (new_n3310_, not_new_n3308_, not_new_n1617__0);
  not g_4286 (not_new_n4123__1, new_n4123_);
  not g_4287 (not_new_n1785_, new_n1785_);
  not g_4288 (not_new_n5674__1, new_n5674_);
  not g_4289 (not_new_n9214_, new_n9214_);
  not g_4290 (not_new_n6884_, new_n6884_);
  not g_4291 (not_pi273_0, pi273);
  not g_4292 (not_new_n7726_, new_n7726_);
  or g_4293 (new_n1164_, not_new_n3858_, not_new_n3857_);
  not g_4294 (not_pi149, pi149);
  not g_4295 (not_new_n5791_, new_n5791_);
  not g_4296 (not_new_n2716_, new_n2716_);
  not g_4297 (not_new_n9682_, new_n9682_);
  not g_4298 (not_new_n8537_, new_n8537_);
  or g_4299 (or_not_new_n2718__not_new_n2717_, not_new_n2718_, not_new_n2717_);
  not g_4300 (not_new_n641__1176490, new_n641_);
  not g_4301 (not_new_n9698_, new_n9698_);
  not g_4302 (not_new_n6922_, new_n6922_);
  or g_4303 (new_n2733_, not_new_n617__2, not_new_n602__0);
  not g_4304 (not_new_n984__332329305696010, new_n984_);
  or g_4305 (new_n6800_, not_new_n6728_, not_new_n6635_);
  or g_4306 (new_n4122_, not_new_n4196_, not_new_n4195_);
  not g_4307 (new_n9078_, new_n8874_);
  or g_4308 (new_n6760_, not_new_n6640__0, not_new_n6719_);
  not g_4309 (not_new_n994__6782230728490, new_n994_);
  not g_4310 (not_new_n666_, new_n666_);
  not g_4311 (not_new_n7016_, new_n7016_);
  or g_4312 (or_not_new_n2246__not_new_n2243_, not_new_n2246_, not_new_n2243_);
  and g_4313 (new_n9483_, new_n9329_, new_n9680_);
  not g_4314 (not_new_n8482_, new_n8482_);
  not g_4315 (not_new_n1289_, new_n1289_);
  not g_4316 (new_n5473_, new_n1011_);
  or g_4317 (new_n2030_, not_new_n593__490, not_new_n643_);
  not g_4318 (not_pi111_0, pi111);
  and g_4319 (new_n1467_, and_and_and_new_n1463__new_n1465__new_n1464__new_n3720_, new_n1462_);
  not g_4320 (new_n4989_, new_n1599_);
  or g_4321 (new_n9240_, not_new_n8849__0, not_new_n1597__332329305696010);
  or g_4322 (new_n3782_, not_new_n642__9, not_new_n1035__6);
  not g_4323 (not_new_n1063__9, new_n1063_);
  or g_4324 (new_n9532_, new_n1045_, new_n635_);
  not g_4325 (not_new_n1395_, new_n1395_);
  not g_4326 (not_new_n7036__1, new_n7036_);
  not g_4327 (not_new_n1613__168070, new_n1613_);
  not g_4328 (new_n7418_, new_n7033_);
  not g_4329 (not_new_n625__5585458640832840070, new_n625_);
  not g_4330 (not_pi261_0, pi261);
  and g_4331 (new_n7091_, new_n7499_, and_new_n7160__new_n7500_);
  not g_4332 (not_new_n9163_, new_n9163_);
  not g_4333 (not_new_n8684_, new_n8684_);
  not g_4334 (not_new_n2616_, new_n2616_);
  not g_4335 (not_new_n4017__1, new_n4017_);
  or g_4336 (new_n7330_, not_new_n7155__0, not_new_n7079_);
  or g_4337 (new_n3755_, not_new_n969_, not_new_n2190_);
  or g_4338 (new_n7425_, not_new_n7123_, not_new_n775__8235430);
  not g_4339 (not_new_n3566_, new_n3566_);
  not g_4340 (not_new_n9441_, new_n9441_);
  or g_4341 (new_n4134_, not_new_n4219_, not_new_n4220_);
  not g_4342 (not_new_n6737__0, new_n6737_);
  not g_4343 (new_n6981_, new_n741_);
  or g_4344 (new_n2058_, not_new_n601__3430, not_new_n643__0);
  or g_4345 (or_not_new_n3116__not_new_n3115_, not_new_n3115_, not_new_n3116_);
  not g_4346 (not_new_n1002__7, new_n1002_);
  and g_4347 (new_n1233_, new_n1813_, new_n1814_);
  not g_4348 (not_new_n6443__57648010, new_n6443_);
  or g_4349 (new_n4567_, not_new_n4498_, not_new_n4566_);
  and g_4350 (new_n1548_, new_n3608_, new_n3609_);
  or g_4351 (new_n3256_, not_new_n624__8, not_new_n3184__4);
  or g_4352 (new_n2289_, not_new_n1584__332329305696010, not_new_n9438_);
  or g_4353 (new_n2603_, not_new_n609__9, not_new_n4453_);
  not g_4354 (not_new_n634__3430, new_n634_);
  or g_4355 (new_n9119_, not_new_n8804_, not_new_n8898_);
  not g_4356 (not_new_n7221_, new_n7221_);
  or g_4357 (new_n8352_, not_new_n8271_, not_new_n8086_);
  not g_4358 (not_new_n2587_, new_n2587_);
  not g_4359 (not_new_n10000_, new_n10000_);
  not g_4360 (not_pi017, pi017);
  not g_4361 (not_new_n4974_, new_n4974_);
  or g_4362 (new_n8071_, not_new_n8069_, not_new_n8070_);
  or g_4363 (new_n7591_, or_not_new_n7908__not_new_n7743_, not_new_n7763_);
  not g_4364 (not_new_n5748__1, new_n5748_);
  not g_4365 (not_new_n7568_, new_n7568_);
  not g_4366 (not_new_n7137_, new_n7137_);
  not g_4367 (not_new_n5491_, new_n5491_);
  not g_4368 (not_new_n1051__24010, new_n1051_);
  not g_4369 (not_new_n7360__0, new_n7360_);
  not g_4370 (not_new_n6176_, new_n6176_);
  not g_4371 (not_new_n4095_, new_n4095_);
  not g_4372 (not_new_n8867_, new_n8867_);
  not g_4373 (not_new_n5036_, new_n5036_);
  buf g_4374 (po013, pi206);
  not g_4375 (not_new_n5670_, new_n5670_);
  not g_4376 (not_new_n7297_, new_n7297_);
  or g_4377 (new_n2759_, not_new_n4129__2, not_new_n3310__1);
  not g_4378 (not_new_n3952_, new_n3952_);
  not g_4379 (not_new_n7291_, new_n7291_);
  or g_4380 (new_n7223_, not_new_n6994_, not_new_n7427_);
  not g_4381 (not_new_n4302_, new_n4302_);
  and g_4382 (new_n1189_, new_n1656_, new_n1658_);
  or g_4383 (new_n2994_, not_new_n1027__4, not_new_n1150_);
  not g_4384 (not_new_n588__3430, new_n588_);
  not g_4385 (not_new_n3415_, new_n3415_);
  not g_4386 (not_new_n9651_, new_n9651_);
  not g_4387 (not_new_n8448_, new_n8448_);
  not g_4388 (new_n6246_, new_n1599_);
  not g_4389 (not_new_n4938__0, new_n4938_);
  not g_4390 (not_new_n5761_, new_n5761_);
  not g_4391 (not_new_n9453_, new_n9453_);
  not g_4392 (new_n7638_, new_n1071_);
  not g_4393 (not_new_n9496_, new_n9496_);
  or g_4394 (new_n3775_, not_new_n3469_, not_new_n2000_);
  or g_4395 (new_n9072_, not_new_n9069_, not_new_n1067__403536070);
  not g_4396 (not_new_n9660_, new_n9660_);
  not g_4397 (not_new_n7158_, new_n7158_);
  not g_4398 (not_new_n6977_, new_n6977_);
  not g_4399 (not_new_n1197_, new_n1197_);
  not g_4400 (not_new_n626__8, new_n626_);
  or g_4401 (new_n682_, not_new_n1494_, not_new_n3011_);
  not g_4402 (not_new_n5512_, new_n5512_);
  not g_4403 (not_new_n1598__168070, new_n1598_);
  not g_4404 (not_new_n4834_, new_n4834_);
  not g_4405 (not_new_n9980_, new_n9980_);
  not g_4406 (not_new_n6076_, new_n6076_);
  not g_4407 (new_n6533_, new_n643_);
  not g_4408 (not_new_n8170__1, new_n8170_);
  not g_4409 (not_new_n7880_, new_n7880_);
  not g_4410 (not_new_n9445_, new_n9445_);
  not g_4411 (not_new_n3717_, new_n3717_);
  not g_4412 (not_new_n3372__1, new_n3372_);
  not g_4413 (not_new_n622__6782230728490, new_n622_);
  not g_4414 (not_new_n2839_, new_n2839_);
  or g_4415 (new_n3127_, not_new_n581__26517308458596534717790233816010, not_new_n629__6);
  and g_4416 (and_new_n4337__new_n4336_, new_n4336_, new_n4337_);
  not g_4417 (not_new_n3104_, new_n3104_);
  or g_4418 (new_n3280_, not_new_n645__8, not_new_n3184__1176490);
  not g_4419 (not_new_n593__5, new_n593_);
  not g_4420 (not_new_n7136_, new_n7136_);
  not g_4421 (not_new_n9222_, new_n9222_);
  not g_4422 (not_new_n1023__2, new_n1023_);
  not g_4423 (not_new_n3372__2, new_n3372_);
  not g_4424 (not_new_n7295_, new_n7295_);
  and g_4425 (new_n1556_, new_n3624_, new_n3625_);
  or g_4426 (new_n8315_, not_new_n8314_, not_new_n8159__0);
  not g_4427 (not_new_n10165__0, new_n10165_);
  not g_4428 (not_new_n591__1176490, new_n591_);
  or g_4429 (new_n7097_, not_new_n7566_, not_new_n7565_);
  not g_4430 (not_pi257_1, pi257);
  not g_4431 (not_new_n3668_, new_n3668_);
  or g_4432 (new_n9791_, not_new_n9383_, not_new_n625__1915812313805664144010);
  or g_4433 (new_n7369_, not_new_n7357__0, not_new_n737__0);
  not g_4434 (not_new_n6552_, new_n6552_);
  not g_4435 (not_new_n1602__47475615099430, new_n1602_);
  or g_4436 (new_n1826_, not_pi133, not_new_n587__3);
  not g_4437 (not_new_n610_, new_n610_);
  not g_4438 (not_new_n1902_, new_n1902_);
  not g_4439 (not_new_n3476_, new_n3476_);
  or g_4440 (new_n638_, not_new_n2036_, or_or_not_new_n2034__not_new_n2035__not_new_n2037_);
  or g_4441 (po221, not_new_n1430_, or_or_not_new_n2577__not_new_n2581__not_new_n1431_);
  not g_4442 (not_new_n3788_, new_n3788_);
  not g_4443 (not_new_n708_, new_n708_);
  or g_4444 (new_n2288_, not_new_n1585__332329305696010, not_new_n5738_);
  not g_4445 (not_new_n608__8235430, new_n608_);
  or g_4446 (new_n4860_, not_new_n4746_, not_new_n1597__7);
  not g_4447 (not_new_n6472_, new_n6472_);
  not g_4448 (not_new_n8673_, new_n8673_);
  not g_4449 (not_new_n1045__57648010, new_n1045_);
  or g_4450 (new_n7670_, not_new_n7632_, not_new_n7875_);
  not g_4451 (not_new_n631__7, new_n631_);
  not g_4452 (not_new_n7025_, new_n7025_);
  not g_4453 (not_new_n1607__1, new_n1607_);
  not g_4454 (not_new_n1043__1, new_n1043_);
  not g_4455 (not_new_n1588__5, new_n1588_);
  not g_4456 (not_new_n1576__2, new_n1576_);
  or g_4457 (new_n9065_, not_new_n638__273687473400809163430, not_new_n1063__2824752490);
  not g_4458 (not_pi040_4, pi040);
  not g_4459 (not_new_n9377_, new_n9377_);
  and g_4460 (new_n1495_, and_new_n3016__new_n998_, new_n3014_);
  not g_4461 (not_new_n5940_, new_n5940_);
  not g_4462 (not_new_n1597__39098210485829880490, new_n1597_);
  not g_4463 (not_new_n4127__2, new_n4127_);
  not g_4464 (new_n5432_, pi130);
  and g_4465 (new_n1437_, new_n2612_, new_n2610_);
  not g_4466 (not_new_n5444_, new_n5444_);
  not g_4467 (not_new_n1043__968890104070, new_n1043_);
  not g_4468 (not_new_n2918_, new_n2918_);
  not g_4469 (not_pi172, pi172);
  or g_4470 (new_n7563_, not_new_n7155__1, not_new_n7154_);
  or g_4471 (new_n7980_, not_new_n7781__0, not_new_n7740_);
  not g_4472 (not_new_n1601__3430, new_n1601_);
  not g_4473 (not_new_n581__113988951853731430, new_n581_);
  not g_4474 (not_new_n4684_, new_n4684_);
  not g_4475 (not_new_n5900_, new_n5900_);
  not g_4476 (not_new_n5971_, new_n5971_);
  not g_4477 (not_new_n9011__0, new_n9011_);
  or g_4478 (new_n4054_, not_new_n3981__0, or_not_pi064_5585458640832840070_not_new_n4019__0);
  not g_4479 (not_new_n6650_, new_n6650_);
  not g_4480 (new_n6975_, new_n737_);
  not g_4481 (new_n4016_, new_n3952_);
  or g_4482 (new_n2721_, not_new_n933_, not_new_n986_);
  or g_4483 (new_n5623_, not_pi133_2, not_new_n5439_);
  or g_4484 (new_n9784_, not_new_n9414_, not_new_n630__16284135979104490);
  not g_4485 (not_new_n1346_, new_n1346_);
  not g_4486 (not_new_n648__138412872010, new_n648_);
  not g_4487 (not_new_n593__57648010, new_n593_);
  or g_4488 (new_n1831_, not_new_n1583__2, not_new_n7592_);
  or g_4489 (new_n2661_, not_new_n606__24010, not_new_n5481__0);
  or g_4490 (or_not_new_n618__19773267430_not_new_n6865_, not_new_n6865_, not_new_n618__19773267430);
  not g_4491 (not_pi255_2, pi255);
  not g_4492 (not_new_n6494_, new_n6494_);
  or g_4493 (new_n2547_, not_new_n2546_, not_new_n611__7);
  not g_4494 (not_new_n2014__0, new_n2014_);
  not g_4495 (not_new_n630__5585458640832840070, new_n630_);
  not g_4496 (not_new_n1728__6, new_n1728_);
  or g_4497 (new_n3427_, not_pi027_0, not_new_n1536__57648010);
  and g_4498 (new_n1503_, new_n998_, new_n3027_);
  or g_4499 (new_n9781_, not_new_n9779_, not_new_n9780_);
  or g_4500 (new_n2127_, not_new_n1588__57648010, not_new_n1069_);
  not g_4501 (not_new_n7855__0, new_n7855_);
  or g_4502 (new_n3943_, not_new_n4014__0, not_new_n3914__0);
  or g_4503 (new_n7995_, not_new_n7663__2, not_new_n1597__403536070);
  or g_4504 (po203, or_or_not_new_n1560__not_new_n2459__not_new_n1389_, not_new_n1390_);
  not g_4505 (not_new_n7676_, new_n7676_);
  not g_4506 (not_new_n585__47475615099430, new_n585_);
  not g_4507 (not_new_n8843_, new_n8843_);
  not g_4508 (not_new_n7168_, new_n7168_);
  and g_4509 (new_n10000_, and_new_n9915__new_n10334_, new_n10333_);
  not g_4510 (not_new_n1616__1176490, new_n1616_);
  or g_4511 (new_n6176_, not_new_n642__168070, not_new_n5898__1);
  not g_4512 (not_new_n2673_, new_n2673_);
  not g_4513 (not_new_n2706_, new_n2706_);
  not g_4514 (not_new_n7932_, new_n7932_);
  or g_4515 (new_n8338_, not_new_n8078_, not_new_n8337_);
  not g_4516 (not_new_n6304_, new_n6304_);
  or g_4517 (new_n2060_, not_new_n1585__24010, not_new_n5834_);
  not g_4518 (not_new_n1172_, new_n1172_);
  or g_4519 (new_n2666_, or_not_new_n2665__not_new_n2664_, not_new_n2663_);
  not g_4520 (not_new_n1613__1176490, new_n1613_);
  or g_4521 (new_n2924_, not_new_n646__3, not_new_n604__2824752490);
  not g_4522 (not_new_n585_, new_n585_);
  or g_4523 (new_n3696_, not_pi234, not_new_n989__2824752490);
  or g_4524 (new_n3443_, not_new_n1003__1, not_new_n1594__7);
  or g_4525 (new_n8024_, not_new_n7636__0, not_new_n640__19773267430);
  not g_4526 (not_new_n4299_, new_n4299_);
  not g_4527 (not_new_n9154_, new_n9154_);
  or g_4528 (new_n7484_, not_new_n7482_, not_new_n7252_);
  or g_4529 (new_n8262_, not_new_n8433_, not_new_n8423_);
  not g_4530 (not_new_n994__968890104070, new_n994_);
  not g_4531 (not_new_n5438_, new_n5438_);
  not g_4532 (not_new_n5518_, new_n5518_);
  and g_4533 (and_new_n2374__new_n2373_, new_n2373_, new_n2374_);
  not g_4534 (not_new_n9427__2, new_n9427_);
  not g_4535 (not_po298_24010, po298);
  not g_4536 (not_pi049_2, pi049);
  and g_4537 (new_n3961_, not_pi041_1, and_and_not_pi040_1_not_pi039_1_not_pi042_1);
  xor g_4538 (key_gate_127, key_127, not_new_n1696_);
  not g_4539 (not_new_n5418_, new_n5418_);
  or g_4540 (new_n3381_, not_new_n1614__0, not_new_n1730_);
  not g_4541 (new_n6276_, new_n648_);
  not g_4542 (new_n4418_, new_n1009_);
  and g_4543 (new_n1349_, new_n2357_, and_new_n2359__new_n2358_);
  or g_4544 (po190, not_new_n1363_, or_not_new_n1547__not_new_n1364_);
  or g_4545 (new_n7247_, not_new_n723_, not_new_n7040_);
  or g_4546 (new_n4695_, not_new_n1017__3, not_new_n4437_);
  or g_4547 (new_n4894_, not_new_n4738_, not_new_n1055__8);
  or g_4548 (new_n2282_, not_new_n587__2326305139872070, not_pi157);
  not g_4549 (not_new_n2489_, new_n2489_);
  not g_4550 (not_new_n936_, new_n936_);
  or g_4551 (new_n5578_, not_new_n1012__5, not_pi146_1);
  not g_4552 (not_new_n5745_, new_n5745_);
  or g_4553 (new_n9767_, not_new_n9376__0, not_new_n617__1915812313805664144010);
  not g_4554 (not_new_n1544_, new_n1544_);
  not g_4555 (not_new_n1039__3430, new_n1039_);
  or g_4556 (new_n5452_, not_new_n5550_, not_new_n5549_);
  or g_4557 (new_n7059_, not_new_n7497_, not_new_n7498_);
  not g_4558 (not_new_n4131__1, new_n4131_);
  not g_4559 (not_new_n4182_, new_n4182_);
  not g_4560 (not_new_n8244__1, new_n8244_);
  and g_4561 (new_n1415_, new_n1414_, and_new_n2513__new_n2512_);
  not g_4562 (not_new_n1053__9, new_n1053_);
  buf g_4563 (po044, pi220);
  not g_4564 (not_new_n643__5, new_n643_);
  or g_4565 (new_n10242_, not_new_n9896_, not_new_n1049__113988951853731430);
  or g_4566 (new_n6869_, not_new_n618__138412872010, not_new_n6540__1);
  not g_4567 (not_new_n3692_, new_n3692_);
  not g_4568 (not_new_n10025_, new_n10025_);
  or g_4569 (new_n9771_, not_new_n9769_, not_new_n9630_);
  or g_4570 (new_n9847_, not_new_n9845_, not_new_n9846_);
  not g_4571 (not_new_n8082__0, new_n8082_);
  not g_4572 (not_pi189_0, pi189);
  or g_4573 (new_n680_, not_new_n3178_, not_new_n3177_);
  not g_4574 (not_new_n9435_, new_n9435_);
  not g_4575 (not_new_n5164_, new_n5164_);
  not g_4576 (new_n8170_, new_n617_);
  or g_4577 (new_n5682_, not_new_n5680__0, not_new_n5681_);
  not g_4578 (not_new_n619__138412872010, new_n619_);
  and g_4579 (new_n4298_, and_new_n4351__new_n4350_, new_n4346_);
  not g_4580 (not_new_n6155_, new_n6155_);
  or g_4581 (new_n2767_, not_new_n3311__2, not_new_n1037__1);
  or g_4582 (new_n4196_, not_new_n4107_, not_new_n4172__0);
  or g_4583 (new_n5109_, not_new_n4945_, not_new_n4900_);
  or g_4584 (new_n9726_, not_new_n1049__2326305139872070, not_new_n9369_);
  or g_4585 (new_n6148_, not_new_n5804__0, not_new_n622__1176490);
  not g_4586 (not_new_n1049__168070, new_n1049_);
  or g_4587 (or_or_not_new_n1552__not_new_n2419__not_new_n1373_, or_not_new_n1552__not_new_n2419_, not_new_n1373_);
  and g_4588 (new_n597_, new_n1586_, new_n1611_);
  not g_4589 (not_new_n1631__19773267430, key_gate_76);
  not g_4590 (not_new_n927__1, new_n927_);
  or g_4591 (new_n4220_, not_new_n4160_, not_new_n4084_);
  not g_4592 (not_new_n593__332329305696010, new_n593_);
  not g_4593 (not_new_n8282__0, new_n8282_);
  not g_4594 (not_pi044_2, pi044);
  not g_4595 (not_new_n2206_, new_n2206_);
  not g_4596 (not_new_n3921_, key_gate_75);
  not g_4597 (not_new_n593__4, new_n593_);
  and g_4598 (new_n8082_, new_n8364_, new_n8365_);
  not g_4599 (not_new_n613__7, new_n613_);
  not g_4600 (not_new_n594__490, new_n594_);
  not g_4601 (not_new_n594__332329305696010, new_n594_);
  and g_4602 (new_n4915_, new_n5228_, new_n5225_);
  or g_4603 (new_n10257_, not_new_n10256_, not_new_n10255_);
  or g_4604 (new_n6432_, or_or_not_new_n6349__not_new_n6373__7_not_new_n1041__490, not_new_n6235__1);
  and g_4605 (new_n8701_, new_n8795_, new_n8700_);
  or g_4606 (or_not_new_n2982__not_new_n2985_, not_new_n2985_, not_new_n2982_);
  or g_4607 (or_not_new_n2899__not_new_n2898_, not_new_n2898_, not_new_n2899_);
  or g_4608 (new_n3687_, not_new_n637__9, not_po298_1176490);
  not g_4609 (not_new_n930_, new_n930_);
  not g_4610 (not_new_n5624_, new_n5624_);
  and g_4611 (new_n1547_, new_n3606_, new_n3607_);
  not g_4612 (not_new_n602__2824752490, new_n602_);
  or g_4613 (po083, key_gate_40, not_new_n1210_);
  not g_4614 (not_new_n618__797922662976120010, new_n618_);
  not g_4615 (not_new_n6105_, new_n6105_);
  or g_4616 (new_n6040_, not_new_n5915__0, not_new_n6039_);
  not g_4617 (not_new_n3318__1, new_n3318_);
  or g_4618 (new_n7055_, not_new_n7472_, not_new_n7471_);
  not g_4619 (not_pi181, pi181);
  not g_4620 (not_new_n4955__0, new_n4955_);
  not g_4621 (not_new_n1581__7, new_n1581_);
  not g_4622 (not_new_n6504_, new_n6504_);
  not g_4623 (not_new_n6079_, new_n6079_);
  or g_4624 (new_n6375_, not_new_n6247_, not_new_n621__57648010);
  not g_4625 (not_new_n2844_, new_n2844_);
  not g_4626 (not_new_n1536__332329305696010, new_n1536_);
  not g_4627 (not_new_n7359_, new_n7359_);
  not g_4628 (not_new_n3315__2, new_n3315_);
  or g_4629 (new_n4850_, not_new_n4752_, not_new_n1049__7);
  not g_4630 (not_new_n1482_, new_n1482_);
  or g_4631 (new_n4701_, not_new_n4553_, not_new_n4699_);
  not g_4632 (not_new_n645__8, new_n645_);
  not g_4633 (not_new_n639__2326305139872070, new_n639_);
  or g_4634 (new_n9265_, not_new_n625__39098210485829880490, not_new_n8855__0);
  not g_4635 (not_new_n9849_, new_n9849_);
  not g_4636 (not_new_n6493_, new_n6493_);
  not g_4637 (not_new_n1069__8235430, new_n1069_);
  not g_4638 (not_new_n7241_, new_n7241_);
  and g_4639 (new_n1181_, key_gate_125, key_gate_44);
  or g_4640 (or_or_not_new_n1558__not_new_n2449__not_new_n1385_, or_not_new_n1558__not_new_n2449_, not_new_n1385_);
  or g_4641 (new_n8258_, not_new_n8435_, not_new_n8425_);
  or g_4642 (new_n3647_, not_new_n1611__2326305139872070, not_new_n980_);
  or g_4643 (new_n4059_, not_pi057_3, not_new_n3943_);
  not g_4644 (not_new_n9491__0, new_n9491_);
  xnor g_4645 (key_gate_112, key_112, not_new_n1534_);
  or g_4646 (new_n3661_, not_new_n628__9, not_po298_3);
  not g_4647 (not_new_n7378_, new_n7378_);
  not g_4648 (not_new_n9864_, new_n9864_);
  not g_4649 (not_new_n601__2824752490, new_n601_);
  not g_4650 (not_new_n1534__1, key_gate_5);
  or g_4651 (new_n4652_, not_new_n4651_, not_new_n4650_);
  or g_4652 (new_n6846_, not_new_n6495__0, not_new_n6699_);
  and g_4653 (and_new_n10212__new_n10211_, new_n10212_, new_n10211_);
  or g_4654 (new_n755_, not_new_n3221_, not_new_n3220_);
  or g_4655 (or_or_not_new_n1319__not_new_n1317__not_new_n2211_, not_new_n2211_, or_not_new_n1319__not_new_n1317_);
  or g_4656 (new_n3448_, not_new_n1002__1, not_new_n1594__8);
  and g_4657 (and_new_n8667__new_n8666_, new_n8667_, new_n8666_);
  not g_4658 (not_new_n1534__2824752490, key_gate_5);
  not g_4659 (not_new_n9524__0, new_n9524_);
  not g_4660 (not_new_n6516__0, new_n6516_);
  not g_4661 (not_new_n5462__0, new_n5462_);
  or g_4662 (new_n1165_, not_new_n3859_, not_new_n3860_);
  and g_4663 (new_n1329_, new_n2270_, new_n2269_);
  not g_4664 (new_n7167_, new_n6987_);
  or g_4665 (new_n1656_, not_po296_7, not_pi024);
  not g_4666 (not_pi103, pi103);
  not g_4667 (not_new_n7610__0, new_n7610_);
  or g_4668 (new_n7399_, not_new_n743__0, not_new_n7354__2);
  not g_4669 (not_new_n5688_, new_n5688_);
  not g_4670 (not_new_n631__57648010, new_n631_);
  not g_4671 (not_new_n7021__1, new_n7021_);
  or g_4672 (new_n2173_, not_new_n1583__2824752490, not_new_n7691_);
  not g_4673 (not_new_n2872_, new_n2872_);
  not g_4674 (not_pi087, pi087);
  not g_4675 (not_new_n1020__4, new_n1020_);
  and g_4676 (new_n8214_, new_n8421_, new_n8356_);
  not g_4677 (not_new_n5040_, new_n5040_);
  not g_4678 (new_n8576_, new_n8239_);
  not g_4679 (not_new_n1055__3430, new_n1055_);
  not g_4680 (not_new_n644__0, new_n644_);
  not g_4681 (not_new_n7614_, new_n7614_);
  and g_4682 (and_new_n2389__new_n2388_, new_n2388_, new_n2389_);
  not g_4683 (not_new_n613__0, new_n613_);
  not g_4684 (not_new_n8978__3, new_n8978_);
  not g_4685 (not_new_n6625__1, new_n6625_);
  not g_4686 (not_new_n5291_, new_n5291_);
  not g_4687 (not_new_n1018__5, new_n1018_);
  or g_4688 (new_n2553_, not_new_n609__4, not_new_n4465_);
  and g_4689 (new_n1323_, new_n2235_, and_new_n1322__new_n2236_);
  or g_4690 (new_n10096_, new_n1057_, new_n636_);
  not g_4691 (not_new_n969_, new_n969_);
  or g_4692 (or_or_or_not_new_n2928__not_new_n2931__not_new_n2930__not_new_n2932_, or_or_not_new_n2928__not_new_n2931__not_new_n2930_, not_new_n2932_);
  not g_4693 (not_new_n606__3, new_n606_);
  not g_4694 (not_new_n9155_, new_n9155_);
  not g_4695 (not_new_n9476_, new_n9476_);
  not g_4696 (not_new_n7026__0, new_n7026_);
  or g_4697 (new_n3244_, not_pi129_0, not_new_n1626__0);
  not g_4698 (not_new_n9625_, new_n9625_);
  not g_4699 (not_new_n8314_, new_n8314_);
  or g_4700 (new_n8898_, not_new_n9117_, not_new_n8878_);
  or g_4701 (new_n9026_, not_new_n8847_, not_new_n8991_);
  or g_4702 (new_n1836_, not_new_n8907_, not_new_n1591__2);
  or g_4703 (new_n1946_, not_new_n5826_, not_new_n1585__8);
  not g_4704 (not_new_n2509_, new_n2509_);
  or g_4705 (new_n6763_, not_new_n6761_, not_new_n6762_);
  not g_4706 (not_new_n5993_, new_n5993_);
  not g_4707 (not_new_n1631__490, key_gate_76);
  or g_4708 (or_not_new_n2803__not_new_n2806_, not_new_n2806_, not_new_n2803_);
  not g_4709 (not_new_n4766__0, new_n4766_);
  not g_4710 (not_new_n6151_, new_n6151_);
  not g_4711 (new_n8160_, new_n636_);
  or g_4712 (new_n9205_, not_new_n1045__113988951853731430, not_new_n8835_);
  and g_4713 (and_new_n1234__new_n1818_, new_n1818_, new_n1234_);
  not g_4714 (not_new_n8162_, new_n8162_);
  not g_4715 (not_new_n2927_, new_n2927_);
  not g_4716 (not_new_n1065__2326305139872070, new_n1065_);
  not g_4717 (new_n6263_, new_n639_);
  or g_4718 (new_n1824_, not_new_n1819_, not_new_n1236_);
  not g_4719 (not_new_n588__8, new_n588_);
  or g_4720 (or_not_new_n6538__1_not_new_n6877_, not_new_n6538__1, not_new_n6877_);
  or g_4721 (new_n8188_, not_new_n8578_, not_new_n8577_);
  not g_4722 (not_new_n7727_, new_n7727_);
  not g_4723 (not_new_n5884_, new_n5884_);
  or g_4724 (new_n8753_, not_new_n8678_, not_new_n8595__3);
  not g_4725 (not_new_n7757_, new_n7757_);
  not g_4726 (not_new_n9939_, new_n9939_);
  not g_4727 (not_new_n1471_, new_n1471_);
  not g_4728 (not_new_n646__6782230728490, new_n646_);
  not g_4729 (not_new_n927__0, new_n927_);
  or g_4730 (new_n9373_, not_new_n9455_, not_new_n9454_);
  not g_4731 (not_new_n1055__168070, new_n1055_);
  not g_4732 (not_new_n5361_, new_n5361_);
  not g_4733 (new_n6498_, new_n1597_);
  or g_4734 (new_n7477_, not_new_n7475_, not_new_n7476_);
  or g_4735 (new_n5703_, not_new_n5517__0, not_new_n5516_);
  not g_4736 (new_n4449_, pi179);
  not g_4737 (not_new_n8044_, new_n8044_);
  not g_4738 (not_pi107_0, pi107);
  not g_4739 (new_n5458_, new_n1017_);
  not g_4740 (not_pi185_0, pi185);
  not g_4741 (not_new_n2464_, new_n2464_);
  not g_4742 (not_new_n1061__5, new_n1061_);
  not g_4743 (not_new_n7043__1, new_n7043_);
  not g_4744 (not_new_n3892_, new_n3892_);
  not g_4745 (not_new_n7631__0, new_n7631_);
  not g_4746 (not_new_n7604_, new_n7604_);
  not g_4747 (not_new_n6626_, new_n6626_);
  not g_4748 (not_new_n9875__0, new_n9875_);
  or g_4749 (new_n2630_, not_new_n1004__0, not_new_n608__70);
  not g_4750 (not_new_n5540_, new_n5540_);
  not g_4751 (new_n4435_, pi172);
  not g_4752 (not_new_n1596__5585458640832840070, new_n1596_);
  not g_4753 (not_new_n587__70, new_n587_);
  or g_4754 (new_n4692_, not_new_n4691_, not_new_n4690_);
  or g_4755 (new_n1992_, not_new_n636_, not_new_n593__10);
  not g_4756 (not_new_n1065__5, new_n1065_);
  not g_4757 (not_new_n7886_, new_n7886_);
  not g_4758 (not_new_n3207_, new_n3207_);
  or g_4759 (new_n8435_, not_new_n8266__1, not_new_n8090_);
  or g_4760 (new_n2417_, not_new_n643__1, not_new_n603__490);
  not g_4761 (not_new_n9415__0, new_n9415_);
  not g_4762 (not_new_n605__5, new_n605_);
  or g_4763 (new_n5530_, pi133, new_n1007_);
  not g_4764 (not_new_n608__5, new_n608_);
  not g_4765 (not_new_n8832_, new_n8832_);
  not g_4766 (not_new_n9118_, new_n9118_);
  or g_4767 (new_n7906_, not_new_n642__19773267430, not_new_n7752__0);
  not g_4768 (not_new_n8128__0, new_n8128_);
  not g_4769 (not_new_n6971_, new_n6971_);
  not g_4770 (new_n6291_, new_n1047_);
  not g_4771 (not_new_n10012_, new_n10012_);
  not g_4772 (new_n4238_, new_n674_);
  not g_4773 (not_new_n1607__4, new_n1607_);
  not g_4774 (not_new_n7014_, new_n7014_);
  not g_4775 (not_new_n617__2824752490, new_n617_);
  and g_4776 (new_n1229_, new_n1794_, new_n1795_);
  and g_4777 (and_new_n1294__new_n2103_, new_n1294_, new_n2103_);
  not g_4778 (not_new_n4418__0, new_n4418_);
  not g_4779 (not_new_n5467_, new_n5467_);
  or g_4780 (new_n9256_, not_new_n630__47475615099430, not_new_n8886_);
  not g_4781 (not_new_n4167_, new_n4167_);
  not g_4782 (new_n6062_, new_n5892_);
  not g_4783 (not_new_n8698_, new_n8698_);
  not g_4784 (new_n4841_, new_n4746_);
  or g_4785 (or_not_new_n6373__9_not_new_n6237_, not_new_n6373__9, not_new_n6237_);
  not g_4786 (not_new_n4626_, new_n4626_);
  and g_4787 (new_n4784_, new_n4874_, new_n4875_);
  not g_4788 (not_new_n586__168070, new_n586_);
  not g_4789 (not_new_n6988__0, new_n6988_);
  not g_4790 (not_new_n8651_, new_n8651_);
  or g_4791 (new_n8020_, not_new_n639__138412872010, not_new_n7633__0);
  not g_4792 (not_new_n7083_, new_n7083_);
  not g_4793 (not_new_n7887__0, new_n7887_);
  and g_4794 (new_n7707_, new_n7580_, new_n7842_);
  not g_4795 (not_new_n984__113988951853731430, new_n984_);
  not g_4796 (new_n8147_, new_n633_);
  not g_4797 (not_new_n6122_, new_n6122_);
  not g_4798 (not_new_n8402_, new_n8402_);
  xnor g_4799 (key_gate_113, key_113, not_new_n1711_);
  not g_4800 (not_new_n1063__3, new_n1063_);
  or g_4801 (new_n2118_, not_new_n9444_, not_new_n1584__8235430);
  not g_4802 (new_n4921_, new_n1037_);
  not g_4803 (not_new_n636__0, new_n636_);
  or g_4804 (new_n2150_, not_pi118, not_new_n588__2824752490);
  or g_4805 (new_n9001_, not_new_n1043__2824752490, not_new_n8981_);
  not g_4806 (not_new_n5810_, new_n5810_);
  and g_4807 (new_n4288_, and_new_n4323__new_n4324_, new_n4325_);
  or g_4808 (new_n5556_, not_new_n5517_, not_new_n5555_);
  not g_4809 (not_new_n617__2, new_n617_);
  or g_4810 (new_n5350_, not_new_n5348_, not_new_n5209__0);
  not g_4811 (not_new_n2576_, new_n2576_);
  or g_4812 (new_n6697_, not_new_n6577_, not_new_n6695_);
  or g_4813 (po183, not_new_n1349_, not_new_n1350_);
  not g_4814 (not_new_n629__113988951853731430, new_n629_);
  not g_4815 (not_new_n4557_, new_n4557_);
  not g_4816 (not_new_n927_, new_n927_);
  or g_4817 (new_n7387_, not_new_n7385_, not_new_n7386_);
  not g_4818 (not_new_n4794_, new_n4794_);
  not g_4819 (not_new_n628__10, new_n628_);
  or g_4820 (new_n5008_, not_new_n5329_, not_new_n5328_);
  or g_4821 (new_n2520_, not_new_n608__0, not_new_n1011_);
  not g_4822 (not_new_n6560_, new_n6560_);
  not g_4823 (not_new_n10034_, new_n10034_);
  not g_4824 (not_new_n7954_, new_n7954_);
  and g_4825 (new_n3922_, new_n4038_, new_n3948_);
  or g_4826 (new_n3183_, not_new_n1624_, not_new_n922__1);
  not g_4827 (not_new_n7770__0, new_n7770_);
  or g_4828 (new_n7962_, not_new_n7600__0, not_new_n635__19773267430);
  not g_4829 (not_new_n10052__0, new_n10052_);
  not g_4830 (not_new_n3981__0, new_n3981_);
  or g_4831 (new_n630_, not_new_n2188_, or_or_not_new_n2189__not_new_n2186__not_new_n2187_);
  not g_4832 (new_n1622_, new_n941_);
  or g_4833 (new_n8461_, not_new_n8244__3, not_new_n8315_);
  or g_4834 (po284, or_or_or_not_new_n2883__not_new_n2886__not_new_n2885__not_new_n2887_, not_new_n2884_);
  not g_4835 (not_new_n601__19773267430, new_n601_);
  or g_4836 (new_n2783_, not_new_n994__7, not_new_n4125__1);
  or g_4837 (new_n4998_, not_new_n4978_, not_new_n5217_);
  not g_4838 (not_new_n589__3788186922656647816827176259430, new_n589_);
  not g_4839 (not_new_n598__332329305696010, new_n598_);
  not g_4840 (not_new_n7621_, new_n7621_);
  or g_4841 (new_n9727_, not_new_n9725_, not_new_n9726_);
  or g_4842 (new_n2944_, not_new_n4137__1, not_new_n994__47475615099430);
  and g_4843 (new_n8228_, new_n8283_, new_n8387_);
  or g_4844 (new_n3858_, not_new_n630__490, not_new_n1576__24010);
  and g_4845 (new_n8658_, new_n1031_, new_n8706_);
  not g_4846 (not_new_n5798_, new_n5798_);
  not g_4847 (not_new_n7239_, new_n7239_);
  or g_4848 (new_n1735_, not_new_n1728__3, not_pi079);
  not g_4849 (not_new_n6343_, new_n6343_);
  or g_4850 (new_n6858_, not_new_n6483__0, not_new_n632__2824752490);
  not g_4851 (not_new_n7750__0, new_n7750_);
  not g_4852 (not_new_n9714__0, new_n9714_);
  not g_4853 (not_new_n641__490, new_n641_);
  not g_4854 (not_new_n3969_, new_n3969_);
  not g_4855 (new_n6262_, new_n640_);
  not g_4856 (not_new_n5718_, new_n5718_);
  not g_4857 (not_new_n632__3430, new_n632_);
  not g_4858 (not_new_n7586_, new_n7586_);
  not g_4859 (not_new_n7745_, new_n7745_);
  not g_4860 (not_new_n9686_, new_n9686_);
  or g_4861 (new_n920_, not_new_n3372_, not_new_n1622_);
  not g_4862 (not_new_n8900_, new_n8900_);
  or g_4863 (new_n4504_, not_new_n4551_, not_new_n4552_);
  or g_4864 (new_n9161_, not_new_n8874__1, not_new_n9131_);
  or g_4865 (new_n1998_, not_new_n588__490, not_pi110);
  not g_4866 (not_new_n9677_, new_n9677_);
  not g_4867 (not_new_n610__3, new_n610_);
  not g_4868 (new_n5196_, new_n5066_);
  not g_4869 (not_pi262_1, pi262);
  not g_4870 (new_n5166_, new_n4999_);
  not g_4871 (not_new_n9918__0, new_n9918_);
  not g_4872 (not_new_n9185_, new_n9185_);
  not g_4873 (new_n6529_, new_n636_);
  not g_4874 (new_n6284_, new_n1055_);
  not g_4875 (not_new_n6064__0, new_n6064_);
  not g_4876 (not_new_n1049__9, new_n1049_);
  not g_4877 (not_new_n6817_, new_n6817_);
  not g_4878 (not_new_n5720_, new_n5720_);
  not g_4879 (not_new_n3192_, new_n3192_);
  and g_4880 (new_n7743_, new_n7986_, new_n7987_);
  not g_4881 (not_new_n1589__10, new_n1589_);
  or g_4882 (or_not_new_n3944__not_new_n3914__1, not_new_n3914__1, not_new_n3944_);
  not g_4883 (not_new_n640__9, new_n640_);
  not g_4884 (not_new_n3112_, new_n3112_);
  or g_4885 (new_n4673_, not_new_n4569_, not_new_n4671_);
  not g_4886 (not_new_n9306_, new_n9306_);
  or g_4887 (new_n5688_, not_new_n5687_, not_new_n5686__0);
  not g_4888 (not_new_n3310__490, new_n3310_);
  or g_4889 (or_not_new_n10210__not_new_n10153_, not_new_n10210_, not_new_n10153_);
  not g_4890 (not_new_n3408_, new_n3408_);
  not g_4891 (not_new_n984__2, new_n984_);
  not g_4892 (not_new_n585__16284135979104490, new_n585_);
  and g_4893 (new_n10027_, new_n3909_, new_n3910_);
  not g_4894 (not_new_n631__273687473400809163430, new_n631_);
  or g_4895 (new_n4656_, not_pi179_4, not_new_n4450__0);
  not g_4896 (not_po298_332329305696010, po298);
  not g_4897 (not_new_n1577_, new_n1577_);
  not g_4898 (not_new_n5909_, new_n5909_);
  or g_4899 (new_n7788_, not_new_n7599_, not_new_n631__6782230728490);
  or g_4900 (new_n3535_, not_new_n1862__0, not_new_n1612__3);
  or g_4901 (new_n9018_, not_new_n9002_, not_new_n8837__0);
  or g_4902 (new_n2545_, not_new_n605__3, not_new_n5487_);
  not g_4903 (not_new_n1580__968890104070, new_n1580_);
  not g_4904 (not_new_n8987__0, new_n8987_);
  not g_4905 (not_new_n1576__332329305696010, new_n1576_);
  not g_4906 (not_pi245, pi245);
  not g_4907 (new_n9063_, new_n8975_);
  not g_4908 (not_new_n6863_, new_n6863_);
  or g_4909 (new_n8190_, not_new_n8462_, not_new_n8461_);
  and g_4910 (new_n1425_, new_n2552_, new_n2550_);
  not g_4911 (new_n7640_, new_n633_);
  not g_4912 (not_new_n1474_, new_n1474_);
  or g_4913 (new_n3957_, not_new_n4066_, not_new_n4065_);
  not g_4914 (new_n8035_, new_n7725_);
  not g_4915 (not_po296_248930711762415449007872216849586085868492917169640490, po296);
  not g_4916 (not_new_n1591__138412872010, new_n1591_);
  or g_4917 (new_n3689_, not_po298_8235430, not_new_n633__9);
  not g_4918 (not_new_n8169__1, new_n8169_);
  or g_4919 (new_n2821_, not_new_n4113__2, not_new_n3310__5);
  not g_4920 (new_n5218_, new_n4998_);
  or g_4921 (new_n7254_, not_new_n7010_, not_new_n7454_);
  not g_4922 (not_new_n8806_, new_n8806_);
  not g_4923 (not_po296_725745515342319093317411710931737859674906464051430, po296);
  not g_4924 (not_new_n5754_, new_n5754_);
  not g_4925 (not_new_n5845_, new_n5845_);
  not g_4926 (not_new_n5173_, new_n5173_);
  or g_4927 (new_n9540_, not_new_n9539_, not_new_n9484_);
  or g_4928 (new_n2488_, not_new_n4120__0, not_new_n600__332329305696010);
  or g_4929 (new_n981_, not_pi003, not_new_n1536__8);
  not g_4930 (not_new_n7118_, new_n7118_);
  not g_4931 (not_new_n5366_, new_n5366_);
  or g_4932 (new_n3169_, not_new_n581__17984650426474121466202803405696493492512490, not_new_n627__6);
  not g_4933 (not_new_n8380_, new_n8380_);
  or g_4934 (new_n7535_, not_new_n7035__1, not_new_n7002__1);
  not g_4935 (not_new_n4898__2, new_n4898_);
  or g_4936 (new_n6906_, not_new_n6630_, not_new_n6803_);
  not g_4937 (not_new_n7262_, new_n7262_);
  or g_4938 (new_n3043_, not_new_n639__4, not_new_n3372__19773267430);
  not g_4939 (not_new_n8715_, new_n8715_);
  not g_4940 (not_new_n5805_, new_n5805_);
  or g_4941 (new_n7514_, not_new_n7005__0, not_new_n7037__0);
  not g_4942 (new_n6475_, new_n1043_);
  or g_4943 (new_n3947_, not_new_n3971_, not_new_n4014__1);
  not g_4944 (not_new_n8253_, new_n8253_);
  not g_4945 (not_new_n635__16284135979104490, new_n635_);
  not g_4946 (new_n4153_, new_n4147_);
  not g_4947 (not_new_n4766_, new_n4766_);
  and g_4948 (new_n1517_, and_new_n3052__new_n998_, new_n3050_);
  or g_4949 (new_n7848_, not_new_n7634_, not_new_n1604__1176490);
  not g_4950 (not_new_n989__968890104070, new_n989_);
  or g_4951 (new_n2627_, not_new_n611__168070, not_new_n2626_);
  not g_4952 (not_new_n625__47475615099430, new_n625_);
  and g_4953 (new_n10014_, new_n10281_, new_n10282_);
  or g_4954 (new_n3016_, not_new_n3372__490, not_new_n628__4);
  not g_4955 (new_n4000_, new_n3939_);
  or g_4956 (new_n5918_, not_new_n5765_, not_new_n1598__70);
  or g_4957 (new_n2854_, not_new_n4117__1, not_new_n994__168070);
  or g_4958 (new_n4884_, not_new_n4795_, not_new_n1065__7);
  not g_4959 (not_new_n4708_, new_n4708_);
  or g_4960 (new_n6674_, not_new_n1045__1176490, not_new_n6487__0);
  and g_4961 (new_n7748_, new_n8016_, new_n8015_);
  not g_4962 (not_new_n585__3430, new_n585_);
  not g_4963 (not_new_n7156_, new_n7156_);
  not g_4964 (new_n5540_, new_n5498_);
  and g_4965 (new_n1400_, new_n2485_, new_n2486_);
  not g_4966 (not_new_n6770_, new_n6770_);
  or g_4967 (new_n3593_, not_new_n944_, not_new_n1611__0);
  not g_4968 (not_new_n1473_, new_n1473_);
  or g_4969 (new_n9406_, not_new_n1069__138412872010, not_new_n646__332329305696010);
  not g_4970 (not_new_n624__8235430, new_n624_);
  and g_4971 (and_and_new_n2067__new_n2070__new_n2068_, and_new_n2067__new_n2070_, new_n2068_);
  not g_4972 (not_new_n692_, new_n692_);
  not g_4973 (not_new_n8409_, new_n8409_);
  not g_4974 (not_pi272_1, pi272);
  or g_4975 (new_n9079_, not_new_n1604__19773267430, not_new_n9078_);
  not g_4976 (not_new_n7633_, new_n7633_);
  not g_4977 (not_new_n8034_, new_n8034_);
  not g_4978 (not_new_n5081_, new_n5081_);
  or g_4979 (new_n3319_, not_new_n1534__2, not_pi059_0);
  not g_4980 (not_new_n7464_, new_n7464_);
  and g_4981 (new_n8811_, new_n9099_, new_n9093_);
  not g_4982 (not_new_n4736_, new_n4736_);
  not g_4983 (not_new_n629__2824752490, new_n629_);
  not g_4984 (new_n9413_, new_n1067_);
  or g_4985 (new_n9632_, not_new_n1597__2326305139872070, not_new_n617__39098210485829880490);
  or g_4986 (new_n4684_, not_new_n4442__0, not_pi175_3);
  not g_4987 (not_new_n589__1915812313805664144010, new_n589_);
  not g_4988 (not_new_n5864_, new_n5864_);
  not g_4989 (new_n3324_, new_n1000_);
  not g_4990 (not_new_n609__70, new_n609_);
  not g_4991 (not_new_n4390_, new_n4390_);
  not g_4992 (not_new_n1591__403536070, new_n1591_);
  not g_4993 (new_n5096_, new_n4930_);
  not g_4994 (not_new_n7260_, new_n7260_);
  not g_4995 (not_new_n2875_, new_n2875_);
  not g_4996 (not_new_n8821_, new_n8821_);
  not g_4997 (not_new_n646__70, new_n646_);
  or g_4998 (new_n8051_, not_new_n7656__0, not_new_n1063__1176490);
  not g_4999 (not_new_n9883_, new_n9883_);
  not g_5000 (not_new_n9872_, new_n9872_);
  or g_5001 (or_not_new_n1996__not_new_n1997_, not_new_n1997_, not_new_n1996_);
  and g_5002 (new_n6623_, new_n6879_, new_n6878_);
  xor g_5003 (key_gate_33, new_n1714_, key_33);
  or g_5004 (new_n3271_, not_new_n1602__5, not_new_n589__1577753820348458066150427430);
  not g_5005 (new_n4439_, pi174);
  or g_5006 (new_n4338_, not_new_n4236_, not_new_n673_);
  or g_5007 (new_n4402_, not_new_n4399_, not_new_n4317_);
  not g_5008 (not_new_n3375__4, new_n3375_);
  not g_5009 (not_new_n619__0, new_n619_);
  not g_5010 (not_new_n1035__0, new_n1035_);
  or g_5011 (new_n3115_, not_new_n618__5, not_new_n581__11044276742439206463052992010);
  not g_5012 (new_n4413_, new_n1020_);
  or g_5013 (new_n7827_, not_new_n7825_, not_new_n7826_);
  or g_5014 (new_n1737_, not_pi081, not_new_n1728__5);
  not g_5015 (not_new_n4750__0, new_n4750_);
  or g_5016 (new_n4062_, not_new_n3988_, not_new_n4034_);
  not g_5017 (new_n4949_, new_n617_);
  not g_5018 (new_n2313_, new_n980_);
  or g_5019 (new_n7517_, not_new_n7234_, not_new_n7515_);
  or g_5020 (new_n10026_, not_new_n9931_, not_new_n10216_);
  not g_5021 (not_new_n8955_, new_n8955_);
  not g_5022 (not_new_n8262__1, new_n8262_);
  not g_5023 (new_n8851_, new_n1598_);
  not g_5024 (not_new_n9111_, new_n9111_);
  or g_5025 (new_n2121_, not_new_n8916_, not_new_n1591__8235430);
  not g_5026 (not_pi037_2, pi037);
  and g_5027 (and_new_n4298__new_n4341_, new_n4341_, new_n4298_);
  and g_5028 (new_n1376_, new_n2426_, new_n2425_);
  and g_5029 (and_new_n4327__new_n4331_, new_n4327_, new_n4331_);
  not g_5030 (not_new_n639_, new_n639_);
  or g_5031 (new_n7545_, not_new_n7543_, not_new_n7331_);
  not g_5032 (new_n7611_, new_n635_);
  not g_5033 (not_new_n5241_, new_n5241_);
  not g_5034 (not_new_n5853_, new_n5853_);
  not g_5035 (not_pi266_2, pi266);
  or g_5036 (or_not_new_n999__1_not_new_n3377_, not_new_n3377_, not_new_n999__1);
  and g_5037 (new_n7147_, new_n7519_, new_n7518_);
  not g_5038 (not_new_n606__1176490, new_n606_);
  and g_5039 (new_n1271_, and_new_n1270__new_n1989_, new_n1988_);
  or g_5040 (new_n3242_, not_new_n1031__7, not_new_n3185__2326305139872070);
  or g_5041 (or_or_or_not_new_n2973__not_new_n2976__not_new_n2975__not_new_n2977_, or_or_not_new_n2973__not_new_n2976__not_new_n2975_, not_new_n2977_);
  not g_5042 (not_new_n605__70, new_n605_);
  or g_5043 (new_n9015_, new_n1045_, new_n635_);
  not g_5044 (not_new_n625__968890104070, new_n625_);
  not g_5045 (not_new_n1591__4, new_n1591_);
  not g_5046 (new_n4786_, new_n1031_);
  not g_5047 (not_new_n5223_, new_n5223_);
  not g_5048 (not_new_n8595__2, new_n8595_);
  or g_5049 (new_n6142_, not_new_n6138__0, not_new_n5912__0);
  not g_5050 (not_pi096, pi096);
  not g_5051 (not_pi064_9, pi064);
  or g_5052 (new_n4039_, not_pi051_3, not_new_n3947_);
  not g_5053 (new_n9927_, new_n1059_);
  not g_5054 (not_new_n581__63668057609090279857414351392240010, new_n581_);
  or g_5055 (new_n5966_, not_new_n5847_, not_new_n6079_);
  not g_5056 (not_new_n8833_, new_n8833_);
  not g_5057 (new_n10061_, new_n9899_);
  or g_5058 (new_n9499_, not_new_n1031__2824752490, not_new_n641__2824752490);
  not g_5059 (not_new_n7639__0, new_n7639_);
  not g_5060 (not_new_n6023__0, new_n6023_);
  or g_5061 (new_n9783_, not_new_n9781_, not_new_n9624_);
  not g_5062 (not_new_n4329_, new_n4329_);
  not g_5063 (not_new_n7649_, new_n7649_);
  not g_5064 (not_new_n1606__3, new_n1606_);
  not g_5065 (not_new_n6606_, new_n6606_);
  or g_5066 (new_n2193_, not_new_n1585__19773267430, not_new_n5832_);
  or g_5067 (or_or_not_new_n1235__not_new_n1233__not_new_n1812_, or_not_new_n1235__not_new_n1233_, not_new_n1812_);
  not g_5068 (not_new_n5542_, new_n5542_);
  not g_5069 (not_new_n1612__19773267430, new_n1612_);
  not g_5070 (not_new_n1584__57648010, new_n1584_);
  and g_5071 (and_new_n2010__new_n2013_, new_n2010_, new_n2013_);
  not g_5072 (not_new_n4249_, new_n4249_);
  not g_5073 (not_new_n637__113988951853731430, new_n637_);
  not g_5074 (not_new_n1043__403536070, new_n1043_);
  not g_5075 (not_new_n617__10, new_n617_);
  not g_5076 (not_new_n1602__968890104070, new_n1602_);
  not g_5077 (not_new_n4363_, new_n4363_);
  not g_5078 (not_new_n9519__0, new_n9519_);
  not g_5079 (not_new_n1004__4, new_n1004_);
  not g_5080 (new_n8652_, new_n1606_);
  and g_5081 (new_n6461_, new_n6896_, new_n6545_);
  not g_5082 (not_new_n3311__1176490, new_n3311_);
  not g_5083 (not_new_n5574_, new_n5574_);
  not g_5084 (not_new_n4605_, new_n4605_);
  not g_5085 (not_new_n5080_, new_n5080_);
  not g_5086 (new_n8882_, new_n637_);
  not g_5087 (not_new_n1067__8235430, new_n1067_);
  not g_5088 (not_pi049_3, pi049);
  not g_5089 (not_new_n4483_, new_n4483_);
  not g_5090 (not_new_n6174_, new_n6174_);
  not g_5091 (not_new_n6949_, new_n6949_);
  not g_5092 (not_po296_490, po296);
  not g_5093 (not_new_n9702_, new_n9702_);
  not g_5094 (not_new_n5866_, new_n5866_);
  and g_5095 (new_n6335_, new_n6232_, new_n6267_);
  not g_5096 (not_new_n8002_, new_n8002_);
  not g_5097 (not_new_n7959_, new_n7959_);
  or g_5098 (new_n2232_, not_new_n9440_, not_new_n1584__968890104070);
  not g_5099 (not_new_n3914_, new_n3914_);
  not g_5100 (not_new_n6976__2, new_n6976_);
  not g_5101 (not_new_n3740_, new_n3740_);
  not g_5102 (not_new_n597__6782230728490, new_n597_);
  or g_5103 (new_n6141_, not_new_n6139_, or_not_new_n5766__1_not_new_n6140_);
  xor g_5104 (key_gate_123, key_123, not_new_n1684_);
  not g_5105 (not_new_n5216_, new_n5216_);
  or g_5106 (new_n10123_, not_new_n9905_, not_new_n9906_);
  not g_5107 (not_po298_113988951853731430, po298);
  not g_5108 (not_new_n6974__24010, new_n6974_);
  not g_5109 (not_pi265_4, pi265);
  not g_5110 (not_new_n5489_, new_n5489_);
  not g_5111 (not_new_n4322_, new_n4322_);
  not g_5112 (not_new_n3911_, new_n3911_);
  not g_5113 (not_new_n7334_, new_n7334_);
  not g_5114 (not_new_n6553_, new_n6553_);
  not g_5115 (not_new_n4086_, new_n4086_);
  not g_5116 (not_new_n6897_, new_n6897_);
  and g_5117 (new_n1368_, new_n2405_, new_n2406_);
  not g_5118 (new_n6133_, new_n5858_);
  not g_5119 (not_new_n7104_, new_n7104_);
  not g_5120 (not_new_n3373_, new_n3373_);
  not g_5121 (not_new_n5171_, new_n5171_);
  not g_5122 (not_new_n5178_, new_n5178_);
  not g_5123 (not_new_n1537__9, new_n1537_);
  or g_5124 (new_n3135_, not_new_n928__1176490, not_new_n1603__3);
  not g_5125 (not_pi163_2, pi163);
  not g_5126 (not_new_n2595_, new_n2595_);
  or g_5127 (new_n4531_, not_new_n4530_, not_new_n4479_);
  not g_5128 (not_new_n9463_, new_n9463_);
  not g_5129 (not_new_n744__1, new_n744_);
  not g_5130 (not_pi064_490, pi064);
  not g_5131 (not_new_n9234_, new_n9234_);
  not g_5132 (not_new_n3313_, new_n3313_);
  or g_5133 (new_n8984_, not_new_n622__6782230728490, not_new_n1599__2824752490);
  or g_5134 (new_n5328_, not_new_n5060_, not_new_n5061_);
  or g_5135 (new_n2070_, not_new_n1588__168070, not_new_n1063_);
  not g_5136 (not_new_n1065__490, new_n1065_);
  and g_5137 (and_new_n5582__new_n5648_, new_n5582_, new_n5648_);
  not g_5138 (not_new_n7961_, new_n7961_);
  not g_5139 (not_new_n8248__1, new_n8248_);
  not g_5140 (not_new_n9989_, new_n9989_);
  not g_5141 (not_new_n994__1176490, new_n994_);
  not g_5142 (not_new_n635__9, new_n635_);
  or g_5143 (new_n1904_, not_new_n585__7, not_new_n4114_);
  or g_5144 (new_n2815_, not_pi255_3, not_po296_17984650426474121466202803405696493492512490);
  not g_5145 (not_pi092, pi092);
  not g_5146 (not_new_n8995_, new_n8995_);
  not g_5147 (not_new_n591__138412872010, new_n591_);
  not g_5148 (not_new_n4465__0, new_n4465_);
  not g_5149 (not_new_n630__8, new_n630_);
  or g_5150 (new_n9503_, not_new_n9399_, not_new_n9701_);
  not g_5151 (not_new_n2883_, new_n2883_);
  not g_5152 (not_new_n9140__0, new_n9140_);
  or g_5153 (new_n3836_, not_new_n631__490, not_new_n1576__3);
  or g_5154 (new_n7269_, not_new_n7010__0, not_new_n7454__0);
  not g_5155 (not_new_n1576__113988951853731430, new_n1576_);
  or g_5156 (new_n3051_, not_new_n1027__968890104070, not_new_n1169_);
  not g_5157 (not_new_n1065__9, new_n1065_);
  not g_5158 (not_new_n1059__9, new_n1059_);
  or g_5159 (new_n2355_, not_new_n1031__2, not_new_n598_);
  not g_5160 (not_new_n4697_, new_n4697_);
  not g_5161 (not_new_n627__1176490, new_n627_);
  or g_5162 (new_n7978_, not_new_n632__138412872010, not_new_n7607__0);
  not g_5163 (not_new_n617__8, new_n617_);
  not g_5164 (not_new_n9283_, new_n9283_);
  not g_5165 (not_new_n6619__0, new_n6619_);
  not g_5166 (not_new_n3346_, new_n3346_);
  or g_5167 (new_n8028_, not_new_n7609_, not_new_n1035__70);
  and g_5168 (and_new_n6385__new_n6386_, new_n6385_, new_n6386_);
  not g_5169 (new_n9877_, new_n635_);
  not g_5170 (not_new_n1585__403536070, new_n1585_);
  or g_5171 (new_n5484_, not_new_n5658_, not_new_n5657_);
  not g_5172 (not_new_n2211_, new_n2211_);
  not g_5173 (not_new_n602__1, new_n602_);
  not g_5174 (not_new_n3153_, new_n3153_);
  not g_5175 (not_new_n1602__57648010, new_n1602_);
  not g_5176 (not_new_n6877_, new_n6877_);
  not g_5177 (not_new_n5181_, new_n5181_);
  not g_5178 (not_new_n5030_, new_n5030_);
  not g_5179 (not_new_n1007__7, new_n1007_);
  not g_5180 (new_n8445_, new_n8273_);
  or g_5181 (or_or_not_new_n3965__not_new_n3966__not_new_n3968_, not_new_n3968_, or_not_new_n3965__not_new_n3966_);
  or g_5182 (new_n7017_, not_new_n7292_, not_new_n6997_);
  not g_5183 (new_n4541_, new_n4473_);
  not g_5184 (not_new_n10156__0, new_n10156_);
  not g_5185 (not_new_n2733_, new_n2733_);
  not g_5186 (not_new_n610__0, new_n610_);
  not g_5187 (not_new_n7322_, new_n7322_);
  not g_5188 (not_new_n2746_, new_n2746_);
  not g_5189 (not_new_n3825_, new_n3825_);
  not g_5190 (not_new_n1631__57648010, key_gate_76);
  or g_5191 (new_n7272_, not_new_n7267__0, not_new_n7089_);
  not g_5192 (new_n7244_, new_n7143_);
  not g_5193 (not_new_n1430_, new_n1430_);
  not g_5194 (not_new_n4795_, new_n4795_);
  not g_5195 (not_new_n8447_, new_n8447_);
  or g_5196 (new_n7408_, not_new_n763_, not_new_n6974__10);
  or g_5197 (new_n5757_, not_new_n624__168070, not_new_n5744_);
  or g_5198 (new_n7949_, not_new_n647__19773267430, not_new_n7616__0);
  not g_5199 (not_new_n6242__0, new_n6242_);
  or g_5200 (or_or_not_new_n1315__not_new_n1313__not_new_n2192_, not_new_n2192_, or_not_new_n1315__not_new_n1313_);
  or g_5201 (or_not_new_n6226__0_not_new_n6336_, not_new_n6336_, not_new_n6226__0);
  or g_5202 (new_n6013_, not_new_n5807_, not_new_n6012_);
  not g_5203 (new_n9591_, new_n9503_);
  not g_5204 (new_n9530_, new_n9373_);
  not g_5205 (not_new_n7791_, new_n7791_);
  not g_5206 (not_new_n8593__0, new_n8593_);
  or g_5207 (new_n3194_, not_new_n3185__3, not_new_n1043__4);
  not g_5208 (not_new_n5073_, new_n5073_);
  not g_5209 (not_new_n2509__6, new_n2509_);
  or g_5210 (new_n6847_, not_new_n6691__0, not_new_n6615_);
  and g_5211 (new_n1227_, new_n1762_, new_n3401_);
  or g_5212 (new_n2157_, not_new_n1581__403536070, not_new_n8183_);
  not g_5213 (not_new_n5450_, new_n5450_);
  not g_5214 (not_new_n7631_, new_n7631_);
  or g_5215 (new_n3057_, not_new_n1171_, not_new_n1027__47475615099430);
  not g_5216 (not_new_n1045__168070, new_n1045_);
  or g_5217 (new_n5425_, not_new_n1031__490, not_new_n4932_);
  or g_5218 (new_n6086_, not_new_n6085_, not_new_n5888_);
  or g_5219 (new_n1853_, not_new_n1581__3, not_new_n8193_);
  or g_5220 (new_n8740_, not_new_n1150__0, not_new_n8603_);
  not g_5221 (not_new_n1583_, new_n1583_);
  not g_5222 (not_pi129_3, pi129);
  and g_5223 (new_n1387_, new_n2452_, new_n2453_);
  and g_5224 (new_n1522_, new_n3065_, and_new_n3067__new_n998_);
  not g_5225 (not_new_n6711_, new_n6711_);
  not g_5226 (new_n9096_, new_n8966_);
  not g_5227 (not_new_n2301_, new_n2301_);
  or g_5228 (new_n4135_, not_new_n4221_, not_new_n4222_);
  not g_5229 (not_new_n8343_, new_n8343_);
  or g_5230 (new_n4045_, not_pi046_2, not_new_n4044_);
  not g_5231 (not_pi054_2, pi054);
  not g_5232 (not_new_n636__24010, new_n636_);
  not g_5233 (not_new_n1203_, new_n1203_);
  not g_5234 (not_new_n622__113988951853731430, new_n622_);
  not g_5235 (not_new_n10061__0, new_n10061_);
  or g_5236 (new_n736_, not_new_n3246_, not_new_n3245_);
  not g_5237 (not_new_n585__10, new_n585_);
  or g_5238 (new_n4096_, not_pi268_1, not_new_n4166_);
  or g_5239 (new_n7935_, not_new_n7579_, not_new_n7735__0);
  not g_5240 (not_new_n5002_, new_n5002_);
  or g_5241 (new_n5121_, new_n1045_, new_n635_);
  not g_5242 (not_new_n9871__0, new_n9871_);
  not g_5243 (not_new_n1186_, new_n1186_);
  not g_5244 (not_new_n9594_, new_n9594_);
  not g_5245 (not_new_n6068_, new_n6068_);
  not g_5246 (not_new_n7720_, new_n7720_);
  not g_5247 (not_new_n1037__332329305696010, new_n1037_);
  xor g_5248 (key_gate_17, key_17, not_new_n3992_);
  not g_5249 (not_new_n3345_, new_n3345_);
  or g_5250 (or_or_or_not_new_n2964__not_new_n2967__not_new_n2966__not_new_n2968_, or_or_not_new_n2964__not_new_n2967__not_new_n2966_, not_new_n2968_);
  or g_5251 (new_n5412_, not_new_n636__168070, not_new_n4962_);
  or g_5252 (new_n2793_, or_not_new_n2792__not_new_n2791_, not_new_n2790_);
  or g_5253 (new_n4346_, not_new_n701_, not_new_n4249_);
  not g_5254 (not_new_n3184__490, new_n3184_);
  not g_5255 (not_new_n9048_, new_n9048_);
  not g_5256 (not_new_n5011_, new_n5011_);
  or g_5257 (new_n5500_, not_new_n5534_, not_new_n5535_);
  not g_5258 (not_new_n1210_, new_n1210_);
  or g_5259 (new_n2683_, not_new_n4411_, not_new_n609__8235430);
  not g_5260 (not_new_n3662_, new_n3662_);
  or g_5261 (po270, not_new_n2759_, or_or_or_not_new_n2758__not_new_n2761__not_new_n2760__not_new_n2762_);
  not g_5262 (not_new_n5730_, new_n5730_);
  not g_5263 (not_new_n629__490, new_n629_);
  and g_5264 (new_n4501_, new_n4689_, new_n4688_);
  or g_5265 (new_n2464_, not_new_n9966__0, not_new_n599__19773267430);
  not g_5266 (not_new_n595__47475615099430, new_n595_);
  not g_5267 (not_new_n3730_, new_n3730_);
  not g_5268 (not_new_n1008__4, new_n1008_);
  not g_5269 (not_new_n7769__0, new_n7769_);
  not g_5270 (not_new_n1024__3, new_n1024_);
  or g_5271 (or_not_new_n2645__not_new_n2644_, not_new_n2645_, not_new_n2644_);
  or g_5272 (or_or_not_new_n2151__not_new_n2148__not_new_n2149_, or_not_new_n2151__not_new_n2148_, not_new_n2149_);
  or g_5273 (new_n2351_, not_new_n2350_, not_new_n985_);
  not g_5274 (not_new_n1584_, new_n1584_);
  not g_5275 (not_new_n591__5, new_n591_);
  not g_5276 (not_new_n3441_, new_n3441_);
  not g_5277 (not_new_n7023__1, new_n7023_);
  or g_5278 (po130, not_new_n3466_, not_new_n3465_);
  not g_5279 (not_new_n5526_, new_n5526_);
  not g_5280 (not_new_n6496_, new_n6496_);
  or g_5281 (or_not_new_n2343__not_new_n2344_, not_new_n2344_, not_new_n2343_);
  not g_5282 (not_new_n5986_, new_n5986_);
  or g_5283 (new_n3383_, not_new_n3922__0, not_pi064_2326305139872070);
  or g_5284 (new_n710_, not_new_n3048_, not_new_n1516_);
  not g_5285 (not_new_n10020_, new_n10020_);
  not g_5286 (not_new_n4121__2, new_n4121_);
  not g_5287 (new_n3494_, new_n1069_);
  not g_5288 (new_n5269_, new_n4939_);
  or g_5289 (new_n1752_, not_new_n1728__2824752490, not_pi095);
  not g_5290 (new_n10110_, new_n9951_);
  or g_5291 (new_n702_, not_new_n3078_, not_new_n1526_);
  not g_5292 (not_new_n6737_, new_n6737_);
  and g_5293 (new_n7149_, new_n7532_, new_n7533_);
  and g_5294 (new_n7570_, new_n7788_, new_n7787_);
  not g_5295 (not_new_n7421__0, new_n7421_);
  not g_5296 (not_new_n3687_, new_n3687_);
  and g_5297 (new_n6332_, new_n6373_, new_n6256_);
  or g_5298 (new_n3292_, not_new_n644__8, not_new_n3184__138412872010);
  not g_5299 (not_new_n1256_, new_n1256_);
  not g_5300 (not_new_n1350_, new_n1350_);
  or g_5301 (new_n5930_, not_new_n5749__0, not_new_n5748_);
  or g_5302 (new_n2186_, not_pi184, not_new_n586__138412872010);
  not g_5303 (not_pi269_4, pi269);
  or g_5304 (new_n7381_, not_new_n6990__0, not_new_n7301_);
  or g_5305 (new_n10159_, not_new_n10158_, not_new_n9995_);
  not g_5306 (not_pi267, pi267);
  not g_5307 (not_new_n4347_, new_n4347_);
  or g_5308 (new_n5661_, not_new_n5470__0, not_new_n1012__7);
  not g_5309 (not_new_n1588__273687473400809163430, new_n1588_);
  or g_5310 (new_n2875_, not_new_n612__3, not_new_n4122__2);
  not g_5311 (not_new_n7598_, new_n7598_);
  and g_5312 (new_n1564_, new_n3640_, new_n3641_);
  not g_5313 (not_pi029, pi029);
  not g_5314 (not_new_n5122_, new_n5122_);
  not g_5315 (not_new_n9428_, new_n9428_);
  or g_5316 (new_n9325_, not_new_n1031__403536070, not_new_n8832_);
  not g_5317 (not_new_n5329_, new_n5329_);
  not g_5318 (not_new_n5801_, new_n5801_);
  not g_5319 (not_new_n8038_, new_n8038_);
  or g_5320 (new_n9613_, not_new_n9610_, or_not_new_n9612__not_new_n9611_);
  not g_5321 (not_new_n1453_, new_n1453_);
  not g_5322 (not_new_n9374__0, new_n9374_);
  not g_5323 (not_new_n626__138412872010, new_n626_);
  not g_5324 (not_new_n9472_, new_n9472_);
  buf g_5325 (po006, pi199);
  and g_5326 (new_n8940_, new_n9091_, new_n9183_);
  or g_5327 (new_n10291_, not_new_n1599__47475615099430, not_new_n9937_);
  not g_5328 (not_new_n984__4, new_n984_);
  or g_5329 (new_n6380_, not_new_n6278_, not_new_n1601__168070);
  not g_5330 (not_new_n6471_, new_n6471_);
  not g_5331 (new_n2199_, new_n968_);
  not g_5332 (not_new_n1153_, new_n1153_);
  or g_5333 (new_n6019_, not_new_n5774__0, not_new_n625__8235430);
  not g_5334 (not_new_n6784_, new_n6784_);
  not g_5335 (not_pi225, pi225);
  not g_5336 (not_new_n625__1915812313805664144010, new_n625_);
  not g_5337 (not_new_n1367_, new_n1367_);
  not g_5338 (not_new_n6980_, new_n6980_);
  not g_5339 (new_n1981_, new_n636_);
  and g_5340 (and_new_n2682__new_n2681_, new_n2682_, new_n2681_);
  and g_5341 (new_n10010_, new_n10268_, new_n10267_);
  not g_5342 (not_new_n2974_, new_n2974_);
  not g_5343 (not_new_n7411_, new_n7411_);
  not g_5344 (not_new_n1537__5, new_n1537_);
  not g_5345 (not_new_n3387__3, new_n3387_);
  not g_5346 (not_new_n1467_, new_n1467_);
  not g_5347 (not_new_n8829__0, new_n8829_);
  not g_5348 (not_new_n5483_, new_n5483_);
  or g_5349 (new_n3100_, not_new_n624__5, not_new_n3315__6);
  not g_5350 (not_po296_3119734822845423713013303218219760490, po296);
  not g_5351 (not_new_n1031__2824752490, new_n1031_);
  or g_5352 (new_n10106_, not_new_n643__273687473400809163430, not_new_n1061__16284135979104490);
  or g_5353 (new_n2758_, not_new_n3311__1, not_new_n1069__1);
  not g_5354 (not_new_n1728__138412872010, new_n1728_);
  not g_5355 (not_pi137_1, pi137);
  not g_5356 (not_new_n626__403536070, new_n626_);
  not g_5357 (not_pi057_2, pi057);
  or g_5358 (new_n9965_, not_new_n10305_, not_new_n10306_);
  or g_5359 (new_n4520_, not_pi164_1, not_new_n1008__2);
  not g_5360 (not_new_n5218__0, new_n5218_);
  not g_5361 (not_pi264_1, pi264);
  not g_5362 (not_new_n2930_, new_n2930_);
  or g_5363 (or_not_new_n1863__not_new_n1864_, not_new_n1864_, not_new_n1863_);
  not g_5364 (not_new_n2780_, new_n2780_);
  or g_5365 (new_n2234_, not_new_n6551_, not_new_n1580__6782230728490);
  not g_5366 (not_new_n645__47475615099430, new_n645_);
  or g_5367 (new_n7873_, not_new_n7872_, not_new_n7717_);
  not g_5368 (not_new_n7060_, new_n7060_);
  not g_5369 (not_new_n587__2824752490, new_n587_);
  and g_5370 (new_n8673_, new_n8592_, new_n8672_);
  not g_5371 (not_new_n639__113988951853731430, new_n639_);
  not g_5372 (not_new_n631__657123623635342801395430, new_n631_);
  not g_5373 (not_new_n5462_, new_n5462_);
  not g_5374 (not_new_n8175__0, new_n8175_);
  not g_5375 (not_new_n5485__0, new_n5485_);
  not g_5376 (not_new_n1401_, new_n1401_);
  and g_5377 (new_n7740_, new_n7978_, new_n7977_);
  or g_5378 (new_n7592_, not_new_n7819_, not_new_n7944_);
  not g_5379 (not_new_n2760_, new_n2760_);
  not g_5380 (not_new_n609__4, new_n609_);
  not g_5381 (not_new_n7213_, new_n7213_);
  not g_5382 (not_new_n7741_, new_n7741_);
  or g_5383 (new_n9763_, not_new_n9490_, not_new_n9491__1);
  not g_5384 (not_pi063, pi063);
  not g_5385 (not_new_n9385_, new_n9385_);
  or g_5386 (new_n3152_, not_new_n3315__138412872010, not_new_n637__5);
  or g_5387 (new_n5361_, not_new_n5067_, not_new_n4988__0);
  not g_5388 (not_new_n632__273687473400809163430, new_n632_);
  or g_5389 (new_n4698_, not_new_n4438__0, not_pi173_3);
  or g_5390 (new_n1747_, not_new_n1728__168070, not_pi091);
  or g_5391 (new_n3232_, not_new_n1059__4, not_new_n3185__138412872010);
  or g_5392 (new_n6083_, not_new_n5720__0, not_new_n5890__1);
  or g_5393 (new_n8099_, not_new_n8453_, not_new_n8332_);
  or g_5394 (new_n3217_, not_new_n640__7, not_new_n589__24010);
  not g_5395 (not_new_n9968_, new_n9968_);
  not g_5396 (not_pi141, pi141);
  not g_5397 (not_new_n7457__0, new_n7457_);
  or g_5398 (new_n5320_, not_new_n5137_, not_new_n5318_);
  not g_5399 (not_new_n3923__0, new_n3923_);
  or g_5400 (new_n9085_, or_not_new_n9084__not_new_n9083_, not_new_n9082_);
  not g_5401 (not_new_n585__19773267430, new_n585_);
  or g_5402 (new_n5629_, not_new_n5435__0, not_pi132_2);
  not g_5403 (not_new_n6572_, new_n6572_);
  not g_5404 (not_new_n7920_, new_n7920_);
  or g_5405 (new_n5936_, not_new_n5920_, not_new_n5924_);
  and g_5406 (and_new_n6251__new_n6371_, new_n6371_, new_n6251_);
  or g_5407 (new_n4657_, not_new_n4656_, not_new_n4655_);
  or g_5408 (new_n2940_, not_new_n595__138412872010, not_new_n6972_);
  not g_5409 (not_new_n1041__6782230728490, new_n1041_);
  not g_5410 (not_new_n1049__3430, new_n1049_);
  not g_5411 (not_new_n4136__2, new_n4136_);
  or g_5412 (new_n2953_, not_new_n4124__1, not_new_n994__332329305696010);
  not g_5413 (not_new_n629__2326305139872070, new_n629_);
  not g_5414 (not_new_n10152_, new_n10152_);
  and g_5415 (new_n4294_, new_n4335_, and_and_new_n4295__new_n4334__new_n4338_);
  not g_5416 (not_new_n6186_, new_n6186_);
  or g_5417 (new_n3398_, not_new_n1024__3, not_new_n3372__93874803376477543056490);
  not g_5418 (not_new_n8125_, new_n8125_);
  not g_5419 (not_new_n9511_, new_n9511_);
  not g_5420 (not_new_n4462_, new_n4462_);
  or g_5421 (new_n10183_, not_new_n10029__1, not_new_n10100_);
  or g_5422 (new_n4846_, new_n1031_, new_n1035_);
  not g_5423 (not_new_n928__19773267430, new_n928_);
  not g_5424 (new_n8133_, new_n1600_);
  not g_5425 (not_new_n6701_, new_n6701_);
  or g_5426 (new_n7845_, not_new_n7639_, not_new_n1069__1176490);
  not g_5427 (not_new_n9142_, new_n9142_);
  or g_5428 (new_n7851_, not_new_n7630_, not_new_n630__2824752490);
  not g_5429 (not_new_n5073__0, new_n5073_);
  not g_5430 (new_n9414_, new_n1601_);
  not g_5431 (not_new_n1059__19773267430, new_n1059_);
  not g_5432 (not_new_n597__0, new_n597_);
  not g_5433 (not_new_n6700_, new_n6700_);
  not g_5434 (not_new_n6545_, new_n6545_);
  or g_5435 (new_n995_, not_new_n590__1, not_new_n582__0);
  not g_5436 (not_new_n588__16284135979104490, new_n588_);
  not g_5437 (not_new_n593__6782230728490, new_n593_);
  not g_5438 (not_new_n10299_, new_n10299_);
  and g_5439 (new_n1459_, new_n3786_, and_and_new_n3780__new_n3783__new_n3789_);
  not g_5440 (not_new_n6159__0, new_n6159_);
  not g_5441 (not_new_n8109__0, new_n8109_);
  not g_5442 (new_n7180_, new_n6980_);
  not g_5443 (not_new_n1596__1176490, new_n1596_);
  or g_5444 (new_n8527_, not_new_n8525_, not_new_n8526_);
  or g_5445 (new_n977_, not_new_n1536__6, not_pi005);
  not g_5446 (not_new_n8979__0, new_n8979_);
  not g_5447 (not_pi042_3, pi042);
  not g_5448 (not_new_n4519_, new_n4519_);
  not g_5449 (not_new_n587__9, new_n587_);
  not g_5450 (not_new_n10326_, new_n10326_);
  not g_5451 (not_new_n10184__0, new_n10184_);
  or g_5452 (new_n5351_, not_new_n629__24010, not_new_n4952_);
  or g_5453 (new_n7438_, not_new_n6974__2824752490, not_new_n754_);
  not g_5454 (not_new_n4350_, new_n4350_);
  or g_5455 (new_n9493_, not_new_n9472_, not_new_n9629_);
  not g_5456 (not_new_n5362_, new_n5362_);
  or g_5457 (new_n2617_, not_new_n611__24010, not_new_n2616_);
  not g_5458 (new_n6648_, new_n6481_);
  or g_5459 (new_n10168_, not_new_n10124__0, not_new_n10166__0);
  or g_5460 (new_n2181_, not_new_n594__2824752490, not_new_n9871_);
  or g_5461 (new_n2091_, not_new_n586__8235430, not_pi179);
  not g_5462 (not_new_n8513_, new_n8513_);
  or g_5463 (new_n10127_, or_not_new_n10126__not_new_n10125_, not_new_n10124_);
  or g_5464 (or_or_not_new_n2883__not_new_n2886__not_new_n2885_, not_new_n2885_, or_not_new_n2883__not_new_n2886_);
  xnor g_5465 (key_gate_24, new_n1702_, key_24);
  or g_5466 (new_n726_, not_new_n3280_, not_new_n3279_);
  not g_5467 (not_new_n1611__5, new_n1611_);
  not g_5468 (not_new_n1065__16284135979104490, new_n1065_);
  or g_5469 (new_n8766_, not_new_n8645_, not_new_n1602__2824752490);
  and g_5470 (new_n4497_, new_n4674_, new_n4675_);
  and g_5471 (new_n8697_, new_n1601_, new_n8646_);
  not g_5472 (not_new_n1626__1, new_n1626_);
  not g_5473 (not_new_n644__70, new_n644_);
  or g_5474 (po129, not_new_n3460_, not_new_n3461_);
  not g_5475 (not_po296_1299348114471230201171721456984490, po296);
  or g_5476 (new_n3161_, not_new_n644__5, not_new_n3315__47475615099430);
  not g_5477 (not_new_n6529__0, new_n6529_);
  or g_5478 (new_n10140_, new_n1599_, new_n622_);
  not g_5479 (not_new_n1405_, new_n1405_);
  not g_5480 (not_new_n3587_, new_n3587_);
  not g_5481 (not_new_n8634_, new_n8634_);
  or g_5482 (new_n2962_, not_new_n4133__1, not_new_n994__2326305139872070);
  or g_5483 (new_n8982_, not_new_n647__6782230728490, not_new_n1051__2824752490);
  or g_5484 (new_n8074_, not_new_n7672__0, not_new_n7904_);
  or g_5485 (or_not_new_n1331__not_new_n1329_, not_new_n1329_, not_new_n1331_);
  not g_5486 (not_pi202, pi202);
  not g_5487 (not_new_n10203_, new_n10203_);
  not g_5488 (not_new_n2509__10, new_n2509_);
  or g_5489 (new_n8348_, not_new_n8079_, not_new_n8288_);
  not g_5490 (not_new_n7647__0, new_n7647_);
  not g_5491 (not_pi272_0, pi272);
  not g_5492 (new_n9606_, new_n9402_);
  not g_5493 (not_new_n1591__8, new_n1591_);
  or g_5494 (new_n2444_, not_new_n599__8235430, not_new_n9968__0);
  and g_5495 (new_n1488_, new_n2993_, and_new_n2995__new_n998_);
  or g_5496 (new_n634_, not_new_n1884_, or_or_not_new_n1882__not_new_n1883__not_new_n1885_);
  and g_5497 (new_n8816_, new_n9120_, new_n9122_);
  and g_5498 (new_n1383_, new_n2443_, new_n2442_);
  or g_5499 (new_n9099_, new_n1600_, new_n629_);
  not g_5500 (not_new_n9990_, new_n9990_);
  or g_5501 (or_not_new_n8221__not_new_n8220_, not_new_n8220_, not_new_n8221_);
  not g_5502 (new_n8622_, new_n1169_);
  not g_5503 (new_n7600_, new_n1045_);
  not g_5504 (not_new_n1594__5, new_n1594_);
  not g_5505 (not_new_n643__6, new_n643_);
  not g_5506 (not_new_n10291_, new_n10291_);
  or g_5507 (new_n1160_, not_new_n3850_, not_new_n3849_);
  not g_5508 (not_new_n7794_, new_n7794_);
  or g_5509 (new_n9623_, not_new_n630__2326305139872070, not_new_n1601__5585458640832840070);
  and g_5510 (new_n614_, new_n922_, new_n3315_);
  not g_5511 (not_new_n3337_, new_n3337_);
  not g_5512 (not_new_n1597__5585458640832840070, new_n1597_);
  not g_5513 (not_new_n7346_, new_n7346_);
  not g_5514 (not_new_n9857_, new_n9857_);
  not g_5515 (not_new_n600__47475615099430, new_n600_);
  not g_5516 (not_new_n8940_, new_n8940_);
  not g_5517 (not_new_n6323_, new_n6323_);
  not g_5518 (not_new_n4428_, new_n4428_);
  and g_5519 (new_n8801_, new_n9044_, new_n9043_);
  not g_5520 (not_new_n8124_, new_n8124_);
  not g_5521 (not_po296_657123623635342801395430, po296);
  and g_5522 (new_n1351_, and_new_n2364__new_n2363_, new_n2362_);
  or g_5523 (new_n7993_, not_new_n7663__1, not_new_n1597__57648010);
  not g_5524 (not_new_n1049__113988951853731430, new_n1049_);
  not g_5525 (not_new_n4775_, new_n4775_);
  or g_5526 (new_n2018_, not_new_n4133_, not_new_n585__3430);
  or g_5527 (new_n665_, not_new_n3156_, or_not_new_n3158__not_new_n3157_);
  not g_5528 (not_new_n5754__0, new_n5754_);
  not g_5529 (new_n7105_, new_n766_);
  not g_5530 (not_new_n9620__0, new_n9620_);
  and g_5531 (new_n1247_, and_new_n1246__new_n1875_, new_n1874_);
  not g_5532 (new_n4932_, new_n641_);
  not g_5533 (not_new_n7302_, new_n7302_);
  not g_5534 (not_new_n1027__10, new_n1027_);
  not g_5535 (not_new_n1585__10, new_n1585_);
  not g_5536 (new_n4088_, pi272);
  not g_5537 (new_n6058_, new_n5897_);
  not g_5538 (not_new_n8461_, new_n8461_);
  or g_5539 (new_n3612_, not_new_n984__10, not_pi172_0);
  not g_5540 (new_n8110_, new_n1049_);
  not g_5541 (not_new_n4444_, new_n4444_);
  not g_5542 (not_new_n5920__1, new_n5920_);
  or g_5543 (new_n9365_, not_new_n635__332329305696010, not_new_n1045__797922662976120010);
  not g_5544 (not_new_n5803_, new_n5803_);
  not g_5545 (not_new_n641__24010, new_n641_);
  or g_5546 (new_n7215_, not_new_n7421_, not_new_n7001_);
  not g_5547 (not_new_n7109_, new_n7109_);
  not g_5548 (not_new_n8332_, new_n8332_);
  not g_5549 (not_new_n7332_, new_n7332_);
  not g_5550 (not_new_n10206_, new_n10206_);
  or g_5551 (new_n9437_, not_new_n9763_, not_new_n9764_);
  not g_5552 (not_new_n1308_, new_n1308_);
  buf g_5553 (po039, pi225);
  or g_5554 (new_n1537_, not_new_n1228_, not_new_n615_);
  or g_5555 (new_n9849_, not_new_n9578_, not_new_n9847_);
  not g_5556 (not_new_n5347_, new_n5347_);
  not g_5557 (not_new_n5342_, new_n5342_);
  or g_5558 (new_n8902_, not_new_n9324_, not_new_n9325_);
  or g_5559 (po283, or_or_or_not_new_n2874__not_new_n2877__not_new_n2876__not_new_n2878_, not_new_n2875_);
  not g_5560 (not_po296_185621159210175743024531636712070, po296);
  not g_5561 (not_new_n630__490, new_n630_);
  not g_5562 (not_new_n2881_, new_n2881_);
  not g_5563 (not_new_n4396_, new_n4396_);
  or g_5564 (new_n6155_, not_new_n6154_, not_new_n6062_);
  not g_5565 (not_new_n1047__2824752490, new_n1047_);
  not g_5566 (not_new_n581__125892552985318850263419623839875454447587430, new_n581_);
  not g_5567 (not_new_n617__657123623635342801395430, new_n617_);
  not g_5568 (new_n9914_, new_n633_);
  not g_5569 (not_new_n6909_, new_n6909_);
  not g_5570 (not_new_n673_, new_n673_);
  and g_5571 (new_n1327_, new_n2254_, and_new_n1326__new_n2255_);
  not g_5572 (new_n4107_, pi262);
  not g_5573 (not_new_n1039__7, new_n1039_);
  or g_5574 (new_n10013_, not_new_n10151_, not_new_n10150_);
  not g_5575 (not_new_n1576__1, new_n1576_);
  not g_5576 (not_new_n3335_, new_n3335_);
  not g_5577 (not_new_n3854_, new_n3854_);
  not g_5578 (not_new_n3544_, new_n3544_);
  not g_5579 (not_new_n588__6782230728490, new_n588_);
  or g_5580 (or_or_not_new_n8781__not_new_n8701__not_new_n8780_, not_new_n8780_, or_not_new_n8781__not_new_n8701_);
  not g_5581 (not_new_n5839_, new_n5839_);
  or g_5582 (new_n2789_, not_pi252, not_po296_52433383167563036344614587188619514555430);
  or g_5583 (new_n10261_, not_new_n1039__273687473400809163430, not_new_n9884_);
  or g_5584 (new_n7785_, not_new_n628__968890104070, not_new_n7766_);
  or g_5585 (new_n5608_, not_new_n5540_, not_new_n5606_);
  or g_5586 (new_n1706_, not_pi057, not_new_n1631__968890104070);
  or g_5587 (new_n5550_, not_pi138_1, not_new_n1002__5);
  not g_5588 (not_new_n3460_, new_n3460_);
  not g_5589 (not_new_n9325_, new_n9325_);
  not g_5590 (not_new_n1604__4, new_n1604_);
  not g_5591 (not_new_n3835_, new_n3835_);
  not g_5592 (not_new_n6344_, new_n6344_);
  not g_5593 (new_n5088_, new_n4959_);
  and g_5594 (new_n9342_, new_n9662_, new_n9665_);
  or g_5595 (new_n7720_, not_new_n8007_, not_new_n8008_);
  not g_5596 (not_new_n1598__113988951853731430, new_n1598_);
  and g_5597 (and_new_n2399__new_n2398_, new_n2398_, new_n2399_);
  or g_5598 (new_n4502_, not_new_n4555_, not_new_n4556_);
  not g_5599 (not_new_n1043__10, new_n1043_);
  or g_5600 (new_n7801_, not_new_n1051__168070, not_new_n7617_);
  not g_5601 (not_new_n5807__0, new_n5807_);
  not g_5602 (new_n5765_, new_n621_);
  or g_5603 (new_n1913_, not_new_n4920_, not_new_n1589__6);
  not g_5604 (not_new_n1537__403536070, new_n1537_);
  xor g_5605 (key_gate_51, key_51, not_new_n1690_);
  or g_5606 (new_n744_, not_new_n3300_, not_new_n3299_);
  not g_5607 (not_new_n1900__0, new_n1900_);
  not g_5608 (not_new_n634__7, new_n634_);
  or g_5609 (new_n2707_, not_new_n1587__0, not_new_n991_);
  or g_5610 (new_n2363_, not_new_n600__1, not_pi250_0);
  or g_5611 (new_n8625_, not_new_n8720_, not_new_n8721_);
  or g_5612 (new_n5955_, not_new_n5938_, not_new_n5882__0);
  or g_5613 (new_n9838_, not_new_n9395_, not_new_n644__5585458640832840070);
  not g_5614 (not_new_n4243_, new_n4243_);
  or g_5615 (new_n5364_, not_new_n4956_, not_new_n1602__9);
  not g_5616 (not_new_n7581_, new_n7581_);
  not g_5617 (not_new_n8708_, new_n8708_);
  or g_5618 (new_n6049_, not_new_n5905__1, not_new_n5849_);
  and g_5619 (new_n1366_, new_n2400_, new_n2401_);
  not g_5620 (not_new_n1613__138412872010, new_n1613_);
  not g_5621 (not_new_n3429_, new_n3429_);
  and g_5622 (new_n7718_, new_n7997_, new_n7771_);
  not g_5623 (not_new_n2594_, new_n2594_);
  or g_5624 (new_n6383_, not_new_n644__403536070, not_new_n6290_);
  not g_5625 (not_new_n9515_, new_n9515_);
  not g_5626 (not_new_n7249_, new_n7249_);
  not g_5627 (not_new_n630__113988951853731430, new_n630_);
  or g_5628 (or_not_new_n8413__not_new_n8252_, not_new_n8413_, not_new_n8252_);
  not g_5629 (not_new_n3555_, new_n3555_);
  not g_5630 (new_n8638_, new_n1177_);
  or g_5631 (new_n10308_, not_new_n1602__113988951853731430, not_new_n9933_);
  not g_5632 (not_new_n8971_, new_n8971_);
  not g_5633 (not_new_n4802__1, new_n4802_);
  not g_5634 (not_new_n1061__57648010, new_n1061_);
  not g_5635 (not_pi274_0, pi274);
  not g_5636 (not_new_n3506_, new_n3506_);
  not g_5637 (not_new_n6811_, new_n6811_);
  and g_5638 (po112, key_gate_101, pi091);
  not g_5639 (not_new_n1728__2824752490, new_n1728_);
  not g_5640 (not_new_n8866__0, new_n8866_);
  not g_5641 (not_new_n6745_, new_n6745_);
  not g_5642 (not_new_n1059__6, new_n1059_);
  not g_5643 (not_new_n1071__8235430, new_n1071_);
  not g_5644 (not_new_n1604__9, new_n1604_);
  and g_5645 (and_new_n3007__new_n998_, new_n998_, new_n3007_);
  not g_5646 (not_new_n598__1, new_n598_);
  or g_5647 (new_n10128_, new_n1069_, new_n646_);
  not g_5648 (not_new_n1538__47475615099430, new_n1538_);
  not g_5649 (not_pi128, pi128);
  not g_5650 (new_n7108_, new_n768_);
  and g_5651 (new_n9339_, new_n9627_, new_n9621_);
  or g_5652 (or_not_new_n4841__not_new_n4762_, not_new_n4841_, not_new_n4762_);
  not g_5653 (not_new_n2341_, new_n2341_);
  not g_5654 (not_new_n632__4, new_n632_);
  not g_5655 (not_new_n5748__0, new_n5748_);
  not g_5656 (not_new_n1047__168070, new_n1047_);
  not g_5657 (not_new_n6651__0, new_n6651_);
  not g_5658 (not_pi040_3, pi040);
  not g_5659 (not_new_n7870_, new_n7870_);
  not g_5660 (not_new_n9059_, new_n9059_);
  not g_5661 (not_new_n1538__10, new_n1538_);
  not g_5662 (not_new_n4499_, new_n4499_);
  or g_5663 (new_n2575_, not_new_n605__6, not_new_n5490_);
  or g_5664 (or_not_new_n5453__not_new_n5706__1, not_new_n5706__1, not_new_n5453_);
  or g_5665 (new_n1174_, not_new_n3877_, not_new_n3878_);
  not g_5666 (not_new_n5499_, new_n5499_);
  not g_5667 (not_new_n2052__0, new_n2052_);
  not g_5668 (not_new_n7090_, new_n7090_);
  or g_5669 (new_n5396_, not_new_n4957_, not_new_n638__24010);
  or g_5670 (new_n1921_, not_pi138, not_new_n587__8);
  not g_5671 (not_new_n9326__0, new_n9326_);
  not g_5672 (new_n8986_, new_n8878_);
  and g_5673 (new_n5037_, new_n5164_, new_n4909_);
  or g_5674 (new_n2083_, not_new_n8917_, not_new_n1591__168070);
  not g_5675 (not_new_n1597__2, new_n1597_);
  not g_5676 (not_new_n8824_, new_n8824_);
  not g_5677 (not_new_n9535_, new_n9535_);
  not g_5678 (not_new_n8857__0, new_n8857_);
  not g_5679 (new_n7650_, new_n1055_);
  not g_5680 (not_pi051_3, pi051);
  not g_5681 (not_new_n8131__0, new_n8131_);
  or g_5682 (new_n3600_, not_new_n984__4, not_pi166_0);
  or g_5683 (new_n5355_, not_new_n5196_, not_new_n5353_);
  not g_5684 (not_new_n7590_, new_n7590_);
  not g_5685 (not_new_n9950_, new_n9950_);
  or g_5686 (new_n9683_, not_new_n9387__0, not_new_n9539__0);
  and g_5687 (new_n6582_, new_n6724_, new_n6455_);
  or g_5688 (new_n10219_, not_new_n9989_, not_new_n10029__3);
  not g_5689 (not_new_n6178_, new_n6178_);
  or g_5690 (new_n9765_, not_new_n9376_, not_new_n617__273687473400809163430);
  not g_5691 (not_new_n8687_, new_n8687_);
  not g_5692 (not_new_n8155_, new_n8155_);
  or g_5693 (new_n3003_, not_new_n1153_, not_new_n1027__7);
  not g_5694 (new_n4797_, new_n1063_);
  not g_5695 (not_new_n3583_, new_n3583_);
  not g_5696 (not_new_n8209_, new_n8209_);
  or g_5697 (new_n2997_, not_new_n1151_, not_new_n1027__5);
  not g_5698 (not_new_n630__797922662976120010, new_n630_);
  not g_5699 (not_new_n3375__0, new_n3375_);
  not g_5700 (not_new_n7597_, new_n7597_);
  or g_5701 (or_not_new_n1247__not_new_n1245_, not_new_n1247_, not_new_n1245_);
  or g_5702 (new_n8493_, not_new_n619__8235430, not_new_n8250_);
  not g_5703 (not_new_n595__1176490, new_n595_);
  not g_5704 (not_new_n9611_, new_n9611_);
  not g_5705 (not_new_n5367_, new_n5367_);
  and g_5706 (new_n7142_, new_n7492_, new_n7493_);
  or g_5707 (new_n5340_, not_new_n4949__0, not_new_n1597__10);
  not g_5708 (not_new_n1190_, new_n1190_);
  not g_5709 (not_new_n648__47475615099430, new_n648_);
  not g_5710 (not_new_n1600__403536070, new_n1600_);
  not g_5711 (not_new_n6771_, new_n6771_);
  not g_5712 (not_new_n6974__1, new_n6974_);
  not g_5713 (not_new_n7735__1, new_n7735_);
  not g_5714 (not_new_n641__57648010, new_n641_);
  not g_5715 (not_new_n8125__0, new_n8125_);
  not g_5716 (not_new_n8027_, new_n8027_);
  or g_5717 (new_n6132_, not_new_n5764__1, not_new_n618__57648010);
  or g_5718 (new_n8721_, not_new_n8623_, not_new_n1170__0);
  and g_5719 (new_n8076_, new_n8301_, new_n8300_);
  not g_5720 (not_new_n1363_, new_n1363_);
  or g_5721 (new_n2598_, not_new_n610__8, not_new_n4469__0);
  or g_5722 (new_n2905_, not_pi265_4, not_po296_5080218607396233653221881976522165017724345248360010);
  not g_5723 (not_new_n6645_, new_n6645_);
  not g_5724 (not_new_n8601_, new_n8601_);
  not g_5725 (not_new_n1065__6782230728490, new_n1065_);
  or g_5726 (new_n9614_, new_n1069_, new_n646_);
  or g_5727 (new_n3657_, not_new_n642__8, not_po298_1);
  not g_5728 (not_new_n7743_, new_n7743_);
  not g_5729 (new_n7867_, new_n7744_);
  not g_5730 (not_new_n1728__968890104070, new_n1728_);
  not g_5731 (not_new_n6842_, new_n6842_);
  not g_5732 (not_new_n5915__0, new_n5915_);
  or g_5733 (new_n4149_, not_new_n4163__0, not_pi261_1);
  not g_5734 (not_pi172_3, pi172);
  not g_5735 (not_new_n5459__1, new_n5459_);
  not g_5736 (not_new_n4333_, new_n4333_);
  not g_5737 (not_new_n1534__2326305139872070, key_gate_5);
  not g_5738 (not_new_n590__1, new_n590_);
  not g_5739 (not_new_n1824__0, new_n1824_);
  not g_5740 (not_new_n5307_, new_n5307_);
  or g_5741 (new_n2326_, not_new_n601__2326305139872070, not_new_n618__0);
  not g_5742 (not_new_n3904_, new_n3904_);
  and g_5743 (new_n5726_, new_n5723_, new_n5975_);
  or g_5744 (new_n3845_, not_new_n6443__8, not_new_n619__6);
  or g_5745 (new_n950_, or_or_not_new_n1255__not_new_n1253__not_new_n1907_, not_new_n1906_);
  not g_5746 (not_new_n10069_, new_n10069_);
  not g_5747 (not_new_n7828_, new_n7828_);
  not g_5748 (not_new_n7107_, new_n7107_);
  not g_5749 (not_new_n8902_, new_n8902_);
  not g_5750 (not_new_n6543_, new_n6543_);
  not g_5751 (not_new_n9830_, new_n9830_);
  not g_5752 (not_new_n3966_, new_n3966_);
  not g_5753 (not_new_n8918_, new_n8918_);
  not g_5754 (not_new_n9467_, new_n9467_);
  or g_5755 (new_n9148_, new_n1051_, new_n647_);
  not g_5756 (not_pi246, pi246);
  not g_5757 (not_new_n4446_, new_n4446_);
  and g_5758 (new_n3970_, not_pi057_2, not_pi058_2);
  and g_5759 (and_not_pi048_2_not_pi047_2, not_pi048_2, not_pi047_2);
  not g_5760 (not_new_n1045__6, new_n1045_);
  or g_5761 (new_n3236_, not_new_n3185__6782230728490, not_new_n1055__4);
  and g_5762 (new_n3920_, new_n3947_, new_n4041_);
  not g_5763 (not_new_n1591__10, new_n1591_);
  or g_5764 (new_n3136_, not_new_n639__6, not_new_n581__9095436801298611408202050198891430);
  not g_5765 (not_new_n3184__6, new_n3184_);
  or g_5766 (new_n10265_, not_new_n9881_, not_new_n632__273687473400809163430);
  not g_5767 (not_new_n6370_, new_n6370_);
  not g_5768 (not_new_n1537__1, new_n1537_);
  or g_5769 (po146, not_new_n3518_, not_new_n3519_);
  or g_5770 (new_n8321_, not_new_n8304_, not_new_n8248__0);
  not g_5771 (not_new_n6009_, new_n6009_);
  not g_5772 (not_new_n943_, new_n943_);
  and g_5773 (new_n5060_, new_n5324_, new_n5323_);
  and g_5774 (new_n1279_, and_new_n1278__new_n2027_, new_n2026_);
  or g_5775 (new_n9669_, new_n1057_, new_n636_);
  not g_5776 (not_new_n8584_, new_n8584_);
  not g_5777 (not_new_n4640_, new_n4640_);
  not g_5778 (not_new_n3477_, new_n3477_);
  not g_5779 (not_new_n1003__6, new_n1003_);
  not g_5780 (not_new_n1601__8, new_n1601_);
  not g_5781 (not_new_n9957_, new_n9957_);
  or g_5782 (new_n9817_, not_new_n633__113988951853731430, not_new_n9413__0);
  not g_5783 (not_new_n1576__968890104070, new_n1576_);
  not g_5784 (not_new_n7025__0, new_n7025_);
  or g_5785 (new_n2913_, not_new_n595__403536070, not_new_n7049_);
  not g_5786 (new_n7183_, new_n6977_);
  not g_5787 (new_n8179_, new_n641_);
  or g_5788 (new_n3952_, not_new_n4014__2, not_new_n3974_);
  not g_5789 (not_new_n8229_, new_n8229_);
  not g_5790 (not_new_n1057_, new_n1057_);
  not g_5791 (not_new_n7847_, new_n7847_);
  not g_5792 (not_new_n635__19773267430, new_n635_);
  not g_5793 (not_new_n6760_, new_n6760_);
  not g_5794 (not_new_n9858_, new_n9858_);
  not g_5795 (not_new_n2523_, new_n2523_);
  not g_5796 (not_new_n3943_, new_n3943_);
  not g_5797 (not_new_n9558_, new_n9558_);
  not g_5798 (not_new_n4286__0, new_n4286_);
  or g_5799 (new_n6409_, not_new_n625__403536070, not_new_n6300_);
  or g_5800 (new_n9198_, not_new_n8841_, not_new_n1049__47475615099430);
  not g_5801 (not_new_n8654_, new_n8654_);
  not g_5802 (not_new_n5875_, new_n5875_);
  or g_5803 (new_n10307_, not_new_n625__657123623635342801395430, not_new_n9932_);
  not g_5804 (new_n5455_, pi140);
  not g_5805 (not_new_n9919__0, new_n9919_);
  not g_5806 (not_new_n977_, new_n977_);
  not g_5807 (not_new_n9812_, new_n9812_);
  not g_5808 (not_new_n9378_, new_n9378_);
  or g_5809 (new_n2260_, not_new_n1588__47475615099430, not_new_n1599_);
  not g_5810 (not_pi028_0, pi028);
  or g_5811 (new_n10206_, not_new_n9909__0, not_new_n10128__0);
  not g_5812 (not_new_n7551_, new_n7551_);
  or g_5813 (new_n8037_, not_new_n7754__4, not_new_n7725_);
  not g_5814 (not_new_n1589__490, new_n1589_);
  not g_5815 (new_n4807_, new_n1055_);
  not g_5816 (not_new_n8066_, new_n8066_);
  not g_5817 (not_new_n623__3, new_n623_);
  not g_5818 (new_n6074_, new_n5905_);
  not g_5819 (not_new_n1581__1, new_n1581_);
  or g_5820 (new_n1045_, not_new_n3432_, not_new_n3433_);
  and g_5821 (and_new_n4351__new_n4350_, new_n4350_, new_n4351_);
  not g_5822 (not_new_n1876_, new_n1876_);
  or g_5823 (or_or_not_new_n2170__not_new_n2167__not_new_n2168_, or_not_new_n2170__not_new_n2167_, not_new_n2168_);
  or g_5824 (new_n7681_, not_new_n8047_, not_new_n8046_);
  not g_5825 (not_new_n9481_, new_n9481_);
  not g_5826 (not_new_n9895_, new_n9895_);
  xor g_5827 (key_gate_6, key_6, new_n3931_);
  not g_5828 (not_new_n4436__0, new_n4436_);
  not g_5829 (not_new_n9200_, new_n9200_);
  or g_5830 (new_n10278_, not_new_n10276_, not_new_n10277_);
  not g_5831 (not_new_n1526_, new_n1526_);
  or g_5832 (new_n6819_, not_new_n6570_, not_new_n6496_);
  not g_5833 (not_new_n2694_, new_n2694_);
  not g_5834 (new_n7567_, new_n7097_);
  xor g_5835 (key_gate_57, key_57, not_new_n3921_);
  or g_5836 (new_n5199_, new_n1600_, new_n629_);
  or g_5837 (new_n10232_, not_new_n10179_, not_new_n9951__0);
  not g_5838 (not_new_n5115_, new_n5115_);
  not g_5839 (not_new_n8837__1, new_n8837_);
  or g_5840 (new_n8068_, not_new_n7761_, not_new_n7731_);
  not g_5841 (not_new_n4598_, new_n4598_);
  not g_5842 (not_new_n637__2326305139872070, new_n637_);
  not g_5843 (not_new_n1591__16284135979104490, new_n1591_);
  not g_5844 (not_new_n2282_, new_n2282_);
  not g_5845 (not_new_n3453_, new_n3453_);
  not g_5846 (not_new_n10116_, new_n10116_);
  and g_5847 (new_n8968_, new_n9263_, new_n9264_);
  or g_5848 (new_n4689_, not_pi174_2, not_new_n4440_);
  not g_5849 (not_new_n2806_, new_n2806_);
  not g_5850 (not_new_n9949__0, new_n9949_);
  not g_5851 (new_n2275_, new_n976_);
  not g_5852 (new_n3363_, new_n1020_);
  not g_5853 (not_new_n984__57648010, new_n984_);
  not g_5854 (not_new_n4740_, new_n4740_);
  or g_5855 (new_n8301_, not_new_n8106_, not_new_n631__16284135979104490);
  and g_5856 (new_n1571_, new_n3653_, new_n3652_);
  not g_5857 (not_new_n1014__4, new_n1014_);
  not g_5858 (not_new_n585__138412872010, new_n585_);
  not g_5859 (not_new_n10217_, new_n10217_);
  not g_5860 (not_new_n1631__8, key_gate_76);
  not g_5861 (not_new_n6001_, new_n6001_);
  or g_5862 (new_n2459_, not_new_n9871__0, not_new_n599__2824752490);
  or g_5863 (new_n1007_, not_new_n3336_, not_new_n3335_);
  not g_5864 (new_n4269_, new_n690_);
  not g_5865 (not_new_n6364_, new_n6364_);
  not g_5866 (not_new_n605__490, new_n605_);
  not g_5867 (not_new_n3861_, new_n3861_);
  not g_5868 (not_new_n1596__47475615099430, new_n1596_);
  not g_5869 (not_new_n5665_, new_n5665_);
  not g_5870 (not_new_n7563_, new_n7563_);
  not g_5871 (not_new_n996_, new_n996_);
  not g_5872 (not_new_n606__4, new_n606_);
  or g_5873 (new_n2596_, or_not_new_n2595__not_new_n2594_, not_new_n2593_);
  not g_5874 (not_new_n4570_, new_n4570_);
  and g_5875 (new_n6961_, new_n7181_, new_n7182_);
  or g_5876 (new_n7522_, not_new_n7521_, not_new_n7520_);
  not g_5877 (not_new_n636__113988951853731430, new_n636_);
  or g_5878 (new_n10016_, not_new_n10136_, not_new_n10137_);
  not g_5879 (not_new_n7355_, new_n7355_);
  or g_5880 (new_n6547_, not_new_n6811_, not_new_n6528_);
  not g_5881 (not_new_n9847_, new_n9847_);
  not g_5882 (not_new_n994__3430, new_n994_);
  not g_5883 (not_new_n7436__0, new_n7436_);
  not g_5884 (not_new_n1619__0, new_n1619_);
  not g_5885 (not_new_n8367_, new_n8367_);
  not g_5886 (not_new_n4442__0, new_n4442_);
  not g_5887 (not_new_n586__4, new_n586_);
  not g_5888 (not_new_n7774_, new_n7774_);
  or g_5889 (new_n8232_, not_new_n8539_, not_new_n8538_);
  not g_5890 (not_new_n1356_, new_n1356_);
  or g_5891 (new_n8575_, not_new_n8153__0, not_new_n644__47475615099430);
  or g_5892 (new_n3639_, not_new_n972_, not_new_n1611__968890104070);
  or g_5893 (new_n5989_, not_new_n5783_, not_new_n1067__70);
  not g_5894 (not_new_n8621_, new_n8621_);
  not g_5895 (not_new_n1628_, new_n1628_);
  or g_5896 (new_n4205_, not_pi254_1, not_new_n4096_);
  not g_5897 (new_n8140_, new_n1603_);
  or g_5898 (new_n8796_, not_new_n8713__2, or_not_new_n1158__1_not_new_n8715__0);
  not g_5899 (not_new_n6983__0, new_n6983_);
  or g_5900 (new_n8884_, not_new_n1065__2326305139872070, not_new_n637__6782230728490);
  or g_5901 (new_n9290_, not_new_n8883_, not_new_n1067__19773267430);
  not g_5902 (new_n4845_, new_n4755_);
  not g_5903 (not_new_n9530_, new_n9530_);
  and g_5904 (new_n1463_, and_new_n3729__new_n3726_, new_n3723_);
  not g_5905 (not_pi263_2, pi263);
  or g_5906 (new_n6426_, not_new_n6234__0, or_or_not_new_n6337__not_new_n6373__6_not_new_n6338_);
  or g_5907 (or_not_new_n6327__not_new_n6373__2, not_new_n6373__2, not_new_n6327_);
  or g_5908 (new_n5566_, not_new_n1015__5, not_new_n5680_);
  not g_5909 (not_new_n775__8235430, new_n775_);
  not g_5910 (not_new_n719__0, new_n719_);
  or g_5911 (or_not_new_n2189__not_new_n2186_, not_new_n2189_, not_new_n2186_);
  not g_5912 (not_new_n761_, new_n761_);
  or g_5913 (new_n6191_, not_new_n633__8235430, not_new_n5784__0);
  not g_5914 (not_new_n9943__0, new_n9943_);
  not g_5915 (not_new_n1926_, new_n1926_);
  or g_5916 (new_n2937_, not_new_n1039__1, not_new_n3311__168070);
  or g_5917 (new_n3496_, not_new_n1613__8235430, not_new_n2128_);
  not g_5918 (not_new_n643__24010, new_n643_);
  and g_5919 (new_n6462_, new_n6862_, new_n6861_);
  or g_5920 (new_n7322_, not_new_n7113__0, not_new_n6967_);
  not g_5921 (not_new_n7611__1, new_n7611_);
  not g_5922 (not_new_n9196_, new_n9196_);
  or g_5923 (new_n2175_, not_new_n9344_, not_new_n1584__2824752490);
  or g_5924 (new_n6378_, not_new_n6246_, not_new_n622__8235430);
  not g_5925 (not_new_n6974__10, new_n6974_);
  not g_5926 (not_new_n4220_, new_n4220_);
  or g_5927 (new_n7426_, not_new_n757_, not_new_n6974__1176490);
  or g_5928 (new_n8553_, not_new_n1069__403536070, not_new_n8146__0);
  not g_5929 (new_n6541_, new_n618_);
  not g_5930 (not_new_n8087_, new_n8087_);
  not g_5931 (not_new_n3539_, new_n3539_);
  not g_5932 (not_new_n6981__1, new_n6981_);
  or g_5933 (new_n4190_, not_new_n4111_, not_new_n4175_);
  not g_5934 (not_new_n4130_, new_n4130_);
  and g_5935 (and_new_n5083__new_n5411_, new_n5411_, new_n5083_);
  not g_5936 (not_new_n1611__9, new_n1611_);
  not g_5937 (not_new_n753_, new_n753_);
  not g_5938 (not_new_n587__1, new_n587_);
  not g_5939 (not_new_n5873_, new_n5873_);
  or g_5940 (or_not_new_n2015__not_new_n2016_, not_new_n2015_, not_new_n2016_);
  not g_5941 (not_new_n10332_, new_n10332_);
  not g_5942 (not_new_n775__19773267430, new_n775_);
  not g_5943 (not_new_n7041__0, new_n7041_);
  or g_5944 (new_n9546_, not_new_n9365__0, not_new_n9530_);
  not g_5945 (not_new_n3181_, new_n3181_);
  or g_5946 (new_n6495_, not_new_n6690_, not_new_n6490_);
  or g_5947 (new_n5114_, new_n1051_, new_n647_);
  not g_5948 (not_new_n6477_, new_n6477_);
  not g_5949 (not_new_n6347_, new_n6347_);
  not g_5950 (not_new_n1067__3, new_n1067_);
  not g_5951 (not_new_n1589__19773267430, new_n1589_);
  or g_5952 (new_n8573_, not_new_n8449_, not_new_n8270_);
  not g_5953 (not_new_n1393_, new_n1393_);
  not g_5954 (not_new_n7039_, new_n7039_);
  and g_5955 (new_n6350_, new_n6401_, and_and_new_n6373__new_n6254__new_n6402_);
  and g_5956 (new_n6451_, new_n6733_, new_n6734_);
  or g_5957 (new_n8578_, not_new_n8272_, not_new_n8239_);
  and g_5958 (new_n3962_, not_pi040_2, not_pi039_2);
  not g_5959 (not_new_n7708_, new_n7708_);
  or g_5960 (new_n3827_, not_new_n6443_, not_new_n647__70);
  not g_5961 (not_new_n8304__0, new_n8304_);
  not g_5962 (new_n9892_, new_n641_);
  not g_5963 (not_new_n3311__6, new_n3311_);
  and g_5964 (new_n1514_, new_n1515_, new_n3046_);
  not g_5965 (not_new_n6539__2, new_n6539_);
  and g_5966 (new_n1293_, new_n2099_, new_n2098_);
  or g_5967 (new_n2015_, not_new_n586__3430, not_pi175);
  not g_5968 (not_new_n1012__7, new_n1012_);
  or g_5969 (new_n3891_, not_new_n626__3430, not_new_n9920_);
  not g_5970 (not_new_n595__9, new_n595_);
  or g_5971 (new_n7899_, not_new_n7733_, not_new_n7898_);
  or g_5972 (or_or_not_new_n2015__not_new_n2016__not_new_n2018_, or_not_new_n2015__not_new_n2016_, not_new_n2018_);
  not g_5973 (not_new_n641__403536070, new_n641_);
  not g_5974 (not_new_n941_, new_n941_);
  or g_5975 (or_not_new_n1920__not_new_n1921_, not_new_n1921_, not_new_n1920_);
  or g_5976 (new_n10304_, not_new_n10303_, not_new_n10302_);
  or g_5977 (new_n7470_, not_new_n7468_, not_new_n7469_);
  and g_5978 (and_new_n2692__new_n2691_, new_n2692_, new_n2691_);
  not g_5979 (not_new_n994__332329305696010, new_n994_);
  not g_5980 (not_po296_32199057558131797268376070, po296);
  not g_5981 (not_new_n5207_, new_n5207_);
  or g_5982 (or_or_not_new_n1303__not_new_n1301__not_new_n2135_, or_not_new_n1303__not_new_n1301_, not_new_n2135_);
  and g_5983 (new_n1453_, new_n2680_, and_new_n2682__new_n2681_);
  or g_5984 (new_n9956_, not_new_n10245_, not_new_n10244_);
  not g_5985 (not_new_n7079_, new_n7079_);
  or g_5986 (new_n7836_, not_new_n7835_, not_new_n7574_);
  or g_5987 (new_n2654_, not_new_n1007_, not_new_n607__490);
  not g_5988 (not_new_n10298_, new_n10298_);
  or g_5989 (new_n1019_, not_new_n3360_, not_new_n3359_);
  or g_5990 (new_n7789_, not_new_n7773_, not_new_n7777_);
  not g_5991 (not_new_n8110__1, new_n8110_);
  not g_5992 (not_new_n6864_, new_n6864_);
  or g_5993 (new_n3748_, not_new_n639__10, not_new_n1603__6);
  not g_5994 (not_new_n9870__0, new_n9870_);
  not g_5995 (not_new_n4950_, new_n4950_);
  not g_5996 (not_new_n1589__4, new_n1589_);
  and g_5997 (po094, pi073, key_gate_101);
  or g_5998 (new_n10331_, not_new_n10024__0, not_new_n10206_);
  or g_5999 (new_n7304_, not_new_n7012__0, not_new_n7258__0);
  not g_6000 (not_new_n1063__6782230728490, new_n1063_);
  or g_6001 (new_n5305_, not_new_n4935_, not_new_n1045__9);
  not g_6002 (not_new_n10082_, new_n10082_);
  not g_6003 (not_new_n4418_, new_n4418_);
  not g_6004 (not_new_n9786_, new_n9786_);
  not g_6005 (not_new_n9945__0, new_n9945_);
  or g_6006 (new_n9777_, not_new_n9422__0, not_new_n9687_);
  or g_6007 (new_n8510_, not_new_n8506_, not_new_n8278__0);
  not g_6008 (not_new_n595__3, new_n595_);
  not g_6009 (not_new_n8282_, new_n8282_);
  not g_6010 (not_new_n4504__0, new_n4504_);
  not g_6011 (not_new_n8933_, new_n8933_);
  not g_6012 (not_new_n4917_, new_n4917_);
  or g_6013 (new_n4357_, not_new_n4354_, not_new_n4302_);
  not g_6014 (not_new_n989__2824752490, new_n989_);
  not g_6015 (new_n8141_, new_n640_);
  or g_6016 (new_n3094_, not_new_n635__5, not_new_n3315__4);
  or g_6017 (new_n2387_, not_new_n648__1, not_new_n603__6);
  not g_6018 (not_new_n9055_, new_n9055_);
  not g_6019 (not_new_n9592_, new_n9592_);
  and g_6020 (new_n10021_, new_n10314_, new_n10315_);
  not g_6021 (not_new_n8863_, new_n8863_);
  not g_6022 (not_new_n4125__1, new_n4125_);
  and g_6023 (new_n1403_, new_n2493_, new_n2492_);
  not g_6024 (not_new_n8925_, new_n8925_);
  or g_6025 (new_n9647_, not_new_n9332_, not_new_n9426_);
  not g_6026 (not_new_n1349_, new_n1349_);
  or g_6027 (new_n3009_, not_new_n581__6, not_new_n1605__1);
  or g_6028 (new_n3821_, not_new_n1581__797922662976120010, not_new_n1574_);
  or g_6029 (new_n7060_, not_new_n7505_, not_new_n7504_);
  not g_6030 (not_new_n5861_, new_n5861_);
  or g_6031 (new_n3613_, not_new_n1611__10, not_new_n954_);
  not g_6032 (new_n9941_, new_n1598_);
  not g_6033 (not_new_n4825__0, new_n4825_);
  not g_6034 (not_new_n3315__0, new_n3315_);
  not g_6035 (not_new_n4344__0, new_n4344_);
  not g_6036 (not_new_n640__3430, new_n640_);
  or g_6037 (po230, not_new_n1450_, not_new_n1449_);
  or g_6038 (new_n8589_, not_new_n8409_, not_new_n8178__0);
  not g_6039 (new_n5093_, new_n5071_);
  not g_6040 (not_new_n3766_, new_n3766_);
  or g_6041 (new_n10312_, not_new_n10020__0, not_new_n10019_);
  or g_6042 (new_n4144_, not_pi266_1, not_new_n4155__0);
  or g_6043 (new_n5171_, not_new_n633__3430, not_new_n5170_);
  not g_6044 (not_new_n3315__332329305696010, new_n3315_);
  not g_6045 (new_n5467_, pi144);
  not g_6046 (not_new_n3351_, new_n3351_);
  or g_6047 (or_or_not_new_n2928__not_new_n2931__not_new_n2930_, not_new_n2930_, or_not_new_n2928__not_new_n2931_);
  or g_6048 (new_n8506_, not_new_n8505_, not_new_n8504_);
  not g_6049 (not_new_n1005__6, new_n1005_);
  not g_6050 (not_new_n10133_, new_n10133_);
  not g_6051 (not_new_n618__57648010, new_n618_);
  not g_6052 (not_new_n4796__0, new_n4796_);
  not g_6053 (not_new_n603__57648010, new_n603_);
  or g_6054 (new_n7000_, not_new_n735_, not_new_n7033_);
  or g_6055 (new_n7497_, not_new_n7143__0, not_new_n7142_);
  or g_6056 (new_n2241_, not_new_n1600_, not_new_n1588__6782230728490);
  not g_6057 (not_new_n7408_, new_n7408_);
  not g_6058 (not_new_n10093_, new_n10093_);
  or g_6059 (new_n681_, not_new_n1493_, not_new_n3008_);
  and g_6060 (new_n1216_, new_n1778_, and_new_n1215__new_n1780_);
  not g_6061 (not_new_n594__70, new_n594_);
  not g_6062 (not_new_n7854_, new_n7854_);
  not g_6063 (not_new_n4694_, new_n4694_);
  and g_6064 (new_n6624_, new_n6881_, new_n6880_);
  not g_6065 (not_new_n7029_, new_n7029_);
  not g_6066 (not_new_n1027__113988951853731430, new_n1027_);
  not g_6067 (not_new_n4227__0, new_n4227_);
  not g_6068 (not_new_n8146_, new_n8146_);
  not g_6069 (not_new_n1629_, new_n1629_);
  or g_6070 (new_n9798_, not_new_n9407_, not_new_n639__113988951853731430);
  not g_6071 (not_new_n1045_, new_n1045_);
  and g_6072 (new_n9989_, new_n9866_, new_n10108_);
  not g_6073 (not_new_n5948__0, new_n5948_);
  not g_6074 (new_n5777_, new_n640_);
  not g_6075 (not_new_n1678_, key_gate_108);
  not g_6076 (not_new_n9089_, new_n9089_);
  not g_6077 (not_new_n3352_, new_n3352_);
  not g_6078 (not_new_n4457__0, new_n4457_);
  not g_6079 (not_new_n1612__16284135979104490, new_n1612_);
  and g_6080 (new_n1223_, and_and_new_n1750__new_n1751__new_n1753_, new_n1752_);
  and g_6081 (new_n1434_, new_n2599_, new_n2598_);
  not g_6082 (not_new_n731__0, new_n731_);
  or g_6083 (new_n3672_, not_pi222, not_new_n989__8);
  not g_6084 (not_new_n1603__138412872010, new_n1603_);
  not g_6085 (not_new_n5439_, new_n5439_);
  not g_6086 (not_new_n6188_, new_n6188_);
  or g_6087 (new_n9200_, not_new_n8956__0, not_new_n9155_);
  not g_6088 (new_n1577_, new_n939_);
  not g_6089 (new_n5754_, new_n635_);
  not g_6090 (not_new_n5661_, new_n5661_);
  not g_6091 (not_new_n8331_, new_n8331_);
  not g_6092 (not_new_n591__332329305696010, new_n591_);
  or g_6093 (new_n6734_, not_new_n625__2824752490, not_new_n6507_);
  not g_6094 (not_po296_4599865365447399609768010, po296);
  or g_6095 (new_n5826_, not_new_n6093_, not_new_n6094_);
  not g_6096 (not_new_n7018__0, new_n7018_);
  xnor g_6097 (key_gate_12, key_12, new_n3987_);
  not g_6098 (not_po296_14811132966169777414641055325137507340304213552070, po296);
  or g_6099 (new_n4721_, not_new_n620__5, not_new_n4718__0);
  or g_6100 (new_n9611_, not_new_n9333_, not_new_n9514_);
  or g_6101 (new_n9070_, not_new_n8885_, not_new_n8884_);
  not g_6102 (not_new_n6947_, new_n6947_);
  or g_6103 (new_n2480_, not_new_n598__6782230728490, not_new_n1599__0);
  not g_6104 (not_new_n6515__0, new_n6515_);
  not g_6105 (not_new_n6139_, new_n6139_);
  not g_6106 (not_new_n3231_, new_n3231_);
  not g_6107 (not_new_n1616__3, new_n1616_);
  not g_6108 (not_new_n6974__19773267430, new_n6974_);
  not g_6109 (not_new_n6190_, new_n6190_);
  or g_6110 (new_n8998_, not_new_n8924_, not_new_n8798__0);
  not g_6111 (not_new_n603__24010, new_n603_);
  not g_6112 (not_new_n2237_, new_n2237_);
  not g_6113 (not_new_n6523__0, new_n6523_);
  or g_6114 (new_n5560_, not_new_n5559_, not_new_n5515_);
  not g_6115 (not_new_n3114_, new_n3114_);
  not g_6116 (not_new_n3171_, new_n3171_);
  not g_6117 (not_new_n8184_, new_n8184_);
  or g_6118 (new_n4805_, not_new_n4825__0, not_new_n4807__0);
  or g_6119 (new_n9358_, not_new_n642__2326305139872070, not_new_n1035__168070);
  or g_6120 (new_n5990_, not_new_n5784_, not_new_n633__1176490);
  not g_6121 (not_new_n5835_, new_n5835_);
  not g_6122 (not_new_n3395_, new_n3395_);
  not g_6123 (not_new_n4312_, new_n4312_);
  or g_6124 (new_n650_, not_new_n3106_, not_new_n3107_);
  and g_6125 (new_n607_, new_n2505_, new_n3366_);
  not g_6126 (not_new_n4603_, new_n4603_);
  not g_6127 (not_new_n619__168070, new_n619_);
  not g_6128 (new_n3401_, new_n1033_);
  not g_6129 (not_new_n3982_, new_n3982_);
  not g_6130 (not_new_n4489_, new_n4489_);
  not g_6131 (not_new_n8466_, new_n8466_);
  or g_6132 (new_n3766_, not_new_n3444_, not_new_n1905_);
  or g_6133 (new_n1033_, not_new_n3399_, not_new_n3400_);
  not g_6134 (new_n7794_, new_n7615_);
  not g_6135 (not_new_n8718_, new_n8718_);
  not g_6136 (not_new_n1332_, new_n1332_);
  not g_6137 (not_new_n7311_, new_n7311_);
  or g_6138 (new_n3857_, not_new_n6443__24010, not_new_n630__70);
  or g_6139 (new_n10162_, not_new_n9996_, not_new_n10160_);
  not g_6140 (not_new_n1035_, new_n1035_);
  not g_6141 (not_new_n3276_, new_n3276_);
  not g_6142 (not_new_n7437_, new_n7437_);
  not g_6143 (not_po296_541169560379521116689596608490, po296);
  not g_6144 (not_new_n8025_, new_n8025_);
  not g_6145 (not_new_n2889_, new_n2889_);
  or g_6146 (new_n5272_, not_new_n4939_, not_new_n4906_);
  or g_6147 (new_n8286_, not_new_n8119_, not_new_n1043__8235430);
  or g_6148 (new_n2769_, not_new_n2766_, not_new_n1616__3);
  not g_6149 (not_new_n8856__0, new_n8856_);
  not g_6150 (not_new_n8385_, new_n8385_);
  and g_6151 (new_n6345_, new_n6225_, new_n1061_);
  or g_6152 (new_n2296_, not_new_n593__332329305696010, not_new_n618_);
  or g_6153 (new_n578_, not_new_n9892_, not_new_n1031_);
  or g_6154 (new_n2982_, not_new_n3311__57648010, not_new_n1047__1);
  not g_6155 (not_new_n5869_, new_n5869_);
  not g_6156 (not_new_n604__1176490, new_n604_);
  not g_6157 (not_new_n1597__797922662976120010, new_n1597_);
  or g_6158 (new_n2166_, not_new_n2161_, not_new_n1308_);
  or g_6159 (new_n2402_, not_new_n603__9, not_new_n627__1);
  not g_6160 (not_new_n10262_, new_n10262_);
  not g_6161 (not_new_n7371_, new_n7371_);
  or g_6162 (new_n9287_, not_new_n8973__0, not_new_n9162_);
  not g_6163 (not_new_n9301_, new_n9301_);
  not g_6164 (new_n6264_, new_n1069_);
  not g_6165 (not_new_n589__9, new_n589_);
  not g_6166 (not_new_n1607__168070, new_n1607_);
  or g_6167 (new_n2788_, not_new_n7059_, not_new_n595__5);
  not g_6168 (not_new_n9356__1, new_n9356_);
  not g_6169 (not_new_n1616__403536070, new_n1616_);
  not g_6170 (not_new_n8339_, new_n8339_);
  not g_6171 (not_new_n1599__47475615099430, new_n1599_);
  not g_6172 (not_new_n1057__19773267430, new_n1057_);
  and g_6173 (and_new_n3792__new_n3795_, new_n3795_, new_n3792_);
  not g_6174 (not_new_n5218_, new_n5218_);
  not g_6175 (not_new_n6974__403536070, new_n6974_);
  and g_6176 (new_n9869_, new_n10181_, new_n10233_);
  or g_6177 (new_n8225_, not_new_n8516_, not_new_n8515_);
  not g_6178 (not_new_n2978_, new_n2978_);
  not g_6179 (not_new_n3311__57648010, new_n3311_);
  or g_6180 (new_n8728_, not_new_n1049__968890104070, not_new_n8635_);
  not g_6181 (not_new_n6655__1, new_n6655_);
  or g_6182 (new_n5919_, not_new_n1037__70, not_new_n5747_);
  not g_6183 (not_new_n2500_, new_n2500_);
  not g_6184 (not_new_n6443__70, new_n6443_);
  or g_6185 (new_n10329_, not_new_n1069__47475615099430, not_new_n9908_);
  or g_6186 (new_n699_, not_new_n1523_, not_new_n3069_);
  not g_6187 (not_pi242, pi242);
  not g_6188 (not_new_n618__1176490, new_n618_);
  or g_6189 (new_n5154_, not_new_n1059__9, not_new_n644__24010);
  xor g_6190 (key_gate_2, key_2, new_n1696_);
  or g_6191 (new_n10258_, not_new_n10201_, not_new_n9901__0);
  not g_6192 (not_new_n4788__0, new_n4788_);
  not g_6193 (not_new_n643__2326305139872070, new_n643_);
  not g_6194 (not_new_n982_, new_n982_);
  or g_6195 (new_n4113_, not_new_n4177_, not_new_n4178_);
  not g_6196 (not_new_n8186_, new_n8186_);
  not g_6197 (not_new_n7639_, new_n7639_);
  not g_6198 (new_n7163_, new_n7006_);
  and g_6199 (new_n3933_, new_n3936_, new_n4007_);
  and g_6200 (and_new_n2335__new_n2336_, new_n2336_, new_n2335_);
  not g_6201 (not_new_n1600__3, new_n1600_);
  not g_6202 (not_new_n634_, new_n634_);
  not g_6203 (not_new_n2645_, new_n2645_);
  not g_6204 (not_new_n4904_, new_n4904_);
  not g_6205 (not_pi025, pi025);
  or g_6206 (or_or_not_new_n2794__not_new_n2797__not_new_n2796_, not_new_n2796_, or_not_new_n2794__not_new_n2797_);
  or g_6207 (new_n9232_, not_new_n618__39098210485829880490, not_new_n8893__0);
  or g_6208 (new_n7849_, not_new_n640__2824752490, not_new_n7636_);
  or g_6209 (new_n4729_, new_n1035_, or_new_n1031__new_n1037_);
  not g_6210 (not_new_n7160_, new_n7160_);
  or g_6211 (or_not_new_n1550__not_new_n1370_, not_new_n1370_, not_new_n1550_);
  not g_6212 (not_new_n4159__0, new_n4159_);
  not g_6213 (not_new_n9996_, new_n9996_);
  not g_6214 (new_n7660_, new_n1069_);
  or g_6215 (new_n4649_, not_pi180_1, not_new_n4490_);
  not g_6216 (not_new_n6874_, new_n6874_);
  or g_6217 (new_n2897_, not_new_n641__1, not_new_n604__8235430);
  not g_6218 (not_new_n4477__0, new_n4477_);
  not g_6219 (not_pi067, pi067);
  and g_6220 (new_n7699_, new_n7910_, new_n7698_);
  not g_6221 (not_new_n591__10, new_n591_);
  or g_6222 (new_n5214_, not_new_n621__3430, not_new_n1598__8);
  not g_6223 (not_new_n635__57648010, new_n635_);
  not g_6224 (new_n6253_, new_n628_);
  or g_6225 (new_n6496_, not_new_n6646_, or_not_new_n6780__not_new_n6662_);
  not g_6226 (not_new_n1625_, new_n1625_);
  not g_6227 (not_new_n606__24010, new_n606_);
  not g_6228 (not_new_n639__9, new_n639_);
  not g_6229 (not_new_n7141_, new_n7141_);
  or g_6230 (po155, not_new_n3536_, not_new_n3537_);
  not g_6231 (not_new_n5634_, new_n5634_);
  not g_6232 (new_n5558_, new_n5515_);
  not g_6233 (not_new_n8888__0, new_n8888_);
  not g_6234 (not_new_n956_, new_n956_);
  not g_6235 (not_new_n7651_, new_n7651_);
  not g_6236 (not_new_n1597__7, new_n1597_);
  not g_6237 (not_new_n5744__0, new_n5744_);
  not g_6238 (not_new_n623__2, new_n623_);
  not g_6239 (not_po298_4, po298);
  not g_6240 (not_new_n6965_, new_n6965_);
  not g_6241 (not_pi137_3, pi137);
  or g_6242 (new_n2776_, not_new_n3311__3, not_new_n1055__1);
  or g_6243 (new_n5010_, not_new_n5342_, not_new_n5343_);
  or g_6244 (new_n9754_, not_new_n9486__0, not_new_n1607__403536070);
  not g_6245 (not_pi150_0, pi150);
  or g_6246 (new_n10273_, not_new_n10271_, not_new_n10154_);
  not g_6247 (new_n7930_, new_n7746_);
  or g_6248 (po141, not_new_n3508_, not_new_n3509_);
  not g_6249 (not_new_n3944_, new_n3944_);
  not g_6250 (new_n1848_, new_n631_);
  not g_6251 (not_pi141_1, pi141);
  not g_6252 (not_new_n3372__6782230728490, new_n3372_);
  and g_6253 (and_new_n1290__new_n2084_, new_n2084_, new_n1290_);
  not g_6254 (new_n4270_, new_n689_);
  not g_6255 (new_n8860_, new_n1053_);
  not g_6256 (not_new_n7705_, new_n7705_);
  not g_6257 (not_new_n5233_, new_n5233_);
  or g_6258 (new_n6467_, not_new_n6645_, or_not_new_n6782__not_new_n6621_);
  not g_6259 (not_new_n593__2824752490, new_n593_);
  not g_6260 (not_new_n6721_, new_n6721_);
  not g_6261 (not_new_n1585__47475615099430, new_n1585_);
  or g_6262 (new_n3270_, not_new_n3184__70, not_new_n630__8);
  not g_6263 (not_new_n9945_, new_n9945_);
  or g_6264 (new_n3628_, not_pi180_0, not_new_n984__57648010);
  not g_6265 (not_new_n928__1, new_n928_);
  not g_6266 (not_new_n3166_, new_n3166_);
  not g_6267 (not_new_n9774_, new_n9774_);
  not g_6268 (not_new_n7019__1, new_n7019_);
  and g_6269 (new_n593_, new_n1609_, new_n3366_);
  not g_6270 (not_new_n8113__1, new_n8113_);
  not g_6271 (not_new_n6549_, new_n6549_);
  not g_6272 (not_new_n6556_, new_n6556_);
  or g_6273 (new_n2441_, not_new_n597__1176490, not_new_n4793__0);
  not g_6274 (not_po296_4183778472590916451475308348590993345191760458870147715430, po296);
  not g_6275 (not_new_n10124__0, new_n10124_);
  not g_6276 (new_n5058_, new_n619_);
  or g_6277 (new_n1670_, not_pi045, not_new_n1631__70);
  or g_6278 (new_n3071_, not_new_n1057__2, not_new_n581__2326305139872070);
  or g_6279 (new_n1912_, not_new_n8820_, not_new_n1591__6);
  not g_6280 (not_new_n594__4, new_n594_);
  not g_6281 (not_new_n9450_, new_n9450_);
  not g_6282 (not_new_n8326_, new_n8326_);
  or g_6283 (new_n7909_, not_new_n7739__1, not_new_n7697_);
  or g_6284 (po123, not_new_n3431_, not_new_n3430_);
  or g_6285 (new_n9022_, not_new_n8996_, not_new_n8992_);
  not g_6286 (not_pi040_0, pi040);
  not g_6287 (not_new_n1181_, key_gate_50);
  or g_6288 (new_n3826_, or_not_new_n3363__not_new_n583__0, not_pi161_1);
  or g_6289 (new_n2374_, not_new_n9958__0, not_new_n599__3);
  not g_6290 (not_new_n2753_, new_n2753_);
  not g_6291 (not_new_n1069_, new_n1069_);
  or g_6292 (new_n2986_, not_po296_205005145156954906122290109080958673914396262484637238056070, not_pi274_0);
  not g_6293 (not_new_n5792_, new_n5792_);
  not g_6294 (new_n6259_, new_n625_);
  or g_6295 (new_n2334_, or_not_new_n1405__not_new_n616_, not_new_n3307_);
  or g_6296 (or_or_not_new_n6328__not_new_n6373__3_not_new_n6329_, or_not_new_n6328__not_new_n6373__3, not_new_n6329_);
  not g_6297 (not_new_n5053_, new_n5053_);
  not g_6298 (not_new_n933_, new_n933_);
  not g_6299 (not_new_n989__16284135979104490, new_n989_);
  not g_6300 (not_new_n5436_, new_n5436_);
  or g_6301 (new_n7250_, not_new_n7141_, not_new_n7249_);
  and g_6302 (and_not_pi044_1_not_pi043_1, not_pi044_1, not_pi043_1);
  not g_6303 (not_new_n639__138412872010, new_n639_);
  not g_6304 (not_new_n5785__0, new_n5785_);
  not g_6305 (not_new_n620__5, new_n620_);
  or g_6306 (new_n2646_, or_not_new_n2645__not_new_n2644_, not_new_n2643_);
  not g_6307 (not_new_n5428_, new_n5428_);
  not g_6308 (not_new_n1585__1, new_n1585_);
  and g_6309 (new_n6337_, new_n6232_, new_n6275_);
  not g_6310 (not_new_n8254_, new_n8254_);
  not g_6311 (not_new_n638__39098210485829880490, new_n638_);
  or g_6312 (new_n4104_, not_new_n4170_, not_pi271_0);
  not g_6313 (not_new_n3119_, new_n3119_);
  not g_6314 (not_new_n3537_, new_n3537_);
  or g_6315 (new_n10237_, not_new_n1051__47475615099430, not_new_n9897_);
  not g_6316 (not_new_n10284_, new_n10284_);
  or g_6317 (new_n6632_, not_new_n6800_, not_new_n6513_);
  not g_6318 (not_new_n619__6782230728490, new_n619_);
  not g_6319 (not_new_n1276_, new_n1276_);
  not g_6320 (new_n6525_, new_n626_);
  not g_6321 (not_new_n2763_, new_n2763_);
  not g_6322 (not_new_n6519__0, new_n6519_);
  not g_6323 (not_new_n2268_, new_n2268_);
  not g_6324 (not_new_n1045__403536070, new_n1045_);
  or g_6325 (or_or_not_new_n1231__not_new_n1229__not_new_n1793_, or_not_new_n1231__not_new_n1229_, not_new_n1793_);
  not g_6326 (not_new_n9937_, new_n9937_);
  not g_6327 (not_new_n8308_, new_n8308_);
  not g_6328 (not_new_n6911_, new_n6911_);
  not g_6329 (not_new_n1611__8, new_n1611_);
  not g_6330 (not_new_n3270_, new_n3270_);
  not g_6331 (not_new_n8491_, new_n8491_);
  or g_6332 (new_n6121_, not_new_n632__8235430, not_new_n5750__0);
  not g_6333 (not_new_n1538__8235430, new_n1538_);
  and g_6334 (new_n8691_, new_n8762_, new_n8763_);
  not g_6335 (not_new_n8486_, new_n8486_);
  not g_6336 (not_new_n1020__3, new_n1020_);
  not g_6337 (not_new_n1007__2, new_n1007_);
  not g_6338 (not_new_n626__5, new_n626_);
  not g_6339 (not_new_n1537__2824752490, new_n1537_);
  not g_6340 (not_new_n636__3430, new_n636_);
  not g_6341 (not_new_n2546_, new_n2546_);
  or g_6342 (new_n6915_, not_new_n6661_, not_new_n6914_);
  or g_6343 (new_n6875_, not_new_n6873_, not_new_n6874_);
  not g_6344 (not_new_n6795_, new_n6795_);
  not g_6345 (not_new_n1214_, new_n1214_);
  not g_6346 (not_new_n6540_, new_n6540_);
  or g_6347 (new_n9580_, new_n1057_, new_n636_);
  not g_6348 (not_new_n7498_, new_n7498_);
  not g_6349 (not_new_n2877_, new_n2877_);
  not g_6350 (not_new_n617__57648010, new_n617_);
  not g_6351 (not_new_n685_, new_n685_);
  and g_6352 (and_new_n9717__new_n9715_, new_n9715_, new_n9717_);
  or g_6353 (new_n9712_, not_new_n621__113988951853731430, not_new_n9625_);
  or g_6354 (new_n7972_, not_new_n1039__403536070, not_new_n7606__1);
  not g_6355 (not_new_n4523_, new_n4523_);
  not g_6356 (not_new_n6719__0, new_n6719_);
  not g_6357 (not_new_n3585_, new_n3585_);
  or g_6358 (new_n2046_, not_new_n5019_, not_new_n1589__3430);
  or g_6359 (new_n9233_, not_new_n1596__2326305139872070, not_new_n8892__0);
  not g_6360 (not_new_n7222_, new_n7222_);
  not g_6361 (not_new_n9016_, new_n9016_);
  not g_6362 (not_new_n626__6782230728490, new_n626_);
  and g_6363 (and_new_n6422__new_n6426_, new_n6426_, new_n6422_);
  or g_6364 (new_n642_, or_or_not_new_n1763__not_new_n1764__not_new_n1766_, not_new_n1765_);
  not g_6365 (not_new_n3674_, new_n3674_);
  not g_6366 (not_new_n1616__138412872010, new_n1616_);
  not g_6367 (new_n6299_, new_n1603_);
  or g_6368 (new_n7937_, not_new_n7735__1, not_new_n7582_);
  not g_6369 (not_new_n4171__0, new_n4171_);
  not g_6370 (not_new_n8939_, new_n8939_);
  not g_6371 (not_new_n9591_, new_n9591_);
  not g_6372 (not_new_n4004__0, new_n4004_);
  and g_6373 (new_n9453_, new_n1031_, new_n641_);
  or g_6374 (new_n7150_, not_new_n7216_, not_new_n7217_);
  or g_6375 (or_not_new_n1275__not_new_n1273_, not_new_n1273_, not_new_n1275_);
  not g_6376 (not_new_n9770_, new_n9770_);
  not g_6377 (not_new_n1576__490, new_n1576_);
  not g_6378 (new_n7430_, new_n7028_);
  and g_6379 (and_new_n4344__new_n4343_, new_n4343_, new_n4344_);
  not g_6380 (not_new_n9485_, new_n9485_);
  or g_6381 (or_not_new_n1303__not_new_n1301_, not_new_n1303_, not_new_n1301_);
  and g_6382 (new_n1435_, new_n2602_, new_n2600_);
  or g_6383 (new_n5388_, not_new_n5386_, not_new_n5174_);
  not g_6384 (not_new_n2735_, new_n2735_);
  not g_6385 (not_new_n6805_, new_n6805_);
  not g_6386 (new_n5779_, new_n1604_);
  and g_6387 (and_not_pi051_1_not_pi050_1, not_pi051_1, not_pi050_1);
  or g_6388 (new_n8795_, not_new_n8655_, not_new_n8716__0);
  not g_6389 (not_new_n5066_, new_n5066_);
  not g_6390 (not_new_n1041__9, new_n1041_);
  or g_6391 (new_n10091_, not_new_n626__225393402906922580878632490, not_new_n1053__2326305139872070);
  not g_6392 (not_new_n4116_, new_n4116_);
  not g_6393 (not_new_n2782_, new_n2782_);
  or g_6394 (new_n1061_, not_new_n3472_, not_new_n3473_);
  or g_6395 (new_n1748_, not_new_n1728__1176490, not_pi092);
  not g_6396 (not_new_n1055__6, new_n1055_);
  or g_6397 (new_n5502_, not_new_n5527_, not_new_n5528_);
  not g_6398 (not_new_n7243_, new_n7243_);
  or g_6399 (new_n2532_, not_new_n2509__1, not_pi195);
  or g_6400 (new_n6719_, not_new_n6533_, not_new_n1061__168070);
  not g_6401 (not_new_n642__10, new_n642_);
  not g_6402 (not_new_n5612_, new_n5612_);
  not g_6403 (not_new_n7425_, new_n7425_);
  not g_6404 (not_new_n4981_, new_n4981_);
  not g_6405 (not_new_n1051__6, new_n1051_);
  or g_6406 (new_n3129_, not_new_n928__24010, not_new_n1601__3);
  not g_6407 (not_new_n5588_, new_n5588_);
  not g_6408 (not_new_n8266__5, new_n8266_);
  not g_6409 (not_pi176, pi176);
  not g_6410 (not_new_n2752_, new_n2752_);
  or g_6411 (new_n9029_, new_n624_, new_n1041_);
  and g_6412 (new_n8669_, and_new_n8731__new_n8730_, new_n8729_);
  not g_6413 (not_new_n622__3, new_n622_);
  not g_6414 (not_new_n5420_, new_n5420_);
  buf g_6415 (po051, pi213);
  and g_6416 (new_n10003_, new_n10189_, new_n9858_);
  not g_6417 (not_new_n594__403536070, new_n594_);
  or g_6418 (new_n2442_, not_new_n603__8235430, not_new_n645__1);
  not g_6419 (not_new_n5320_, new_n5320_);
  or g_6420 (new_n7349_, not_new_n775__4, not_new_n7103_);
  or g_6421 (new_n4375_, not_new_n4308_, not_new_n4372_);
  not g_6422 (not_pi050, pi050);
  not g_6423 (not_new_n7779_, new_n7779_);
  not g_6424 (not_new_n2873_, new_n2873_);
  not g_6425 (not_new_n6102_, new_n6102_);
  not g_6426 (new_n8264_, new_n1035_);
  or g_6427 (new_n7797_, not_new_n7598__0, not_new_n7597_);
  not g_6428 (not_new_n9332_, new_n9332_);
  not g_6429 (not_new_n1723_, key_gate_120);
  not g_6430 (new_n9369_, new_n648_);
  and g_6431 (new_n5042_, and_new_n5289__new_n5287_, new_n5204_);
  not g_6432 (not_new_n7505_, new_n7505_);
  and g_6433 (new_n1182_, new_n1637_, new_n1635_);
  or g_6434 (po062, key_gate_82, not_new_n1189_);
  or g_6435 (new_n9160_, not_new_n8854__0, not_new_n9099__0);
  or g_6436 (new_n7243_, not_new_n7239_, not_new_n7241_);
  not g_6437 (not_new_n1598__16284135979104490, new_n1598_);
  and g_6438 (new_n7738_, new_n7968_, new_n7969_);
  not g_6439 (not_new_n1805__0, new_n1805_);
  not g_6440 (not_new_n1576__138412872010, new_n1576_);
  not g_6441 (not_new_n7448__1, new_n7448_);
  or g_6442 (new_n7033_, not_new_n7417_, not_new_n7416_);
  not g_6443 (not_new_n8830_, new_n8830_);
  not g_6444 (not_new_n631__24010, new_n631_);
  not g_6445 (not_new_n928__0, new_n928_);
  not g_6446 (not_new_n5394_, new_n5394_);
  not g_6447 (not_new_n2090_, new_n2090_);
  not g_6448 (not_new_n593__19773267430, new_n593_);
  or g_6449 (new_n8464_, not_new_n8110__0, not_new_n648__332329305696010);
  or g_6450 (new_n10179_, new_n637_, new_n1065_);
  not g_6451 (not_new_n4980_, new_n4980_);
  or g_6452 (new_n668_, or_not_new_n3167__not_new_n3166_, not_new_n3165_);
  or g_6453 (new_n9805_, not_new_n9521_, not_new_n9500_);
  or g_6454 (new_n6686_, not_new_n6576_, not_new_n6685_);
  not g_6455 (not_new_n621__138412872010, new_n621_);
  not g_6456 (not_new_n7150_, new_n7150_);
  or g_6457 (new_n4627_, not_new_n4482_, not_new_n4483__0);
  not g_6458 (new_n8707_, new_n1607_);
  or g_6459 (new_n2874_, not_new_n1599__1, not_new_n613__3);
  or g_6460 (new_n3522_, not_new_n1537__113988951853731430, not_pi127_0);
  not g_6461 (not_new_n1179_, new_n1179_);
  not g_6462 (not_new_n7166_, new_n7166_);
  or g_6463 (new_n9566_, not_new_n1039__113988951853731430, not_new_n628__273687473400809163430);
  not g_6464 (not_new_n7734_, new_n7734_);
  not g_6465 (not_pi199, pi199);
  not g_6466 (not_new_n4718_, new_n4718_);
  not g_6467 (not_new_n1059__2824752490, new_n1059_);
  not g_6468 (not_new_n8555_, new_n8555_);
  not g_6469 (not_new_n4186_, new_n4186_);
  not g_6470 (not_new_n2014_, new_n2014_);
  not g_6471 (not_new_n1055__332329305696010, new_n1055_);
  not g_6472 (not_new_n601__24010, new_n601_);
  or g_6473 (new_n5103_, new_n1047_, new_n634_);
  or g_6474 (or_or_not_new_n1920__not_new_n1921__not_new_n1923_, not_new_n1923_, or_not_new_n1920__not_new_n1921_);
  not g_6475 (not_new_n1788_, new_n1788_);
  or g_6476 (new_n5983_, not_new_n5982_, not_new_n5717_);
  not g_6477 (not_new_n7634_, new_n7634_);
  not g_6478 (not_new_n3381_, new_n3381_);
  or g_6479 (new_n6556_, not_new_n6930_, not_new_n6931_);
  not g_6480 (not_new_n1045__113988951853731430, new_n1045_);
  or g_6481 (new_n6565_, not_new_n6902_, not_new_n6901_);
  not g_6482 (not_pi156, pi156);
  not g_6483 (not_new_n1065__2824752490, new_n1065_);
  not g_6484 (new_n9092_, new_n8888_);
  not g_6485 (not_new_n608__1176490, new_n608_);
  or g_6486 (new_n5479_, not_new_n5615_, not_new_n5614_);
  or g_6487 (new_n2040_, not_new_n7693_, not_new_n1583__3430);
  and g_6488 (new_n8592_, new_n8591_, new_n8669_);
  or g_6489 (new_n10054_, new_n1045_, new_n635_);
  not g_6490 (not_new_n6109_, new_n6109_);
  not g_6491 (not_new_n7317_, new_n7317_);
  not g_6492 (not_new_n4531_, new_n4531_);
  not g_6493 (not_new_n2305_, new_n2305_);
  not g_6494 (new_n4987_, new_n630_);
  or g_6495 (new_n9769_, not_new_n9768_, not_new_n9767_);
  or g_6496 (new_n3726_, not_new_n3724_, not_new_n3725_);
  not g_6497 (not_new_n4925_, new_n4925_);
  and g_6498 (new_n5723_, new_n5714_, new_n5948_);
  not g_6499 (not_new_n8029_, new_n8029_);
  or g_6500 (po247, not_new_n3680_, not_new_n3681_);
  not g_6501 (not_new_n8519_, new_n8519_);
  or g_6502 (new_n5357_, not_new_n4987_, not_new_n1601__9);
  not g_6503 (not_new_n3310__168070, new_n3310_);
  not g_6504 (not_new_n4311_, new_n4311_);
  or g_6505 (new_n8521_, not_new_n8133__0, not_new_n629__968890104070);
  not g_6506 (not_new_n5475_, new_n5475_);
  or g_6507 (new_n6990_, not_new_n7320_, not_new_n6980_);
  or g_6508 (new_n10221_, not_new_n9948_, not_new_n9865_);
  not g_6509 (not_new_n766_, new_n766_);
  not g_6510 (not_new_n640__6782230728490, new_n640_);
  not g_6511 (new_n3444_, new_n1049_);
  and g_6512 (new_n8923_, new_n1037_, new_n632_);
  or g_6513 (new_n5119_, not_new_n1047__9, not_new_n634__24010);
  and g_6514 (and_and_new_n1735__new_n1736__new_n1738_, and_new_n1735__new_n1736_, new_n1738_);
  or g_6515 (new_n2041_, not_new_n5835_, not_new_n1585__3430);
  not g_6516 (not_new_n4831_, new_n4831_);
  not g_6517 (not_new_n743_, new_n743_);
  not g_6518 (new_n5790_, new_n1057_);
  not g_6519 (not_new_n9916_, new_n9916_);
  not g_6520 (not_new_n2055_, new_n2055_);
  or g_6521 (new_n1170_, not_new_n3869_, not_new_n3870_);
  not g_6522 (not_new_n8274_, new_n8274_);
  not g_6523 (not_new_n1047__57648010, new_n1047_);
  not g_6524 (not_new_n4211_, new_n4211_);
  and g_6525 (new_n6614_, new_n6837_, new_n6838_);
  or g_6526 (new_n8344_, not_new_n8153_, not_new_n644__6782230728490);
  or g_6527 (new_n5615_, not_new_n5536_, not_new_n5613_);
  not g_6528 (not_new_n10045__1, new_n10045_);
  not g_6529 (not_new_n6443__138412872010, new_n6443_);
  not g_6530 (not_new_n8648_, new_n8648_);
  or g_6531 (or_not_new_n3128__not_new_n3127_, not_new_n3127_, not_new_n3128_);
  not g_6532 (not_new_n9274_, new_n9274_);
  or g_6533 (new_n5482_, not_new_n5633_, not_new_n5634_);
  not g_6534 (not_new_n621__0, new_n621_);
  or g_6535 (new_n9527_, not_new_n9356_, not_new_n9357_);
  not g_6536 (not_new_n8944_, new_n8944_);
  not g_6537 (not_new_n598__7, new_n598_);
  not g_6538 (not_new_n7885_, new_n7885_);
  not g_6539 (not_new_n1325_, new_n1325_);
  not g_6540 (not_new_n617__968890104070, new_n617_);
  not g_6541 (not_new_n8716_, new_n8716_);
  not g_6542 (not_new_n1035__490, new_n1035_);
  not g_6543 (not_new_n10014_, new_n10014_);
  or g_6544 (new_n5588_, not_new_n5644_, not_new_n5432__0);
  and g_6545 (new_n8941_, new_n8979_, new_n9103_);
  or g_6546 (or_not_new_n2908__not_new_n2907_, not_new_n2907_, not_new_n2908_);
  not g_6547 (not_new_n3118_, new_n3118_);
  or g_6548 (new_n9879_, not_new_n635__16284135979104490, not_new_n1045__39098210485829880490);
  and g_6549 (new_n5506_, new_n5645_, new_n5646_);
  or g_6550 (new_n6394_, not_new_n6270_, not_new_n1057__3430);
  not g_6551 (not_new_n7029__1, new_n7029_);
  not g_6552 (not_new_n5756_, new_n5756_);
  not g_6553 (not_new_n733_, new_n733_);
  not g_6554 (not_new_n601_, new_n601_);
  and g_6555 (new_n8933_, new_n8992_, new_n9041_);
  not g_6556 (not_new_n3987_, key_gate_12);
  not g_6557 (not_new_n9780_, new_n9780_);
  not g_6558 (new_n8030_, new_n7724_);
  and g_6559 (and_new_n8664__new_n8663_, new_n8663_, new_n8664_);
  not g_6560 (new_n9024_, new_n8847_);
  or g_6561 (new_n3358_, not_new_n3916__0, not_pi064_2824752490);
  not g_6562 (not_new_n8415_, new_n8415_);
  or g_6563 (or_not_new_n3143__not_new_n3142_, not_new_n3142_, not_new_n3143_);
  not g_6564 (not_new_n1065__8, new_n1065_);
  not g_6565 (not_new_n7875_, new_n7875_);
  not g_6566 (not_new_n7624_, new_n7624_);
  not g_6567 (new_n2209_, new_n629_);
  not g_6568 (not_new_n6724_, new_n6724_);
  not g_6569 (not_new_n3370_, new_n3370_);
  not g_6570 (not_new_n935_, new_n935_);
  or g_6571 (new_n5491_, not_new_n5703_, not_new_n5704_);
  or g_6572 (new_n2856_, not_new_n1043__1, not_new_n3311__9);
  or g_6573 (new_n7799_, not_new_n7767_, not_new_n648__138412872010);
  not g_6574 (not_new_n8838__0, new_n8838_);
  or g_6575 (new_n4635_, not_new_n4517_, not_new_n4633_);
  not g_6576 (new_n8626_, new_n1067_);
  not g_6577 (not_new_n4115__0, new_n4115_);
  or g_6578 (new_n3320_, not_new_n3926__0, not_pi064_2);
  not g_6579 (not_new_n9808_, new_n9808_);
  not g_6580 (not_new_n1067__9, new_n1067_);
  and g_6581 (new_n1500_, new_n1501_, new_n3025_);
  or g_6582 (new_n9710_, not_new_n9467_, not_new_n9427__2);
  not g_6583 (not_new_n5849_, new_n5849_);
  not g_6584 (not_new_n4165__0, new_n4165_);
  not g_6585 (not_new_n3937_, new_n3937_);
  not g_6586 (not_new_n618__657123623635342801395430, new_n618_);
  or g_6587 (new_n7353_, not_new_n772_, not_new_n6974__4);
  not g_6588 (not_new_n984__24010, new_n984_);
  or g_6589 (new_n2967_, not_new_n7066_, not_new_n595__47475615099430);
  not g_6590 (not_new_n3926__0, new_n3926_);
  and g_6591 (new_n8215_, new_n8091_, new_n8373_);
  not g_6592 (not_new_n7876__0, new_n7876_);
  not g_6593 (not_new_n5219__0, new_n5219_);
  not g_6594 (not_new_n599__9, new_n599_);
  not g_6595 (not_new_n7686_, new_n7686_);
  or g_6596 (new_n5279_, not_new_n4908_, not_new_n4996_);
  not g_6597 (not_new_n9843_, new_n9843_);
  or g_6598 (po128, not_new_n3455_, not_new_n3456_);
  or g_6599 (new_n4217_, not_pi272_2, not_new_n4086_);
  or g_6600 (new_n5675_, not_new_n5465__1, not_pi144_3);
  or g_6601 (new_n7939_, not_new_n7706_, not_new_n7735__2);
  or g_6602 (new_n5286_, not_new_n5192_, not_new_n5195__0);
  or g_6603 (new_n5902_, not_new_n5802_, not_new_n5986_);
  not g_6604 (not_new_n7760_, new_n7760_);
  or g_6605 (new_n9278_, not_new_n9130_, not_new_n8971_);
  not g_6606 (not_new_n5226_, new_n5226_);
  not g_6607 (not_new_n9504_, new_n9504_);
  not g_6608 (not_new_n1500_, new_n1500_);
  not g_6609 (not_new_n598__47475615099430, new_n598_);
  or g_6610 (new_n5235_, not_new_n4984__0, not_new_n5166_);
  or g_6611 (new_n2594_, not_new_n607__6, not_new_n1019_);
  not g_6612 (not_new_n9287_, new_n9287_);
  not g_6613 (not_po296_7490483309651862334944941026945644936490, po296);
  or g_6614 (new_n3772_, not_new_n3494_, not_new_n2095_);
  not g_6615 (not_new_n637__1176490, new_n637_);
  and g_6616 (new_n8216_, new_n8374_, new_n8428_);
  not g_6617 (not_new_n4131__0, new_n4131_);
  not g_6618 (not_new_n7659_, new_n7659_);
  not g_6619 (not_new_n4454__0, new_n4454_);
  or g_6620 (new_n2315_, not_new_n593__2326305139872070, not_new_n619_);
  or g_6621 (new_n5090_, new_n624_, new_n1041_);
  not g_6622 (not_new_n4517_, new_n4517_);
  or g_6623 (new_n10254_, not_new_n1043__16284135979104490, not_new_n9887_);
  not g_6624 (not_new_n601__1, new_n601_);
  or g_6625 (new_n9824_, not_new_n9385_, not_new_n638__657123623635342801395430);
  not g_6626 (not_pi034_3, pi034);
  not g_6627 (not_pi044, pi044);
  not g_6628 (not_new_n2020_, new_n2020_);
  or g_6629 (new_n1055_, not_new_n3457_, not_new_n3458_);
  not g_6630 (not_new_n640__138412872010, new_n640_);
  not g_6631 (new_n5781_, new_n1071_);
  or g_6632 (new_n5690_, not_new_n5688_, not_new_n1016__6);
  not g_6633 (not_new_n3184__4, new_n3184_);
  not g_6634 (not_new_n2256_, new_n2256_);
  not g_6635 (not_new_n986__0, new_n986_);
  not g_6636 (not_new_n1360_, new_n1360_);
  not g_6637 (not_new_n4436_, new_n4436_);
  or g_6638 (new_n1910_, not_new_n8191_, not_new_n1581__6);
  not g_6639 (not_new_n627__4, new_n627_);
  and g_6640 (new_n7713_, new_n7868_, new_n7985_);
  not g_6641 (not_new_n6519__2, new_n6519_);
  not g_6642 (new_n4832_, new_n4790_);
  not g_6643 (not_new_n1389_, new_n1389_);
  or g_6644 (new_n2570_, not_new_n608__5, not_new_n1016__0);
  not g_6645 (not_new_n5174_, new_n5174_);
  not g_6646 (new_n1599_, new_n973_);
  or g_6647 (new_n3421_, not_new_n1843_, not_new_n1613__2);
  or g_6648 (new_n975_, not_pi006, not_new_n1536__5);
  not g_6649 (new_n9936_, new_n1599_);
  or g_6650 (new_n2807_, not_pi254, not_po296_2569235775210588780886114772242356213216070);
  not g_6651 (new_n4274_, new_n687_);
  not g_6652 (not_new_n2092_, new_n2092_);
  not g_6653 (not_new_n9973_, new_n9973_);
  not g_6654 (not_new_n1049__4, new_n1049_);
  or g_6655 (new_n2360_, not_new_n1035__0, not_new_n598__0);
  not g_6656 (not_new_n8095_, new_n8095_);
  or g_6657 (po118, not_new_n3406_, not_new_n3405_);
  not g_6658 (not_new_n5311_, new_n5311_);
  not g_6659 (new_n7629_, new_n639_);
  not g_6660 (new_n5445_, pi136);
  not g_6661 (not_new_n1307_, new_n1307_);
  not g_6662 (new_n5110_, new_n5056_);
  or g_6663 (new_n4867_, not_new_n4838_, not_new_n4772__0);
  not g_6664 (new_n9521_, new_n9499_);
  or g_6665 (new_n9704_, not_new_n9465_, not_new_n9506__2);
  or g_6666 (new_n7301_, not_new_n6977__1, not_new_n7195_);
  not g_6667 (not_new_n7160__0, new_n7160_);
  or g_6668 (new_n7231_, not_new_n7003_, not_new_n7433_);
  or g_6669 (po148, not_new_n3523_, not_new_n3522_);
  and g_6670 (new_n8810_, new_n8808_, new_n8803_);
  or g_6671 (new_n2544_, not_new_n1014_, not_new_n607__1);
  not g_6672 (not_new_n9993_, new_n9993_);
  or g_6673 (new_n712_, not_new_n1528_, not_new_n3084_);
  not g_6674 (not_new_n10331_, new_n10331_);
  not g_6675 (not_new_n622__4, new_n622_);
  not g_6676 (not_new_n8263_, new_n8263_);
  or g_6677 (new_n4643_, not_pi162_2, not_new_n4415__0);
  not g_6678 (not_new_n9178_, new_n9178_);
  not g_6679 (not_new_n4000_, new_n4000_);
  not g_6680 (not_new_n7916_, new_n7916_);
  or g_6681 (new_n949_, or_or_not_new_n1251__not_new_n1249__not_new_n1888_, not_new_n1887_);
  not g_6682 (not_new_n595__138412872010, new_n595_);
  or g_6683 (new_n3060_, not_new_n1027__332329305696010, not_new_n1172_);
  or g_6684 (new_n5401_, not_new_n5075_, not_new_n5074_);
  not g_6685 (not_new_n5676_, new_n5676_);
  and g_6686 (new_n1476_, new_n1477_, new_n2767_);
  not g_6687 (not_new_n588__47475615099430, new_n588_);
  not g_6688 (not_new_n1027__3, new_n1027_);
  or g_6689 (new_n3034_, not_new_n629__4, not_new_n3372__57648010);
  not g_6690 (not_new_n5492_, new_n5492_);
  or g_6691 (new_n7069_, not_new_n7564_, not_new_n7563_);
  not g_6692 (not_new_n6749_, new_n6749_);
  not g_6693 (not_new_n9952_, new_n9952_);
  not g_6694 (not_new_n1027__24010, new_n1027_);
  or g_6695 (new_n7198_, not_new_n7197_, not_new_n7076_);
  and g_6696 (and_new_n6227__new_n6232_, new_n6232_, new_n6227_);
  not g_6697 (not_new_n1604__24010, new_n1604_);
  or g_6698 (new_n7941_, not_new_n7620_, not_new_n7695_);
  not g_6699 (not_new_n6682_, new_n6682_);
  not g_6700 (not_new_n3315__3, new_n3315_);
  not g_6701 (not_new_n602__490, new_n602_);
  and g_6702 (new_n3934_, new_n3954_, new_n4006_);
  and g_6703 (new_n4290_, new_n4229_, new_n709_);
  not g_6704 (not_new_n4288_, new_n4288_);
  not g_6705 (not_new_n9564_, new_n9564_);
  not g_6706 (not_pi246_0, pi246);
  not g_6707 (not_new_n1613__403536070, new_n1613_);
  or g_6708 (new_n6602_, not_new_n6913_, not_new_n6912_);
  not g_6709 (not_pi143_0, pi143);
  not g_6710 (not_new_n7754__1, new_n7754_);
  not g_6711 (not_new_n7478_, new_n7478_);
  and g_6712 (new_n6313_, new_n6385_, new_n6386_);
  not g_6713 (not_new_n9030_, new_n9030_);
  not g_6714 (not_new_n1009__3, new_n1009_);
  or g_6715 (new_n7029_, not_new_n7425_, not_new_n7426_);
  not g_6716 (not_new_n1612__1, new_n1612_);
  not g_6717 (not_new_n5900__3, new_n5900_);
  or g_6718 (new_n1868_, not_new_n624__0, not_new_n601__3);
  not g_6719 (not_new_n6512_, new_n6512_);
  and g_6720 (new_n1559_, new_n3630_, new_n3631_);
  or g_6721 (new_n6513_, not_new_n645__57648010, not_new_n6514_);
  not g_6722 (not_new_n619__3430, new_n619_);
  not g_6723 (not_new_n4792_, new_n4792_);
  xor g_6724 (key_gate_95, not_new_n1726_, key_95);
  not g_6725 (not_new_n5878__1, new_n5878_);
  or g_6726 (new_n3802_, not_new_n3489_, not_new_n2076_);
  or g_6727 (new_n5555_, new_n1018_, pi140);
  or g_6728 (new_n7587_, not_new_n7899_, not_new_n7902_);
  or g_6729 (new_n2344_, not_new_n1606_, not_new_n1588__797922662976120010);
  not g_6730 (new_n1587_, new_n985_);
  or g_6731 (new_n5447_, not_new_n5543_, not_new_n5542_);
  not g_6732 (not_new_n5904_, new_n5904_);
  or g_6733 (new_n4392_, not_new_n4279_, not_new_n685_);
  not g_6734 (not_new_n639__0, new_n639_);
  not g_6735 (not_new_n646__332329305696010, new_n646_);
  or g_6736 (new_n9740_, not_new_n9354_, not_new_n1041__968890104070);
  not g_6737 (new_n1609_, new_n940_);
  or g_6738 (new_n7807_, not_new_n7774__0, not_new_n7597__1);
  or g_6739 (new_n3592_, not_pi162_0, not_new_n984__0);
  not g_6740 (not_new_n9840_, new_n9840_);
  or g_6741 (new_n2474_, not_new_n9964__0, not_new_n599__968890104070);
  not g_6742 (not_new_n1063__403536070, new_n1063_);
  not g_6743 (not_new_n1657_, key_gate_22);
  not g_6744 (not_new_n1589__2824752490, new_n1589_);
  not g_6745 (not_new_n5545_, new_n5545_);
  not g_6746 (not_new_n9898_, new_n9898_);
  not g_6747 (not_new_n9936_, new_n9936_);
  and g_6748 (and_new_n7605__new_n7973_, new_n7605_, new_n7973_);
  or g_6749 (or_not_new_n1548__not_new_n1366_, not_new_n1366_, not_new_n1548_);
  buf g_6750 (po019, pi212);
  not g_6751 (new_n6208_, new_n5873_);
  or g_6752 (new_n9570_, not_new_n9568_, not_new_n9461_);
  not g_6753 (new_n10045_, new_n9893_);
  not g_6754 (not_new_n635__8, new_n635_);
  not g_6755 (not_pi152, pi152);
  or g_6756 (new_n5164_, new_n1063_, new_n638_);
  or g_6757 (new_n3771_, not_new_n3770_, not_new_n3769_);
  or g_6758 (new_n4813_, not_new_n4737__0, not_new_n4812__0);
  or g_6759 (new_n5069_, not_new_n5278_, not_new_n5280_);
  or g_6760 (new_n8126_, not_new_n8321_, not_new_n8121_);
  not g_6761 (not_new_n602__47475615099430, new_n602_);
  not g_6762 (not_new_n6069_, new_n6069_);
  or g_6763 (new_n9931_, not_new_n10217_, not_new_n10105_);
  and g_6764 (new_n8804_, new_n9075_, new_n9076_);
  or g_6765 (new_n5981_, not_new_n5786_, not_new_n638__1176490);
  not g_6766 (not_new_n5860_, new_n5860_);
  xnor g_6767 (key_gate_87, key_87, not_new_n1636_);
  or g_6768 (new_n8568_, not_new_n8400_, not_new_n8177__0);
  not g_6769 (not_new_n3247_, new_n3247_);
  not g_6770 (not_new_n5565_, new_n5565_);
  or g_6771 (new_n7063_, not_new_n7523_, not_new_n7524_);
  not g_6772 (not_new_n998__0, new_n998_);
  not g_6773 (not_new_n1402_, new_n1402_);
  not g_6774 (not_new_n9727_, new_n9727_);
  not g_6775 (not_pi032_0, pi032);
  not g_6776 (not_new_n5078__0, new_n5078_);
  and g_6777 (and_new_n1302__new_n2141_, new_n1302_, new_n2141_);
  and g_6778 (new_n1396_, new_n2476_, new_n2475_);
  not g_6779 (not_new_n1028__1, new_n1028_);
  or g_6780 (new_n2167_, not_pi183, not_new_n586__19773267430);
  not g_6781 (not_new_n4074_, new_n4074_);
  not g_6782 (new_n4789_, new_n1069_);
  not g_6783 (not_new_n7040__0, new_n7040_);
  not g_6784 (not_new_n1059__113988951853731430, new_n1059_);
  not g_6785 (not_new_n3992_, key_gate_56);
  not g_6786 (not_new_n618__1915812313805664144010, new_n618_);
  not g_6787 (new_n5787_, new_n1061_);
  not g_6788 (not_new_n10059_, new_n10059_);
  and g_6789 (new_n1267_, new_n1969_, and_new_n1266__new_n1970_);
  or g_6790 (new_n9787_, not_new_n9415__0, not_new_n1601__273687473400809163430);
  not g_6791 (not_new_n602__403536070, new_n602_);
  or g_6792 (or_or_or_not_new_n6363__not_new_n6358__not_new_n6361__not_new_n6366_, or_or_not_new_n6363__not_new_n6358__not_new_n6361_, not_new_n6366_);
  not g_6793 (not_new_n1002__0, new_n1002_);
  not g_6794 (not_new_n1049__8, new_n1049_);
  not g_6795 (not_new_n3222_, new_n3222_);
  and g_6796 (new_n1470_, pi275, new_n923_);
  and g_6797 (and_new_n7159__new_n7547_, new_n7159_, new_n7547_);
  not g_6798 (not_new_n3316_, new_n3316_);
  not g_6799 (not_new_n6443__797922662976120010, new_n6443_);
  not g_6800 (not_new_n1063__490, new_n1063_);
  not g_6801 (not_new_n8874__0, new_n8874_);
  not g_6802 (not_new_n2248_, new_n2248_);
  not g_6803 (not_new_n644__8, new_n644_);
  or g_6804 (new_n1982_, not_new_n626__0, not_new_n601__9);
  not g_6805 (not_new_n648__19773267430, new_n648_);
  not g_6806 (not_new_n7220_, new_n7220_);
  or g_6807 (new_n2339_, not_pi192, not_new_n586__797922662976120010);
  and g_6808 (po106, key_gate_101, pi085);
  not g_6809 (not_new_n1604__47475615099430, new_n1604_);
  or g_6810 (new_n7386_, not_new_n6979__1, not_new_n7022__1);
  not g_6811 (not_new_n3483_, new_n3483_);
  or g_6812 (new_n2799_, not_new_n604__7, not_new_n645__3);
  not g_6813 (not_new_n1011__6, new_n1011_);
  not g_6814 (new_n4162_, new_n4150_);
  not g_6815 (not_new_n1631__7, key_gate_76);
  or g_6816 (new_n6845_, not_new_n631__968890104070, not_new_n6475__2);
  or g_6817 (new_n10270_, not_new_n10008__0, not_new_n1607__19773267430);
  or g_6818 (new_n2320_, not_new_n587__113988951853731430, not_pi159);
  not g_6819 (not_new_n5927_, new_n5927_);
  and g_6820 (and_and_new_n1460__new_n1466__new_n1458_, and_new_n1460__new_n1466_, new_n1458_);
  not g_6821 (new_n3951_, pi051);
  or g_6822 (new_n674_, not_new_n3095_, or_not_new_n3097__not_new_n3096_);
  or g_6823 (new_n3466_, not_new_n1613__70, not_new_n2014_);
  not g_6824 (not_new_n7439__0, new_n7439_);
  not g_6825 (not_new_n622__2, new_n622_);
  or g_6826 (new_n3239_, not_new_n589__47475615099430, not_new_n626__7);
  or g_6827 (new_n7946_, not_new_n7755_, not_new_n7845_);
  not g_6828 (not_new_n9181_, new_n9181_);
  not g_6829 (not_new_n3449_, new_n3449_);
  not g_6830 (not_new_n7003__0, new_n7003_);
  not g_6831 (not_new_n10277_, new_n10277_);
  not g_6832 (not_new_n1041__57648010, new_n1041_);
  or g_6833 (new_n8310_, not_new_n8104_, not_new_n8105__0);
  or g_6834 (new_n5992_, not_new_n5782_, not_new_n1069__10);
  and g_6835 (new_n4493_, new_n4660_, new_n4661_);
  or g_6836 (new_n7959_, not_new_n7807_, not_new_n7618__0);
  and g_6837 (new_n1509_, new_n998_, new_n3036_);
  or g_6838 (new_n6912_, not_new_n6485_, not_new_n1035__10);
  not g_6839 (new_n7218_, new_n7150_);
  not g_6840 (not_new_n4116__0, new_n4116_);
  not g_6841 (not_new_n8170__0, new_n8170_);
  not g_6842 (not_pi052_2, pi052);
  not g_6843 (not_new_n9086__0, new_n9086_);
  not g_6844 (not_new_n721_, new_n721_);
  not g_6845 (new_n7648_, new_n627_);
  not g_6846 (not_new_n5075_, new_n5075_);
  not g_6847 (not_pi234, pi234);
  not g_6848 (not_new_n3066_, new_n3066_);
  not g_6849 (not_new_n585__5, new_n585_);
  not g_6850 (not_new_n1581__797922662976120010, new_n1581_);
  not g_6851 (not_pi165_3, pi165);
  not g_6852 (not_new_n8966__0, new_n8966_);
  or g_6853 (new_n9251_, not_new_n8852_, not_new_n629__47475615099430);
  not g_6854 (not_new_n7803_, new_n7803_);
  or g_6855 (new_n3895_, not_new_n9925_, not_new_n1055__7);
  or g_6856 (new_n1667_, not_new_n1631__10, not_pi044);
  and g_6857 (and_new_n8082__new_n8430_, new_n8082_, new_n8430_);
  not g_6858 (new_n2133_, new_n640_);
  not g_6859 (not_new_n3704_, new_n3704_);
  or g_6860 (new_n10199_, not_new_n9919__0, not_new_n10059__0);
  or g_6861 (new_n7382_, not_new_n7321__0, not_new_n7380_);
  not g_6862 (not_new_n609__8235430, new_n609_);
  or g_6863 (new_n2515_, or_not_new_n4461__not_new_n609__0, not_new_n611__2);
  not g_6864 (not_new_n7356_, new_n7356_);
  or g_6865 (new_n4018_, not_new_n3913__0, or_or_not_new_n3944__not_new_n3914__1_not_new_n4014__4);
  not g_6866 (not_new_n2555_, new_n2555_);
  or g_6867 (new_n7461_, not_new_n7460_, not_new_n746_);
  not g_6868 (not_new_n6831_, new_n6831_);
  not g_6869 (not_new_n638__490, new_n638_);
  or g_6870 (new_n6027_, not_new_n5916_, not_new_n5813_);
  not g_6871 (not_new_n10272_, new_n10272_);
  not g_6872 (not_new_n5059_, new_n5059_);
  not g_6873 (not_new_n1195_, new_n1195_);
  or g_6874 (new_n2551_, not_new_n606__3, not_new_n5487__0);
  or g_6875 (new_n5802_, not_new_n5985_, not_new_n5983_);
  and g_6876 (new_n6454_, new_n6446_, new_n6683_);
  not g_6877 (not_new_n628__24010, new_n628_);
  or g_6878 (po205, not_new_n1394_, or_or_not_new_n1562__not_new_n2469__not_new_n1393_);
  or g_6879 (new_n990_, not_new_n582_, not_new_n583_);
  or g_6880 (new_n2244_, not_pi155, not_new_n587__47475615099430);
  not g_6881 (not_pi080, pi080);
  or g_6882 (new_n3912_, not_new_n10026_, not_new_n10025_);
  not g_6883 (not_new_n8096_, new_n8096_);
  not g_6884 (new_n8162_, new_n637_);
  not g_6885 (not_new_n4463_, new_n4463_);
  or g_6886 (new_n3268_, not_new_n3184__10, not_new_n629__8);
  or g_6887 (new_n3536_, not_new_n1538__4, not_pi134_0);
  not g_6888 (new_n4809_, new_n1053_);
  not g_6889 (not_new_n8978__1, new_n8978_);
  not g_6890 (not_new_n7456_, new_n7456_);
  or g_6891 (new_n10245_, not_new_n10243_, not_new_n10224_);
  not g_6892 (not_new_n3385_, new_n3385_);
  not g_6893 (not_new_n4998__1, new_n4998_);
  not g_6894 (new_n1791_, new_n641_);
  not g_6895 (not_new_n5708_, new_n5708_);
  or g_6896 (or_not_new_n2794__not_new_n2797_, not_new_n2794_, not_new_n2797_);
  or g_6897 (new_n3649_, not_new_n2334_, not_new_n1611__16284135979104490);
  not g_6898 (not_new_n2933_, new_n2933_);
  or g_6899 (new_n7662_, not_new_n621__19773267430, not_new_n7621_);
  not g_6900 (not_new_n1765_, new_n1765_);
  not g_6901 (not_new_n5159_, new_n5159_);
  and g_6902 (new_n4905_, new_n5177_, new_n4904_);
  or g_6903 (new_n2137_, not_new_n9443_, not_new_n1584__57648010);
  or g_6904 (new_n3540_, not_pi136_0, not_new_n1538__6);
  or g_6905 (new_n2976_, not_new_n595__332329305696010, not_new_n7055_);
  not g_6906 (not_new_n6905_, new_n6905_);
  not g_6907 (new_n7616_, new_n1051_);
  or g_6908 (new_n6032_, not_new_n5801__0, not_new_n5984__0);
  or g_6909 (new_n3676_, not_pi224, not_new_n989__10);
  not g_6910 (not_new_n6373__9, new_n6373_);
  or g_6911 (new_n8369_, not_new_n1601__47475615099430, not_new_n8134__0);
  not g_6912 (not_new_n6527__1, new_n6527_);
  not g_6913 (new_n1810_, new_n628_);
  not g_6914 (new_n6507_, new_n1602_);
  or g_6915 (new_n6637_, not_new_n6535_, not_new_n6721_);
  not g_6916 (not_new_n3758_, new_n3758_);
  or g_6917 (new_n7956_, not_new_n7955_, not_new_n7954_);
  not g_6918 (not_new_n1049__5, new_n1049_);
  not g_6919 (not_new_n1043__6, new_n1043_);
  not g_6920 (not_new_n1588__490, new_n1588_);
  not g_6921 (not_new_n8319_, new_n8319_);
  not g_6922 (not_new_n4464__0, new_n4464_);
  or g_6923 (new_n2572_, not_pi199, not_new_n2509__5);
  not g_6924 (not_new_n1043__168070, new_n1043_);
  or g_6925 (new_n10015_, not_new_n10146_, not_new_n10147_);
  not g_6926 (not_new_n6330_, new_n6330_);
  or g_6927 (new_n9032_, not_new_n8828__0, not_new_n9028_);
  not g_6928 (new_n1572_, new_n6243_);
  not g_6929 (not_new_n5655_, new_n5655_);
  not g_6930 (not_new_n7139_, new_n7139_);
  not g_6931 (not_new_n5669_, new_n5669_);
  not g_6932 (not_new_n4372_, new_n4372_);
  not g_6933 (not_new_n628__93874803376477543056490, new_n628_);
  or g_6934 (new_n7273_, not_new_n719__0, not_new_n7043__0);
  not g_6935 (not_new_n5919_, new_n5919_);
  not g_6936 (not_new_n6930_, new_n6930_);
  not g_6937 (not_new_n4411_, new_n4411_);
  not g_6938 (not_new_n6998__1, new_n6998_);
  not g_6939 (not_new_n5764_, new_n5764_);
  not g_6940 (not_new_n6813_, new_n6813_);
  not g_6941 (not_new_n6597_, new_n6597_);
  not g_6942 (not_new_n3514_, new_n3514_);
  or g_6943 (new_n1004_, not_new_n3330_, not_new_n3329_);
  or g_6944 (new_n6798_, not_new_n6596_, not_new_n6631__0);
  not g_6945 (not_new_n646_, new_n646_);
  not g_6946 (not_new_n629__24010, new_n629_);
  or g_6947 (new_n5960_, not_new_n5920__0, not_new_n5762_);
  not g_6948 (not_pi254_1, pi254);
  not g_6949 (not_new_n1585__6, new_n1585_);
  not g_6950 (not_new_n632__5, new_n632_);
  or g_6951 (new_n7727_, not_new_n8044_, not_new_n8043_);
  and g_6952 (new_n1389_, new_n2457_, new_n2458_);
  not g_6953 (not_new_n1538__968890104070, new_n1538_);
  or g_6954 (new_n4680_, not_new_n4678_, not_new_n4565_);
  not g_6955 (not_new_n7150__0, new_n7150_);
  not g_6956 (not_new_n1021_, new_n1021_);
  not g_6957 (not_new_n627__57648010, new_n627_);
  not g_6958 (not_new_n8138__1, new_n8138_);
  or g_6959 (new_n8878_, not_new_n646__6782230728490, not_new_n1069__2824752490);
  or g_6960 (or_not_new_n1556__not_new_n2439_, not_new_n2439_, not_new_n1556_);
  or g_6961 (new_n4152_, not_new_n4157__0, not_pi270_1);
  not g_6962 (not_new_n7357_, new_n7357_);
  or g_6963 (new_n9853_, not_new_n9360_, not_new_n1031__19773267430);
  not g_6964 (not_new_n620__6, new_n620_);
  not g_6965 (not_new_n6070_, new_n6070_);
  not g_6966 (not_new_n8550_, new_n8550_);
  not g_6967 (not_new_n6824_, new_n6824_);
  not g_6968 (not_new_n10179_, new_n10179_);
  not g_6969 (new_n8427_, new_n8173_);
  not g_6970 (not_new_n6338_, new_n6338_);
  or g_6971 (new_n3053_, not_new_n1069__2, not_new_n581__19773267430);
  not g_6972 (not_new_n955_, new_n955_);
  not g_6973 (not_new_n1696_, key_gate_2);
  not g_6974 (not_new_n6042_, new_n6042_);
  not g_6975 (not_new_n5244_, new_n5244_);
  not g_6976 (not_new_n1616__0, new_n1616_);
  not g_6977 (new_n8987_, new_n8854_);
  and g_6978 (new_n8939_, new_n8810_, new_n9090_);
  not g_6979 (not_new_n3561_, new_n3561_);
  not g_6980 (not_new_n3387__4, new_n3387_);
  or g_6981 (new_n4647_, not_new_n4509_, not_pi162_3);
  and g_6982 (new_n9330_, new_n9580_, new_n9579_);
  or g_6983 (new_n9133_, not_new_n8899__0, not_new_n9132_);
  not g_6984 (new_n8156_, new_n626_);
  not g_6985 (not_new_n7119_, new_n7119_);
  not g_6986 (not_new_n1604__2824752490, new_n1604_);
  not g_6987 (not_new_n5105_, new_n5105_);
  or g_6988 (new_n2682_, not_new_n2509__1176490, not_pi210);
  not g_6989 (not_new_n2745_, new_n2745_);
  not g_6990 (not_new_n2821_, new_n2821_);
  not g_6991 (new_n5772_, new_n639_);
  or g_6992 (or_not_new_n2339__not_new_n2340_, not_new_n2339_, not_new_n2340_);
  and g_6993 (new_n6460_, new_n6459_, new_n6740_);
  or g_6994 (new_n7471_, not_new_n7137__0, not_new_n7136_);
  not g_6995 (not_new_n5779__0, new_n5779_);
  not g_6996 (not_new_n1039__168070, new_n1039_);
  or g_6997 (new_n8567_, not_new_n638__39098210485829880490, not_new_n8150__2);
  not g_6998 (new_n4938_, new_n1047_);
  or g_6999 (new_n4123_, not_new_n4198_, not_new_n4197_);
  or g_7000 (new_n3569_, not_new_n2185__0, not_new_n1612__2824752490);
  not g_7001 (new_n3484_, new_n1065_);
  or g_7002 (new_n9125_, not_new_n9124_, not_new_n8948_);
  or g_7003 (po127, not_new_n3451_, not_new_n3450_);
  not g_7004 (not_new_n1065__403536070, new_n1065_);
  not g_7005 (not_new_n604__490, new_n604_);
  not g_7006 (new_n6282_, new_n642_);
  not g_7007 (new_n9392_, new_n1055_);
  not g_7008 (not_new_n9427__0, new_n9427_);
  xnor g_7009 (key_gate_121, not_new_n3933_, key_121);
  or g_7010 (new_n2847_, not_new_n1067__1, not_new_n3311__8);
  or g_7011 (new_n10335_, not_new_n9912_, not_new_n637__113988951853731430);
  not g_7012 (not_new_n8117__1, new_n8117_);
  and g_7013 (new_n5067_, new_n5357_, new_n5356_);
  and g_7014 (new_n1356_, new_n2375_, and_new_n1543__new_n2376_);
  not g_7015 (not_new_n622__9, new_n622_);
  not g_7016 (not_new_n8362_, new_n8362_);
  not g_7017 (not_new_n5703_, new_n5703_);
  not g_7018 (not_new_n5445__0, new_n5445_);
  not g_7019 (not_new_n9802_, new_n9802_);
  not g_7020 (not_new_n7217_, new_n7217_);
  not g_7021 (not_new_n5026_, new_n5026_);
  not g_7022 (not_new_n8744_, new_n8744_);
  or g_7023 (new_n3077_, not_new_n1053__3, not_new_n581__113988951853731430);
  not g_7024 (not_new_n3507_, new_n3507_);
  not g_7025 (not_new_n732__0, new_n732_);
  not g_7026 (not_new_n1059__3430, new_n1059_);
  not g_7027 (not_new_n8017_, new_n8017_);
  not g_7028 (not_new_n6786_, new_n6786_);
  not g_7029 (not_new_n643__4, new_n643_);
  not g_7030 (not_pi249_0, pi249);
  not g_7031 (not_new_n9617_, new_n9617_);
  or g_7032 (new_n9947_, not_new_n10155_, not_new_n9940_);
  and g_7033 (new_n3924_, new_n3989_, new_n4035_);
  not g_7034 (not_new_n622__2824752490, new_n622_);
  and g_7035 (new_n8596_, new_n8768_, and_new_n8664__new_n8663_);
  not g_7036 (new_n9385_, new_n1063_);
  not g_7037 (not_new_n1059__6782230728490, new_n1059_);
  not g_7038 (new_n4014_, new_n3941_);
  or g_7039 (new_n6020_, not_new_n6019_, not_new_n5893_);
  and g_7040 (new_n7711_, new_n7771_, new_n7862_);
  not g_7041 (not_new_n5530_, new_n5530_);
  not g_7042 (new_n8517_, new_n8225_);
  not g_7043 (not_new_n1354_, new_n1354_);
  or g_7044 (po169, not_new_n3564_, not_new_n3565_);
  not g_7045 (not_pi008_0, pi008);
  not g_7046 (not_new_n5056_, new_n5056_);
  not g_7047 (new_n6287_, new_n1043_);
  not g_7048 (not_new_n1602__10, new_n1602_);
  or g_7049 (new_n7420_, not_new_n6974__24010, not_new_n760_);
  and g_7050 (new_n1490_, new_n2999_, and_new_n3001__new_n998_);
  not g_7051 (new_n8855_, new_n1602_);
  not g_7052 (new_n9698_, new_n9424_);
  not g_7053 (not_new_n6565_, new_n6565_);
  and g_7054 (new_n1185_, new_n1644_, new_n1646_);
  not g_7055 (not_new_n3315__403536070, new_n3315_);
  not g_7056 (not_new_n7247_, new_n7247_);
  or g_7057 (new_n5952_, not_new_n5921_, not_new_n5761_);
  not g_7058 (not_new_n8121__0, new_n8121_);
  not g_7059 (new_n4941_, new_n648_);
  and g_7060 (new_n1255_, and_new_n1254__new_n1913_, new_n1912_);
  not g_7061 (not_new_n7306_, new_n7306_);
  not g_7062 (not_new_n1006__5, new_n1006_);
  not g_7063 (not_new_n2501_, new_n2501_);
  or g_7064 (new_n3810_, not_new_n3809_, not_new_n3808_);
  or g_7065 (new_n3650_, not_new_n984__113988951853731430, not_pi191_0);
  not g_7066 (new_n1631_, key_gate_77);
  not g_7067 (not_new_n7418__0, new_n7418_);
  not g_7068 (not_new_n6311_, new_n6311_);
  not g_7069 (new_n5430_, new_n1010_);
  not g_7070 (not_new_n1063__57648010, new_n1063_);
  not g_7071 (not_new_n4564_, new_n4564_);
  not g_7072 (not_new_n9073_, new_n9073_);
  not g_7073 (not_new_n8287_, new_n8287_);
  not g_7074 (not_new_n5771__0, new_n5771_);
  or g_7075 (or_not_new_n1283__not_new_n1281_, not_new_n1281_, not_new_n1283_);
  not g_7076 (not_new_n5856_, new_n5856_);
  or g_7077 (new_n4115_, not_new_n4181_, not_new_n4182_);
  not g_7078 (not_new_n5885__0, new_n5885_);
  or g_7079 (new_n3506_, not_new_n1537__19773267430, not_pi119_0);
  not g_7080 (not_new_n7161_, new_n7161_);
  or g_7081 (new_n5643_, not_new_n5519__0, not_new_n5430_);
  and g_7082 (new_n5728_, new_n5725_, new_n5727_);
  not g_7083 (not_new_n6216_, new_n6216_);
  or g_7084 (new_n8776_, or_or_not_new_n8696__not_new_n8690__not_new_n8689_, not_new_n8688_);
  or g_7085 (new_n6425_, or_or_or_not_new_n6226__0_not_new_n6336__not_new_n6373__5_not_new_n6242__2, not_new_n1059__24010);
  not g_7086 (new_n6066_, new_n5891_);
  not g_7087 (not_new_n1011__2, new_n1011_);
  or g_7088 (new_n8197_, not_new_n8537_, not_new_n8536_);
  not g_7089 (not_new_n608__0, new_n608_);
  not g_7090 (not_new_n8192_, new_n8192_);
  not g_7091 (not_new_n8286__0, new_n8286_);
  not g_7092 (new_n6658_, new_n6508_);
  or g_7093 (new_n3512_, not_new_n1537__6782230728490, not_pi122_0);
  or g_7094 (new_n8957_, not_new_n9024_, not_new_n9036_);
  or g_7095 (new_n2540_, not_new_n608__2, not_new_n1013__0);
  not g_7096 (not_new_n4018_, new_n4018_);
  and g_7097 (new_n8812_, new_n9150_, new_n9153_);
  not g_7098 (not_new_n5763__0, new_n5763_);
  not g_7099 (not_new_n4835__0, new_n4835_);
  not g_7100 (not_new_n634__19773267430, new_n634_);
  or g_7101 (new_n2183_, not_new_n591__19773267430, not_new_n4781_);
  not g_7102 (not_new_n9718_, new_n9718_);
  not g_7103 (not_new_n6125_, new_n6125_);
  or g_7104 (new_n7911_, not_new_n7829_, not_new_n7827__0);
  or g_7105 (new_n3418_, not_new_n1008__1, not_new_n1594__2);
  not g_7106 (new_n5102_, new_n4945_);
  and g_7107 (new_n1343_, and_new_n2335__new_n2336_, new_n2337_);
  or g_7108 (new_n2471_, not_new_n597__138412872010, not_new_n4776__0);
  not g_7109 (new_n8550_, new_n8234_);
  not g_7110 (not_new_n7199_, new_n7199_);
  not g_7111 (new_n5519_, new_n5431_);
  or g_7112 (po204, not_new_n1392_, or_or_not_new_n1561__not_new_n2464__not_new_n1391_);
  not g_7113 (not_new_n4747_, new_n4747_);
  not g_7114 (not_new_n661_, new_n661_);
  and g_7115 (new_n4907_, new_n5156_, new_n4902_);
  or g_7116 (new_n10063_, new_n1045_, new_n635_);
  not g_7117 (not_new_n3291_, new_n3291_);
  not g_7118 (new_n5784_, new_n1067_);
  not g_7119 (not_new_n5431_, new_n5431_);
  not g_7120 (not_new_n6376_, new_n6376_);
  not g_7121 (not_new_n3185__490, new_n3185_);
  not g_7122 (not_new_n9326__2, new_n9326_);
  or g_7123 (new_n5296_, not_new_n5113__0, not_new_n5294_);
  or g_7124 (new_n2586_, or_not_new_n2585__not_new_n2584_, not_new_n2583_);
  not g_7125 (not_new_n9232_, new_n9232_);
  or g_7126 (new_n9595_, new_n1067_, new_n633_);
  and g_7127 (new_n4913_, new_n5246_, new_n5243_);
  not g_7128 (not_new_n6759_, new_n6759_);
  not g_7129 (not_new_n4591_, new_n4591_);
  or g_7130 (new_n7372_, not_new_n7019__1, not_new_n6975__1);
  not g_7131 (not_new_n585__8235430, new_n585_);
  not g_7132 (not_new_n599__3430, new_n599_);
  not g_7133 (not_new_n9734_, new_n9734_);
  not g_7134 (not_new_n3676_, new_n3676_);
  or g_7135 (new_n7854_, not_new_n7576_, not_new_n7853_);
  not g_7136 (not_pi204, pi204);
  not g_7137 (not_new_n5838_, new_n5838_);
  not g_7138 (not_new_n6518_, new_n6518_);
  or g_7139 (new_n7771_, not_new_n1598__1176490, not_new_n7661_);
  and g_7140 (new_n8814_, new_n9134_, new_n9137_);
  and g_7141 (and_new_n4928__new_n5310_, new_n5310_, new_n4928_);
  not g_7142 (not_new_n641__2, new_n641_);
  or g_7143 (new_n6923_, not_new_n6536__0, not_new_n646__403536070);
  or g_7144 (new_n683_, not_new_n1496_, not_new_n3017_);
  not g_7145 (not_new_n637__24010, new_n637_);
  not g_7146 (new_n5536_, new_n5500_);
  not g_7147 (not_new_n7616_, new_n7616_);
  not g_7148 (not_new_n1581__47475615099430, new_n1581_);
  or g_7149 (new_n2635_, not_new_n605__490, not_new_n5479_);
  not g_7150 (not_new_n2223_, new_n2223_);
  or g_7151 (new_n7723_, not_new_n8023_, not_new_n8024_);
  not g_7152 (not_new_n10296_, new_n10296_);
  or g_7153 (new_n2618_, not_new_n4454__0, not_new_n610__10);
  or g_7154 (new_n6713_, not_new_n644__2824752490, not_new_n6522_);
  and g_7155 (and_and_new_n1731__new_n1732__new_n1734_, new_n1734_, and_new_n1731__new_n1732_);
  not g_7156 (not_new_n695_, new_n695_);
  not g_7157 (not_new_n3234_, new_n3234_);
  not g_7158 (not_new_n6931_, new_n6931_);
  not g_7159 (not_new_n1612__6, new_n1612_);
  or g_7160 (new_n3787_, not_new_n2038_, not_new_n3479_);
  or g_7161 (new_n6788_, not_new_n6787_, not_new_n6712_);
  not g_7162 (new_n9938_, new_n1600_);
  or g_7163 (new_n8714_, not_new_n8707_, or_not_new_n8713__not_new_n8715_);
  not g_7164 (not_pi164_3, pi164);
  not g_7165 (new_n4839_, new_n4745_);
  not g_7166 (not_new_n5462__1, new_n5462_);
  or g_7167 (new_n1903_, not_new_n588__7, not_pi105);
  not g_7168 (not_new_n1057__7, new_n1057_);
  not g_7169 (not_new_n7010__1, new_n7010_);
  or g_7170 (new_n4369_, not_new_n4306_, not_new_n4366_);
  not g_7171 (not_new_n1020_, new_n1020_);
  not g_7172 (not_new_n6961_, new_n6961_);
  not g_7173 (not_new_n5197_, new_n5197_);
  not g_7174 (not_new_n2729_, new_n2729_);
  or g_7175 (new_n10105_, new_n643_, new_n1061_);
  not g_7176 (new_n5551_, new_n5452_);
  not g_7177 (not_new_n3310__3430, new_n3310_);
  and g_7178 (new_n1541_, new_n3594_, new_n3595_);
  not g_7179 (not_new_n4495_, new_n4495_);
  not g_7180 (not_new_n7619__0, new_n7619_);
  not g_7181 (not_new_n4995_, new_n4995_);
  not g_7182 (not_new_n4513_, new_n4513_);
  not g_7183 (not_new_n5951_, new_n5951_);
  or g_7184 (new_n4678_, not_new_n4677_, not_new_n4676_);
  or g_7185 (new_n5299_, not_new_n5297_, not_new_n5298_);
  not g_7186 (not_new_n2798_, new_n2798_);
  and g_7187 (new_n9472_, new_n9419_, new_n9626_);
  not g_7188 (not_new_n9629_, new_n9629_);
  or g_7189 (new_n8486_, not_new_n628__16284135979104490, not_new_n8117__1);
  and g_7190 (and_new_n3004__new_n998_, new_n3004_, new_n998_);
  not g_7191 (not_pi166_3, pi166);
  not g_7192 (not_new_n1065__10, new_n1065_);
  not g_7193 (not_new_n628__57648010, new_n628_);
  not g_7194 (new_n9646_, new_n9426_);
  not g_7195 (not_new_n8341_, new_n8341_);
  not g_7196 (not_new_n775__70, new_n775_);
  not g_7197 (not_new_n1252_, new_n1252_);
  xor g_7198 (key_gate_5, key_5, new_n1534_);
  not g_7199 (not_new_n648__403536070, new_n648_);
  or g_7200 (new_n7343_, not_new_n7101_, not_new_n775__2);
  not g_7201 (not_new_n3271_, new_n3271_);
  not g_7202 (not_new_n586__5, new_n586_);
  or g_7203 (new_n931_, or_not_new_n1027__0_not_new_n3384_, not_new_n1023__1);
  and g_7204 (new_n5044_, new_n4991_, new_n5198_);
  not g_7205 (not_new_n1583__7, new_n1583_);
  or g_7206 (new_n7859_, not_new_n629__2824752490, not_new_n7626_);
  not g_7207 (not_new_n8404_, new_n8404_);
  or g_7208 (new_n9550_, not_new_n9520_, not_new_n9524_);
  not g_7209 (not_new_n3372__19773267430, new_n3372_);
  or g_7210 (new_n6397_, not_new_n6291_, not_new_n634__57648010);
  not g_7211 (not_new_n638__1577753820348458066150427430, new_n638_);
  not g_7212 (not_new_n4787_, new_n4787_);
  not g_7213 (not_new_n2666_, new_n2666_);
  not g_7214 (not_new_n1601__70, new_n1601_);
  not g_7215 (not_new_n9420__0, new_n9420_);
  or g_7216 (new_n6934_, not_new_n6933_, not_new_n6932_);
  not g_7217 (not_new_n6521__0, new_n6521_);
  and g_7218 (new_n6233_, new_n6382_, and_and_and_new_n6385__new_n6386__new_n6241__new_n6375_);
  not g_7219 (not_new_n5797_, new_n5797_);
  or g_7220 (or_not_new_n9166__not_new_n9106_, not_new_n9106_, not_new_n9166_);
  not g_7221 (new_n7664_, new_n1596_);
  not g_7222 (not_new_n10166__0, new_n10166_);
  or g_7223 (new_n8536_, not_new_n8390_, not_new_n8262__1);
  or g_7224 (new_n3679_, not_new_n636__9, not_po298_490);
  and g_7225 (new_n4914_, new_n5234_, new_n5237_);
  or g_7226 (new_n3305_, not_new_n1581__113988951853731430, not_new_n8098__0);
  or g_7227 (or_not_new_n4227__not_new_n1608_, not_new_n1608_, not_new_n4227_);
  not g_7228 (not_new_n9913_, new_n9913_);
  and g_7229 (new_n1334_, new_n2290_, new_n2291_);
  not g_7230 (not_new_n1011__7, new_n1011_);
  not g_7231 (not_new_n594__6782230728490, new_n594_);
  and g_7232 (and_new_n2364__new_n2363_, new_n2364_, new_n2363_);
  not g_7233 (not_new_n8614_, new_n8614_);
  and g_7234 (new_n1300_, and_and_new_n2124__new_n2127__new_n2125_, new_n2126_);
  not g_7235 (not_new_n5095__1, new_n5095_);
  or g_7236 (new_n4035_, not_pi055_2, not_new_n3949_);
  not g_7237 (not_new_n925_, new_n925_);
  not g_7238 (not_new_n8756_, new_n8756_);
  not g_7239 (not_new_n8170__2, new_n8170_);
  or g_7240 (new_n9785_, not_new_n1601__39098210485829880490, not_new_n9415_);
  or g_7241 (new_n1947_, not_new_n9431_, not_new_n1584__8);
  or g_7242 (or_or_or_not_new_n6239__not_new_n6350__not_new_n6232__3_not_new_n6317__0, not_new_n6317__0, or_or_not_new_n6239__not_new_n6350__not_new_n6232__3);
  not g_7243 (not_new_n7754__4, new_n7754_);
  not g_7244 (not_new_n4432__0, new_n4432_);
  or g_7245 (or_not_new_n1028__8_not_new_n1622__1, not_new_n1028__8, not_new_n1622__1);
  and g_7246 (new_n6586_, new_n6653_, new_n6744_);
  or g_7247 (or_not_new_n1551__not_new_n1372_, not_new_n1551_, not_new_n1372_);
  not g_7248 (not_new_n7664__1, new_n7664_);
  or g_7249 (new_n6717_, not_new_n6657_, not_new_n6448_);
  not g_7250 (not_new_n6738_, new_n6738_);
  not g_7251 (not_new_n7838_, new_n7838_);
  not g_7252 (not_new_n2093_, new_n2093_);
  not g_7253 (not_new_n6501_, new_n6501_);
  or g_7254 (new_n9263_, not_new_n8855_, not_new_n625__5585458640832840070);
  not g_7255 (not_new_n1536__7, new_n1536_);
  not g_7256 (not_new_n646__3430, new_n646_);
  not g_7257 (not_new_n1589__168070, new_n1589_);
  not g_7258 (not_new_n4537_, new_n4537_);
  not g_7259 (not_new_n9375_, new_n9375_);
  not g_7260 (not_new_n6612_, new_n6612_);
  or g_7261 (new_n5143_, new_n1051_, new_n647_);
  not g_7262 (not_new_n587__6782230728490, new_n587_);
  not g_7263 (not_new_n8961_, new_n8961_);
  not g_7264 (not_new_n1583__2, new_n1583_);
  and g_7265 (new_n5862_, new_n625_, new_n5774_);
  not g_7266 (not_new_n9247_, new_n9247_);
  not g_7267 (not_new_n581__5, new_n581_);
  not g_7268 (not_new_n643__490, new_n643_);
  not g_7269 (not_new_n994__7, new_n994_);
  or g_7270 (new_n9100_, new_n621_, new_n1598_);
  not g_7271 (not_new_n4075_, new_n4075_);
  not g_7272 (not_pi031, pi031);
  not g_7273 (not_new_n1017__6, new_n1017_);
  and g_7274 (new_n8597_, new_n8794_, new_n8717_);
  or g_7275 (new_n4395_, not_new_n4281_, not_new_n652_);
  or g_7276 (new_n9281_, not_new_n9279_, not_new_n9280_);
  not g_7277 (not_new_n1055__968890104070, new_n1055_);
  and g_7278 (and_and_new_n1915__new_n1918__new_n1916_, and_new_n1915__new_n1918_, new_n1916_);
  or g_7279 (new_n648_, not_new_n1903_, or_or_not_new_n1901__not_new_n1902__not_new_n1904_);
  not g_7280 (not_new_n4023_, new_n4023_);
  or g_7281 (new_n6008_, not_new_n6007_, not_new_n5891_);
  and g_7282 (new_n1558_, new_n3629_, new_n3628_);
  or g_7283 (new_n1016_, not_new_n3353_, not_new_n3354_);
  or g_7284 (new_n6205_, not_new_n6074_, not_new_n5904_);
  or g_7285 (new_n6832_, not_new_n6474__1, not_new_n1049__168070);
  or g_7286 (new_n2376_, not_new_n4725__0, not_new_n597__3);
  not g_7287 (not_new_n4832_, new_n4832_);
  not g_7288 (not_new_n7400_, new_n7400_);
  not g_7289 (not_new_n1065__332329305696010, new_n1065_);
  or g_7290 (new_n5627_, not_new_n5501_, not_new_n5502__0);
  not g_7291 (not_new_n7009__1, new_n7009_);
  or g_7292 (new_n1063_, not_new_n3477_, not_new_n3478_);
  not g_7293 (not_new_n4357_, new_n4357_);
  not g_7294 (not_new_n631_, new_n631_);
  or g_7295 (new_n3635_, not_new_n1611__19773267430, not_new_n968_);
  not g_7296 (not_new_n588__332329305696010, new_n588_);
  not g_7297 (not_new_n1800_, new_n1800_);
  not g_7298 (not_new_n3567_, new_n3567_);
  and g_7299 (new_n1448_, new_n2660_, and_new_n2662__new_n2661_);
  not g_7300 (not_new_n637__0, new_n637_);
  not g_7301 (not_new_n2907_, new_n2907_);
  not g_7302 (not_new_n9753_, new_n9753_);
  or g_7303 (new_n7279_, not_new_n7015_, not_new_n7278_);
  and g_7304 (new_n1471_, new_n2715_, new_n2713_);
  not g_7305 (not_pi263_0, pi263);
  and g_7306 (new_n1319_, new_n2216_, and_new_n1318__new_n2217_);
  not g_7307 (new_n9513_, new_n9394_);
  not g_7308 (not_new_n4005_, new_n4005_);
  not g_7309 (not_new_n4093_, new_n4093_);
  not g_7310 (not_new_n3421_, new_n3421_);
  and g_7311 (new_n8944_, new_n9098_, new_n8891_);
  or g_7312 (or_not_new_n2300__not_new_n2301_, not_new_n2300_, not_new_n2301_);
  not g_7313 (not_new_n10033_, new_n10033_);
  or g_7314 (new_n2851_, not_pi259_0, not_po296_43181145673964365640352930977077280875522488490);
  or g_7315 (new_n6609_, not_new_n6949_, not_new_n6948_);
  not g_7316 (not_new_n613__1, new_n613_);
  not g_7317 (not_new_n4814_, new_n4814_);
  or g_7318 (new_n9322_, not_new_n626__93874803376477543056490, not_new_n8860_);
  not g_7319 (not_new_n7733_, new_n7733_);
  not g_7320 (not_new_n10143_, new_n10143_);
  or g_7321 (new_n2029_, not_new_n9868_, not_new_n594__490);
  or g_7322 (new_n7113_, not_new_n7326_, not_new_n7310_);
  not g_7323 (not_new_n7407_, new_n7407_);
  or g_7324 (or_not_new_n3149__not_new_n3148_, not_new_n3149_, not_new_n3148_);
  not g_7325 (new_n6524_, new_n627_);
  not g_7326 (not_new_n5258_, new_n5258_);
  or g_7327 (new_n7858_, not_new_n1600__1176490, not_new_n7625_);
  not g_7328 (not_new_n1057__8, new_n1057_);
  not g_7329 (new_n6064_, new_n5811_);
  not g_7330 (not_new_n1027__19773267430, new_n1027_);
  or g_7331 (new_n1889_, not_new_n1585__5, not_new_n5735_);
  and g_7332 (new_n4803_, new_n4890_, new_n4891_);
  not g_7333 (not_pi060, pi060);
  not g_7334 (new_n5776_, new_n1603_);
  not g_7335 (not_new_n9355_, new_n9355_);
  not g_7336 (new_n4993_, new_n1596_);
  not g_7337 (not_new_n2509__3, new_n2509_);
  not g_7338 (not_new_n7666__0, new_n7666_);
  not g_7339 (not_new_n984__6782230728490, new_n984_);
  not g_7340 (not_new_n3445_, new_n3445_);
  or g_7341 (new_n8426_, not_new_n8371_, not_new_n8174_);
  not g_7342 (not_new_n9736_, new_n9736_);
  not g_7343 (not_new_n1067__968890104070, new_n1067_);
  or g_7344 (new_n2743_, not_new_n595__0, not_new_n6971_);
  not g_7345 (not_new_n1454_, new_n1454_);
  not g_7346 (not_new_n1528_, new_n1528_);
  not g_7347 (not_new_n1037__2, new_n1037_);
  not g_7348 (not_new_n6451__0, new_n6451_);
  not g_7349 (not_po296_9, po296);
  not g_7350 (not_new_n1285_, new_n1285_);
  not g_7351 (not_new_n6508_, new_n6508_);
  not g_7352 (not_new_n4508_, new_n4508_);
  not g_7353 (not_new_n2218_, new_n2218_);
  not g_7354 (not_new_n1600__57648010, new_n1600_);
  or g_7355 (new_n7175_, not_new_n7158_, not_new_n742_);
  or g_7356 (new_n3248_, not_new_n3184__0, not_new_n648__8);
  not g_7357 (not_new_n7345_, new_n7345_);
  or g_7358 (or_not_new_n7311__not_new_n7203_, not_new_n7311_, not_new_n7203_);
  not g_7359 (not_new_n5473_, new_n5473_);
  or g_7360 (new_n5349_, not_new_n5259_, not_new_n4994__0);
  and g_7361 (new_n7728_, new_n7574_, new_n7892_);
  not g_7362 (not_new_n7063_, new_n7063_);
  not g_7363 (not_new_n7075_, new_n7075_);
  not g_7364 (not_new_n6522_, new_n6522_);
  not g_7365 (not_new_n7017_, new_n7017_);
  not g_7366 (new_n4926_, new_n624_);
  and g_7367 (new_n8209_, new_n8474_, new_n8286_);
  not g_7368 (not_pi062_2, pi062);
  not g_7369 (new_n9697_, new_n9367_);
  not g_7370 (new_n4924_, new_n628_);
  not g_7371 (not_new_n3249_, new_n3249_);
  not g_7372 (not_new_n4803_, new_n4803_);
  or g_7373 (new_n3869_, not_new_n646__70, not_new_n6443__2824752490);
  or g_7374 (new_n2792_, not_new_n4134__1, not_new_n994__8);
  not g_7375 (not_new_n4978_, new_n4978_);
  not g_7376 (new_n10235_, new_n10020_);
  and g_7377 (new_n9334_, new_n9329_, new_n9539_);
  not g_7378 (new_n7613_, new_n624_);
  not g_7379 (not_new_n8631_, new_n8631_);
  not g_7380 (not_new_n3534_, new_n3534_);
  or g_7381 (new_n3106_, not_new_n928__6, not_new_n1606__2);
  not g_7382 (not_new_n2585_, new_n2585_);
  not g_7383 (not_new_n1616__19773267430, new_n1616_);
  not g_7384 (not_new_n4642_, new_n4642_);
  or g_7385 (new_n9778_, not_new_n9637__0, not_new_n9776_);
  or g_7386 (new_n2556_, not_new_n2553_, or_not_new_n2555__not_new_n2554_);
  not g_7387 (not_new_n617__0, new_n617_);
  not g_7388 (not_new_n6995_, new_n6995_);
  and g_7389 (new_n4307_, new_n4370_, new_n4371_);
  not g_7390 (not_new_n581__77309937197074445241370944070, new_n581_);
  not g_7391 (not_new_n2343_, new_n2343_);
  or g_7392 (new_n1934_, not_new_n9956_, not_new_n594__7);
  not g_7393 (not_new_n1581__3, new_n1581_);
  not g_7394 (not_new_n4213_, new_n4213_);
  and g_7395 (new_n9479_, new_n9331_, new_n9664_);
  not g_7396 (not_new_n4734_, new_n4734_);
  not g_7397 (not_new_n8840_, new_n8840_);
  not g_7398 (not_new_n9160_, new_n9160_);
  or g_7399 (new_n7812_, not_new_n7811_, not_new_n7703_);
  or g_7400 (or_not_new_n2836__not_new_n2835_, not_new_n2836_, not_new_n2835_);
  not g_7401 (not_new_n603__6782230728490, new_n603_);
  not g_7402 (not_new_n4960_, new_n4960_);
  and g_7403 (new_n1283_, and_new_n1282__new_n2046_, new_n2045_);
  not g_7404 (not_new_n641__8235430, new_n641_);
  not g_7405 (not_new_n1599__9, new_n1599_);
  not g_7406 (not_new_n8398_, new_n8398_);
  or g_7407 (new_n7058_, not_new_n7491_, not_new_n7490_);
  not g_7408 (not_new_n4478_, new_n4478_);
  or g_7409 (new_n2368_, not_new_n600__2, not_new_n4071__0);
  or g_7410 (or_or_or_not_new_n6240__not_new_n6330__not_new_n6331__not_new_n6242__1, or_or_not_new_n6240__not_new_n6330__not_new_n6331_, not_new_n6242__1);
  not g_7411 (not_pi068, pi068);
  not g_7412 (not_new_n1047__1176490, new_n1047_);
  not g_7413 (not_new_n3971_, new_n3971_);
  or g_7414 (new_n4790_, not_new_n4792__0, not_new_n4831__0);
  not g_7415 (not_new_n10013__0, new_n10013_);
  not g_7416 (not_new_n1015__5, new_n1015_);
  or g_7417 (new_n1766_, not_new_n585_, not_pi265);
  not g_7418 (not_new_n1055__8235430, new_n1055_);
  not g_7419 (not_new_n646__47475615099430, new_n646_);
  not g_7420 (not_new_n6237_, new_n6237_);
  and g_7421 (and_new_n4323__new_n4324_, new_n4323_, new_n4324_);
  not g_7422 (not_new_n609_, new_n609_);
  not g_7423 (not_new_n9021_, new_n9021_);
  not g_7424 (not_new_n8289_, new_n8289_);
  or g_7425 (new_n8236_, not_new_n8559_, not_new_n8558_);
  not g_7426 (not_new_n5472_, new_n5472_);
  not g_7427 (not_new_n7566_, new_n7566_);
  or g_7428 (new_n9121_, not_new_n9119__0, not_new_n9082__0);
  or g_7429 (new_n3636_, not_new_n984__138412872010, not_pi184_0);
  not g_7430 (not_new_n626__6, new_n626_);
  not g_7431 (not_new_n8305_, new_n8305_);
  not g_7432 (new_n7800_, new_n7735_);
  or g_7433 (po261, not_new_n3709_, not_new_n3708_);
  and g_7434 (and_new_n8750__new_n8736_, new_n8750_, new_n8736_);
  not g_7435 (not_new_n1173_, new_n1173_);
  not g_7436 (not_new_n1043__70, new_n1043_);
  not g_7437 (new_n6269_, new_n643_);
  or g_7438 (new_n2253_, not_new_n6550_, not_new_n1580__47475615099430);
  not g_7439 (not_po296_8, po296);
  not g_7440 (not_new_n5616_, new_n5616_);
  or g_7441 (or_or_not_new_n1267__not_new_n1265__not_new_n1964_, or_not_new_n1267__not_new_n1265_, not_new_n1964_);
  or g_7442 (new_n10253_, not_new_n631__225393402906922580878632490, not_new_n9889__0);
  not g_7443 (not_new_n4199_, new_n4199_);
  and g_7444 (new_n5045_, and_new_n5084__new_n5345_, new_n5344_);
  not g_7445 (not_new_n1037__10, new_n1037_);
  or g_7446 (new_n7316_, not_new_n7180_, not_new_n6961_);
  not g_7447 (new_n6477_, new_n1041_);
  or g_7448 (new_n2227_, not_new_n4122_, not_new_n585__6782230728490);
  not g_7449 (not_new_n4014__1, new_n4014_);
  not g_7450 (not_new_n599__0, new_n599_);
  not g_7451 (not_new_n622__403536070, new_n622_);
  and g_7452 (new_n7088_, and_new_n7161__new_n7474_, new_n7473_);
  or g_7453 (new_n7249_, not_new_n7009_, not_new_n7448_);
  not g_7454 (not_new_n1598__2824752490, new_n1598_);
  or g_7455 (new_n6834_, not_new_n1049__1176490, not_new_n6474__2);
  or g_7456 (new_n3651_, not_new_n1615_, not_new_n1611__113988951853731430);
  and g_7457 (new_n10001_, new_n9859_, new_n10180_);
  not g_7458 (not_new_n1028__6, new_n1028_);
  not g_7459 (new_n9037_, new_n8957_);
  or g_7460 (or_not_new_n8995__1_not_new_n8799__1, not_new_n8799__1, not_new_n8995__1);
  not g_7461 (not_new_n619__5, new_n619_);
  not g_7462 (not_new_n4244_, new_n4244_);
  not g_7463 (not_new_n4542_, new_n4542_);
  and g_7464 (new_n6458_, new_n6730_, new_n6728_);
  not g_7465 (not_new_n599__8235430, new_n599_);
  or g_7466 (new_n1813_, not_new_n1585__1, not_new_n5830_);
  or g_7467 (new_n9760_, not_new_n618__93874803376477543056490, not_new_n9421__0);
  not g_7468 (not_new_n5639_, new_n5639_);
  and g_7469 (new_n3963_, not_pi047_1, and_and_and_not_pi051_1_not_pi050_1_not_pi049_1_not_pi048_1);
  not g_7470 (new_n6816_, new_n6641_);
  or g_7471 (or_not_new_n2769__not_new_n1476_, not_new_n2769_, not_new_n1476_);
  or g_7472 (new_n10072_, not_new_n1039__5585458640832840070, not_new_n628__13410686196639649008070);
  not g_7473 (not_new_n1071__6, new_n1071_);
  not g_7474 (not_new_n10344_, new_n10344_);
  not g_7475 (not_new_n581__2, new_n581_);
  not g_7476 (not_pi137_2, pi137);
  or g_7477 (new_n3884_, not_new_n1576__2326305139872070, not_new_n627__490);
  or g_7478 (new_n2999_, not_new_n581__3, not_new_n1045__2);
  or g_7479 (or_not_new_n4827__not_new_n4799_, not_new_n4827_, not_new_n4799_);
  not g_7480 (not_new_n7631__1, new_n7631_);
  or g_7481 (new_n6754_, not_new_n6631_, not_new_n6737_);
  not g_7482 (not_new_n10297_, new_n10297_);
  and g_7483 (and_new_n6440__new_n6441_, new_n6441_, new_n6440_);
  not g_7484 (not_new_n1940_, new_n1940_);
  or g_7485 (new_n8244_, not_new_n8205_, not_new_n8415_);
  not g_7486 (not_new_n1047__10, new_n1047_);
  or g_7487 (new_n3187_, not_new_n647__7, not_new_n589_);
  not g_7488 (not_new_n5232_, new_n5232_);
  not g_7489 (not_new_n994__797922662976120010, new_n994_);
  not g_7490 (not_new_n7523_, new_n7523_);
  not g_7491 (not_new_n1534__19773267430, key_gate_5);
  or g_7492 (new_n3350_, not_new_n3919__0, not_pi064_1176490);
  not g_7493 (not_new_n5517_, new_n5517_);
  not g_7494 (not_new_n6587_, new_n6587_);
  not g_7495 (not_new_n620__1, new_n620_);
  not g_7496 (not_new_n629__3430, new_n629_);
  not g_7497 (not_new_n4399_, new_n4399_);
  not g_7498 (not_new_n1596__3430, new_n1596_);
  not g_7499 (not_new_n4678_, new_n4678_);
  not g_7500 (not_new_n3310__8235430, new_n3310_);
  not g_7501 (not_new_n1613__3, new_n1613_);
  not g_7502 (not_new_n9294_, new_n9294_);
  not g_7503 (new_n6177_, new_n5867_);
  or g_7504 (new_n1804_, not_new_n1588__1, not_new_n1035_);
  not g_7505 (not_new_n9273_, new_n9273_);
  or g_7506 (new_n4386_, not_new_n4275_, not_new_n687_);
  or g_7507 (or_or_or_not_new_n2785__not_new_n2788__not_new_n2787__not_new_n2789_, or_or_not_new_n2785__not_new_n2788__not_new_n2787_, not_new_n2789_);
  not g_7508 (not_new_n6605_, new_n6605_);
  not g_7509 (not_new_n3051_, new_n3051_);
  not g_7510 (not_new_n5899__2, new_n5899_);
  and g_7511 (and_and_new_n6388__new_n6313__new_n6224_, and_new_n6388__new_n6313_, new_n6224_);
  not g_7512 (not_new_n2249_, new_n2249_);
  or g_7513 (new_n7233_, not_new_n7036_, not_new_n727_);
  or g_7514 (new_n2428_, not_new_n4132__0, not_new_n600__24010);
  not g_7515 (not_new_n3922_, new_n3922_);
  not g_7516 (not_new_n8494_, new_n8494_);
  or g_7517 (new_n5731_, not_new_n6026_, not_new_n6029_);
  or g_7518 (or_or_not_new_n2053__not_new_n2054__not_new_n2056_, or_not_new_n2053__not_new_n2054_, not_new_n2056_);
  not g_7519 (not_new_n8167__0, new_n8167_);
  not g_7520 (new_n4164_, new_n4149_);
  not g_7521 (not_new_n639__6, new_n639_);
  not g_7522 (not_new_n1031__3, new_n1031_);
  or g_7523 (new_n10200_, not_new_n10066_, not_new_n9879__0);
  not g_7524 (not_new_n6547__0, new_n6547_);
  and g_7525 (and_new_n2632__new_n2631_, new_n2631_, new_n2632_);
  not g_7526 (not_new_n4255_, new_n4255_);
  not g_7527 (not_new_n6370__0, new_n6370_);
  not g_7528 (not_new_n2097_, new_n2097_);
  not g_7529 (not_new_n8006_, new_n8006_);
  or g_7530 (new_n3015_, not_new_n1157_, not_new_n1027__70);
  not g_7531 (new_n9407_, new_n1603_);
  not g_7532 (not_new_n629__6782230728490, new_n629_);
  not g_7533 (not_new_n9427_, new_n9427_);
  not g_7534 (not_new_n8129__1, new_n8129_);
  or g_7535 (new_n1719_, not_po296_16284135979104490, not_pi003_0);
  or g_7536 (new_n2566_, not_new_n2563_, or_not_new_n2565__not_new_n2564_);
  not g_7537 (not_pi148_2, pi148);
  or g_7538 (new_n6408_, new_n1031_, new_n714_);
  or g_7539 (new_n4382_, not_new_n4270_, not_new_n657_);
  or g_7540 (new_n7337_, not_new_n7334__0, not_new_n736__2);
  not g_7541 (not_new_n631__0, new_n631_);
  or g_7542 (new_n8859_, not_new_n1049__6782230728490, not_new_n648__16284135979104490);
  or g_7543 (new_n7910_, not_new_n7794_, not_new_n7578_);
  not g_7544 (not_new_n6741_, new_n6741_);
  not g_7545 (not_new_n8060_, new_n8060_);
  not g_7546 (not_pi213, pi213);
  not g_7547 (not_pi050_0, pi050);
  and g_7548 (and_new_n1575__new_n938_, new_n1575_, new_n938_);
  not g_7549 (not_new_n4837_, new_n4837_);
  not g_7550 (not_new_n4497_, new_n4497_);
  not g_7551 (not_new_n9855_, new_n9855_);
  not g_7552 (not_new_n7795_, new_n7795_);
  and g_7553 (new_n5847_, new_n6119_, new_n5919_);
  not g_7554 (not_new_n9449_, new_n9449_);
  or g_7555 (or_or_not_new_n4234__not_new_n4336__not_new_n675_, or_not_new_n4234__not_new_n4336_, not_new_n675_);
  not g_7556 (not_new_n4899__1, new_n4899_);
  not g_7557 (new_n1576_, new_n6443_);
  or g_7558 (new_n1817_, not_new_n1591__1, not_new_n8818_);
  not g_7559 (not_new_n9349_, new_n9349_);
  or g_7560 (new_n6369_, not_new_n6368_, not_new_n6309_);
  not g_7561 (not_new_n8922_, new_n8922_);
  not g_7562 (not_new_n7246_, new_n7246_);
  not g_7563 (not_new_n7805_, new_n7805_);
  not g_7564 (not_new_n4428__0, new_n4428_);
  or g_7565 (new_n6077_, not_new_n5919__0, not_new_n5763__0);
  not g_7566 (not_new_n1057__6782230728490, new_n1057_);
  or g_7567 (new_n6422_, not_new_n6332_, not_new_n6333_);
  not g_7568 (not_new_n3262_, new_n3262_);
  not g_7569 (not_new_n3339_, new_n3339_);
  not g_7570 (not_new_n2879_, new_n2879_);
  not g_7571 (not_new_n589__8, new_n589_);
  or g_7572 (new_n6110_, not_new_n5956__0, not_new_n5880_);
  not g_7573 (not_new_n8237_, new_n8237_);
  or g_7574 (new_n8379_, not_new_n617__332329305696010, not_new_n8278_);
  or g_7575 (new_n3887_, not_new_n6443__113988951853731430, not_new_n642__10);
  not g_7576 (not_new_n5942_, new_n5942_);
  or g_7577 (new_n7404_, not_new_n775__10, not_new_n7116_);
  not g_7578 (new_n2095_, new_n646_);
  or g_7579 (new_n6384_, not_new_n6286_, not_new_n638__2824752490);
  and g_7580 (new_n8591_, and_and_new_n8724__new_n8726__new_n8728_, new_n8727_);
  not g_7581 (not_new_n4262_, new_n4262_);
  or g_7582 (new_n9230_, not_new_n618__5585458640832840070, not_new_n8893_);
  not g_7583 (not_new_n4643_, new_n4643_);
  not g_7584 (not_new_n5166__0, new_n5166_);
  and g_7585 (and_not_pi034_1_not_pi033_3, not_pi033_3, not_pi034_1);
  and g_7586 (new_n8598_, new_n8703_, new_n8783_);
  not g_7587 (not_new_n8433_, new_n8433_);
  or g_7588 (new_n2310_, not_new_n6549_, not_new_n1580__16284135979104490);
  or g_7589 (new_n7654_, not_new_n7828_, not_new_n7911_);
  not g_7590 (not_new_n4505_, new_n4505_);
  not g_7591 (not_new_n9638_, new_n9638_);
  not g_7592 (not_new_n10223_, new_n10223_);
  not g_7593 (not_new_n1177_, new_n1177_);
  not g_7594 (not_new_n1616__8235430, new_n1616_);
  or g_7595 (new_n4547_, not_new_n4508_, not_new_n4546_);
  not g_7596 (not_new_n7689_, new_n7689_);
  or g_7597 (new_n1745_, not_new_n1728__3430, not_pi089);
  or g_7598 (new_n7869_, not_new_n618__968890104070, not_new_n7664_);
  not g_7599 (not_new_n586__2326305139872070, new_n586_);
  not g_7600 (not_new_n6640_, new_n6640_);
  not g_7601 (not_new_n3494_, new_n3494_);
  or g_7602 (or_or_not_new_n6318__not_new_n6373__0_not_new_n6319_, not_new_n6319_, or_not_new_n6318__not_new_n6373__0);
  not g_7603 (not_new_n1037__2824752490, new_n1037_);
  not g_7604 (not_new_n989__10, new_n989_);
  or g_7605 (new_n9816_, not_new_n9814_, not_new_n9602_);
  not g_7606 (not_new_n9394__0, new_n9394_);
  not g_7607 (not_pi252, pi252);
  not g_7608 (new_n7633_, new_n1603_);
  and g_7609 (new_n3990_, new_n4061_, new_n4062_);
  not g_7610 (not_new_n3357_, new_n3357_);
  not g_7611 (new_n1608_, new_n990_);
  not g_7612 (not_new_n4639_, new_n4639_);
  or g_7613 (new_n3989_, not_new_n4033_, not_new_n3950_);
  not g_7614 (not_new_n2915_, new_n2915_);
  or g_7615 (new_n9651_, new_n645_, new_n1071_);
  not g_7616 (not_new_n620_, new_n620_);
  or g_7617 (new_n3317_, not_pi064_1, not_new_n3987__0);
  not g_7618 (not_new_n3547_, new_n3547_);
  not g_7619 (not_new_n1006__3, new_n1006_);
  not g_7620 (not_new_n1613__10, new_n1613_);
  or g_7621 (new_n5276_, not_new_n5078__2, not_new_n5037_);
  and g_7622 (po101, key_gate_101, pi080);
  or g_7623 (or_not_new_n5426__not_new_n605_, not_new_n5426_, not_new_n605_);
  not g_7624 (not_new_n8444_, new_n8444_);
  not g_7625 (not_pi186_0, pi186);
  not g_7626 (not_new_n3185__6, new_n3185_);
  not g_7627 (not_new_n7027_, new_n7027_);
  not g_7628 (not_new_n637__138412872010, new_n637_);
  or g_7629 (new_n6772_, not_new_n6812_, not_new_n6771_);
  not g_7630 (not_new_n7744__0, new_n7744_);
  not g_7631 (not_new_n3509_, new_n3509_);
  or g_7632 (new_n2410_, not_new_n1055__0, not_new_n598__10);
  not g_7633 (not_new_n662_, new_n662_);
  not g_7634 (not_new_n9647_, new_n9647_);
  not g_7635 (not_po298_490, po298);
  or g_7636 (new_n5931_, not_new_n5753_, not_new_n5930_);
  not g_7637 (not_new_n1059__1, new_n1059_);
  not g_7638 (not_new_n598__24010, new_n598_);
  or g_7639 (new_n3481_, not_new_n2071_, not_new_n1613__24010);
  not g_7640 (new_n5178_, new_n4974_);
  or g_7641 (new_n8267_, not_new_n8420_, not_new_n8214_);
  or g_7642 (new_n8008_, not_new_n629__19773267430, not_new_n7626__0);
  or g_7643 (new_n8973_, not_new_n9170_, not_new_n9073_);
  not g_7644 (not_new_n4624_, new_n4624_);
  or g_7645 (new_n9795_, not_new_n9793_, not_new_n9794_);
  or g_7646 (new_n9276_, not_new_n8897__0, not_new_n1604__968890104070);
  not g_7647 (not_new_n9639_, new_n9639_);
  not g_7648 (not_new_n589__10, new_n589_);
  or g_7649 (new_n8414_, not_new_n8254_, not_new_n8275__0);
  not g_7650 (not_new_n586__6782230728490, new_n586_);
  not g_7651 (not_new_n3124_, new_n3124_);
  not g_7652 (not_new_n1043__3, new_n1043_);
  not g_7653 (not_new_n7627_, new_n7627_);
  or g_7654 (new_n6937_, not_new_n6546__0, not_new_n6769_);
  not g_7655 (not_new_n8145__0, new_n8145_);
  and g_7656 (new_n8949_, new_n8804_, new_n9127_);
  not g_7657 (not_new_n6487__1, new_n6487_);
  not g_7658 (not_new_n1534__113988951853731430, key_gate_5);
  not g_7659 (not_new_n7416_, new_n7416_);
  or g_7660 (new_n5694_, not_new_n5458__0, not_pi141_3);
  or g_7661 (or_not_new_n1596__3430_not_new_n5729_, not_new_n1596__3430, not_new_n5729_);
  or g_7662 (new_n618_, not_new_n2283_, or_or_not_new_n2284__not_new_n2281__not_new_n2282_);
  or g_7663 (po231, not_new_n1453_, not_new_n1452_);
  and g_7664 (and_new_n2029__new_n2032_, new_n2029_, new_n2032_);
  not g_7665 (not_new_n4205_, new_n4205_);
  not g_7666 (new_n10154_, new_n10011_);
  or g_7667 (or_not_new_n2783__not_new_n2782_, not_new_n2783_, not_new_n2782_);
  not g_7668 (new_n7421_, new_n7034_);
  not g_7669 (not_new_n1059__70, new_n1059_);
  not g_7670 (not_new_n1602__9, new_n1602_);
  not g_7671 (not_new_n3134_, new_n3134_);
  or g_7672 (new_n5620_, not_new_n5616_, or_not_new_n5441__not_new_n5617__1);
  not g_7673 (not_new_n1304_, new_n1304_);
  or g_7674 (new_n4409_, or_not_new_n649__0_not_new_n4287_, not_new_n4286__0);
  not g_7675 (not_new_n600__6782230728490, new_n600_);
  not g_7676 (not_new_n9064_, new_n9064_);
  not g_7677 (not_new_n7484_, new_n7484_);
  not g_7678 (not_new_n633__332329305696010, new_n633_);
  not g_7679 (new_n5942_, new_n5761_);
  not g_7680 (not_new_n5508__0, new_n5508_);
  not g_7681 (new_n7775_, new_n7658_);
  not g_7682 (not_new_n1007__5, new_n1007_);
  not g_7683 (not_new_n3354_, new_n3354_);
  or g_7684 (new_n5817_, not_new_n6151_, not_new_n6150_);
  not g_7685 (not_new_n9334_, new_n9334_);
  not g_7686 (not_new_n5021_, new_n5021_);
  not g_7687 (not_new_n3315__19773267430, new_n3315_);
  or g_7688 (new_n9562_, not_new_n9560_, not_new_n9460_);
  not g_7689 (not_pi131, pi131);
  or g_7690 (new_n10170_, new_n645_, new_n1071_);
  not g_7691 (not_new_n625_, new_n625_);
  not g_7692 (not_new_n5029_, new_n5029_);
  not g_7693 (not_new_n3400_, new_n3400_);
  xor g_7694 (key_gate_52, new_n1693_, key_52);
  or g_7695 (new_n3001_, not_new_n3372__7, not_new_n635__4);
  or g_7696 (new_n4219_, not_new_n4151_, not_pi253_1);
  or g_7697 (new_n5797_, not_new_n5975_, not_new_n6046_);
  not g_7698 (not_new_n611__6, new_n611_);
  not g_7699 (not_new_n7354__2, new_n7354_);
  or g_7700 (new_n2063_, not_new_n6567_, not_new_n1580__168070);
  not g_7701 (not_new_n1606__1, new_n1606_);
  or g_7702 (new_n3739_, not_new_n3499_, not_new_n2114_);
  not g_7703 (not_new_n5113_, new_n5113_);
  not g_7704 (not_new_n628__490, new_n628_);
  not g_7705 (not_new_n9462_, new_n9462_);
  not g_7706 (not_new_n6494__0, new_n6494_);
  not g_7707 (not_new_n7121_, new_n7121_);
  or g_7708 (new_n1710_, not_po296_47475615099430, not_pi006_0);
  not g_7709 (not_new_n1603__113988951853731430, new_n1603_);
  not g_7710 (not_new_n1534__47475615099430, key_gate_5);
  not g_7711 (not_new_n4369_, new_n4369_);
  and g_7712 (new_n4793_, new_n4883_, new_n4882_);
  not g_7713 (not_new_n6657_, new_n6657_);
  not g_7714 (not_new_n9281_, new_n9281_);
  not g_7715 (not_new_n4127_, new_n4127_);
  not g_7716 (not_new_n4496__0, new_n4496_);
  not g_7717 (not_new_n593__70, new_n593_);
  not g_7718 (not_new_n9442_, new_n9442_);
  not g_7719 (not_new_n585__3, new_n585_);
  or g_7720 (new_n2629_, not_pi274, not_po296_77309937197074445241370944070);
  not g_7721 (not_new_n9856_, new_n9856_);
  not g_7722 (not_new_n4785_, new_n4785_);
  not g_7723 (not_new_n1537__24010, new_n1537_);
  not g_7724 (not_new_n4971_, new_n4971_);
  not g_7725 (not_new_n6613__2, new_n6613_);
  not g_7726 (not_new_n7430_, new_n7430_);
  and g_7727 (new_n1543_, new_n3598_, new_n3599_);
  not g_7728 (not_new_n3328_, new_n3328_);
  not g_7729 (new_n5562_, new_n5459_);
  and g_7730 (new_n1226_, and_and_new_n1222__new_n1223__new_n1225_, new_n1224_);
  or g_7731 (new_n9596_, new_n637_, new_n1065_);
  or g_7732 (new_n5537_, pi135, new_n1005_);
  not g_7733 (not_new_n9456_, new_n9456_);
  not g_7734 (new_n7928_, new_n7747_);
  or g_7735 (new_n2737_, not_new_n2726_, not_new_n2736_);
  not g_7736 (not_new_n3375_, new_n3375_);
  or g_7737 (new_n7367_, not_new_n7099_, not_new_n7109__1);
  not g_7738 (not_new_n632__19773267430, new_n632_);
  not g_7739 (not_new_n2192_, new_n2192_);
  or g_7740 (new_n3200_, not_new_n1596__4, not_new_n3185__6);
  not g_7741 (not_new_n9175_, new_n9175_);
  or g_7742 (new_n3834_, not_new_n635__490, not_new_n1576__2);
  and g_7743 (new_n5031_, and_new_n4928__new_n5310_, new_n5309_);
  or g_7744 (new_n9782_, not_new_n9494__0, not_new_n9688_);
  or g_7745 (or_not_new_n9191__not_new_n9190_, not_new_n9190_, not_new_n9191_);
  and g_7746 (new_n6236_, new_n6382_, new_n6227_);
  not g_7747 (not_new_n5464_, new_n5464_);
  not g_7748 (new_n9180_, new_n8895_);
  or g_7749 (new_n4870_, not_new_n1602__7, not_new_n4778_);
  not g_7750 (not_new_n7045__0, new_n7045_);
  or g_7751 (new_n6829_, not_new_n6492__0, not_new_n647__403536070);
  not g_7752 (not_new_n5872_, new_n5872_);
  or g_7753 (new_n5248_, new_n1051_, new_n647_);
  or g_7754 (new_n3159_, not_new_n1061__3, not_new_n928__6782230728490);
  not g_7755 (not_new_n1596_, new_n1596_);
  not g_7756 (not_new_n1884_, new_n1884_);
  not g_7757 (not_new_n9094_, new_n9094_);
  or g_7758 (new_n3637_, not_new_n1611__138412872010, not_new_n970_);
  not g_7759 (not_new_n628__1915812313805664144010, new_n628_);
  or g_7760 (new_n8410_, not_new_n8115_, not_new_n641__8235430);
  not g_7761 (not_new_n1027__6782230728490, new_n1027_);
  not g_7762 (new_n7131_, new_n748_);
  or g_7763 (po249, not_new_n3684_, not_new_n3685_);
  or g_7764 (new_n1983_, not_new_n7587_, not_new_n1583__10);
  not g_7765 (not_new_n4774__0, new_n4774_);
  or g_7766 (new_n2400_, not_new_n598__8, not_new_n1051__0);
  or g_7767 (new_n6029_, not_new_n5871_, not_new_n6027_);
  or g_7768 (new_n4519_, not_new_n4518_, not_new_n4485_);
  not g_7769 (new_n4266_, new_n691_);
  not g_7770 (not_new_n1576__797922662976120010, new_n1576_);
  not g_7771 (not_new_n4133_, new_n4133_);
  not g_7772 (not_new_n8045_, new_n8045_);
  not g_7773 (not_new_n7120_, new_n7120_);
  not g_7774 (not_new_n9820_, new_n9820_);
  not g_7775 (not_new_n994__2, new_n994_);
  or g_7776 (new_n5380_, not_new_n1071__9, not_new_n4973_);
  not g_7777 (not_new_n6235__1, new_n6235_);
  not g_7778 (new_n4085_, pi263);
  or g_7779 (new_n1970_, not_new_n1589__9, not_new_n4912_);
  not g_7780 (not_new_n599__4, new_n599_);
  not g_7781 (not_new_n3755_, new_n3755_);
  not g_7782 (not_new_n5783__0, new_n5783_);
  or g_7783 (new_n7971_, not_new_n7942_, not_new_n7738_);
  or g_7784 (or_or_not_new_n1825__not_new_n1826__not_new_n1828_, or_not_new_n1825__not_new_n1826_, not_new_n1828_);
  or g_7785 (new_n2283_, not_pi125, not_new_n588__2326305139872070);
  not g_7786 (not_new_n4195_, new_n4195_);
  not g_7787 (not_new_n5774__1, new_n5774_);
  or g_7788 (new_n6742_, not_new_n1599__490, not_new_n6499_);
  not g_7789 (not_new_n7668_, new_n7668_);
  or g_7790 (new_n9558_, not_new_n9374_, not_new_n9557_);
  not g_7791 (not_new_n3372__13410686196639649008070, new_n3372_);
  and g_7792 (new_n1478_, new_n642_, new_n1616_);
  not g_7793 (not_new_n643__47475615099430, new_n643_);
  or g_7794 (new_n752_, not_new_n3213_, not_new_n3212_);
  not g_7795 (not_new_n624__403536070, new_n624_);
  not g_7796 (not_new_n1053__4, new_n1053_);
  not g_7797 (not_new_n4459__0, new_n4459_);
  not g_7798 (not_new_n611__168070, new_n611_);
  not g_7799 (not_new_n1020__1, new_n1020_);
  or g_7800 (new_n6021_, not_new_n5775_, not_new_n6002_);
  not g_7801 (not_new_n5757__0, new_n5757_);
  or g_7802 (new_n2179_, not_new_n4916_, not_new_n1589__2824752490);
  not g_7803 (new_n4282_, new_n683_);
  not g_7804 (not_new_n8390_, new_n8390_);
  or g_7805 (new_n2669_, not_po296_185621159210175743024531636712070, not_pi269);
  not g_7806 (not_new_n595__24010, new_n595_);
  not g_7807 (not_new_n1170__0, new_n1170_);
  not g_7808 (new_n3469_, new_n1059_);
  or g_7809 (new_n2332_, not_new_n8908_, not_new_n1591__16284135979104490);
  not g_7810 (not_pi148, pi148);
  or g_7811 (new_n2056_, not_new_n585__168070, not_new_n4131_);
  not g_7812 (not_new_n9841_, new_n9841_);
  not g_7813 (new_n6500_, new_n1599_);
  not g_7814 (not_new_n629__6, new_n629_);
  not g_7815 (not_new_n1055__16284135979104490, new_n1055_);
  not g_7816 (not_new_n9997_, new_n9997_);
  not g_7817 (not_new_n9295_, new_n9295_);
  or g_7818 (new_n9222_, not_new_n8822_, not_new_n1037__968890104070);
  not g_7819 (not_new_n9074_, new_n9074_);
  not g_7820 (not_new_n3403_, new_n3403_);
  not g_7821 (not_new_n1055__3, new_n1055_);
  not g_7822 (new_n4095_, pi268);
  not g_7823 (not_new_n8224_, new_n8224_);
  or g_7824 (new_n5933_, not_new_n1045__10, not_new_n5754_);
  not g_7825 (not_new_n646__9, new_n646_);
  or g_7826 (new_n3185_, not_new_n1531_, not_new_n3182__0);
  not g_7827 (new_n3489_, new_n1067_);
  or g_7828 (new_n7067_, not_new_n7551_, not_new_n7552_);
  not g_7829 (not_new_n9206_, new_n9206_);
  not g_7830 (not_new_n9407__0, new_n9407_);
  and g_7831 (new_n609_, new_n2505_, new_n583_);
  not g_7832 (not_new_n984__16284135979104490, new_n984_);
  or g_7833 (new_n3769_, not_new_n1924_, not_new_n3449_);
  or g_7834 (new_n6219_, not_new_n1053__3430, not_new_n5792__0);
  or g_7835 (new_n5291_, not_new_n4950_, not_new_n5084__2);
  and g_7836 (new_n5727_, new_n5995_, new_n5993_);
  not g_7837 (not_new_n8220_, new_n8220_);
  or g_7838 (new_n2738_, not_new_n1588__273687473400809163430, not_new_n1595_);
  not g_7839 (not_new_n1335_, new_n1335_);
  or g_7840 (or_not_new_n4837__not_new_n4772_, not_new_n4772_, not_new_n4837_);
  not g_7841 (not_pi060_0, pi060);
  not g_7842 (not_new_n9627__0, new_n9627_);
  not g_7843 (not_new_n7068_, new_n7068_);
  or g_7844 (new_n2610_, not_new_n1002__0, not_new_n608__9);
  not g_7845 (not_new_n1015__1, new_n1015_);
  not g_7846 (not_new_n1866_, new_n1866_);
  and g_7847 (new_n8078_, new_n8335_, new_n8336_);
  or g_7848 (new_n3081_, not_new_n1179_, not_new_n1027__273687473400809163430);
  not g_7849 (not_new_n625__0, new_n625_);
  not g_7850 (not_new_n1596__3, new_n1596_);
  not g_7851 (not_new_n1600__8235430, new_n1600_);
  and g_7852 (and_new_n9511__new_n9839_, new_n9511_, new_n9839_);
  or g_7853 (new_n3442_, not_new_n1536__19773267430, not_pi024_0);
  not g_7854 (not_new_n1612__24010, new_n1612_);
  not g_7855 (new_n9415_, new_n630_);
  not g_7856 (not_new_n644__2326305139872070, new_n644_);
  not g_7857 (not_new_n2223__0, new_n2223_);
  not g_7858 (not_new_n8172__0, new_n8172_);
  not g_7859 (not_new_n1067__3430, new_n1067_);
  or g_7860 (or_not_new_n2749__not_new_n2752_, not_new_n2752_, not_new_n2749_);
  not g_7861 (not_new_n640__6, new_n640_);
  not g_7862 (not_new_n4724_, new_n4724_);
  not g_7863 (not_new_n4812__0, new_n4812_);
  not g_7864 (not_new_n631__3, new_n631_);
  not g_7865 (new_n8152_, new_n644_);
  not g_7866 (not_new_n8517_, new_n8517_);
  not g_7867 (not_new_n5989_, new_n5989_);
  and g_7868 (new_n4318_, and_new_n4403__new_n4407_, new_n4406_);
  or g_7869 (new_n7365_, not_new_n768_, not_new_n6974__8);
  and g_7870 (new_n1431_, new_n2580_, new_n2582_);
  not g_7871 (not_new_n2226_, new_n2226_);
  or g_7872 (new_n5406_, not_new_n1061__490, not_new_n4970__0);
  or g_7873 (or_or_not_new_n1279__not_new_n1277__not_new_n2021_, not_new_n2021_, or_not_new_n1279__not_new_n1277_);
  or g_7874 (new_n2062_, not_new_n1581__24010, not_new_n8198_);
  or g_7875 (new_n7324_, not_new_n7113__1, not_new_n7072_);
  not g_7876 (not_new_n6892_, new_n6892_);
  not g_7877 (not_new_n2983_, new_n2983_);
  not g_7878 (not_new_n1263_, new_n1263_);
  or g_7879 (new_n9968_, not_new_n10332_, not_new_n10331_);
  or g_7880 (new_n3832_, not_new_n634__490, not_new_n1576__1);
  or g_7881 (new_n2068_, not_new_n593__24010, not_new_n637_);
  or g_7882 (new_n2299_, not_new_n2294_, not_new_n1336_);
  not g_7883 (not_new_n2977_, new_n2977_);
  not g_7884 (not_new_n1011_, new_n1011_);
  and g_7885 (new_n1261_, new_n1946_, new_n1947_);
  not g_7886 (not_new_n8127__1, new_n8127_);
  not g_7887 (new_n5771_, new_n625_);
  or g_7888 (new_n2271_, not_new_n8195_, not_new_n1581__47475615099430);
  not g_7889 (not_new_n5671_, new_n5671_);
  or g_7890 (new_n2272_, not_new_n6564_, not_new_n1580__332329305696010);
  not g_7891 (not_new_n590__0, new_n590_);
  or g_7892 (new_n9039_, or_or_not_new_n8833__not_new_n8830__0_not_new_n9222_, not_new_n9221_);
  not g_7893 (not_new_n6622__0, new_n6622_);
  not g_7894 (not_pi081, pi081);
  or g_7895 (new_n9548_, not_new_n9457_, not_new_n9546_);
  not g_7896 (not_new_n7404_, new_n7404_);
  not g_7897 (not_new_n9002__0, new_n9002_);
  not g_7898 (not_new_n6542_, new_n6542_);
  not g_7899 (not_new_n3945_, new_n3945_);
  not g_7900 (not_new_n8643_, new_n8643_);
  or g_7901 (new_n5652_, not_new_n1011__7, not_new_n5472_);
  or g_7902 (new_n3330_, not_new_n3933__0, not_pi064_6);
  or g_7903 (new_n9173_, not_new_n8978__1, not_new_n8809_);
  not g_7904 (not_new_n5504__0, new_n5504_);
  not g_7905 (not_new_n6540__0, new_n6540_);
  or g_7906 (new_n688_, not_new_n1506_, not_new_n3032_);
  not g_7907 (not_new_n596__70, key_gate_88);
  not g_7908 (not_new_n9066_, new_n9066_);
  not g_7909 (not_new_n1502_, new_n1502_);
  not g_7910 (not_pi269_3, pi269);
  not g_7911 (not_new_n3289_, new_n3289_);
  not g_7912 (not_new_n8079_, new_n8079_);
  not g_7913 (not_new_n608__57648010, new_n608_);
  and g_7914 (po103, key_gate_101, pi082);
  not g_7915 (not_new_n2980_, new_n2980_);
  not g_7916 (not_new_n1039__16284135979104490, new_n1039_);
  not g_7917 (not_new_n1487_, new_n1487_);
  or g_7918 (new_n5475_, not_new_n5712_, not_new_n5711_);
  not g_7919 (not_new_n5926_, new_n5926_);
  or g_7920 (new_n7895_, not_new_n7894_, not_new_n7769__0);
  or g_7921 (new_n4857_, not_new_n4760__1, not_new_n4843__1);
  not g_7922 (not_new_n1525_, new_n1525_);
  or g_7923 (new_n6951_, not_new_n6950_, not_new_n6814_);
  and g_7924 (new_n1570_, new_n3650_, new_n3651_);
  not g_7925 (not_new_n1071__47475615099430, new_n1071_);
  not g_7926 (not_new_n618__225393402906922580878632490, new_n618_);
  not g_7927 (not_new_n1051__968890104070, new_n1051_);
  not g_7928 (not_new_n7979_, new_n7979_);
  not g_7929 (not_new_n647__6, new_n647_);
  or g_7930 (new_n2925_, not_new_n640__3, not_new_n602__19773267430);
  not g_7931 (new_n4770_, new_n1599_);
  not g_7932 (not_new_n4606_, new_n4606_);
  not g_7933 (not_new_n602__4, new_n602_);
  not g_7934 (new_n8822_, new_n632_);
  not g_7935 (new_n5923_, new_n5775_);
  not g_7936 (not_new_n7944_, new_n7944_);
  not g_7937 (not_new_n586__3430, new_n586_);
  not g_7938 (not_new_n2947_, new_n2947_);
  or g_7939 (new_n9642_, not_new_n621__16284135979104490, not_new_n1598__6782230728490);
  or g_7940 (new_n3800_, not_new_n634__10, not_new_n1047__6);
  or g_7941 (new_n3523_, not_new_n1613__113988951853731430, not_new_n2345_);
  and g_7942 (and_new_n2359__new_n2358_, new_n2359_, new_n2358_);
  or g_7943 (new_n2954_, or_not_new_n2953__not_new_n2952_, not_new_n2951_);
  not g_7944 (not_new_n9641_, new_n9641_);
  not g_7945 (not_new_n3893_, new_n3893_);
  not g_7946 (not_new_n635__47475615099430, new_n635_);
  or g_7947 (new_n2347_, not_new_n1588__5585458640832840070, not_new_n1605_);
  or g_7948 (new_n1671_, not_po296_490, not_pi019);
  not g_7949 (not_pi044_0, pi044);
  or g_7950 (new_n8328_, not_new_n8326_, not_new_n8208_);
  not g_7951 (not_new_n7222__0, new_n7222_);
  and g_7952 (new_n1395_, new_n2473_, new_n2472_);
  and g_7953 (new_n9861_, new_n10119_, new_n9860_);
  not g_7954 (not_new_n3575_, new_n3575_);
  or g_7955 (new_n9522_, new_n642_, new_n1035_);
  or g_7956 (new_n2648_, not_new_n610__3430, not_new_n4457__0);
  not g_7957 (not_new_n1559_, new_n1559_);
  not g_7958 (not_pi124, pi124);
  not g_7959 (not_new_n4483__0, new_n4483_);
  not g_7960 (not_new_n649__0, new_n649_);
  not g_7961 (not_new_n6453_, new_n6453_);
  not g_7962 (not_new_n7023__0, new_n7023_);
  not g_7963 (not_new_n6292_, new_n6292_);
  not g_7964 (new_n3994_, pi033);
  not g_7965 (new_n6539_, new_n617_);
  not g_7966 (not_new_n1604__1176490, new_n1604_);
  not g_7967 (not_new_n3979__0, new_n3979_);
  or g_7968 (new_n4036_, not_new_n3991_, not_new_n4032__0);
  not g_7969 (new_n6805_, new_n6627_);
  or g_7970 (new_n6655_, not_new_n6488_, not_new_n1043__3430);
  or g_7971 (new_n6730_, not_new_n6510_, not_new_n1604__24010);
  not g_7972 (not_new_n4799_, new_n4799_);
  or g_7973 (new_n9604_, new_n645_, new_n1071_);
  not g_7974 (not_new_n624__138412872010, new_n624_);
  not g_7975 (not_new_n8126__0, new_n8126_);
  not g_7976 (not_new_n1493_, new_n1493_);
  or g_7977 (new_n5063_, not_new_n5288_, not_new_n5042_);
  not g_7978 (not_new_n7015__0, new_n7015_);
  not g_7979 (not_new_n4134__2, new_n4134_);
  or g_7980 (new_n3278_, not_new_n3184__168070, not_new_n632__8);
  not g_7981 (new_n7234_, new_n7146_);
  or g_7982 (new_n1742_, not_new_n1728__10, not_pi086);
  not g_7983 (not_new_n4445_, new_n4445_);
  not g_7984 (not_new_n989__3, new_n989_);
  or g_7985 (new_n7967_, not_new_n7809__0, not_new_n7737_);
  not g_7986 (not_new_n585__403536070, new_n585_);
  not g_7987 (not_new_n8171__0, new_n8171_);
  not g_7988 (new_n5453_, new_n1019_);
  not g_7989 (not_new_n5035_, new_n5035_);
  not g_7990 (not_new_n8551_, new_n8551_);
  or g_7991 (new_n4823_, not_new_n4729_, not_new_n1039__7);
  buf g_7992 (po033, pi231);
  not g_7993 (not_new_n2944_, new_n2944_);
  not g_7994 (not_new_n772_, new_n772_);
  not g_7995 (not_new_n5673_, new_n5673_);
  not g_7996 (not_new_n4632_, new_n4632_);
  not g_7997 (not_new_n9631__0, new_n9631_);
  or g_7998 (new_n964_, or_or_not_new_n1307__not_new_n1305__not_new_n2154_, not_new_n2153_);
  not g_7999 (not_new_n1631__1, key_gate_76);
  not g_8000 (not_new_n1728__797922662976120010, new_n1728_);
  and g_8001 (new_n583_, new_n1022_, new_n1021_);
  or g_8002 (or_or_not_new_n1406__not_new_n1407__not_new_n1410_, or_not_new_n1406__not_new_n1407_, not_new_n1410_);
  not g_8003 (not_new_n1027__6, new_n1027_);
  not g_8004 (not_new_n596__403536070, key_gate_88);
  not g_8005 (not_new_n4555_, new_n4555_);
  buf g_8006 (po021, pi243);
  not g_8007 (not_new_n8352_, new_n8352_);
  or g_8008 (new_n5378_, not_new_n5230_, not_new_n5071_);
  or g_8009 (new_n8047_, not_new_n7727_, not_new_n7756_);
  or g_8010 (new_n8565_, not_new_n8564_, not_new_n8563_);
  or g_8011 (new_n7968_, not_new_n7613__0, not_new_n1041__1176490);
  not g_8012 (not_new_n596__16284135979104490, key_gate_88);
  not g_8013 (not_new_n8440_, new_n8440_);
  and g_8014 (new_n9450_, new_n9451_, new_n9519_);
  or g_8015 (new_n1693_, not_new_n596__403536070, key_gate_17);
  not g_8016 (not_new_n1699_, key_gate_8);
  or g_8017 (new_n7479_, not_new_n7268_, not_new_n7477_);
  not g_8018 (not_new_n604__5, new_n604_);
  not g_8019 (not_new_n2837_, new_n2837_);
  not g_8020 (not_pi047, pi047);
  or g_8021 (new_n9208_, not_new_n9206_, not_new_n9002__0);
  not g_8022 (not_new_n636__2326305139872070, new_n636_);
  or g_8023 (new_n647_, not_new_n1922_, or_or_not_new_n1920__not_new_n1921__not_new_n1923_);
  not g_8024 (not_new_n6794_, new_n6794_);
  not g_8025 (new_n8150_, new_n1063_);
  or g_8026 (new_n3863_, not_new_n640__70, not_new_n6443__8235430);
  not g_8027 (new_n2237_, new_n972_);
  or g_8028 (new_n7431_, not_new_n775__403536070, not_new_n7125_);
  not g_8029 (not_po296_39098210485829880490, po296);
  not g_8030 (new_n7345_, new_n7026_);
  or g_8031 (new_n8720_, not_new_n1169__0, not_new_n8627_);
  and g_8032 (and_new_n2672__new_n2671_, new_n2671_, new_n2672_);
  not g_8033 (not_new_n5091_, new_n5091_);
  not g_8034 (new_n8650_, new_n1597_);
  not g_8035 (not_new_n8264__1, new_n8264_);
  not g_8036 (not_new_n3557_, new_n3557_);
  not g_8037 (not_new_n5628_, new_n5628_);
  not g_8038 (not_new_n4449_, new_n4449_);
  not g_8039 (not_new_n7366__2, new_n7366_);
  and g_8040 (and_and_new_n2295__new_n2298__new_n2296_, and_new_n2295__new_n2298_, new_n2296_);
  not g_8041 (not_new_n1057__10, new_n1057_);
  not g_8042 (not_new_n608__6, new_n608_);
  or g_8043 (new_n7414_, not_new_n6974__490, not_new_n762_);
  not g_8044 (not_new_n4561_, new_n4561_);
  or g_8045 (new_n2489_, not_new_n599__332329305696010, not_new_n9962__0);
  not g_8046 (new_n5922_, new_n5801_);
  not g_8047 (not_new_n4166__0, new_n4166_);
  not g_8048 (not_new_n2705_, new_n2705_);
  or g_8049 (new_n9843_, not_new_n9428__0, not_new_n9692_);
  or g_8050 (new_n10089_, new_n626_, new_n1053_);
  or g_8051 (new_n4532_, not_new_n1005__2, not_pi167_1);
  and g_8052 (new_n5888_, new_n6141_, new_n6142_);
  not g_8053 (not_new_n5607_, new_n5607_);
  not g_8054 (not_new_n1031__57648010, new_n1031_);
  not g_8055 (not_new_n1005__1, new_n1005_);
  not g_8056 (not_new_n8142__0, new_n8142_);
  and g_8057 (and_and_new_n1750__new_n1751__new_n1753_, new_n1753_, and_new_n1750__new_n1751_);
  and g_8058 (new_n4727_, new_n4820_, new_n4731_);
  not g_8059 (not_new_n4492_, new_n4492_);
  or g_8060 (new_n2884_, not_new_n4135__2, not_new_n3310__10);
  or g_8061 (new_n3844_, not_new_n1576__7, not_new_n628__490);
  not g_8062 (not_new_n9539_, new_n9539_);
  and g_8063 (new_n1516_, new_n3047_, and_new_n3049__new_n998_);
  not g_8064 (not_new_n4196_, new_n4196_);
  not g_8065 (not_new_n1616__6782230728490, new_n1616_);
  not g_8066 (not_new_n7365_, new_n7365_);
  not g_8067 (not_new_n1005__5, new_n1005_);
  not g_8068 (not_new_n9827_, new_n9827_);
  not g_8069 (not_new_n4980__0, new_n4980_);
  and g_8070 (new_n3968_, not_pi042_2, and_not_pi040_3_not_pi041_2);
  not g_8071 (new_n4279_, new_n653_);
  not g_8072 (not_new_n5830_, new_n5830_);
  not g_8073 (not_new_n8136__0, new_n8136_);
  not g_8074 (not_new_n4977_, new_n4977_);
  xor g_8075 (key_gate_41, not_new_n3977_, key_41);
  not g_8076 (new_n8540_, new_n8232_);
  or g_8077 (po223, or_or_not_new_n2597__not_new_n2601__not_new_n1435_, not_new_n1434_);
  or g_8078 (new_n3408_, not_new_n1594__0, not_new_n1010__1);
  or g_8079 (or_or_not_new_n1291__not_new_n1289__not_new_n2078_, or_not_new_n1291__not_new_n1289_, not_new_n2078_);
  or g_8080 (new_n3407_, not_pi031_0, not_new_n1536__24010);
  or g_8081 (new_n972_, or_or_not_new_n1323__not_new_n1321__not_new_n2230_, not_new_n2229_);
  and g_8082 (and_new_n6373__new_n6401_, new_n6373_, new_n6401_);
  or g_8083 (new_n6400_, not_new_n6255_, not_new_n635__8235430);
  not g_8084 (new_n8289_, new_n8139_);
  or g_8085 (new_n7347_, not_new_n6974__2, not_new_n774_);
  not g_8086 (not_new_n8623_, new_n8623_);
  not g_8087 (not_new_n10285_, new_n10285_);
  not g_8088 (not_new_n5955_, new_n5955_);
  or g_8089 (new_n2567_, not_new_n611__9, not_new_n2566_);
  or g_8090 (new_n2869_, not_po296_2115876138024253916377293617876786762900601936010, not_pi261_0);
  or g_8091 (new_n2255_, not_new_n5011_, not_new_n1589__6782230728490);
  and g_8092 (new_n8689_, new_n8751_, new_n8752_);
  not g_8093 (not_new_n621__5, new_n621_);
  or g_8094 (new_n6549_, not_new_n6871_, not_new_n6872_);
  not g_8095 (not_new_n1400_, new_n1400_);
  not g_8096 (not_new_n5962_, new_n5962_);
  not g_8097 (not_new_n984__797922662976120010, new_n984_);
  not g_8098 (not_new_n6443__2, new_n6443_);
  or g_8099 (new_n3334_, not_new_n3931__0, not_pi064_8);
  not g_8100 (not_pi233, pi233);
  not g_8101 (not_new_n6508__1, new_n6508_);
  not g_8102 (not_new_n6236_, new_n6236_);
  not g_8103 (not_new_n6800_, new_n6800_);
  not g_8104 (not_new_n9006_, new_n9006_);
  not g_8105 (not_new_n7399_, new_n7399_);
  or g_8106 (new_n7784_, not_new_n7610_, not_new_n7783_);
  not g_8107 (not_new_n6563_, new_n6563_);
  not g_8108 (not_new_n3113_, new_n3113_);
  not g_8109 (not_new_n597__3430, new_n597_);
  or g_8110 (new_n5021_, not_new_n5421_, not_new_n5420_);
  not g_8111 (not_pi038_2, pi038);
  not g_8112 (new_n9887_, new_n631_);
  not g_8113 (not_new_n619__70, new_n619_);
  not g_8114 (not_new_n4273_, new_n4273_);
  or g_8115 (new_n8323_, not_new_n631__113988951853731430, not_new_n8106__0);
  not g_8116 (not_new_n3815_, new_n3815_);
  or g_8117 (new_n4674_, not_new_n1014__3, not_new_n4443_);
  not g_8118 (not_new_n648__2326305139872070, new_n648_);
  or g_8119 (po082, key_gate_69, not_new_n1209_);
  not g_8120 (not_new_n7035_, new_n7035_);
  not g_8121 (not_new_n4429_, new_n4429_);
  not g_8122 (not_new_n5249_, new_n5249_);
  or g_8123 (new_n6741_, not_new_n629__57648010, not_new_n6502_);
  or g_8124 (new_n3145_, not_new_n645__6, not_new_n581__3119734822845423713013303218219760490);
  not g_8125 (not_new_n1538__57648010, new_n1538_);
  or g_8126 (new_n5780_, not_new_n5781_, not_new_n645__168070);
  not g_8127 (not_new_n2965_, new_n2965_);
  not g_8128 (not_new_n7909_, new_n7909_);
  or g_8129 (new_n2203_, not_new_n1602_, not_new_n1588__138412872010);
  not g_8130 (not_new_n6514_, new_n6514_);
  not g_8131 (not_new_n9361_, new_n9361_);
  or g_8132 (new_n9245_, not_new_n8850__0, not_new_n1598__968890104070);
  or g_8133 (new_n1006_, not_new_n3333_, not_new_n3334_);
  or g_8134 (or_or_not_new_n1564__not_new_n2479__not_new_n1397_, or_not_new_n1564__not_new_n2479_, not_new_n1397_);
  not g_8135 (not_new_n8977_, new_n8977_);
  and g_8136 (new_n5034_, new_n5146_, new_n5082_);
  and g_8137 (new_n9992_, new_n10130_, new_n10221_);
  not g_8138 (not_new_n643__403536070, new_n643_);
  not g_8139 (not_new_n5203_, new_n5203_);
  or g_8140 (new_n7401_, not_new_n7400_, not_new_n7399_);
  not g_8141 (not_new_n5325_, new_n5325_);
  not g_8142 (not_new_n6487__0, new_n6487_);
  not g_8143 (not_new_n9916__0, new_n9916_);
  not g_8144 (not_new_n622__6, new_n622_);
  or g_8145 (new_n5284_, not_new_n5197_, not_new_n621__24010);
  not g_8146 (not_new_n1603__16284135979104490, new_n1603_);
  not g_8147 (not_new_n8505_, new_n8505_);
  not g_8148 (not_new_n604__2824752490, new_n604_);
  not g_8149 (not_new_n3375__2, new_n3375_);
  or g_8150 (new_n2184_, not_new_n1603_, not_new_n1588__19773267430);
  or g_8151 (new_n3575_, not_new_n2242__0, not_new_n1612__968890104070);
  not g_8152 (not_new_n7769_, new_n7769_);
  not g_8153 (not_new_n1041__2, new_n1041_);
  and g_8154 (and_new_n1306__new_n2160_, new_n2160_, new_n1306_);
  not g_8155 (not_new_n9252_, new_n9252_);
  not g_8156 (not_new_n8636_, new_n8636_);
  and g_8157 (and_new_n3067__new_n998_, new_n3067_, new_n998_);
  or g_8158 (new_n2956_, not_new_n4124__2, not_new_n612__6);
  not g_8159 (not_new_n581__185621159210175743024531636712070, new_n581_);
  or g_8160 (or_not_new_n4322__0_not_new_n680__0, not_new_n4322__0, not_new_n680__0);
  or g_8161 (new_n5264_, not_new_n5083__0, not_new_n5247_);
  not g_8162 (new_n5448_, new_n1003_);
  not g_8163 (not_new_n7353_, new_n7353_);
  not g_8164 (not_new_n598__3, new_n598_);
  or g_8165 (new_n8413_, or_not_new_n8221__not_new_n8220_, not_new_n8376__0);
  not g_8166 (not_new_n1185_, new_n1185_);
  not g_8167 (not_new_n8880_, new_n8880_);
  or g_8168 (new_n7890_, not_new_n7729_, not_new_n7889_);
  not g_8169 (not_new_n5010_, new_n5010_);
  not g_8170 (not_new_n6574_, new_n6574_);
  or g_8171 (new_n1907_, not_new_n1583__6, not_new_n7685_);
  not g_8172 (not_new_n647__16284135979104490, new_n647_);
  or g_8173 (or_not_new_n1482__not_new_n2858_, not_new_n1482_, not_new_n2858_);
  not g_8174 (not_new_n5065_, new_n5065_);
  or g_8175 (new_n3910_, not_new_n643__24010, not_new_n9929__0);
  not g_8176 (not_new_n632__0, new_n632_);
  or g_8177 (new_n2784_, or_not_new_n2783__not_new_n2782_, not_new_n2781_);
  not g_8178 (not_new_n1382_, new_n1382_);
  or g_8179 (new_n9808_, not_new_n9401_, not_new_n1071__968890104070);
  not g_8180 (not_new_n3468_, new_n3468_);
  or g_8181 (new_n2409_, not_new_n599__10, not_new_n9973__0);
  or g_8182 (new_n6130_, not_new_n5808__0, or_not_new_n1596__3430_not_new_n5729_);
  not g_8183 (not_new_n1594__57648010, new_n1594_);
  or g_8184 (new_n3104_, not_new_n928__5, not_new_n1605__2);
  and g_8185 (new_n4310_, new_n4380_, new_n4379_);
  or g_8186 (new_n2882_, or_not_new_n2881__not_new_n2880_, not_new_n2879_);
  not g_8187 (not_new_n5898_, new_n5898_);
  not g_8188 (not_new_n1537__138412872010, new_n1537_);
  not g_8189 (not_new_n608__3430, new_n608_);
  not g_8190 (not_new_n3571_, new_n3571_);
  not g_8191 (new_n4812_, new_n4729_);
  or g_8192 (new_n9239_, not_new_n617__5585458640832840070, not_new_n8848__0);
  or g_8193 (new_n1877_, not_new_n9874_, not_new_n594__4);
  not g_8194 (not_new_n3995_, new_n3995_);
  or g_8195 (new_n6179_, not_new_n5899__2, not_new_n5867_);
  not g_8196 (not_new_n10270_, new_n10270_);
  not g_8197 (not_new_n2914_, new_n2914_);
  not g_8198 (not_new_n3487_, new_n3487_);
  xnor g_8199 (key_gate_106, not_new_n1714_, key_106);
  not g_8200 (not_new_n8226_, new_n8226_);
  or g_8201 (new_n3828_, not_new_n647__490, not_new_n1576_);
  not g_8202 (not_new_n5533_, new_n5533_);
  not g_8203 (not_new_n6213_, new_n6213_);
  not g_8204 (not_new_n636__332329305696010, new_n636_);
  not g_8205 (not_new_n1039_, new_n1039_);
  not g_8206 (not_new_n2603_, new_n2603_);
  not g_8207 (not_new_n3478_, new_n3478_);
  or g_8208 (new_n2932_, not_pi268_0, not_po296_1742514982336908143055105517947102601079450420187483430);
  or g_8209 (new_n731_, not_new_n3289_, not_new_n3290_);
  or g_8210 (or_or_not_new_n1556__not_new_n2439__not_new_n1381_, or_not_new_n1556__not_new_n2439_, not_new_n1381_);
  not g_8211 (not_new_n10230_, new_n10230_);
  or g_8212 (new_n2531_, not_new_n5485__0, not_new_n606__1);
  not g_8213 (not_new_n5391_, new_n5391_);
  not g_8214 (not_new_n3533_, new_n3533_);
  or g_8215 (or_or_not_new_n2955__not_new_n2958__not_new_n2957_, not_new_n2957_, or_not_new_n2955__not_new_n2958_);
  not g_8216 (new_n2342_, new_n620_);
  not g_8217 (not_new_n1394_, new_n1394_);
  and g_8218 (new_n8679_, new_n8600_, new_n1178_);
  or g_8219 (new_n2819_, not_new_n2816_, or_not_new_n2818__not_new_n2817_);
  or g_8220 (new_n5610_, not_pi135_2, not_new_n5444_);
  not g_8221 (not_new_n1933_, new_n1933_);
  not g_8222 (not_new_n8171__1, new_n8171_);
  or g_8223 (new_n8293_, not_new_n642__968890104070, not_new_n8265__1);
  not g_8224 (new_n3375_, new_n1024_);
  or g_8225 (new_n7659_, not_new_n7836_, not_new_n7838_);
  not g_8226 (not_new_n2551_, new_n2551_);
  or g_8227 (new_n10030_, not_new_n618__657123623635342801395430, not_new_n10013_);
  not g_8228 (not_new_n4019__0, new_n4019_);
  not g_8229 (not_pi169_2, pi169);
  not g_8230 (not_new_n3365_, new_n3365_);
  or g_8231 (new_n9621_, new_n630_, new_n1601_);
  not g_8232 (not_new_n3935_, new_n3935_);
  not g_8233 (not_new_n4938_, new_n4938_);
  not g_8234 (not_new_n9396_, new_n9396_);
  or g_8235 (new_n1178_, not_new_n3886_, not_new_n3885_);
  not g_8236 (not_pi192, pi192);
  not g_8237 (not_new_n2973_, new_n2973_);
  xnor g_8238 (key_gate_72, key_72, new_n1681_);
  not g_8239 (not_new_n2928_, new_n2928_);
  not g_8240 (not_pi146_1, pi146);
  not g_8241 (not_new_n1612__5, new_n1612_);
  or g_8242 (new_n3809_, not_new_n1043__6, not_new_n631__10);
  not g_8243 (not_new_n587__0, new_n587_);
  not g_8244 (not_new_n9483_, new_n9483_);
  not g_8245 (not_new_n594__2824752490, new_n594_);
  not g_8246 (new_n5443_, pi135);
  or g_8247 (new_n3120_, not_new_n928__70, not_new_n1598__3);
  not g_8248 (not_new_n667_, new_n667_);
  or g_8249 (new_n6091_, not_new_n1051__70, not_new_n5760__0);
  or g_8250 (new_n8488_, not_new_n8111__0, not_new_n1037__403536070);
  or g_8251 (new_n1784_, not_pi099, not_new_n588__0);
  not g_8252 (not_new_n622__24010, new_n622_);
  not g_8253 (not_new_n1597__332329305696010, new_n1597_);
  or g_8254 (new_n5173_, not_new_n4903_, not_new_n4999_);
  or g_8255 (new_n5534_, not_new_n1006__5, not_new_n5617_);
  or g_8256 (new_n2744_, not_po296_3119734822845423713013303218219760490, not_pi247);
  not g_8257 (not_new_n5239_, new_n5239_);
  and g_8258 (new_n1422_, new_n2538_, new_n2539_);
  not g_8259 (not_new_n8395_, new_n8395_);
  and g_8260 (new_n1563_, new_n3638_, new_n3639_);
  or g_8261 (new_n10075_, not_new_n9901_, not_new_n10074_);
  or g_8262 (new_n3193_, not_new_n635__7, not_new_n589__2);
  not g_8263 (not_new_n1174_, new_n1174_);
  not g_8264 (not_new_n7202_, new_n7202_);
  not g_8265 (not_new_n6065_, new_n6065_);
  or g_8266 (new_n4856_, not_new_n4747_, not_new_n1607__4);
  not g_8267 (not_new_n9524_, new_n9524_);
  not g_8268 (not_new_n774_, new_n774_);
  not g_8269 (not_new_n6695_, new_n6695_);
  not g_8270 (not_new_n6654__0, new_n6654_);
  not g_8271 (not_new_n7651__0, new_n7651_);
  not g_8272 (not_new_n3410_, new_n3410_);
  not g_8273 (not_new_n1155_, new_n1155_);
  not g_8274 (not_new_n7502_, new_n7502_);
  not g_8275 (not_new_n718__2, new_n718_);
  not g_8276 (not_new_n1037__16284135979104490, new_n1037_);
  not g_8277 (new_n9668_, new_n9428_);
  or g_8278 (new_n4722_, not_new_n623__5, not_new_n4719_);
  or g_8279 (po065, key_gate_64, not_new_n1192_);
  not g_8280 (not_new_n5897_, new_n5897_);
  not g_8281 (not_new_n3589_, new_n3589_);
  not g_8282 (not_new_n1404_, new_n1404_);
  not g_8283 (not_new_n634__403536070, new_n634_);
  or g_8284 (new_n9636_, not_new_n9494_, not_new_n9627_);
  not g_8285 (not_new_n6907_, new_n6907_);
  not g_8286 (not_new_n9308_, new_n9308_);
  not g_8287 (not_new_n3523_, new_n3523_);
  not g_8288 (not_new_n1261_, new_n1261_);
  or g_8289 (new_n2516_, not_new_n1416_, not_new_n611__3);
  not g_8290 (new_n7655_, new_n637_);
  not g_8291 (not_new_n5160_, new_n5160_);
  or g_8292 (new_n5637_, not_new_n5433__0, not_new_n1009__7);
  or g_8293 (new_n7021_, not_new_n7362_, not_new_n7361_);
  not g_8294 (not_new_n10202_, new_n10202_);
  or g_8295 (new_n2650_, not_new_n1006__0, not_new_n608__3430);
  not g_8296 (not_new_n600_, new_n600_);
  not g_8297 (not_new_n3465_, new_n3465_);
  not g_8298 (not_new_n2016_, new_n2016_);
  not g_8299 (not_new_n4943_, new_n4943_);
  or g_8300 (new_n4864_, not_new_n1599__7, not_new_n4745_);
  or g_8301 (new_n5065_, not_new_n5201_, not_new_n5044_);
  and g_8302 (new_n1250_, new_n1891_, new_n1892_);
  not g_8303 (not_new_n8709_, new_n8709_);
  not g_8304 (not_new_n8164__0, new_n8164_);
  not g_8305 (not_new_n648__16284135979104490, new_n648_);
  or g_8306 (new_n5644_, not_new_n5642_, not_new_n5643_);
  buf g_8307 (po012, pi205);
  not g_8308 (not_new_n9722_, new_n9722_);
  and g_8309 (new_n6242_, new_n6382_, new_n6317_);
  or g_8310 (new_n9320_, not_new_n8978__3, not_new_n9165_);
  or g_8311 (new_n6728_, not_new_n6511_, not_new_n1071__3430);
  not g_8312 (not_new_n619__4, new_n619_);
  not g_8313 (not_new_n7839_, new_n7839_);
  not g_8314 (not_new_n1537__0, new_n1537_);
  and g_8315 (new_n6331_, new_n6232_, new_n1045_);
  not g_8316 (not_new_n7081_, new_n7081_);
  not g_8317 (not_new_n4586_, new_n4586_);
  or g_8318 (new_n5814_, not_new_n6067_, not_new_n5795_);
  not g_8319 (new_n10037_, new_n9940_);
  or g_8320 (new_n3309_, not_new_n1619__0, not_new_n1595__0);
  or g_8321 (new_n3428_, not_new_n1594__4, not_new_n1006__1);
  not g_8322 (not_new_n608__1, new_n608_);
  not g_8323 (not_new_n645__7, new_n645_);
  or g_8324 (new_n6194_, not_new_n5902_, not_new_n5870_);
  not g_8325 (not_new_n1537__6, new_n1537_);
  or g_8326 (new_n6085_, not_new_n5890__2, not_new_n5909_);
  not g_8327 (not_new_n8394_, new_n8394_);
  not g_8328 (not_new_n1498_, new_n1498_);
  not g_8329 (not_new_n9985_, new_n9985_);
  and g_8330 (new_n7732_, new_n7901_, new_n7572_);
  not g_8331 (not_new_n6233__1, new_n6233_);
  or g_8332 (new_n677_, or_not_new_n3110__not_new_n3109_, not_new_n3108_);
  or g_8333 (new_n9201_, not_new_n9199_, not_new_n9010_);
  not g_8334 (not_new_n7864_, new_n7864_);
  or g_8335 (new_n7352_, not_new_n775__5, not_new_n7104_);
  or g_8336 (new_n6196_, not_new_n5785__0, not_new_n637__1176490);
  or g_8337 (new_n9894_, not_new_n10057_, not_new_n10058_);
  not g_8338 (not_new_n3185_, new_n3185_);
  not g_8339 (new_n4816_, new_n4731_);
  not g_8340 (not_new_n9779_, new_n9779_);
  not g_8341 (not_new_n3536_, new_n3536_);
  not g_8342 (not_new_n1005__7, new_n1005_);
  not g_8343 (not_new_n8069_, new_n8069_);
  not g_8344 (not_new_n634__16284135979104490, new_n634_);
  not g_8345 (not_new_n4193_, new_n4193_);
  or g_8346 (new_n3770_, not_new_n1051__6, not_new_n647__10);
  not g_8347 (not_new_n1580__8, new_n1580_);
  not g_8348 (not_new_n6232__3, new_n6232_);
  or g_8349 (new_n10287_, not_new_n10148_, not_new_n10285_);
  not g_8350 (not_pi008, pi008);
  not g_8351 (new_n9351_, new_n1039_);
  not g_8352 (not_new_n6633_, new_n6633_);
  not g_8353 (not_new_n959_, new_n959_);
  not g_8354 (not_new_n4279_, new_n4279_);
  not g_8355 (not_new_n5939_, new_n5939_);
  not g_8356 (not_po298_47475615099430, po298);
  not g_8357 (not_new_n4475__0, new_n4475_);
  not g_8358 (not_new_n1041__8, new_n1041_);
  and g_8359 (new_n1523_, new_n3068_, and_new_n3070__new_n998_);
  or g_8360 (or_or_not_new_n1567__not_new_n2494__not_new_n1403_, not_new_n1403_, or_not_new_n1567__not_new_n2494_);
  not g_8361 (not_new_n4164_, new_n4164_);
  not g_8362 (not_new_n1602__8, new_n1602_);
  or g_8363 (new_n8907_, not_new_n9219_, not_new_n9220_);
  or g_8364 (new_n6879_, not_new_n6875_, not_new_n6647__0);
  or g_8365 (new_n6568_, not_new_n6942_, not_new_n6941_);
  not g_8366 (not_new_n600__332329305696010, new_n600_);
  and g_8367 (new_n6336_, new_n6232_, new_n6260_);
  or g_8368 (new_n8039_, not_new_n7660__0, not_new_n646__19773267430);
  or g_8369 (new_n7536_, not_new_n7534_, not_new_n7535_);
  not g_8370 (not_new_n1388_, new_n1388_);
  and g_8371 (new_n4908_, new_n4905_, new_n5186_);
  not g_8372 (not_new_n9102_, new_n9102_);
  not g_8373 (not_new_n3372__3430, new_n3372_);
  not g_8374 (not_new_n5741__0, new_n5741_);
  or g_8375 (new_n10316_, not_new_n9910__0, not_new_n639__273687473400809163430);
  xor g_8376 (key_gate_9, key_9, not_new_n1183_);
  not g_8377 (not_new_n605__3430, new_n605_);
  or g_8378 (po176, not_new_n3578_, not_new_n3579_);
  not g_8379 (not_new_n8861_, new_n8861_);
  or g_8380 (new_n10230_, not_new_n9951_, not_new_n9859_);
  not g_8381 (new_n6982_, new_n743_);
  not g_8382 (new_n8360_, new_n8144_);
  or g_8383 (new_n4355_, not_new_n698_, not_new_n4252_);
  not g_8384 (not_new_n8556_, new_n8556_);
  not g_8385 (not_new_n5770__1, new_n5770_);
  xor g_8386 (key_gate_23, key_23, new_n1726_);
  not g_8387 (not_new_n599__2, new_n599_);
  or g_8388 (new_n9184_, not_new_n9097_, not_new_n621__332329305696010);
  or g_8389 (or_not_new_n4234__not_new_n4336_, not_new_n4336_, not_new_n4234_);
  not g_8390 (not_new_n1059__8, new_n1059_);
  not g_8391 (not_new_n1051__3, new_n1051_);
  not g_8392 (not_new_n6997__0, new_n6997_);
  or g_8393 (new_n3335_, not_pi037_0, not_new_n1534__9);
  not g_8394 (not_new_n10128_, new_n10128_);
  not g_8395 (not_pi219, pi219);
  not g_8396 (not_pi041_0, pi041);
  not g_8397 (not_po296_5, po296);
  not g_8398 (not_new_n1159__1, new_n1159_);
  not g_8399 (not_new_n1481_, new_n1481_);
  not g_8400 (not_pi171_0, pi171);
  not g_8401 (not_new_n597__490, new_n597_);
  and g_8402 (new_n5025_, new_n1031_, new_n641_);
  not g_8403 (not_new_n627__3430, new_n627_);
  not g_8404 (not_new_n1005__0, new_n1005_);
  or g_8405 (new_n5234_, not_new_n5050_, not_new_n5233_);
  and g_8406 (new_n9991_, new_n9859_, new_n9865_);
  or g_8407 (new_n1961_, not_new_n4136_, not_new_n585__10);
  not g_8408 (new_n6796_, new_n6542_);
  or g_8409 (new_n1180_, not_new_n3889_, not_new_n3890_);
  not g_8410 (not_new_n7251_, new_n7251_);
  not g_8411 (not_new_n1622__0, new_n1622_);
  not g_8412 (not_new_n8391_, new_n8391_);
  or g_8413 (new_n6201_, not_new_n6023__0, not_new_n5903_);
  or g_8414 (new_n7889_, not_new_n7887_, not_new_n7888_);
  not g_8415 (not_new_n4103_, new_n4103_);
  not g_8416 (not_new_n7047__0, new_n7047_);
  not g_8417 (not_new_n5760__0, new_n5760_);
  not g_8418 (not_new_n3957_, new_n3957_);
  or g_8419 (new_n1633_, key_gate_78, key_gate_63);
  or g_8420 (or_not_new_n5460__not_new_n5686__1, not_new_n5460_, not_new_n5686__1);
  not g_8421 (not_new_n6887_, new_n6887_);
  or g_8422 (new_n5097_, not_new_n5022_, not_new_n4898_);
  or g_8423 (new_n5485_, not_new_n5665_, not_new_n5664_);
  not g_8424 (not_new_n8995__1, new_n8995_);
  not g_8425 (new_n4491_, pi180);
  or g_8426 (new_n6128_, not_new_n5884__0, not_new_n619__70);
  and g_8427 (new_n6334_, and_new_n6373__new_n6401_, new_n6253_);
  not g_8428 (not_new_n621__273687473400809163430, new_n621_);
  or g_8429 (new_n3529_, not_new_n1805__0, not_new_n1612__0);
  or g_8430 (new_n4372_, not_new_n4369_, not_new_n4307_);
  or g_8431 (new_n9314_, not_new_n9312_, not_new_n9313_);
  or g_8432 (new_n756_, not_new_n3223_, not_new_n3222_);
  not g_8433 (not_new_n8969_, new_n8969_);
  not g_8434 (not_new_n10255_, new_n10255_);
  and g_8435 (new_n1568_, new_n3649_, new_n3648_);
  not g_8436 (not_new_n8680_, new_n8680_);
  or g_8437 (new_n3332_, not_new_n3932__0, not_pi064_7);
  not g_8438 (not_pi064_797922662976120010, pi064);
  not g_8439 (not_new_n3310__24010, new_n3310_);
  not g_8440 (not_new_n7071_, new_n7071_);
  or g_8441 (new_n8583_, not_new_n8240_, not_new_n8273_);
  or g_8442 (new_n7300_, not_new_n7415__1, not_new_n6995__1);
  not g_8443 (not_new_n9408_, new_n9408_);
  not g_8444 (not_new_n9116_, new_n9116_);
  not g_8445 (not_new_n5754__1, new_n5754_);
  not g_8446 (not_new_n4978__0, new_n4978_);
  or g_8447 (new_n8544_, not_new_n8264__1, not_new_n642__47475615099430);
  not g_8448 (not_new_n645__138412872010, new_n645_);
  not g_8449 (not_new_n4787__0, new_n4787_);
  not g_8450 (not_new_n6855_, new_n6855_);
  and g_8451 (new_n1200_, new_n1689_, new_n1691_);
  not g_8452 (not_new_n2938_, new_n2938_);
  not g_8453 (not_new_n7601__0, new_n7601_);
  not g_8454 (not_new_n619__3, new_n619_);
  not g_8455 (not_new_n5254_, new_n5254_);
  not g_8456 (not_new_n928_, new_n928_);
  not g_8457 (not_new_n9060_, new_n9060_);
  not g_8458 (not_new_n4096_, new_n4096_);
  not g_8459 (not_pi167, pi167);
  not g_8460 (not_new_n5912__0, new_n5912_);
  xnor g_8461 (key_gate_69, key_69, not_new_n1717_);
  not g_8462 (new_n7445_, new_n7040_);
  or g_8463 (new_n1734_, not_pi078, not_new_n1728__2);
  not g_8464 (not_new_n7937_, new_n7937_);
  not g_8465 (not_new_n984__70, new_n984_);
  and g_8466 (and_new_n2238__new_n2241_, new_n2241_, new_n2238_);
  or g_8467 (new_n1047_, not_new_n3438_, not_new_n3437_);
  or g_8468 (new_n2466_, not_new_n597__19773267430, not_new_n4779__0);
  or g_8469 (new_n7364_, not_new_n7108_, not_new_n775__9);
  not g_8470 (not_new_n6487_, new_n6487_);
  or g_8471 (new_n2923_, not_pi267, not_po296_248930711762415449007872216849586085868492917169640490);
  and g_8472 (new_n1375_, new_n2422_, and_new_n2424__new_n2423_);
  not g_8473 (not_new_n6373__1, new_n6373_);
  not g_8474 (not_pi088, pi088);
  not g_8475 (new_n8958_, new_n619_);
  not g_8476 (not_new_n9253_, new_n9253_);
  or g_8477 (new_n4690_, not_new_n4439__0, not_new_n1016__4);
  not g_8478 (not_new_n1055__4, new_n1055_);
  not g_8479 (not_new_n5136_, new_n5136_);
  not g_8480 (not_new_n2601_, new_n2601_);
  or g_8481 (new_n6905_, not_new_n6631__1, not_new_n6759_);
  not g_8482 (not_new_n3700_, new_n3700_);
  not g_8483 (not_new_n4019__1, new_n4019_);
  not g_8484 (not_pi206, pi206);
  not g_8485 (not_pi130_1, pi130);
  not g_8486 (not_new_n638__403536070, new_n638_);
  or g_8487 (new_n695_, not_new_n3057_, not_new_n1519_);
  not g_8488 (not_new_n8707__0, new_n8707_);
  or g_8489 (new_n5986_, not_new_n5905_, not_new_n5724_);
  or g_8490 (or_not_new_n2585__not_new_n2584_, not_new_n2585_, not_new_n2584_);
  or g_8491 (new_n6075_, not_new_n5763_, not_new_n5837_);
  not g_8492 (not_new_n5251_, new_n5251_);
  or g_8493 (new_n1001_, not_new_n3317_, not_new_n3316_);
  not g_8494 (not_new_n1863_, new_n1863_);
  not g_8495 (not_new_n3444_, new_n3444_);
  not g_8496 (new_n9945_, new_n618_);
  not g_8497 (not_pi047_1, pi047);
  not g_8498 (not_new_n7338_, new_n7338_);
  or g_8499 (new_n6736_, not_new_n6735_, not_new_n6451_);
  not g_8500 (not_pi133_2, pi133);
  not g_8501 (new_n6548_, new_n641_);
  or g_8502 (new_n10149_, new_n617_, new_n1597_);
  not g_8503 (not_new_n7767_, new_n7767_);
  or g_8504 (new_n2504_, not_new_n4756__0, not_new_n597__797922662976120010);
  not g_8505 (not_new_n1047__24010, new_n1047_);
  or g_8506 (new_n4094_, not_new_n4165_, not_pi249_1);
  or g_8507 (new_n7524_, not_new_n7230_, not_new_n7522_);
  not g_8508 (new_n4983_, new_n633_);
  not g_8509 (not_new_n6239_, new_n6239_);
  not g_8510 (not_new_n2841_, new_n2841_);
  or g_8511 (new_n10155_, not_new_n10016__0, not_new_n10144_);
  or g_8512 (new_n1717_, not_new_n596__2326305139872070, key_gate_119);
  not g_8513 (not_new_n611__490, new_n611_);
  or g_8514 (new_n3498_, not_new_n1028__7, not_new_n1594__57648010);
  not g_8515 (not_new_n1606__0, new_n1606_);
  not g_8516 (new_n9524_, new_n9358_);
  or g_8517 (new_n5609_, not_new_n5443_, not_new_n1005__6);
  not g_8518 (not_new_n1603__168070, new_n1603_);
  not g_8519 (not_new_n4768_, new_n4768_);
  not g_8520 (not_new_n597__2, new_n597_);
  not g_8521 (not_new_n5617_, new_n5617_);
  or g_8522 (new_n2845_, not_new_n994__24010, not_new_n4130__1);
  not g_8523 (not_new_n2509__24010, new_n2509_);
  or g_8524 (new_n2415_, not_new_n598__70, not_new_n1057__0);
  or g_8525 (new_n2858_, not_new_n1616__490, not_new_n2855_);
  not g_8526 (not_new_n1057__1, new_n1057_);
  or g_8527 (new_n7384_, not_new_n6979__0, not_new_n7022__0);
  not g_8528 (not_new_n1599__168070, new_n1599_);
  not g_8529 (not_new_n1601__1915812313805664144010, new_n1601_);
  not g_8530 (not_new_n4774_, new_n4774_);
  or g_8531 (new_n6795_, not_new_n6543_, not_new_n6740_);
  not g_8532 (not_new_n10220_, new_n10220_);
  not g_8533 (not_new_n3552_, new_n3552_);
  not g_8534 (not_new_n611__2824752490, new_n611_);
  not g_8535 (not_new_n630__3, new_n630_);
  and g_8536 (new_n1207_, new_n1710_, new_n1712_);
  not g_8537 (not_new_n7504_, new_n7504_);
  not g_8538 (not_new_n2188_, new_n2188_);
  or g_8539 (new_n9821_, not_new_n9820_, not_new_n9819_);
  or g_8540 (new_n6853_, not_new_n6486__0, not_new_n628__19773267430);
  not g_8541 (not_new_n596__4, key_gate_88);
  not g_8542 (not_new_n4315_, new_n4315_);
  or g_8543 (new_n7888_, not_new_n638__332329305696010, not_new_n7643__0);
  and g_8544 (new_n1420_, new_n2529_, new_n2528_);
  not g_8545 (not_new_n595_, new_n595_);
  not g_8546 (not_new_n5788__0, new_n5788_);
  and g_8547 (new_n1315_, and_new_n1314__new_n2198_, new_n2197_);
  or g_8548 (new_n8751_, not_new_n8595__1, not_new_n8673_);
  and g_8549 (new_n5856_, and_new_n6016__new_n5855_, new_n6013_);
  not g_8550 (new_n1905_, new_n648_);
  not g_8551 (not_new_n1599__5, new_n1599_);
  not g_8552 (not_new_n8232_, new_n8232_);
  or g_8553 (new_n7020_, not_new_n7365_, not_new_n7364_);
  not g_8554 (not_new_n4556_, new_n4556_);
  or g_8555 (new_n3298_, not_new_n626__8, not_new_n3184__47475615099430);
  not g_8556 (not_new_n644__2, new_n644_);
  not g_8557 (not_pi260_1, pi260);
  not g_8558 (new_n1612_, new_n1538_);
  not g_8559 (not_new_n8793_, new_n8793_);
  not g_8560 (not_new_n634__968890104070, new_n634_);
  not g_8561 (not_new_n9672_, new_n9672_);
  not g_8562 (not_new_n10232_, new_n10232_);
  and g_8563 (new_n1493_, new_n3009_, new_n3010_);
  not g_8564 (not_new_n5863_, new_n5863_);
  not g_8565 (not_new_n3866_, new_n3866_);
  not g_8566 (not_new_n1605__0, new_n1605_);
  not g_8567 (not_pi250_0, pi250);
  or g_8568 (new_n6000_, not_new_n5923_, not_new_n5718_);
  or g_8569 (new_n2633_, not_new_n609__490, not_new_n4456_);
  not g_8570 (new_n9381_, new_n629_);
  and g_8571 (new_n3919_, new_n3952_, new_n4042_);
  not g_8572 (new_n9880_, new_n1047_);
  not g_8573 (not_new_n5511__0, new_n5511_);
  not g_8574 (not_new_n2169_, new_n2169_);
  or g_8575 (new_n6554_, not_new_n6920_, not_new_n6921_);
  not g_8576 (not_new_n1613__5, new_n1613_);
  not g_8577 (not_new_n5916_, new_n5916_);
  or g_8578 (new_n8775_, not_new_n8647_, not_new_n1164__0);
  not g_8579 (not_new_n7663__0, new_n7663_);
  not g_8580 (not_new_n1049__47475615099430, new_n1049_);
  not g_8581 (not_new_n643_, new_n643_);
  and g_8582 (new_n7745_, new_n7998_, new_n7999_);
  not g_8583 (not_new_n1611__70, new_n1611_);
  not g_8584 (not_pi232, pi232);
  not g_8585 (not_new_n7644_, new_n7644_);
  or g_8586 (new_n7378_, not_new_n739__0, not_new_n7366__2);
  not g_8587 (not_new_n4128__2, new_n4128_);
  not g_8588 (not_new_n5749_, new_n5749_);
  not g_8589 (not_new_n623__0, new_n623_);
  not g_8590 (not_new_n3689_, new_n3689_);
  not g_8591 (not_new_n598__19773267430, new_n598_);
  not g_8592 (not_new_n604__47475615099430, new_n604_);
  not g_8593 (not_new_n8462_, new_n8462_);
  not g_8594 (not_new_n7293__0, new_n7293_);
  or g_8595 (new_n9229_, not_new_n9227_, not_new_n9107_);
  or g_8596 (new_n6126_, not_new_n6124_, not_new_n6125_);
  not g_8597 (new_n5547_, new_n5496_);
  not g_8598 (not_new_n4150_, new_n4150_);
  not g_8599 (not_new_n7003__1, new_n7003_);
  or g_8600 (new_n2652_, not_new_n2509__3430, not_pi207);
  not g_8601 (not_new_n9703_, new_n9703_);
  not g_8602 (not_new_n9747_, new_n9747_);
  not g_8603 (not_new_n5553_, new_n5553_);
  not g_8604 (not_new_n637__6782230728490, new_n637_);
  not g_8605 (not_pi134_1, pi134);
  and g_8606 (new_n4776_, new_n4868_, new_n4869_);
  or g_8607 (new_n3524_, not_new_n1537__797922662976120010, not_pi128_0);
  not g_8608 (not_new_n7334__0, new_n7334_);
  not g_8609 (not_new_n6132_, new_n6132_);
  not g_8610 (not_new_n7855_, new_n7855_);
  or g_8611 (or_not_new_n5764__0_not_new_n618__8235430, not_new_n618__8235430, not_new_n5764__0);
  not g_8612 (not_new_n611__3, new_n611_);
  not g_8613 (not_new_n625__24010, new_n625_);
  not g_8614 (not_new_n1532_, new_n1532_);
  not g_8615 (not_new_n966_, new_n966_);
  or g_8616 (new_n1151_, not_new_n3832_, not_new_n3831_);
  not g_8617 (not_new_n1059__3, new_n1059_);
  not g_8618 (not_new_n5901_, new_n5901_);
  not g_8619 (new_n3944_, pi061);
  not g_8620 (not_new_n1602__3, new_n1602_);
  not g_8621 (not_new_n7567_, new_n7567_);
  not g_8622 (not_new_n8106_, new_n8106_);
  or g_8623 (new_n10269_, not_new_n619__6782230728490, not_new_n10009__0);
  and g_8624 (new_n8097_, new_n8414_, new_n8383_);
  not g_8625 (not_new_n1385_, new_n1385_);
  not g_8626 (not_new_n8575_, new_n8575_);
  or g_8627 (new_n3814_, not_new_n1609__0, not_new_n991__0);
  or g_8628 (new_n4849_, not_new_n4818__1, not_new_n4749__1);
  not g_8629 (not_new_n1612__8235430, new_n1612_);
  not g_8630 (not_new_n7991_, new_n7991_);
  and g_8631 (new_n601_, new_n1021_, new_n1609_);
  and g_8632 (and_new_n2647__new_n2648_, new_n2647_, new_n2648_);
  or g_8633 (new_n9293_, not_new_n9292_, not_new_n9291_);
  or g_8634 (new_n3013_, not_new_n623__0, not_new_n3372__70);
  not g_8635 (not_pi144_3, pi144);
  not g_8636 (not_new_n3464_, new_n3464_);
  not g_8637 (not_new_n9610_, new_n9610_);
  not g_8638 (not_new_n2845_, new_n2845_);
  or g_8639 (new_n1812_, not_new_n7688_, not_new_n1583__1);
  or g_8640 (new_n9608_, not_new_n9607_, not_new_n9425_);
  or g_8641 (po126, not_new_n3446_, not_new_n3445_);
  not g_8642 (not_new_n2787_, new_n2787_);
  or g_8643 (new_n7062_, not_new_n7517_, not_new_n7516_);
  or g_8644 (new_n2371_, not_new_n597__2, not_new_n4724__0);
  not g_8645 (not_new_n8984_, new_n8984_);
  or g_8646 (po238, not_new_n3662_, not_new_n3663_);
  not g_8647 (not_new_n6854_, new_n6854_);
  not g_8648 (not_new_n3950_, new_n3950_);
  not g_8649 (not_new_n9427__3, new_n9427_);
  not g_8650 (not_new_n620__2, new_n620_);
  and g_8651 (new_n8806_, new_n8801_, new_n9011_);
  or g_8652 (new_n6078_, not_new_n5846_, not_new_n6077_);
  not g_8653 (not_new_n2299_, new_n2299_);
  not g_8654 (not_new_n5159__0, new_n5159_);
  not g_8655 (not_pi142_1, pi142);
  not g_8656 (not_new_n7517_, new_n7517_);
  not g_8657 (not_new_n7612__0, new_n7612_);
  not g_8658 (not_new_n8804_, new_n8804_);
  not g_8659 (not_new_n5388_, new_n5388_);
  or g_8660 (new_n3354_, not_pi064_57648010, not_new_n3917__0);
  or g_8661 (new_n9599_, not_new_n633__2326305139872070, not_new_n9598_);
  not g_8662 (not_new_n1609__1, new_n1609_);
  not g_8663 (new_n4420_, new_n1008_);
  or g_8664 (new_n5733_, not_new_n5910_, not_new_n5857_);
  or g_8665 (new_n5421_, not_new_n5150_, not_new_n5419_);
  and g_8666 (new_n1427_, new_n2560_, new_n2562_);
  not g_8667 (new_n7100_, new_n770_);
  not g_8668 (not_new_n1589__6782230728490, new_n1589_);
  not g_8669 (not_new_n640__2824752490, new_n640_);
  not g_8670 (not_new_n2848_, new_n2848_);
  not g_8671 (not_new_n624__2824752490, new_n624_);
  not g_8672 (not_new_n3722_, new_n3722_);
  not g_8673 (not_new_n6982_, new_n6982_);
  not g_8674 (new_n8386_, new_n8260_);
  and g_8675 (new_n1241_, new_n1852_, new_n1851_);
  or g_8676 (new_n2141_, not_new_n1589__57648010, not_new_n5015_);
  not g_8677 (not_new_n3372__9, new_n3372_);
  not g_8678 (not_new_n7646__0, new_n7646_);
  not g_8679 (not_new_n636__403536070, new_n636_);
  not g_8680 (not_new_n5771_, new_n5771_);
  not g_8681 (not_new_n1594__1176490, new_n1594_);
  not g_8682 (not_new_n4167__0, new_n4167_);
  or g_8683 (new_n5984_, not_new_n1061__3430, not_new_n5800_);
  or g_8684 (or_not_new_n2535__not_new_n2534_, not_new_n2534_, not_new_n2535_);
  not g_8685 (not_new_n9888__1, new_n9888_);
  and g_8686 (new_n9326_, new_n9518_, new_n9517_);
  or g_8687 (new_n3160_, not_new_n643__6, not_new_n581__52433383167563036344614587188619514555430);
  not g_8688 (not_pi166_2, pi166);
  or g_8689 (new_n1538_, not_new_n615__0, not_new_n1345_);
  not g_8690 (not_new_n4749__0, new_n4749_);
  or g_8691 (or_not_new_n8139__1_not_new_n8231_, not_new_n8231_, not_new_n8139__1);
  not g_8692 (not_new_n10102_, new_n10102_);
  xnor g_8693 (key_gate_111, key_111, new_n1708_);
  or g_8694 (new_n8193_, not_new_n8481_, not_new_n8482_);
  not g_8695 (not_new_n5535_, new_n5535_);
  not g_8696 (not_new_n9783_, new_n9783_);
  or g_8697 (or_not_new_n1027__0_not_new_n3384_, not_new_n3384_, not_new_n1027__0);
  not g_8698 (not_new_n686_, new_n686_);
  not g_8699 (not_new_n3664_, new_n3664_);
  or g_8700 (new_n5423_, not_new_n1053__70, not_new_n4961_);
  not g_8701 (not_new_n4628_, new_n4628_);
  or g_8702 (new_n6892_, not_new_n6805_, not_new_n6891_);
  not g_8703 (not_new_n628__8235430, new_n628_);
  not g_8704 (not_new_n597__16284135979104490, new_n597_);
  not g_8705 (not_new_n8262_, new_n8262_);
  or g_8706 (new_n10011_, or_not_new_n10210__not_new_n10153_, not_new_n10030_);
  not g_8707 (not_new_n8557_, new_n8557_);
  and g_8708 (new_n8221_, new_n8382_, new_n8093_);
  not g_8709 (not_new_n621__6782230728490, new_n621_);
  not g_8710 (not_new_n1037__490, new_n1037_);
  not g_8711 (not_new_n1157_, new_n1157_);
  or g_8712 (new_n5938_, not_new_n1041__10, not_new_n5756_);
  or g_8713 (new_n7289_, not_new_n7029__0, not_new_n728__0);
  not g_8714 (not_new_n6502_, new_n6502_);
  not g_8715 (not_new_n624__332329305696010, new_n624_);
  or g_8716 (new_n3228_, not_new_n1063__4, not_new_n3185__2824752490);
  not g_8717 (not_new_n4294_, new_n4294_);
  and g_8718 (new_n9872_, new_n10159_, new_n10162_);
  not g_8719 (not_new_n9341_, new_n9341_);
  not g_8720 (not_new_n7759__0, new_n7759_);
  not g_8721 (not_new_n587__4, new_n587_);
  not g_8722 (not_new_n9045_, new_n9045_);
  not g_8723 (new_n4171_, new_n4104_);
  not g_8724 (not_new_n617__5, new_n617_);
  not g_8725 (not_new_n5680__1, new_n5680_);
  or g_8726 (new_n5543_, not_new_n1004__5, not_pi136_1);
  not g_8727 (not_new_n5129_, new_n5129_);
  not g_8728 (new_n8130_, new_n622_);
  or g_8729 (new_n5882_, not_new_n6075_, not_new_n5838_);
  or g_8730 (or_or_or_not_new_n2838__not_new_n2841__not_new_n2840__not_new_n2842_, or_or_not_new_n2838__not_new_n2841__not_new_n2840_, not_new_n2842_);
  not g_8731 (not_new_n644__1176490, new_n644_);
  not g_8732 (not_new_n626__9, new_n626_);
  or g_8733 (new_n757_, not_new_n3224_, not_new_n3225_);
  not g_8734 (not_new_n7183_, new_n7183_);
  not g_8735 (not_new_n1476_, new_n1476_);
  not g_8736 (not_new_n621__2, new_n621_);
  or g_8737 (new_n6153_, not_new_n5769__0, not_new_n629__1176490);
  not g_8738 (not_new_n5753_, new_n5753_);
  not g_8739 (not_new_n10241_, new_n10241_);
  or g_8740 (new_n7146_, not_new_n7232_, not_new_n7233_);
  not g_8741 (not_new_n1581__4, new_n1581_);
  or g_8742 (new_n1775_, not_new_n1589_, not_new_n5002_);
  or g_8743 (new_n8073_, not_new_n626__113988951853731430, not_new_n7651__2);
  not g_8744 (not_new_n4071__1, new_n4071_);
  or g_8745 (new_n4374_, not_new_n4267_, not_new_n691_);
  not g_8746 (new_n4099_, pi264);
  or g_8747 (new_n7798_, not_new_n7603_, not_new_n7797_);
  not g_8748 (not_new_n9890__0, new_n9890_);
  not g_8749 (not_new_n1057__0, new_n1057_);
  not g_8750 (not_new_n1776_, new_n1776_);
  not g_8751 (not_new_n10156_, new_n10156_);
  not g_8752 (not_new_n644__57648010, new_n644_);
  not g_8753 (not_new_n6443__168070, new_n6443_);
  not g_8754 (not_new_n1043_, new_n1043_);
  or g_8755 (or_or_not_new_n2831__not_new_n1481__not_new_n2830_, not_new_n2830_, or_not_new_n2831__not_new_n1481_);
  or g_8756 (new_n2212_, not_new_n1585__138412872010, not_new_n5732_);
  or g_8757 (po215, not_new_n1417_, not_new_n1419_);
  not g_8758 (not_new_n4198_, new_n4198_);
  and g_8759 (new_n6966_, new_n7212_, new_n6962_);
  and g_8760 (new_n5857_, new_n5886_, new_n6082_);
  not g_8761 (not_new_n7406__0, new_n7406_);
  not g_8762 (not_new_n6318_, new_n6318_);
  or g_8763 (new_n7024_, not_new_n7352_, not_new_n7353_);
  not g_8764 (not_new_n5484__0, new_n5484_);
  and g_8765 (and_new_n2162__new_n2165_, new_n2162_, new_n2165_);
  not g_8766 (not_new_n1585__19773267430, new_n1585_);
  not g_8767 (not_new_n603__3430, new_n603_);
  not g_8768 (not_new_n617__6, new_n617_);
  not g_8769 (not_new_n1152_, new_n1152_);
  not g_8770 (not_new_n2287_, new_n2287_);
  or g_8771 (new_n6555_, not_new_n6926_, not_new_n6925_);
  not g_8772 (not_new_n4183_, new_n4183_);
  or g_8773 (po163, not_new_n3553_, not_new_n3552_);
  or g_8774 (new_n9446_, not_new_n9829_, not_new_n9830_);
  not g_8775 (not_new_n3311__490, new_n3311_);
  or g_8776 (new_n5193_, new_n630_, new_n1601_);
  and g_8777 (and_new_n6316__new_n6227_, new_n6316_, new_n6227_);
  not g_8778 (new_n6998_, new_n732_);
  not g_8779 (not_new_n5016_, new_n5016_);
  or g_8780 (new_n9794_, not_new_n9384__0, not_new_n1602__2326305139872070);
  or g_8781 (new_n4628_, not_new_n4521_, not_new_n4626_);
  not g_8782 (not_new_n621__7, new_n621_);
  or g_8783 (po254, not_new_n3695_, not_new_n3694_);
  or g_8784 (or_not_new_n9855__0_not_new_n10046__0, not_new_n10046__0, not_new_n9855__0);
  not g_8785 (not_new_n8003_, new_n8003_);
  not g_8786 (not_new_n1162_, new_n1162_);
  or g_8787 (new_n7560_, not_new_n735__1, not_new_n7418__1);
  not g_8788 (not_new_n1236_, new_n1236_);
  not g_8789 (not_new_n8091_, new_n8091_);
  not g_8790 (not_new_n6690_, new_n6690_);
  not g_8791 (not_new_n6084_, new_n6084_);
  not g_8792 (not_pi038_0, pi038);
  not g_8793 (not_new_n589__24010, new_n589_);
  not g_8794 (not_new_n599__2824752490, new_n599_);
  not g_8795 (not_new_n9066__0, new_n9066_);
  not g_8796 (not_new_n6974__332329305696010, new_n6974_);
  and g_8797 (new_n1288_, new_n2069_, and_and_new_n2067__new_n2070__new_n2068_);
  not g_8798 (not_new_n646__6, new_n646_);
  not g_8799 (not_pi147_1, pi147);
  and g_8800 (and_and_and_new_n6385__new_n6386__new_n6241__new_n6375_, new_n6375_, and_and_new_n6385__new_n6386__new_n6241_);
  not g_8801 (not_new_n2909_, new_n2909_);
  not g_8802 (not_new_n9123_, new_n9123_);
  not g_8803 (not_new_n2900_, new_n2900_);
  or g_8804 (new_n5288_, not_new_n5286__0, or_not_new_n5041__not_new_n4911_);
  not g_8805 (not_pi039_0, pi039);
  or g_8806 (new_n7881_, not_new_n1601__138412872010, not_new_n7627__1);
  not g_8807 (not_new_n6336_, new_n6336_);
  not g_8808 (not_new_n5051_, new_n5051_);
  or g_8809 (new_n9268_, not_new_n8969_, not_new_n8968_);
  not g_8810 (not_new_n9649_, new_n9649_);
  or g_8811 (new_n3630_, not_pi181_0, not_new_n984__403536070);
  or g_8812 (new_n8178_, not_new_n8159_, not_new_n8442_);
  not g_8813 (not_new_n643__138412872010, new_n643_);
  not g_8814 (not_new_n3225_, new_n3225_);
  not g_8815 (not_new_n6590_, new_n6590_);
  and g_8816 (new_n4292_, and_new_n4337__new_n4336_, new_n4332_);
  not g_8817 (not_new_n1198_, new_n1198_);
  not g_8818 (not_new_n1906_, new_n1906_);
  buf g_8819 (po029, pi235);
  not g_8820 (not_new_n4152_, new_n4152_);
  not g_8821 (not_new_n588__2, new_n588_);
  or g_8822 (new_n9165_, not_new_n9056__0, not_new_n8866__0);
  not g_8823 (not_new_n10292_, new_n10292_);
  not g_8824 (not_new_n718__1, new_n718_);
  not g_8825 (not_new_n8210_, new_n8210_);
  or g_8826 (new_n3694_, not_pi233, not_new_n989__403536070);
  or g_8827 (new_n10053_, new_n1047_, new_n634_);
  not g_8828 (not_new_n630__168070, new_n630_);
  and g_8829 (new_n1505_, new_n998_, new_n3030_);
  not g_8830 (not_new_n5209_, new_n5209_);
  or g_8831 (or_not_new_n4899__0_not_new_n5096__0, not_new_n5096__0, not_new_n4899__0);
  not g_8832 (not_new_n4833__0, new_n4833_);
  not g_8833 (not_new_n4992_, new_n4992_);
  not g_8834 (not_new_n8401_, new_n8401_);
  or g_8835 (new_n9553_, not_new_n9523_, not_new_n9327_);
  not g_8836 (not_new_n639__57648010, new_n639_);
  xnor g_8837 (key_gate_88, new_n596_, key_88);
  not g_8838 (not_new_n637__3430, new_n637_);
  and g_8839 (new_n1447_, and_new_n1446__new_n2659_, new_n2658_);
  not g_8840 (new_n6472_, new_n634_);
  not g_8841 (not_new_n7684_, new_n7684_);
  not g_8842 (not_new_n1057__1176490, new_n1057_);
  or g_8843 (new_n2667_, not_new_n2666_, not_new_n611__403536070);
  not g_8844 (not_new_n8850__0, new_n8850_);
  or g_8845 (new_n3665_, not_po298_5, not_new_n631__9);
  not g_8846 (not_pi180_2, pi180);
  or g_8847 (or_or_not_new_n2497__not_new_n1568__not_new_n2498_, or_not_new_n2497__not_new_n1568_, not_new_n2498_);
  and g_8848 (new_n1539_, new_n3591_, new_n3590_);
  not g_8849 (not_new_n5773__0, new_n5773_);
  not g_8850 (not_new_n5882__2, new_n5882_);
  not g_8851 (not_new_n581__8235430, new_n581_);
  not g_8852 (not_new_n6655_, new_n6655_);
  not g_8853 (not_new_n4473_, new_n4473_);
  not g_8854 (not_new_n588__10, new_n588_);
  not g_8855 (new_n1615_, new_n1569_);
  or g_8856 (new_n2222_, not_new_n1601_, not_new_n1588__968890104070);
  or g_8857 (new_n8065_, not_new_n636__138412872010, not_new_n7647__0);
  not g_8858 (not_new_n1065__3430, new_n1065_);
  not g_8859 (not_new_n1508_, new_n1508_);
  not g_8860 (not_new_n5770__2, new_n5770_);
  not g_8861 (not_new_n3358_, new_n3358_);
  not g_8862 (not_new_n1607__10, new_n1607_);
  or g_8863 (or_not_new_n2525__not_new_n2524_, not_new_n2525_, not_new_n2524_);
  or g_8864 (new_n8006_, not_new_n7746_, not_new_n7719_);
  or g_8865 (new_n1930_, not_new_n6470_, not_new_n1580__8);
  not g_8866 (not_new_n1369_, new_n1369_);
  not g_8867 (not_new_n1534__57648010, key_gate_5);
  not g_8868 (not_new_n1069__9, new_n1069_);
  or g_8869 (new_n2888_, not_new_n640__2, not_new_n604__1176490);
  not g_8870 (not_new_n1581__8235430, new_n1581_);
  not g_8871 (not_new_n4941_, new_n4941_);
  or g_8872 (new_n8474_, not_new_n8472_, not_new_n8473_);
  not g_8873 (not_new_n7451_, new_n7451_);
  or g_8874 (new_n5971_, not_new_n5925_, not_new_n5714_);
  not g_8875 (not_new_n643__16284135979104490, new_n643_);
  not g_8876 (not_new_n1037__1, new_n1037_);
  or g_8877 (new_n2446_, not_new_n597__8235430, not_new_n4791__0);
  or g_8878 (or_not_new_n6339__not_new_n6232__1, not_new_n6339_, not_new_n6232__1);
  not g_8879 (not_new_n9416_, new_n9416_);
  not g_8880 (not_new_n9174_, new_n9174_);
  not g_8881 (not_new_n7737_, new_n7737_);
  not g_8882 (not_new_n8040_, new_n8040_);
  not g_8883 (not_po298_16284135979104490, po298);
  or g_8884 (new_n6956_, not_new_n1053__168070, not_new_n6525__0);
  not g_8885 (not_new_n9778_, new_n9778_);
  not g_8886 (not_new_n3894_, new_n3894_);
  not g_8887 (not_new_n581__11044276742439206463052992010, new_n581_);
  or g_8888 (new_n5483_, not_new_n5641_, not_new_n5640_);
  or g_8889 (new_n9274_, not_new_n9273_, not_new_n9272_);
  not g_8890 (not_new_n4491__0, new_n4491_);
  not g_8891 (not_new_n3701_, new_n3701_);
  or g_8892 (new_n5492_, not_new_n5709_, not_new_n5710_);
  not g_8893 (not_new_n4437_, new_n4437_);
  and g_8894 (and_new_n2702__new_n2701_, new_n2701_, new_n2702_);
  not g_8895 (not_new_n1063__2824752490, new_n1063_);
  and g_8896 (new_n1238_, new_n1834_, new_n1835_);
  not g_8897 (not_new_n598__8235430, new_n598_);
  not g_8898 (not_new_n5918__0, new_n5918_);
  and g_8899 (new_n6584_, new_n6742_, new_n6460_);
  not g_8900 (not_new_n4536_, new_n4536_);
  not g_8901 (not_new_n7542_, new_n7542_);
  not g_8902 (not_new_n642__0, new_n642_);
  not g_8903 (not_po296_24010, po296);
  or g_8904 (or_not_new_n2919__not_new_n2922_, not_new_n2919_, not_new_n2922_);
  not g_8905 (not_new_n8953_, new_n8953_);
  not g_8906 (not_new_n2547_, new_n2547_);
  not g_8907 (not_new_n638__4, new_n638_);
  not g_8908 (not_new_n6319_, new_n6319_);
  or g_8909 (new_n3885_, not_new_n6443__16284135979104490, not_new_n626__70);
  not g_8910 (new_n8657_, new_n1161_);
  or g_8911 (new_n6685_, not_new_n6473__0, not_new_n6677_);
  not g_8912 (not_new_n7815_, new_n7815_);
  or g_8913 (new_n3880_, not_new_n644__490, not_new_n1576__47475615099430);
  or g_8914 (new_n2604_, not_new_n1002_, not_new_n607__7);
  or g_8915 (new_n6724_, not_new_n6516_, not_new_n1067__3430);
  not g_8916 (not_new_n636_, new_n636_);
  not g_8917 (not_new_n4493_, new_n4493_);
  not g_8918 (not_pi049, pi049);
  not g_8919 (not_pi227, pi227);
  not g_8920 (not_new_n7898_, new_n7898_);
  or g_8921 (new_n7182_, not_new_n7366_, not_new_n6976_);
  not g_8922 (new_n8581_, new_n8240_);
  not g_8923 (not_new_n3155_, new_n3155_);
  or g_8924 (new_n5906_, not_new_n5797_, not_new_n6071_);
  or g_8925 (new_n10198_, not_new_n10032__0, not_new_n10062_);
  and g_8926 (new_n8927_, and_new_n9168__new_n9167_, new_n9001_);
  and g_8927 (and_new_n2384__new_n2383_, new_n2384_, new_n2383_);
  not g_8928 (not_new_n638__32199057558131797268376070, new_n638_);
  not g_8929 (not_new_n589__7, new_n589_);
  not g_8930 (not_new_n5902_, new_n5902_);
  not g_8931 (new_n8113_, new_n628_);
  or g_8932 (new_n3714_, not_new_n989__113988951853731430, not_pi243);
  not g_8933 (new_n7844_, new_n7755_);
  not g_8934 (not_new_n3184__2326305139872070, new_n3184_);
  not g_8935 (not_new_n646__8, new_n646_);
  not g_8936 (not_new_n5584_, new_n5584_);
  or g_8937 (new_n5961_, not_new_n1045__490, not_new_n5754__1);
  or g_8938 (or_not_new_n2740__not_new_n2743_, not_new_n2740_, not_new_n2743_);
  or g_8939 (new_n4405_, or_not_new_n4322__0_not_new_n680__0, not_new_n679__0);
  not g_8940 (not_new_n941__0, new_n941_);
  not g_8941 (not_new_n8389_, new_n8389_);
  not g_8942 (new_n7126_, new_n753_);
  not g_8943 (not_new_n4490__0, new_n4490_);
  not g_8944 (not_new_n5974_, new_n5974_);
  not g_8945 (not_new_n1604__70, new_n1604_);
  not g_8946 (not_new_n6496__0, new_n6496_);
  or g_8947 (new_n764_, not_new_n3239_, not_new_n3238_);
  not g_8948 (not_new_n1601__8235430, new_n1601_);
  not g_8949 (not_new_n1342_, new_n1342_);
  not g_8950 (not_new_n581__657123623635342801395430, new_n581_);
  or g_8951 (new_n8295_, not_new_n8113_, not_new_n1039__19773267430);
  not g_8952 (not_pi105, pi105);
  not g_8953 (not_new_n5783_, new_n5783_);
  not g_8954 (not_new_n7270_, new_n7270_);
  not g_8955 (not_new_n8278_, new_n8278_);
  not g_8956 (not_new_n1591__19773267430, new_n1591_);
  not g_8957 (not_new_n586__47475615099430, new_n586_);
  and g_8958 (and_new_n934__new_n986_, new_n934_, new_n986_);
  not g_8959 (not_new_n1843_, new_n1843_);
  not g_8960 (not_new_n1599__1, new_n1599_);
  not g_8961 (not_new_n8372_, new_n8372_);
  not g_8962 (new_n4525_, new_n4481_);
  not g_8963 (new_n9624_, new_n9494_);
  not g_8964 (not_new_n3380_, new_n3380_);
  not g_8965 (not_new_n1585__332329305696010, new_n1585_);
  not g_8966 (new_n6149_, new_n5860_);
  or g_8967 (or_not_new_n6335__not_new_n6373__4, not_new_n6373__4, not_new_n6335_);
  not g_8968 (not_new_n8712_, new_n8712_);
  not g_8969 (not_pi269_1, pi269);
  or g_8970 (new_n655_, not_new_n3123_, or_not_new_n3124__not_new_n3125_);
  not g_8971 (not_new_n4132__2, new_n4132_);
  or g_8972 (new_n10153_, not_new_n1596__39098210485829880490, not_new_n10013__0);
  not g_8973 (not_new_n6085_, new_n6085_);
  or g_8974 (new_n626_, or_or_not_new_n1939__not_new_n1940__not_new_n1942_, not_new_n1941_);
  not g_8975 (not_new_n6674_, new_n6674_);
  or g_8976 (new_n988_, not_new_n1630_, not_new_n923_);
  not g_8977 (not_new_n642__57648010, new_n642_);
  not g_8978 (not_new_n4945__0, new_n4945_);
  not g_8979 (not_new_n5382_, new_n5382_);
  not g_8980 (not_new_n8622_, new_n8622_);
  not g_8981 (not_new_n7001__0, new_n7001_);
  not g_8982 (not_pi054_3, pi054);
  or g_8983 (new_n8586_, not_new_n8584_, not_new_n8585_);
  or g_8984 (new_n8554_, not_new_n8167__0, not_new_n646__968890104070);
  or g_8985 (new_n4851_, not_new_n4817_, not_new_n4751__0);
  not g_8986 (not_new_n5155_, new_n5155_);
  not g_8987 (new_n4267_, new_n659_);
  or g_8988 (new_n5624_, not_new_n1007__7, not_new_n5438__0);
  not g_8989 (new_n9556_, new_n9374_);
  not g_8990 (not_pi161_3, pi161);
  not g_8991 (new_n7331_, new_n7152_);
  not g_8992 (not_new_n994__6, new_n994_);
  or g_8993 (new_n4875_, not_new_n4782__0, not_new_n4834_);
  or g_8994 (po063, key_gate_107, not_new_n1190_);
  or g_8995 (new_n8033_, not_new_n7635__0, not_new_n1071__1176490);
  or g_8996 (new_n4391_, not_new_n686_, not_new_n4276_);
  or g_8997 (new_n2109_, not_new_n2104_, not_new_n1296_);
  or g_8998 (new_n2715_, not_pi245, not_new_n2703_);
  not g_8999 (not_new_n4014__0, new_n4014_);
  or g_9000 (new_n1159_, not_new_n3848_, not_new_n3847_);
  not g_9001 (not_new_n8111_, new_n8111_);
  or g_9002 (new_n2043_, not_new_n8199_, not_new_n1581__3430);
  not g_9003 (not_new_n9197_, new_n9197_);
  not g_9004 (not_new_n5766__1, new_n5766_);
  or g_9005 (new_n2513_, not_new_n606_, not_new_n5426__0);
  not g_9006 (not_new_n2761_, new_n2761_);
  not g_9007 (not_new_n8814_, new_n8814_);
  or g_9008 (new_n1645_, not_new_n596__3, key_gate_27);
  or g_9009 (new_n8917_, not_new_n9294_, not_new_n9295_);
  or g_9010 (new_n6668_, not_new_n1045__168070, not_new_n6487_);
  not g_9011 (not_new_n6647_, new_n6647_);
  not g_9012 (not_new_n9307_, new_n9307_);
  or g_9013 (or_not_new_n2227__not_new_n2224_, not_new_n2227_, not_new_n2224_);
  not g_9014 (not_new_n643__1176490, new_n643_);
  not g_9015 (not_new_n6707_, new_n6707_);
  or g_9016 (new_n1890_, not_new_n1584__5, not_new_n9433_);
  or g_9017 (new_n4659_, not_new_n4577__0, not_new_n4657_);
  or g_9018 (new_n2591_, not_new_n606__7, not_new_n5491__0);
  not g_9019 (not_new_n5922_, new_n5922_);
  not g_9020 (not_new_n8247_, new_n8247_);
  not g_9021 (not_new_n6489_, new_n6489_);
  not g_9022 (new_n9393_, new_n627_);
  not g_9023 (new_n4804_, new_n1057_);
  not g_9024 (not_new_n7225_, new_n7225_);
  or g_9025 (or_not_new_n6349__not_new_n6373__7, not_new_n6373__7, not_new_n6349_);
  not g_9026 (not_new_n4634_, new_n4634_);
  or g_9027 (new_n5129_, new_n624_, new_n1041_);
  not g_9028 (new_n9620_, new_n9416_);
  or g_9029 (or_not_new_n8411__not_new_n8293_, not_new_n8293_, not_new_n8411_);
  not g_9030 (not_new_n8155__1, new_n8155_);
  not g_9031 (not_new_n1027__797922662976120010, new_n1027_);
  not g_9032 (not_new_n1550_, new_n1550_);
  not g_9033 (not_new_n7595_, new_n7595_);
  not g_9034 (not_new_n6527__2, new_n6527_);
  or g_9035 (new_n6594_, not_new_n6884_, not_new_n6885_);
  or g_9036 (new_n5398_, not_new_n638__168070, not_new_n4957__0);
  not g_9037 (not_new_n4085_, new_n4085_);
  not g_9038 (not_new_n6327_, new_n6327_);
  not g_9039 (not_new_n7117_, new_n7117_);
  not g_9040 (not_new_n1728__1, new_n1728_);
  or g_9041 (new_n3938_, or_pi033_pi035, pi034);
  or g_9042 (new_n7012_, not_new_n721_, not_new_n7042_);
  not g_9043 (not_pi248, pi248);
  not g_9044 (not_pi010_0, pi010);
  or g_9045 (new_n2169_, not_pi119, not_new_n588__19773267430);
  not g_9046 (new_n6247_, new_n1598_);
  not g_9047 (not_new_n1517_, new_n1517_);
  not g_9048 (not_po296_152867006319425761937651857692768264010, po296);
  not g_9049 (not_po296_225393402906922580878632490, po296);
  not g_9050 (new_n4422_, new_n1007_);
  and g_9051 (new_n8210_, new_n8483_, and_new_n8112__new_n8484_);
  or g_9052 (new_n5332_, not_new_n4993__0, not_new_n618__168070);
  not g_9053 (not_new_n7618_, new_n7618_);
  not g_9054 (not_new_n10099_, new_n10099_);
  not g_9055 (not_new_n4945__2, new_n4945_);
  not g_9056 (not_new_n1538__490, new_n1538_);
  not g_9057 (not_new_n4108_, new_n4108_);
  not g_9058 (not_new_n4738_, new_n4738_);
  or g_9059 (new_n3229_, not_new_n638__7, not_new_n589__2824752490);
  not g_9060 (not_new_n635__1, new_n635_);
  not g_9061 (not_new_n9706_, new_n9706_);
  and g_9062 (and_new_n5748__new_n6116_, new_n6116_, new_n5748_);
  not g_9063 (not_new_n7902_, new_n7902_);
  and g_9064 (new_n1456_, new_n2699_, and_new_n2697__new_n2698_);
  or g_9065 (new_n6094_, not_new_n5877_, not_new_n5947_);
  not g_9066 (not_new_n4915_, new_n4915_);
  not g_9067 (not_new_n637__19773267430, new_n637_);
  or g_9068 (new_n5973_, not_new_n5791__0, not_new_n1055__490);
  not g_9069 (not_pi035_0, pi035);
  not g_9070 (not_new_n6982__0, new_n6982_);
  not g_9071 (not_new_n2786_, new_n2786_);
  and g_9072 (new_n5024_, new_n628_, new_n1039_);
  not g_9073 (not_new_n1601__113988951853731430, new_n1601_);
  or g_9074 (po061, key_gate_1, not_new_n1188_);
  or g_9075 (new_n1850_, not_new_n7687_, not_new_n1583__3);
  not g_9076 (not_new_n3859_, new_n3859_);
  or g_9077 (new_n1749_, not_pi093, not_new_n1728__8235430);
  not g_9078 (not_new_n4212_, new_n4212_);
  or g_9079 (new_n10132_, not_new_n10020_, not_new_n10131_);
  not g_9080 (not_new_n581__541169560379521116689596608490, new_n581_);
  or g_9081 (new_n3531_, not_new_n1824__0, not_new_n1612__1);
  or g_9082 (or_not_new_n2537__not_new_n2541_, not_new_n2541_, not_new_n2537_);
  not g_9083 (not_new_n601__70, new_n601_);
  or g_9084 (new_n7829_, not_new_n7647_, not_new_n636__19773267430);
  not g_9085 (not_new_n606__8, new_n606_);
  and g_9086 (po117, key_gate_101, pi096);
  not g_9087 (not_new_n595__8, new_n595_);
  not g_9088 (not_new_n5286_, new_n5286_);
  or g_9089 (new_n6566_, not_new_n6906_, not_new_n6905_);
  or g_9090 (new_n676_, or_not_new_n3103__not_new_n3102_, not_new_n3101_);
  or g_9091 (new_n9571_, new_n1051_, new_n647_);
  not g_9092 (not_new_n989__47475615099430, new_n989_);
  not g_9093 (not_new_n3851_, new_n3851_);
  not g_9094 (not_new_n8165_, new_n8165_);
  or g_9095 (new_n9629_, not_new_n9471_, not_new_n9714_);
  not g_9096 (new_n926_, pi245);
  not g_9097 (not_new_n8031_, new_n8031_);
  and g_9098 (new_n5724_, new_n5716_, new_n5984_);
  not g_9099 (not_new_n5784_, new_n5784_);
  or g_9100 (new_n2625_, not_new_n605__70, not_new_n5478_);
  not g_9101 (not_new_n589__9095436801298611408202050198891430, new_n589_);
  not g_9102 (not_new_n7001__1, new_n7001_);
  not g_9103 (new_n1611_, new_n984_);
  not g_9104 (new_n5137_, new_n5057_);
  or g_9105 (new_n6767_, not_new_n6606_, not_new_n6765_);
  not g_9106 (not_new_n2285_, new_n2285_);
  not g_9107 (not_new_n3063_, new_n3063_);
  or g_9108 (new_n4132_, not_new_n4216_, not_new_n4215_);
  not g_9109 (not_new_n637__4, new_n637_);
  not g_9110 (not_new_n6981_, new_n6981_);
  not g_9111 (not_new_n7021_, new_n7021_);
  and g_9112 (and_new_n7161__new_n7474_, new_n7161_, new_n7474_);
  xnor g_9113 (key_gate_28, not_new_n1182_, key_28);
  not g_9114 (not_new_n4831__0, new_n4831_);
  not g_9115 (not_new_n6507__0, new_n6507_);
  or g_9116 (new_n3110_, not_new_n632__5, not_new_n3315__8);
  not g_9117 (not_new_n8948_, new_n8948_);
  and g_9118 (new_n1385_, new_n2448_, new_n2447_);
  or g_9119 (new_n3267_, not_new_n1600__5, not_new_n589__32199057558131797268376070);
  not g_9120 (not_new_n9384_, new_n9384_);
  not g_9121 (not_new_n775__2326305139872070, new_n775_);
  not g_9122 (not_new_n4423_, new_n4423_);
  not g_9123 (not_new_n7145_, new_n7145_);
  not g_9124 (new_n7639_, new_n646_);
  not g_9125 (not_new_n3986_, new_n3986_);
  not g_9126 (not_new_n648__113988951853731430, new_n648_);
  or g_9127 (new_n2599_, not_po296_225393402906922580878632490, not_pi270);
  not g_9128 (not_new_n8887_, new_n8887_);
  not g_9129 (new_n7327_, new_n7113_);
  not g_9130 (not_new_n9581_, new_n9581_);
  or g_9131 (new_n7920_, not_new_n7668_, not_new_n7858_);
  not g_9132 (not_new_n3102_, new_n3102_);
  not g_9133 (not_new_n9309_, new_n9309_);
  not g_9134 (not_new_n3967_, new_n3967_);
  not g_9135 (new_n9105_, new_n8963_);
  not g_9136 (not_new_n1730_, new_n1730_);
  not g_9137 (not_new_n7323_, new_n7323_);
  not g_9138 (not_new_n626__3, new_n626_);
  and g_9139 (new_n1263_, and_new_n1262__new_n1951_, new_n1950_);
  not g_9140 (not_new_n4985_, new_n4985_);
  not g_9141 (not_new_n3812_, new_n3812_);
  not g_9142 (not_new_n3185__8235430, new_n3185_);
  or g_9143 (new_n7615_, not_new_n7790_, not_new_n7792_);
  not g_9144 (not_new_n2066_, new_n2066_);
  not g_9145 (not_new_n1612__2824752490, new_n1612_);
  not g_9146 (not_pi139_0, pi139);
  not g_9147 (not_new_n3185__0, new_n3185_);
  or g_9148 (new_n9806_, not_new_n9658_, not_new_n9499_);
  not g_9149 (not_new_n8895_, new_n8895_);
  or g_9150 (new_n8339_, not_new_n1055__47475615099430, not_new_n8155__0);
  not g_9151 (not_new_n994__24010, new_n994_);
  or g_9152 (new_n7511_, not_new_n7144_, not_new_n7145_);
  and g_9153 (new_n1221_, new_n1219_, and_and_new_n1217__new_n1218__new_n1220_);
  and g_9154 (new_n6588_, new_n6865_, new_n6750_);
  not g_9155 (not_new_n8228_, new_n8228_);
  not g_9156 (not_new_n1582_, new_n1582_);
  not g_9157 (not_new_n5437_, new_n5437_);
  xnor g_9158 (key_gate_101, key_101, new_n1535_);
  not g_9159 (not_new_n5077_, new_n5077_);
  not g_9160 (not_new_n7237_, new_n7237_);
  or g_9161 (new_n5677_, or_not_new_n5466__not_new_n5674__1, not_new_n5673_);
  not g_9162 (not_new_n6658__0, new_n6658_);
  not g_9163 (not_new_n5083_, new_n5083_);
  and g_9164 (and_and_new_n2105__new_n2108__new_n2106_, new_n2106_, and_new_n2105__new_n2108_);
  or g_9165 (or_not_new_n9719__not_new_n9718_, not_new_n9719_, not_new_n9718_);
  not g_9166 (not_new_n1014__0, new_n1014_);
  not g_9167 (not_new_n6536_, new_n6536_);
  not g_9168 (not_new_n4423__0, new_n4423_);
  or g_9169 (new_n7341_, not_new_n6974__0, not_new_n770_);
  not g_9170 (not_new_n1865_, new_n1865_);
  or g_9171 (or_or_not_new_n934__not_new_n933__0_not_new_n941__0, not_new_n941__0, or_not_new_n934__not_new_n933__0);
  not g_9172 (not_new_n629__332329305696010, new_n629_);
  and g_9173 (new_n6443_, new_n623_, new_n6444_);
  not g_9174 (not_new_n3372_, new_n3372_);
  or g_9175 (new_n4715_, not_new_n4713_, not_new_n4545_);
  or g_9176 (new_n10084_, not_new_n10265_, or_or_not_new_n9893__not_new_n9890__0_not_new_n10266_);
  and g_9177 (new_n1418_, new_n2519_, new_n2522_);
  not g_9178 (new_n9379_, new_n1598_);
  not g_9179 (not_new_n8548_, new_n8548_);
  or g_9180 (new_n5411_, not_new_n1059__70, not_new_n4968_);
  not g_9181 (not_new_n9474_, new_n9474_);
  or g_9182 (new_n3341_, not_new_n1534__490, not_pi034_0);
  not g_9183 (not_new_n4420_, new_n4420_);
  not g_9184 (not_new_n1631__2, key_gate_76);
  or g_9185 (new_n7544_, not_new_n7151_, not_new_n7152__0);
  not g_9186 (not_pi162_3, pi162);
  not g_9187 (not_new_n5650_, new_n5650_);
  not g_9188 (not_new_n4360_, new_n4360_);
  not g_9189 (not_pi166, pi166);
  not g_9190 (new_n4718_, new_n623_);
  not g_9191 (not_new_n1583__4, new_n1583_);
  not g_9192 (new_n5460_, new_n1016_);
  not g_9193 (not_new_n4066_, new_n4066_);
  not g_9194 (not_new_n1035__1, new_n1035_);
  not g_9195 (not_po296_205005145156954906122290109080958673914396262484637238056070, po296);
  not g_9196 (not_new_n585__9, new_n585_);
  not g_9197 (not_new_n1059__1176490, new_n1059_);
  or g_9198 (new_n8329_, not_new_n8106__1, not_new_n631__797922662976120010);
  not g_9199 (not_new_n3154_, new_n3154_);
  not g_9200 (not_new_n1886_, new_n1886_);
  not g_9201 (not_new_n1602__1, new_n1602_);
  not g_9202 (not_new_n9854_, new_n9854_);
  not g_9203 (not_new_n8848_, new_n8848_);
  or g_9204 (new_n5618_, not_pi134_3, not_new_n5440__1);
  not g_9205 (not_new_n1427_, new_n1427_);
  not g_9206 (not_new_n1603__1176490, new_n1603_);
  not g_9207 (not_new_n5937_, new_n5937_);
  not g_9208 (not_new_n6943_, new_n6943_);
  not g_9209 (not_new_n5217_, new_n5217_);
  not g_9210 (not_new_n3922__0, new_n3922_);
  not g_9211 (not_new_n7635_, new_n7635_);
  not g_9212 (not_pi029_0, pi029);
  or g_9213 (new_n4539_, not_new_n4538_, not_new_n4475_);
  not g_9214 (not_new_n7471_, new_n7471_);
  not g_9215 (not_new_n8102_, new_n8102_);
  not g_9216 (not_new_n7888_, new_n7888_);
  or g_9217 (new_n7449_, not_new_n775__47475615099430, not_new_n7131_);
  not g_9218 (not_new_n5469_, new_n5469_);
  or g_9219 (new_n2918_, not_new_n2915_, or_not_new_n2917__not_new_n2916_);
  not g_9220 (not_new_n8198_, new_n8198_);
  not g_9221 (not_new_n4924_, new_n4924_);
  not g_9222 (new_n7122_, new_n759_);
  not g_9223 (not_new_n8157_, new_n8157_);
  not g_9224 (not_new_n8110__0, new_n8110_);
  and g_9225 (and_and_new_n6395__new_n6396__new_n6228_, new_n6228_, and_new_n6395__new_n6396_);
  not g_9226 (not_new_n628__403536070, new_n628_);
  not g_9227 (not_new_n2723_, new_n2723_);
  not g_9228 (not_new_n1536__24010, new_n1536_);
  or g_9229 (new_n9764_, not_new_n9633_, not_new_n9762_);
  or g_9230 (new_n8903_, not_new_n9195_, not_new_n9196_);
  not g_9231 (not_pi136_2, pi136);
  not g_9232 (not_new_n630__9, new_n630_);
  or g_9233 (new_n4660_, not_new_n1012__3, not_new_n4447_);
  and g_9234 (new_n1305_, new_n2155_, new_n2156_);
  or g_9235 (new_n9497_, not_new_n9708_, not_new_n9706_);
  not g_9236 (not_new_n9520__0, new_n9520_);
  not g_9237 (not_pi019_0, pi019);
  not g_9238 (not_new_n6387_, new_n6387_);
  not g_9239 (not_new_n9370_, new_n9370_);
  or g_9240 (new_n9216_, not_new_n628__5585458640832840070, not_new_n8823_);
  or g_9241 (new_n2418_, not_new_n600__490, not_new_n4134__0);
  not g_9242 (new_n1580_, new_n934_);
  not g_9243 (not_new_n624__490, new_n624_);
  not g_9244 (not_new_n4437__0, new_n4437_);
  or g_9245 (new_n7190_, not_new_n7189_, not_new_n6990_);
  not g_9246 (not_new_n3793_, new_n3793_);
  not g_9247 (not_new_n9007_, new_n9007_);
  not g_9248 (new_n6076_, new_n5882_);
  not g_9249 (not_new_n1065__1, new_n1065_);
  or g_9250 (new_n8452_, not_new_n8285__0, not_new_n8127__0);
  or g_9251 (new_n6180_, not_new_n5778__0, not_new_n1071__70);
  not g_9252 (not_new_n8779__0, new_n8779_);
  not g_9253 (not_new_n3997__0, new_n3997_);
  not g_9254 (not_new_n743__0, new_n743_);
  not g_9255 (not_new_n588__70, new_n588_);
  or g_9256 (new_n5531_, not_new_n5502_, not_new_n5530_);
  not g_9257 (new_n7603_, new_n1049_);
  not g_9258 (not_new_n3847_, new_n3847_);
  not g_9259 (not_new_n9413__0, new_n9413_);
  not g_9260 (not_new_n7159__0, new_n7159_);
  not g_9261 (not_pi175_1, pi175);
  or g_9262 (or_not_new_n1470__not_new_n3824_, not_new_n1470_, not_new_n3824_);
  not g_9263 (not_new_n8163__0, new_n8163_);
  not g_9264 (not_new_n4174_, new_n4174_);
  not g_9265 (new_n7460_, new_n7087_);
  or g_9266 (new_n9762_, not_new_n9760_, not_new_n9761_);
  or g_9267 (new_n7872_, not_new_n7666__0, not_new_n7771_);
  or g_9268 (po159, not_new_n3545_, not_new_n3544_);
  not g_9269 (not_new_n9776_, new_n9776_);
  or g_9270 (new_n10282_, not_new_n9944_, not_new_n1597__5585458640832840070);
  not g_9271 (not_new_n725__0, new_n725_);
  not g_9272 (not_new_n4001__0, new_n4001_);
  not g_9273 (not_new_n8151__0, new_n8151_);
  not g_9274 (not_new_n1958_, new_n1958_);
  not g_9275 (not_new_n7537_, new_n7537_);
  or g_9276 (new_n5900_, not_new_n6087_, not_new_n6043_);
  not g_9277 (not_new_n6635__0, new_n6635_);
  or g_9278 (new_n7332_, not_new_n7098_, not_new_n775__0);
  not g_9279 (not_new_n595__6782230728490, new_n595_);
  or g_9280 (new_n4192_, not_new_n4112_, not_new_n4174__0);
  not g_9281 (not_new_n2597_, new_n2597_);
  not g_9282 (not_new_n8559_, new_n8559_);
  or g_9283 (or_not_new_n3130__not_new_n3131_, not_new_n3130_, not_new_n3131_);
  not g_9284 (not_new_n7755_, new_n7755_);
  not g_9285 (not_new_n7819_, new_n7819_);
  or g_9286 (new_n5517_, not_new_n5553_, not_new_n5552_);
  not g_9287 (not_new_n6692_, new_n6692_);
  or g_9288 (new_n9095_, not_new_n1601__16284135979104490, not_new_n630__6782230728490);
  not g_9289 (not_new_n1588__8, new_n1588_);
  not g_9290 (not_new_n1495_, new_n1495_);
  not g_9291 (not_new_n588__138412872010, new_n588_);
  or g_9292 (new_n5195_, not_new_n1601__8, not_new_n630__3430);
  or g_9293 (new_n7456_, not_new_n750_, not_new_n6974__332329305696010);
  not g_9294 (not_new_n7047_, new_n7047_);
  not g_9295 (not_new_n3294_, new_n3294_);
  not g_9296 (not_new_n1588__797922662976120010, new_n1588_);
  or g_9297 (new_n7751_, not_new_n7923_, not_new_n7637_);
  not g_9298 (not_new_n8408_, new_n8408_);
  not g_9299 (not_new_n4781_, new_n4781_);
  not g_9300 (not_new_n601__4, new_n601_);
  or g_9301 (or_not_new_n1335__not_new_n1333_, not_new_n1333_, not_new_n1335_);
  not g_9302 (not_new_n9709_, new_n9709_);
  not g_9303 (not_new_n636__490, new_n636_);
  not g_9304 (not_new_n626__113988951853731430, new_n626_);
  not g_9305 (new_n4001_, new_n3935_);
  not g_9306 (not_new_n2459_, new_n2459_);
  or g_9307 (new_n7516_, not_new_n7146__1, not_new_n7306_);
  not g_9308 (not_new_n1600__138412872010, new_n1600_);
  or g_9309 (new_n5663_, not_new_n5661_, not_new_n5662_);
  not g_9310 (not_new_n7259_, new_n7259_);
  and g_9311 (new_n5876_, new_n6218_, new_n5915_);
  and g_9312 (new_n10002_, and_new_n10033__new_n3902_, new_n3903_);
  or g_9313 (new_n669_, or_not_new_n3170__not_new_n3169_, not_new_n3168_);
  or g_9314 (new_n5125_, not_new_n5095_, not_new_n4899_);
  not g_9315 (not_new_n7923_, new_n7923_);
  not g_9316 (not_new_n9113_, new_n9113_);
  not g_9317 (not_new_n978_, new_n978_);
  or g_9318 (new_n8253_, not_new_n8218_, not_new_n8376_);
  or g_9319 (po246, not_new_n3679_, not_new_n3678_);
  not g_9320 (not_new_n6443__968890104070, new_n6443_);
  and g_9321 (and_new_n5740__new_n6096_, new_n5740_, new_n6096_);
  not g_9322 (not_new_n628__19773267430, new_n628_);
  not g_9323 (not_new_n8894__0, new_n8894_);
  not g_9324 (not_new_n984_, new_n984_);
  not g_9325 (not_new_n4769__0, new_n4769_);
  or g_9326 (new_n2477_, not_new_n603__6782230728490, not_new_n621__1);
  or g_9327 (new_n7255_, not_new_n7164_, not_new_n6965_);
  not g_9328 (not_new_n8432_, new_n8432_);
  or g_9329 (new_n8298_, not_new_n8279_, not_new_n628__332329305696010);
  and g_9330 (new_n7083_, new_n7160_, new_n7238_);
  or g_9331 (po217, or_or_not_new_n2537__not_new_n2541__not_new_n1423_, not_new_n1422_);
  not g_9332 (not_new_n3908_, new_n3908_);
  not g_9333 (new_n8114_, new_n1037_);
  not g_9334 (not_new_n4202_, new_n4202_);
  not g_9335 (not_new_n9887_, new_n9887_);
  not g_9336 (not_new_n9735_, new_n9735_);
  not g_9337 (not_new_n596__6782230728490, key_gate_88);
  not g_9338 (not_new_n6454_, new_n6454_);
  not g_9339 (not_new_n6551_, new_n6551_);
  not g_9340 (new_n6303_, new_n1596_);
  or g_9341 (new_n7999_, not_new_n7621__0, not_new_n621__138412872010);
  not g_9342 (not_new_n1598__6, new_n1598_);
  not g_9343 (not_new_n7800_, new_n7800_);
  or g_9344 (new_n2348_, or_not_new_n2346__not_new_n2347_, not_new_n1569__0);
  not g_9345 (not_pi250_4, pi250);
  not g_9346 (not_new_n3527_, new_n3527_);
  and g_9347 (new_n1316_, and_and_new_n2200__new_n2203__new_n2201_, new_n2202_);
  not g_9348 (not_new_n8709__0, new_n8709_);
  not g_9349 (not_new_n9502_, new_n9502_);
  not g_9350 (not_new_n6524_, new_n6524_);
  not g_9351 (not_new_n1580__113988951853731430, new_n1580_);
  or g_9352 (new_n3903_, not_new_n9927_, not_new_n644__3430);
  not g_9353 (not_new_n10251_, new_n10251_);
  or g_9354 (new_n5266_, not_new_n1596__9, not_new_n618__3430);
  and g_9355 (new_n3967_, not_pi038_2, and_and_not_pi037_2_not_pi036_2_not_pi039_3);
  and g_9356 (po099, key_gate_101, pi078);
  not g_9357 (not_new_n5529_, new_n5529_);
  not g_9358 (new_n8654_, new_n1605_);
  not g_9359 (new_n4948_, new_n1597_);
  not g_9360 (not_new_n586__8, new_n586_);
  or g_9361 (new_n6921_, not_new_n6603_, not_new_n6635__5);
  or g_9362 (new_n1940_, not_new_n587__9, not_pi139);
  or g_9363 (or_not_new_n4933__not_new_n4930__0, not_new_n4930__0, not_new_n4933_);
  not g_9364 (not_new_n5525_, new_n5525_);
  not g_9365 (not_new_n989__0, new_n989_);
  or g_9366 (or_or_not_new_n2803__not_new_n2806__not_new_n2805_, not_new_n2805_, or_not_new_n2803__not_new_n2806_);
  or g_9367 (new_n9500_, not_new_n9358_, not_new_n9657_);
  not g_9368 (not_new_n10188_, new_n10188_);
  not g_9369 (not_new_n9131_, new_n9131_);
  not g_9370 (new_n5433_, pi131);
  not g_9371 (not_new_n7469_, new_n7469_);
  or g_9372 (new_n4216_, not_new_n4162_, not_new_n4087_);
  not g_9373 (not_new_n605__1176490, new_n605_);
  not g_9374 (not_new_n1417_, new_n1417_);
  not g_9375 (not_new_n10310_, new_n10310_);
  not g_9376 (not_new_n3163_, new_n3163_);
  not g_9377 (not_new_n4482_, new_n4482_);
  or g_9378 (new_n5673_, not_pi144_2, not_new_n5465__0);
  not g_9379 (not_pi064_8235430, pi064);
  or g_9380 (new_n4603_, not_new_n4427__0, not_new_n1004__4);
  not g_9381 (not_new_n8078_, new_n8078_);
  xnor g_9382 (key_gate_90, not_po296, key_90);
  or g_9383 (new_n4129_, not_new_n4210_, not_new_n4209_);
  not g_9384 (not_pi150, pi150);
  not g_9385 (new_n7106_, new_n769_);
  not g_9386 (not_new_n4425_, new_n4425_);
  or g_9387 (new_n2140_, not_new_n1591__57648010, not_new_n8915_);
  not g_9388 (not_pi055_0, pi055);
  or g_9389 (new_n3936_, not_new_n4001_, not_new_n3962_);
  not g_9390 (not_new_n7062_, new_n7062_);
  not g_9391 (not_new_n1604__8, new_n1604_);
  not g_9392 (not_new_n8962_, new_n8962_);
  not g_9393 (not_new_n6255_, new_n6255_);
  not g_9394 (not_new_n6617__0, new_n6617_);
  not g_9395 (not_new_n630__3430, new_n630_);
  and g_9396 (new_n10017_, new_n10301_, new_n10300_);
  or g_9397 (new_n3686_, not_pi229, not_new_n989__168070);
  not g_9398 (not_pi079, pi079);
  or g_9399 (or_or_not_new_n2265__not_new_n2262__not_new_n2263_, or_not_new_n2265__not_new_n2262_, not_new_n2263_);
  not g_9400 (new_n5086_, new_n4978_);
  and g_9401 (new_n6231_, and_and_new_n6369__new_n6320__new_n6230_, new_n6408_);
  not g_9402 (new_n6285_, new_n1051_);
  or g_9403 (new_n8874_, not_new_n1071__2824752490, not_new_n645__6782230728490);
  not g_9404 (not_new_n4415__1, new_n4415_);
  not g_9405 (not_new_n9972_, new_n9972_);
  and g_9406 (new_n1192_, new_n1667_, new_n1665_);
  not g_9407 (not_new_n601__47475615099430, new_n601_);
  not g_9408 (not_new_n638__657123623635342801395430, new_n638_);
  and g_9409 (and_and_new_n6374__new_n6372__new_n6371_, new_n6371_, and_new_n6374__new_n6372_);
  not g_9410 (not_new_n5765_, new_n5765_);
  not g_9411 (not_pi236, pi236);
  or g_9412 (new_n3294_, not_new_n3184__968890104070, not_new_n636__8);
  not g_9413 (not_new_n7093_, new_n7093_);
  or g_9414 (new_n1039_, not_new_n3418_, not_new_n3417_);
  or g_9415 (or_not_new_n2820__not_new_n2823_, not_new_n2820_, not_new_n2823_);
  or g_9416 (new_n6220_, not_new_n5794__2, not_new_n626__2824752490);
  or g_9417 (new_n8745_, not_new_n8744_, not_new_n8743_);
  or g_9418 (new_n2093_, not_pi115, not_new_n588__8235430);
  not g_9419 (not_new_n7827_, new_n7827_);
  or g_9420 (new_n2760_, not_new_n2757_, not_new_n1616__2);
  not g_9421 (not_new_n1596__490, new_n1596_);
  not g_9422 (not_new_n1901_, new_n1901_);
  not g_9423 (not_new_n2554_, new_n2554_);
  not g_9424 (not_new_n5063__0, new_n5063_);
  not g_9425 (not_new_n1035__3430, new_n1035_);
  or g_9426 (new_n2929_, not_new_n3310__3430, not_new_n4128__2);
  not g_9427 (not_new_n8042_, new_n8042_);
  not g_9428 (not_new_n622_, new_n622_);
  and g_9429 (new_n5851_, new_n6005_, new_n5728_);
  not g_9430 (not_pi074, pi074);
  or g_9431 (or_not_new_n1977__not_new_n1978_, not_new_n1978_, not_new_n1977_);
  not g_9432 (not_new_n1598__4, new_n1598_);
  not g_9433 (not_new_n4780__1, new_n4780_);
  not g_9434 (not_pi172_1, pi172);
  not g_9435 (new_n8283_, new_n8176_);
  or g_9436 (po199, or_or_not_new_n1556__not_new_n2439__not_new_n1381_, not_new_n1382_);
  not g_9437 (not_new_n596__2, key_gate_88);
  or g_9438 (new_n3316_, not_pi057_0, not_new_n1534__1);
  not g_9439 (not_new_n8974_, new_n8974_);
  or g_9440 (new_n7486_, not_new_n7041__0, not_new_n7009__0);
  not g_9441 (not_new_n5465__1, new_n5465_);
  not g_9442 (not_new_n5723_, new_n5723_);
  or g_9443 (new_n3643_, not_new_n976_, not_new_n1611__47475615099430);
  and g_9444 (and_new_n1262__new_n1951_, new_n1951_, new_n1262_);
  or g_9445 (new_n7826_, not_new_n7648__0, not_new_n1055__19773267430);
  not g_9446 (not_new_n9974_, new_n9974_);
  or g_9447 (new_n9262_, not_new_n9260_, not_new_n9092__0);
  not g_9448 (not_new_n9658_, new_n9658_);
  not g_9449 (new_n5575_, new_n5511_);
  not g_9450 (not_new_n9258_, new_n9258_);
  not g_9451 (not_new_n585__332329305696010, new_n585_);
  or g_9452 (new_n2356_, not_new_n1031__3, not_new_n597_);
  not g_9453 (new_n8821_, new_n1037_);
  or g_9454 (new_n6904_, not_new_n6509__0, not_new_n639__2824752490);
  not g_9455 (not_new_n648__8, new_n648_);
  not g_9456 (not_new_n5235_, new_n5235_);
  not g_9457 (not_new_n6989_, new_n6989_);
  or g_9458 (new_n8402_, not_new_n8158__0, not_new_n626__5585458640832840070);
  or g_9459 (new_n5156_, new_n627_, new_n1055_);
  not g_9460 (not_new_n8893__0, new_n8893_);
  not g_9461 (new_n4441_, pi175);
  not g_9462 (not_new_n638__9, new_n638_);
  not g_9463 (not_new_n1055__70, new_n1055_);
  not g_9464 (not_pi033_1, pi033);
  or g_9465 (new_n6897_, or_not_new_n6508__1_not_new_n6600_, not_new_n6808_);
  not g_9466 (not_new_n3526_, new_n3526_);
  not g_9467 (not_new_n2148_, new_n2148_);
  not g_9468 (not_new_n7337_, new_n7337_);
  not g_9469 (not_new_n9918_, new_n9918_);
  or g_9470 (po236, not_new_n3658_, not_new_n3659_);
  not g_9471 (not_new_n1039__24010, new_n1039_);
  or g_9472 (new_n8013_, not_new_n7630__0, not_new_n630__19773267430);
  not g_9473 (not_new_n994__3, new_n994_);
  or g_9474 (new_n4800_, not_new_n4802__0, not_new_n4827__0);
  not g_9475 (not_new_n984__8, new_n984_);
  not g_9476 (not_new_n7095_, new_n7095_);
  or g_9477 (po162, not_new_n3550_, not_new_n3551_);
  not g_9478 (new_n10035_, new_n9926_);
  not g_9479 (not_pi261, pi261);
  not g_9480 (new_n7124_, new_n758_);
  not g_9481 (not_new_n8932_, new_n8932_);
  not g_9482 (not_new_n727__0, new_n727_);
  not g_9483 (new_n8611_, new_n1065_);
  not g_9484 (not_new_n8024_, new_n8024_);
  not g_9485 (not_new_n1596__70, new_n1596_);
  or g_9486 (new_n8791_, not_new_n8596__3, not_new_n8625_);
  or g_9487 (new_n2457_, not_new_n603__2824752490, not_new_n625__1);
  not g_9488 (new_n8637_, new_n1178_);
  not g_9489 (not_new_n1039__0, new_n1039_);
  not g_9490 (not_new_n5925_, new_n5925_);
  or g_9491 (new_n9549_, new_n1045_, new_n635_);
  not g_9492 (not_new_n1420_, new_n1420_);
  or g_9493 (new_n8972_, not_new_n8830_, not_new_n9129_);
  not g_9494 (not_new_n4972_, new_n4972_);
  or g_9495 (new_n8468_, not_new_n8103__0, not_new_n1047__57648010);
  not g_9496 (new_n3315_, new_n998_);
  not g_9497 (not_new_n6851_, new_n6851_);
  not g_9498 (not_new_n9469_, new_n9469_);
  or g_9499 (new_n8416_, not_new_n8307_, not_new_n8084_);
  not g_9500 (not_new_n1384_, new_n1384_);
  or g_9501 (new_n8382_, not_new_n618__332329305696010, not_new_n8171_);
  not g_9502 (not_new_n5709_, new_n5709_);
  not g_9503 (not_new_n6570_, new_n6570_);
  not g_9504 (not_new_n8075_, new_n8075_);
  not g_9505 (not_new_n4770__1, new_n4770_);
  not g_9506 (not_new_n1728__8, new_n1728_);
  or g_9507 (new_n7790_, not_new_n7789_, not_new_n7570_);
  not g_9508 (not_new_n1053__1176490, new_n1053_);
  or g_9509 (new_n2680_, not_new_n608__1176490, not_new_n1009__0);
  not g_9510 (not_pi274, pi274);
  not g_9511 (not_new_n7946_, new_n7946_);
  or g_9512 (or_not_new_n2587__not_new_n2591_, not_new_n2591_, not_new_n2587_);
  not g_9513 (not_new_n1055__2326305139872070, new_n1055_);
  and g_9514 (new_n4774_, new_n4867_, new_n4866_);
  or g_9515 (new_n2961_, not_new_n602__47475615099430, not_new_n638__3);
  and g_9516 (and_new_n9189__new_n9187_, new_n9187_, new_n9189_);
  not g_9517 (not_new_n624__6782230728490, new_n624_);
  not g_9518 (not_new_n4937__0, new_n4937_);
  not g_9519 (not_new_n9834_, new_n9834_);
  or g_9520 (new_n3520_, not_new_n1537__16284135979104490, not_pi126_0);
  not g_9521 (not_new_n8585_, new_n8585_);
  or g_9522 (new_n4560_, not_new_n1016__2, not_pi174_1);
  or g_9523 (new_n8483_, not_new_n1039__138412872010, not_new_n8113__1);
  not g_9524 (new_n8291_, new_n8159_);
  not g_9525 (new_n4958_, new_n638_);
  not g_9526 (not_new_n1020__0, new_n1020_);
  and g_9527 (and_new_n8789__new_n8784_, new_n8784_, new_n8789_);
  or g_9528 (new_n2462_, not_new_n603__19773267430, not_new_n630__1);
  and g_9529 (new_n6225_, new_n6391_, and_and_new_n6388__new_n6313__new_n6224_);
  or g_9530 (new_n1640_, not_pi035, not_new_n1631__1);
  not g_9531 (not_new_n7037__0, new_n7037_);
  not g_9532 (not_new_n6523_, new_n6523_);
  or g_9533 (po185, not_new_n1353_, not_new_n1354_);
  not g_9534 (not_new_n9412__0, new_n9412_);
  not g_9535 (not_new_n9865_, new_n9865_);
  not g_9536 (not_new_n648__2824752490, new_n648_);
  not g_9537 (not_new_n1604__57648010, new_n1604_);
  not g_9538 (not_pi179_2, pi179);
  and g_9539 (new_n7762_, new_n8072_, new_n8073_);
  or g_9540 (new_n2003_, not_new_n1585__70, not_new_n5825_);
  not g_9541 (not_new_n5273_, new_n5273_);
  not g_9542 (not_new_n10108_, new_n10108_);
  not g_9543 (not_pi056, pi056);
  or g_9544 (new_n9033_, not_new_n1043__19773267430, not_new_n631__273687473400809163430);
  or g_9545 (new_n2964_, not_new_n1061__1, not_new_n3311__8235430);
  not g_9546 (not_new_n3311__7, new_n3311_);
  or g_9547 (new_n3463_, not_new_n1017__1, not_new_n1594__70);
  or g_9548 (new_n7694_, not_new_n8074_, not_new_n8075_);
  or g_9549 (new_n6033_, not_new_n626__57648010, not_new_n5794__0);
  not g_9550 (not_new_n1591__70, new_n1591_);
  not g_9551 (not_new_n1534__8, key_gate_5);
  or g_9552 (new_n705_, not_new_n2997_, not_new_n1489_);
  or g_9553 (new_n10167_, not_new_n10166_, not_new_n9997_);
  not g_9554 (not_new_n8839_, new_n8839_);
  or g_9555 (new_n6835_, not_new_n6479__1, not_new_n648__19773267430);
  not g_9556 (not_new_n586__332329305696010, new_n586_);
  or g_9557 (new_n4744_, not_new_n4780_, or_not_new_n4835__not_new_n4777_);
  not g_9558 (not_new_n9328_, new_n9328_);
  not g_9559 (not_new_n3977__0, key_gate_37);
  or g_9560 (new_n4589_, not_new_n4432__0, not_new_n1002__4);
  not g_9561 (not_new_n1037__6, new_n1037_);
  not g_9562 (new_n8641_, new_n1172_);
  and g_9563 (new_n5501_, new_n5623_, new_n5622_);
  not g_9564 (not_new_n595__490, new_n595_);
  or g_9565 (new_n5676_, not_new_n5675_, not_new_n5674__0);
  or g_9566 (new_n1010_, not_new_n3341_, not_new_n3342_);
  or g_9567 (new_n6442_, not_new_n6370__1, not_new_n6306_);
  and g_9568 (new_n9331_, new_n9596_, new_n9595_);
  or g_9569 (new_n7839_, not_new_n7580_, not_new_n7759_);
  or g_9570 (new_n4089_, not_new_n4161_, not_new_n4141_);
  or g_9571 (new_n1830_, not_new_n632__0, not_new_n601__1);
  or g_9572 (new_n4617_, not_new_n4423__0, not_new_n1006__4);
  not g_9573 (not_new_n5965_, new_n5965_);
  not g_9574 (not_new_n7908_, new_n7908_);
  not g_9575 (not_new_n8129_, new_n8129_);
  or g_9576 (new_n6218_, not_new_n6217_, not_new_n6216_);
  or g_9577 (new_n7236_, not_new_n7439_, not_new_n7004_);
  not g_9578 (not_new_n4378_, new_n4378_);
  not g_9579 (not_new_n7165_, new_n7165_);
  not g_9580 (not_new_n2762_, new_n2762_);
  not g_9581 (not_new_n10033__0, new_n10033_);
  or g_9582 (new_n5431_, not_new_n1020__6, not_pi129_2);
  not g_9583 (not_new_n994__113988951853731430, new_n994_);
  not g_9584 (not_new_n596__9, key_gate_88);
  not g_9585 (not_new_n7548_, new_n7548_);
  or g_9586 (new_n3205_, not_new_n621__7, not_new_n589__8);
  not g_9587 (not_new_n644__968890104070, new_n644_);
  not g_9588 (not_new_n581__403536070, new_n581_);
  or g_9589 (new_n9739_, not_new_n9353_, not_new_n624__2326305139872070);
  not g_9590 (not_new_n1065__797922662976120010, new_n1065_);
  not g_9591 (not_new_n3990_, new_n3990_);
  not g_9592 (not_new_n8898__0, new_n8898_);
  not g_9593 (not_new_n8960_, new_n8960_);
  not g_9594 (not_new_n6164_, new_n6164_);
  not g_9595 (not_new_n1584__490, new_n1584_);
  not g_9596 (not_new_n626__0, new_n626_);
  or g_9597 (new_n5474_, not_new_n5577_, not_new_n5578_);
  not g_9598 (not_new_n7366_, new_n7366_);
  not g_9599 (not_new_n603__2326305139872070, new_n603_);
  not g_9600 (not_new_n1047__2, new_n1047_);
  not g_9601 (not_new_n8093_, new_n8093_);
  not g_9602 (not_new_n1599__24010, new_n1599_);
  or g_9603 (new_n8475_, not_new_n8119__0, not_new_n1043__57648010);
  not g_9604 (not_new_n599__5, new_n599_);
  not g_9605 (not_new_n5854_, new_n5854_);
  or g_9606 (new_n2694_, not_new_n607__1176490, not_new_n1020_);
  or g_9607 (new_n2023_, not_new_n1584__490, not_new_n9341_);
  not g_9608 (not_new_n6675_, new_n6675_);
  not g_9609 (not_new_n1728__2326305139872070, new_n1728_);
  or g_9610 (new_n9962_, not_new_n10287_, not_new_n10286_);
  not g_9611 (not_new_n588__113988951853731430, new_n588_);
  not g_9612 (not_new_n8018_, new_n8018_);
  not g_9613 (not_new_n6746_, new_n6746_);
  or g_9614 (new_n7187_, not_new_n6975_, not_new_n7357_);
  not g_9615 (not_new_n1151__0, new_n1151_);
  not g_9616 (not_new_n634__797922662976120010, new_n634_);
  not g_9617 (not_new_n9047_, new_n9047_);
  not g_9618 (not_new_n8657_, new_n8657_);
  not g_9619 (not_new_n1589__7, new_n1589_);
  not g_9620 (not_new_n1019_, new_n1019_);
  or g_9621 (new_n3351_, not_pi047_0, not_new_n1534__8235430);
  or g_9622 (new_n3288_, not_new_n638__8, not_new_n3184__2824752490);
  or g_9623 (new_n2938_, not_new_n3310__24010, not_new_n4071__2);
  not g_9624 (not_new_n5378_, new_n5378_);
  not g_9625 (not_new_n5944_, new_n5944_);
  not g_9626 (not_new_n1537__8, new_n1537_);
  or g_9627 (new_n7287_, not_new_n7286_, not_new_n7093_);
  not g_9628 (not_new_n9438_, new_n9438_);
  not g_9629 (not_new_n642__168070, new_n642_);
  not g_9630 (not_new_n1995_, new_n1995_);
  or g_9631 (new_n9172_, not_new_n8839_, not_new_n8806_);
  not g_9632 (not_pi047_0, pi047);
  not g_9633 (not_new_n10074_, new_n10074_);
  not g_9634 (not_new_n581__3788186922656647816827176259430, new_n581_);
  not g_9635 (not_po298_5, po298);
  or g_9636 (new_n3182_, not_new_n922__0, not_new_n3181_);
  or g_9637 (new_n3553_, not_new_n1612__490, not_new_n2033__0);
  not g_9638 (new_n1990_, new_n954_);
  not g_9639 (not_new_n2625_, new_n2625_);
  not g_9640 (new_n3999_, new_n3938_);
  not g_9641 (not_new_n598__797922662976120010, new_n598_);
  or g_9642 (new_n7994_, not_new_n617__6782230728490, not_new_n7622__0);
  not g_9643 (not_new_n6984_, new_n6984_);
  not g_9644 (not_new_n8310_, new_n8310_);
  or g_9645 (new_n9827_, not_new_n1063__47475615099430, not_new_n9386__0);
  not g_9646 (not_new_n8152__0, new_n8152_);
  or g_9647 (new_n8374_, not_new_n622__138412872010, not_new_n8131_);
  xnor g_9648 (key_gate_66, key_66, new_n3915_);
  not g_9649 (not_new_n3117_, new_n3117_);
  not g_9650 (new_n4757_, new_n1606_);
  not g_9651 (not_new_n4949__0, new_n4949_);
  and g_9652 (and_new_n8112__new_n8484_, new_n8484_, new_n8112_);
  and g_9653 (new_n5050_, new_n5389_, and_new_n4984__new_n5390_);
  not g_9654 (not_new_n1035__3, new_n1035_);
  not g_9655 (not_new_n635__8235430, new_n635_);
  not g_9656 (not_new_n2871_, new_n2871_);
  and g_9657 (new_n4766_, new_n4860_, new_n4861_);
  or g_9658 (new_n5094_, new_n642_, new_n1035_);
  or g_9659 (new_n5157_, new_n644_, new_n1059_);
  not g_9660 (not_new_n631__1915812313805664144010, new_n631_);
  or g_9661 (new_n8844_, not_new_n8859_, not_new_n9012_);
  or g_9662 (new_n2205_, not_pi185, not_new_n586__968890104070);
  not g_9663 (not_new_n6295_, new_n6295_);
  not g_9664 (not_new_n9342_, new_n9342_);
  not g_9665 (not_new_n4657_, new_n4657_);
  not g_9666 (not_new_n642__3430, new_n642_);
  and g_9667 (and_not_pi036_1_not_pi037_1, not_pi037_1, not_pi036_1);
  not g_9668 (not_new_n994__57648010, new_n994_);
  not g_9669 (not_new_n7163_, new_n7163_);
  or g_9670 (new_n9559_, not_new_n9558_, not_new_n9459_);
  not g_9671 (not_new_n3985__0, new_n3985_);
  or g_9672 (new_n5225_, not_new_n5224_, not_new_n5048_);
  not g_9673 (not_new_n7099_, new_n7099_);
  not g_9674 (not_new_n7051_, new_n7051_);
  or g_9675 (new_n8547_, not_new_n8233_, not_new_n8265__2);
  not g_9676 (new_n4787_, new_n1071_);
  not g_9677 (not_pi140_0, pi140);
  not g_9678 (not_pi054, pi054);
  not g_9679 (not_new_n2823_, new_n2823_);
  not g_9680 (not_new_n5630__1, new_n5630_);
  or g_9681 (new_n7512_, not_new_n7510_, not_new_n7168_);
  or g_9682 (new_n3728_, not_new_n2133_, not_new_n963_);
  or g_9683 (new_n739_, not_new_n3252_, not_new_n3251_);
  not g_9684 (not_new_n8882_, new_n8882_);
  not g_9685 (not_new_n2984_, new_n2984_);
  or g_9686 (new_n5301_, not_new_n5110_, not_new_n5299_);
  not g_9687 (not_new_n4120__0, new_n4120_);
  not g_9688 (not_new_n1169__0, new_n1169_);
  not g_9689 (not_new_n5461_, new_n5461_);
  or g_9690 (new_n6941_, not_new_n6770_, not_new_n6640__2);
  or g_9691 (or_not_new_n1231__not_new_n1229_, not_new_n1229_, not_new_n1231_);
  or g_9692 (new_n2328_, not_new_n1585__16284135979104490, not_new_n5733_);
  not g_9693 (not_new_n1053__2, new_n1053_);
  or g_9694 (new_n3139_, not_new_n581__63668057609090279857414351392240010, not_new_n640__6);
  or g_9695 (new_n2713_, not_new_n590__4, or_not_new_n4227__not_new_n1608_);
  not g_9696 (new_n8880_, new_n639_);
  or g_9697 (new_n4465_, not_new_n4687_, not_new_n4686_);
  or g_9698 (new_n1928_, not_new_n1584__7, not_new_n9432_);
  not g_9699 (not_new_n1012__0, new_n1012_);
  or g_9700 (new_n971_, not_pi008, not_new_n1536__3);
  not g_9701 (not_new_n3857_, new_n3857_);
  or g_9702 (new_n5504_, not_new_n5505_, not_new_n5521_);
  not g_9703 (not_new_n2208_, new_n2208_);
  or g_9704 (new_n6948_, not_new_n6529__0, not_new_n1057__1176490);
  not g_9705 (not_new_n9621_, new_n9621_);
  or g_9706 (new_n4058_, not_new_n3983_, not_new_n4026_);
  not g_9707 (new_n7636_, new_n1604_);
  not g_9708 (not_new_n5722_, new_n5722_);
  or g_9709 (new_n6204_, not_new_n5905__2, not_new_n6032_);
  not g_9710 (not_new_n6974__9, new_n6974_);
  or g_9711 (new_n7389_, not_new_n7387_, not_new_n7327_);
  not g_9712 (not_new_n3150_, new_n3150_);
  or g_9713 (new_n8839_, not_new_n9007_, not_new_n9008_);
  not g_9714 (not_new_n5804_, new_n5804_);
  not g_9715 (not_new_n1612__6782230728490, new_n1612_);
  not g_9716 (new_n8148_, new_n1067_);
  not g_9717 (not_new_n4453__0, new_n4453_);
  or g_9718 (or_not_new_n1559__not_new_n2454_, not_new_n2454_, not_new_n1559_);
  or g_9719 (new_n1718_, not_new_n1631__2326305139872070, not_pi061);
  or g_9720 (new_n7521_, not_new_n7036__1, not_new_n7003__1);
  or g_9721 (new_n3101_, not_new_n928__4, not_new_n1041__3);
  not g_9722 (not_new_n7591__0, new_n7591_);
  or g_9723 (new_n7880_, not_new_n7770_, not_new_n7670_);
  not g_9724 (new_n6516_, new_n633_);
  not g_9725 (not_new_n8269_, new_n8269_);
  not g_9726 (not_new_n5507_, new_n5507_);
  not g_9727 (not_new_n597__403536070, new_n597_);
  or g_9728 (new_n6862_, not_new_n6619_, not_new_n619__3430);
  or g_9729 (or_not_new_n1027__13410686196639649008070_not_new_n4227__0, not_new_n1027__13410686196639649008070, not_new_n4227__0);
  not g_9730 (not_new_n7190_, new_n7190_);
  or g_9731 (new_n2581_, not_new_n606__6, not_new_n5490__0);
  not g_9732 (not_new_n8105__2, new_n8105_);
  or g_9733 (new_n8530_, not_new_n8135__0, not_new_n1602__403536070);
  or g_9734 (new_n5353_, not_new_n5351_, not_new_n5352_);
  not g_9735 (not_new_n6481_, new_n6481_);
  xor g_9736 (key_gate_68, key_68, not_new_n1181_);
  not g_9737 (not_new_n1596__138412872010, new_n1596_);
  not g_9738 (new_n4749_, new_n1051_);
  not g_9739 (not_pi253, pi253);
  not g_9740 (not_new_n654_, new_n654_);
  not g_9741 (new_n5791_, new_n627_);
  not g_9742 (not_new_n3095_, new_n3095_);
  or g_9743 (new_n8556_, not_new_n8357_, not_new_n8555_);
  or g_9744 (new_n6781_, not_new_n646__57648010, not_new_n6536_);
  or g_9745 (new_n10064_, not_new_n634__39098210485829880490, not_new_n1047__2326305139872070);
  or g_9746 (new_n7566_, not_new_n775__113988951853731430, not_new_n6986_);
  not g_9747 (not_new_n2509__1, new_n2509_);
  not g_9748 (not_new_n3384__5, new_n3384_);
  or g_9749 (new_n6419_, not_new_n6234_, or_or_not_new_n6327__not_new_n6373__2_not_new_n1051__490);
  not g_9750 (not_new_n1612__168070, new_n1612_);
  not g_9751 (not_new_n3353_, new_n3353_);
  not g_9752 (not_new_n2932_, new_n2932_);
  not g_9753 (not_new_n8100_, new_n8100_);
  not g_9754 (not_new_n624__47475615099430, new_n624_);
  not g_9755 (new_n8313_, new_n8244_);
  and g_9756 (new_n4724_, new_n4823_, new_n4813_);
  or g_9757 (new_n6011_, not_new_n1597__70, not_new_n5767_);
  not g_9758 (not_new_n2189_, new_n2189_);
  or g_9759 (new_n3669_, not_po298_7, not_new_n634__9);
  not g_9760 (not_new_n6589_, new_n6589_);
  not g_9761 (not_new_n6974__16284135979104490, new_n6974_);
  or g_9762 (new_n8905_, not_new_n9208_, not_new_n9207_);
  or g_9763 (new_n1697_, not_new_n1631__2824752490, not_pi054);
  not g_9764 (new_n9005_, new_n8837_);
  not g_9765 (not_new_n8302_, new_n8302_);
  not g_9766 (not_new_n10080_, new_n10080_);
  not g_9767 (not_new_n644__797922662976120010, new_n644_);
  not g_9768 (not_new_n9413_, new_n9413_);
  not g_9769 (new_n8292_, new_n8265_);
  not g_9770 (not_new_n1053__70, new_n1053_);
  or g_9771 (new_n5702_, not_new_n5701_, not_new_n5700_);
  not g_9772 (not_new_n596__6, key_gate_88);
  or g_9773 (new_n1856_, not_new_n5006_, not_new_n1589__3);
  and g_9774 (new_n5717_, new_n5980_, new_n5981_);
  not g_9775 (not_new_n598__490, new_n598_);
  not g_9776 (not_new_n2935_, new_n2935_);
  not g_9777 (not_new_n633__2, new_n633_);
  not g_9778 (not_new_n6634__1, new_n6634_);
  or g_9779 (new_n5194_, not_new_n4988_, not_new_n5193_);
  not g_9780 (not_new_n9103_, new_n9103_);
  not g_9781 (not_pi036, pi036);
  or g_9782 (new_n3889_, not_new_n641__9, not_new_n6443__797922662976120010);
  or g_9783 (new_n3544_, not_new_n1538__8, not_pi138_0);
  or g_9784 (new_n4351_, not_new_n4251_, not_new_n699_);
  not g_9785 (not_new_n7765_, new_n7765_);
  and g_9786 (new_n8662_, new_n8642_, new_n1067_);
  or g_9787 (new_n8997_, not_new_n8798_, not_new_n8922_);
  and g_9788 (new_n4320_, new_n4409_, new_n4408_);
  or g_9789 (new_n3286_, not_new_n3184__403536070, not_new_n637__8);
  not g_9790 (not_new_n10059__0, new_n10059_);
  not g_9791 (not_new_n1536__797922662976120010, new_n1536_);
  not g_9792 (not_new_n1613__9, new_n1613_);
  or g_9793 (new_n2092_, not_pi147, not_new_n587__8235430);
  not g_9794 (new_n9882_, new_n632_);
  not g_9795 (not_new_n10271_, new_n10271_);
  not g_9796 (not_new_n5076_, new_n5076_);
  not g_9797 (not_new_n5498_, new_n5498_);
  not g_9798 (not_new_n7028_, new_n7028_);
  or g_9799 (new_n2440_, not_new_n1067__0, not_new_n598__1176490);
  not g_9800 (new_n4557_, new_n4502_);
  not g_9801 (not_new_n3372__403536070, new_n3372_);
  and g_9802 (new_n3960_, and_not_pi036_1_not_pi037_1, not_pi038_1);
  not g_9803 (not_new_n7042_, new_n7042_);
  or g_9804 (or_not_new_n5484__not_new_n605__0, not_new_n605__0, not_new_n5484_);
  or g_9805 (new_n928_, not_new_n3387_, not_new_n1023_);
  or g_9806 (new_n8564_, not_new_n637__968890104070, not_new_n8149__0);
  not g_9807 (not_new_n7413_, new_n7413_);
  not g_9808 (not_new_n8456_, new_n8456_);
  not g_9809 (not_new_n1538_, new_n1538_);
  not g_9810 (not_new_n1442_, new_n1442_);
  or g_9811 (new_n1727_, not_new_n1631__797922662976120010, not_pi064);
  not g_9812 (not_new_n1047__332329305696010, new_n1047_);
  not g_9813 (not_new_n1600__2824752490, new_n1600_);
  not g_9814 (not_new_n5585_, new_n5585_);
  or g_9815 (new_n3166_, not_new_n581__2569235775210588780886114772242356213216070, not_new_n636__6);
  not g_9816 (not_new_n7878_, new_n7878_);
  or g_9817 (new_n1687_, key_gate_57, not_new_n596__8235430);
  not g_9818 (not_new_n1057__138412872010, new_n1057_);
  not g_9819 (not_new_n7756_, new_n7756_);
  not g_9820 (not_new_n5685_, new_n5685_);
  or g_9821 (po286, or_not_new_n2903__not_new_n1483_, not_new_n2902_);
  not g_9822 (not_new_n3965_, new_n3965_);
  or g_9823 (new_n2426_, not_new_n4801__0, not_new_n597__3430);
  not g_9824 (not_new_n4610_, new_n4610_);
  not g_9825 (new_n4844_, new_n4758_);
  not g_9826 (not_new_n6991__1, new_n6991_);
  not g_9827 (not_pi172_0, pi172);
  not g_9828 (not_new_n1031__8235430, new_n1031_);
  not g_9829 (not_new_n7508_, new_n7508_);
  not g_9830 (not_new_n6335_, new_n6335_);
  not g_9831 (not_new_n8171_, new_n8171_);
  or g_9832 (new_n3172_, not_new_n581__125892552985318850263419623839875454447587430, not_new_n626__6);
  or g_9833 (new_n7716_, not_new_n7988_, not_new_n7989_);
  not g_9834 (not_new_n637__57648010, new_n637_);
  or g_9835 (or_not_new_n1001__not_new_n1000_, not_new_n1001_, not_new_n1000_);
  or g_9836 (new_n9756_, not_new_n9489_, not_new_n9488_);
  or g_9837 (new_n3024_, not_new_n581__70, not_new_n1597__2);
  not g_9838 (not_new_n989__7, new_n989_);
  not g_9839 (not_new_n3868_, new_n3868_);
  not g_9840 (not_new_n5736_, new_n5736_);
  not g_9841 (not_new_n9623_, new_n9623_);
  or g_9842 (new_n7986_, or_not_new_n7664__0_not_new_n618__6782230728490, not_new_n7985_);
  and g_9843 (new_n6607_, new_n6934_, new_n6651_);
  or g_9844 (new_n7792_, not_new_n1045__2824752490, not_new_n7611__0);
  not g_9845 (not_new_n1791_, new_n1791_);
  not g_9846 (not_new_n2204__0, new_n2204_);
  or g_9847 (new_n8539_, not_new_n640__968890104070, not_new_n8143__0);
  not g_9848 (not_new_n5340_, new_n5340_);
  and g_9849 (new_n1281_, new_n2042_, new_n2041_);
  not g_9850 (not_new_n1031__1, new_n1031_);
  not g_9851 (new_n8835_, new_n635_);
  or g_9852 (or_not_new_n5466__not_new_n5674__1, not_new_n5466_, not_new_n5674__1);
  not g_9853 (not_po298_2326305139872070, po298);
  not g_9854 (not_new_n9329_, new_n9329_);
  or g_9855 (new_n9543_, new_n1045_, new_n635_);
  not g_9856 (not_new_n1047__8, new_n1047_);
  not g_9857 (not_new_n5571_, new_n5571_);
  not g_9858 (not_new_n6730_, new_n6730_);
  not g_9859 (not_new_n636__968890104070, new_n636_);
  or g_9860 (new_n3849_, not_new_n6443__10, not_new_n617__70);
  and g_9861 (new_n8953_, new_n8802_, new_n9145_);
  not g_9862 (not_new_n9366__0, new_n9366_);
  not g_9863 (not_new_n8982_, new_n8982_);
  or g_9864 (new_n6874_, not_new_n617__19773267430, not_new_n6498__0);
  or g_9865 (new_n4711_, not_new_n4433__0, not_new_n1019__4);
  not g_9866 (new_n5507_, new_n1028_);
  or g_9867 (new_n9759_, not_new_n1596__797922662976120010, not_new_n9420_);
  not g_9868 (not_new_n587__24010, new_n587_);
  not g_9869 (not_new_n1047__4, new_n1047_);
  not g_9870 (not_new_n7674_, new_n7674_);
  and g_9871 (and_and_new_n2314__new_n2317__new_n2315_, new_n2315_, and_new_n2314__new_n2317_);
  not g_9872 (not_new_n8914_, new_n8914_);
  not g_9873 (not_new_n5642_, new_n5642_);
  or g_9874 (new_n10039_, new_n631_, new_n1043_);
  not g_9875 (not_new_n1028__2, new_n1028_);
  not g_9876 (not_new_n9286_, new_n9286_);
  not g_9877 (not_new_n1600__968890104070, new_n1600_);
  not g_9878 (not_new_n4118__0, new_n4118_);
  not g_9879 (not_new_n1728__47475615099430, new_n1728_);
  not g_9880 (not_new_n7738_, new_n7738_);
  not g_9881 (new_n6497_, new_n1598_);
  or g_9882 (new_n3471_, not_new_n2033_, not_new_n1613__490);
  not g_9883 (not_new_n5034_, new_n5034_);
  or g_9884 (new_n2020_, not_new_n636__0, not_new_n601__70);
  not g_9885 (not_new_n8890_, new_n8890_);
  or g_9886 (or_not_new_n2053__not_new_n2054_, not_new_n2053_, not_new_n2054_);
  or g_9887 (new_n9192_, not_new_n647__47475615099430, not_new_n8843_);
  not g_9888 (not_new_n4773_, new_n4773_);
  not g_9889 (not_new_n6031_, new_n6031_);
  and g_9890 (new_n5516_, new_n5699_, new_n5698_);
  or g_9891 (new_n645_, or_or_not_new_n2110__not_new_n2111__not_new_n2113_, not_new_n2112_);
  not g_9892 (not_new_n3953_, new_n3953_);
  or g_9893 (po134, not_new_n3485_, not_new_n3486_);
  not g_9894 (not_new_n5355_, new_n5355_);
  xor g_9895 (key_gate_7, key_7, not_new_n3926_);
  not g_9896 (not_pi251_0, pi251);
  or g_9897 (new_n6082_, not_new_n6081_, not_new_n5856_);
  and g_9898 (and_new_n1750__new_n1751_, new_n1750_, new_n1751_);
  not g_9899 (not_new_n8885_, new_n8885_);
  not g_9900 (not_pi035, pi035);
  not g_9901 (not_new_n644__168070, new_n644_);
  or g_9902 (new_n2434_, not_new_n9969__0, not_new_n599__168070);
  or g_9903 (new_n8509_, or_not_new_n8169__1_not_new_n8508_, not_new_n8507_);
  or g_9904 (new_n7209_, not_new_n6962_, not_new_n7162_);
  or g_9905 (new_n6162_, not_new_n5771__0, not_new_n1602__490);
  or g_9906 (new_n7819_, not_new_n7945_, not_new_n7705_);
  and g_9907 (and_not_pi060_1_not_pi059_1, not_pi060_1, not_pi059_1);
  not g_9908 (not_new_n1580__16284135979104490, new_n1580_);
  not g_9909 (not_new_n1728__4, new_n1728_);
  not g_9910 (new_n6531_, new_n637_);
  and g_9911 (and_new_n7160__new_n7500_, new_n7160_, new_n7500_);
  not g_9912 (not_new_n1584__2326305139872070, new_n1584_);
  not g_9913 (new_n4075_, pi260);
  not g_9914 (not_new_n5918_, new_n5918_);
  or g_9915 (new_n4587_, not_new_n4432_, not_new_n1002__3);
  or g_9916 (new_n4506_, not_new_n4547_, not_new_n4548_);
  not g_9917 (not_new_n1611__4, new_n1611_);
  xor g_9918 (key_gate_8, new_n1699_, key_8);
  not g_9919 (not_new_n6735_, new_n6735_);
  not g_9920 (not_pi168_2, pi168);
  or g_9921 (or_not_new_n6328__not_new_n6373__3, not_new_n6373__3, not_new_n6328_);
  or g_9922 (new_n7197_, not_new_n7196_, not_new_n6991__0);
  not g_9923 (not_new_n3372__10, new_n3372_);
  not g_9924 (not_new_n1331_, new_n1331_);
  not g_9925 (not_new_n7033_, new_n7033_);
  not g_9926 (not_new_n7010__2, new_n7010_);
  not g_9927 (not_new_n2756_, new_n2756_);
  or g_9928 (new_n3073_, not_new_n636__4, not_new_n3372__5585458640832840070);
  not g_9929 (not_new_n775__113988951853731430, new_n775_);
  not g_9930 (new_n5778_, new_n645_);
  not g_9931 (not_new_n3518_, new_n3518_);
  not g_9932 (not_new_n8251__0, new_n8251_);
  or g_9933 (new_n2910_, not_new_n3311__3430, not_new_n1049__1);
  not g_9934 (new_n4923_, new_n1039_);
  not g_9935 (not_new_n1014__1, new_n1014_);
  not g_9936 (not_new_n762_, new_n762_);
  or g_9937 (new_n1976_, not_new_n1268_, not_new_n1971_);
  not g_9938 (not_new_n1633_, key_gate_3);
  and g_9939 (new_n6592_, new_n6653_, new_n6875_);
  or g_9940 (new_n10272_, not_new_n10010_, not_new_n10011_);
  not g_9941 (not_new_n6234_, new_n6234_);
  not g_9942 (not_new_n8605_, new_n8605_);
  not g_9943 (not_new_n7004_, new_n7004_);
  or g_9944 (new_n8585_, not_new_n8157__0, not_new_n627__968890104070);
  not g_9945 (not_new_n1063__8, new_n1063_);
  not g_9946 (not_new_n5315_, new_n5315_);
  or g_9947 (or_not_new_n2734__not_new_n2733_, not_new_n2734_, not_new_n2733_);
  not g_9948 (not_new_n625__8, new_n625_);
  not g_9949 (not_new_n5711_, new_n5711_);
  not g_9950 (not_new_n9440_, new_n9440_);
  or g_9951 (new_n9114_, not_new_n1598__19773267430, not_new_n621__47475615099430);
  not g_9952 (new_n9074_, new_n8973_);
  not g_9953 (not_new_n3348_, new_n3348_);
  not g_9954 (new_n1594_, new_n1536_);
  not g_9955 (not_new_n5745__0, new_n5745_);
  not g_9956 (not_new_n2191_, new_n2191_);
  not g_9957 (not_new_n2085_, new_n2085_);
  not g_9958 (not_new_n607__8, new_n607_);
  not g_9959 (not_new_n3315__1, new_n3315_);
  not g_9960 (not_new_n5184_, new_n5184_);
  not g_9961 (not_new_n3411_, new_n3411_);
  not g_9962 (not_new_n1591__1176490, new_n1591_);
  not g_9963 (not_pi064_8, pi064);
  and g_9964 (new_n592_, new_n1412_, new_n988_);
  or g_9965 (new_n8391_, not_new_n8350_, not_new_n8271__0);
  or g_9966 (new_n9742_, not_new_n9374__0, not_new_n9685_);
  not g_9967 (not_new_n7423_, new_n7423_);
  or g_9968 (new_n3606_, not_new_n984__7, not_pi169_0);
  and g_9969 (and_new_n1760__new_n1759_, new_n1759_, new_n1760_);
  not g_9970 (not_new_n6968_, new_n6968_);
  not g_9971 (not_new_n8919_, new_n8919_);
  and g_9972 (new_n1527_, new_n3080_, and_new_n3082__new_n998_);
  not g_9973 (not_new_n2544_, new_n2544_);
  or g_9974 (new_n2681_, not_new_n606__1176490, not_new_n5483__0);
  not g_9975 (not_new_n5755_, new_n5755_);
  not g_9976 (not_new_n634__39098210485829880490, new_n634_);
  not g_9977 (not_new_n2829_, new_n2829_);
  not g_9978 (not_new_n611__24010, new_n611_);
  not g_9979 (not_new_n8160__0, new_n8160_);
  not g_9980 (new_n6519_, new_n1063_);
  and g_9981 (new_n1350_, and_new_n1540__new_n2361_, new_n2360_);
  not g_9982 (not_new_n3152_, new_n3152_);
  not g_9983 (not_new_n5627_, new_n5627_);
  or g_9984 (new_n2210_, not_new_n625__0, not_new_n601__19773267430);
  not g_9985 (not_new_n4949_, new_n4949_);
  and g_9986 (new_n1499_, new_n998_, new_n3021_);
  or g_9987 (new_n5935_, not_new_n5742_, not_new_n631__1176490);
  not g_9988 (not_new_n5746_, new_n5746_);
  not g_9989 (not_new_n2864_, new_n2864_);
  and g_9990 (and_new_n1282__new_n2046_, new_n2046_, new_n1282_);
  or g_9991 (new_n5585_, not_new_n5584_, not_new_n5579_);
  not g_9992 (not_new_n9999_, new_n9999_);
  or g_9993 (new_n9677_, not_new_n9676_, not_new_n9372_);
  or g_9994 (new_n9306_, not_new_n8870__0, not_new_n1061__6782230728490);
  or g_9995 (new_n6739_, not_new_n6738_, not_new_n6736_);
  or g_9996 (new_n9068_, new_n637_, new_n1065_);
  not g_9997 (not_new_n4781__0, new_n4781_);
  not g_9998 (not_new_n6548_, new_n6548_);
  and g_9999 (new_n4764_, new_n4858_, new_n4859_);
  not g_10000 (not_new_n10323_, new_n10323_);
  or g_10001 (new_n1166_, not_new_n3862_, not_new_n3861_);
  not g_10002 (not_new_n4270_, new_n4270_);
  not g_10003 (not_new_n1584__8235430, new_n1584_);
  not g_10004 (not_pi175_0, pi175);
  not g_10005 (new_n4161_, new_n4086_);
  not g_10006 (not_new_n7147_, new_n7147_);
  not g_10007 (not_new_n4485_, new_n4485_);
  not g_10008 (not_new_n5497_, new_n5497_);
  not g_10009 (not_new_n7267__0, new_n7267_);
  not g_10010 (not_new_n1067__8, new_n1067_);
  not g_10011 (not_new_n1600__5, new_n1600_);
  or g_10012 (new_n5001_, not_new_n5377_, not_new_n5378_);
  not g_10013 (not_new_n8172__1, new_n8172_);
  not g_10014 (not_new_n6994_, new_n6994_);
  not g_10015 (not_new_n10311_, new_n10311_);
  not g_10016 (not_pi104, pi104);
  not g_10017 (not_new_n6532_, new_n6532_);
  or g_10018 (new_n8912_, not_new_n9255_, not_new_n9254_);
  or g_10019 (new_n5867_, not_new_n6176_, not_new_n6175_);
  not g_10020 (not_po296_6168735096280623662907561568153897267931784070, po296);
  and g_10021 (and_and_not_pi051_1_not_pi050_1_not_pi049_1, not_pi049_1, and_not_pi051_1_not_pi050_1);
  and g_10022 (and_new_n3079__new_n998_, new_n998_, new_n3079_);
  or g_10023 (new_n3353_, not_pi046_0, not_new_n1534__57648010);
  or g_10024 (new_n7240_, not_new_n7442_, not_new_n7005_);
  not g_10025 (not_new_n6246_, new_n6246_);
  not g_10026 (not_new_n7026__1, new_n7026_);
  not g_10027 (not_pi057, pi057);
  not g_10028 (not_new_n6263_, new_n6263_);
  not g_10029 (not_new_n1045__6782230728490, new_n1045_);
  and g_10030 (new_n1231_, and_new_n1230__new_n1799_, new_n1798_);
  or g_10031 (new_n1020_, not_new_n3362_, not_new_n3361_);
  not g_10032 (new_n4076_, pi257);
  not g_10033 (not_pi072, pi072);
  not g_10034 (not_new_n1603__19773267430, new_n1603_);
  not g_10035 (not_new_n1581__2326305139872070, new_n1581_);
  not g_10036 (new_n2218_, new_n970_);
  not g_10037 (not_new_n1039__39098210485829880490, new_n1039_);
  or g_10038 (or_not_new_n4825__not_new_n4804_, not_new_n4825_, not_new_n4804_);
  or g_10039 (new_n5227_, not_new_n640__3430, not_new_n1604__9);
  not g_10040 (not_new_n1045__19773267430, new_n1045_);
  or g_10041 (new_n2878_, not_po296_14811132966169777414641055325137507340304213552070, not_pi262);
  or g_10042 (new_n740_, not_new_n3254_, not_new_n3253_);
  or g_10043 (new_n960_, or_or_not_new_n1295__not_new_n1293__not_new_n2097_, not_new_n2096_);
  or g_10044 (or_not_new_n1782__not_new_n1783_, not_new_n1783_, not_new_n1782_);
  not g_10045 (not_new_n9086_, new_n9086_);
  xnor g_10046 (key_gate_35, new_n1711_, key_35);
  not g_10047 (not_new_n1580__19773267430, new_n1580_);
  or g_10048 (new_n2468_, not_new_n600__138412872010, not_new_n4124__0);
  not g_10049 (not_new_n9093_, new_n9093_);
  not g_10050 (not_new_n718__0, new_n718_);
  not g_10051 (not_new_n5185_, new_n5185_);
  or g_10052 (new_n8222_, not_new_n8500_, not_new_n8499_);
  or g_10053 (or_not_new_n5436__not_new_n5630__1, not_new_n5630__1, not_new_n5436_);
  or g_10054 (new_n5962_, not_new_n5844_, not_new_n5960_);
  or g_10055 (new_n4783_, not_new_n4833__0, not_new_n4787__0);
  not g_10056 (not_new_n1603__490, new_n1603_);
  not g_10057 (not_new_n610__168070, new_n610_);
  or g_10058 (new_n4601_, not_new_n1004__3, not_new_n4427_);
  or g_10059 (new_n9659_, new_n645_, new_n1071_);
  xor g_10060 (key_gate_71, new_n1636_, key_71);
  or g_10061 (new_n7452_, not_new_n775__332329305696010, not_new_n7132_);
  not g_10062 (not_new_n1584__6782230728490, new_n1584_);
  not g_10063 (not_new_n7315__0, new_n7315_);
  or g_10064 (new_n7046_, not_new_n7462_, not_new_n7461_);
  or g_10065 (new_n3314_, not_new_n3990__0, not_pi064_0);
  not g_10066 (not_new_n5705_, new_n5705_);
  or g_10067 (new_n4868_, not_new_n4744_, not_new_n1601__7);
  or g_10068 (new_n3730_, not_new_n3459_, not_new_n1962_);
  or g_10069 (new_n5945_, not_new_n5944_, not_new_n5746_);
  or g_10070 (new_n8104_, not_new_n634__968890104070, not_new_n8109_);
  not g_10071 (not_new_n7438_, new_n7438_);
  not g_10072 (not_new_n2230_, new_n2230_);
  not g_10073 (not_new_n8178_, new_n8178_);
  not g_10074 (not_new_n7116_, new_n7116_);
  not g_10075 (not_new_n3939_, new_n3939_);
  not g_10076 (not_new_n617__47475615099430, new_n617_);
  not g_10077 (not_new_n9510_, new_n9510_);
  or g_10078 (new_n9732_, not_new_n9362_, not_new_n635__2326305139872070);
  not g_10079 (not_new_n5957_, new_n5957_);
  not g_10080 (not_new_n2827_, new_n2827_);
  not g_10081 (not_new_n8978__2, new_n8978_);
  not g_10082 (new_n3953_, pi047);
  or g_10083 (or_not_new_n2597__not_new_n2601_, not_new_n2597_, not_new_n2601_);
  or g_10084 (new_n6569_, not_new_n6958_, not_new_n6959_);
  not g_10085 (not_new_n3165_, new_n3165_);
  not g_10086 (not_new_n4138_, new_n4138_);
  or g_10087 (new_n3230_, not_new_n3185__19773267430, not_new_n1061__4);
  and g_10088 (and_and_new_n8753__new_n8754__new_n8761_, new_n8761_, and_new_n8753__new_n8754_);
  not g_10089 (not_new_n7642_, new_n7642_);
  not g_10090 (not_new_n1613__24010, new_n1613_);
  or g_10091 (new_n10336_, not_new_n1065__39098210485829880490, not_new_n9913_);
  not g_10092 (not_pi064_332329305696010, pi064);
  not g_10093 (new_n6504_, new_n625_);
  or g_10094 (new_n4592_, not_new_n4473__0, not_new_n4472_);
  not g_10095 (not_new_n7442_, new_n7442_);
  not g_10096 (not_new_n10100_, new_n10100_);
  or g_10097 (new_n2552_, not_new_n2509__3, not_pi197);
  not g_10098 (not_new_n9724_, new_n9724_);
  not g_10099 (not_new_n1017__1, new_n1017_);
  not g_10100 (not_new_n4099_, new_n4099_);
  not g_10101 (not_pi069, pi069);
  not g_10102 (not_pi182, pi182);
  or g_10103 (new_n5079_, not_new_n5285_, not_new_n5284_);
  not g_10104 (not_new_n2130_, new_n2130_);
  not g_10105 (not_new_n2545_, new_n2545_);
  not g_10106 (not_new_n639__168070, new_n639_);
  not g_10107 (not_new_n9748_, new_n9748_);
  not g_10108 (new_n6945_, new_n6608_);
  not g_10109 (not_new_n7966_, new_n7966_);
  not g_10110 (not_new_n707_, new_n707_);
  or g_10111 (new_n10059_, new_n1049_, new_n648_);
  or g_10112 (new_n9426_, not_new_n9645_, not_new_n9406_);
  or g_10113 (new_n2706_, not_new_n2705_, not_new_n1573_);
  and g_10114 (and_and_new_n2238__new_n2241__new_n2239_, new_n2239_, and_new_n2238__new_n2241_);
  not g_10115 (not_new_n4701_, new_n4701_);
  not g_10116 (not_new_n2509__0, new_n2509_);
  not g_10117 (not_new_n1622__1, new_n1622_);
  not g_10118 (not_new_n10265_, new_n10265_);
  not g_10119 (not_new_n10182_, new_n10182_);
  not g_10120 (not_new_n3256_, new_n3256_);
  or g_10121 (new_n5685_, not_pi142_2, not_new_n5459__0);
  not g_10122 (not_new_n1578_, new_n1578_);
  not g_10123 (not_new_n7783_, new_n7783_);
  not g_10124 (not_pi001_0, pi001);
  and g_10125 (new_n1560_, new_n3632_, new_n3633_);
  not g_10126 (new_n6255_, new_n1045_);
  not g_10127 (not_new_n2987_, new_n2987_);
  or g_10128 (new_n5964_, not_new_n5920__1, not_new_n5963_);
  not g_10129 (not_new_n5487_, new_n5487_);
  not g_10130 (not_new_n3311__10, new_n3311_);
  or g_10131 (new_n7422_, not_new_n7122_, not_new_n775__1176490);
  or g_10132 (new_n5400_, not_new_n5399_, not_new_n5398_);
  or g_10133 (new_n7314_, not_new_n7315__0, not_new_n7167_);
  not g_10134 (not_pi163_3, pi163);
  not g_10135 (not_new_n2153_, new_n2153_);
  or g_10136 (new_n2770_, not_new_n595__3, not_new_n7053_);
  not g_10137 (not_new_n3311__9, new_n3311_);
  not g_10138 (not_new_n4441__0, new_n4441_);
  or g_10139 (or_or_not_new_n6353__not_new_n6232__5_not_new_n1069__3430, not_new_n1069__3430, or_not_new_n6353__not_new_n6232__5);
  or g_10140 (new_n5978_, not_new_n644__8235430, not_new_n5789_);
  or g_10141 (new_n3731_, not_new_n627__10, not_new_n1055__6);
  or g_10142 (new_n5480_, not_new_n5620_, not_new_n5621_);
  not g_10143 (not_new_n3218_, new_n3218_);
  and g_10144 (new_n4906_, new_n4901_, new_n5111_);
  not g_10145 (not_new_n4803__0, new_n4803_);
  or g_10146 (new_n6732_, not_new_n1601__1176490, not_new_n6503_);
  or g_10147 (new_n6712_, not_new_n6521_, not_new_n1059__168070);
  not g_10148 (not_new_n5247_, new_n5247_);
  not g_10149 (not_new_n8070_, new_n8070_);
  not g_10150 (not_new_n648__5585458640832840070, new_n648_);
  or g_10151 (new_n3052_, not_new_n3372__6782230728490, not_new_n645__4);
  and g_10152 (new_n1551_, new_n3614_, new_n3615_);
  not g_10153 (not_new_n596__57648010, key_gate_88);
  not g_10154 (not_new_n5358_, new_n5358_);
  not g_10155 (not_new_n1537__3430, new_n1537_);
  not g_10156 (not_new_n7636__0, new_n7636_);
  not g_10157 (not_new_n9745_, new_n9745_);
  not g_10158 (not_new_n648__1, new_n648_);
  or g_10159 (new_n5183_, not_new_n5086_, not_new_n4905_);
  not g_10160 (not_new_n625__93874803376477543056490, new_n625_);
  or g_10161 (new_n6093_, not_new_n5878__3, not_new_n5949_);
  not g_10162 (not_new_n9924_, new_n9924_);
  not g_10163 (new_n6984_, new_n742_);
  not g_10164 (not_new_n729_, new_n729_);
  not g_10165 (not_new_n4948__0, new_n4948_);
  not g_10166 (not_new_n1057__403536070, new_n1057_);
  or g_10167 (or_not_new_n1939__not_new_n1940_, not_new_n1939_, not_new_n1940_);
  not g_10168 (not_new_n642__2, new_n642_);
  not g_10169 (not_new_n5123_, new_n5123_);
  not g_10170 (not_new_n4137__0, new_n4137_);
  not g_10171 (not_new_n4071_, new_n4071_);
  not g_10172 (not_new_n1439_, new_n1439_);
  or g_10173 (new_n4343_, not_new_n671_, not_new_n4244_);
  not g_10174 (not_new_n1585__113988951853731430, new_n1585_);
  or g_10175 (new_n3275_, not_new_n589__77309937197074445241370944070, not_new_n1604__5);
  not g_10176 (not_new_n7111_, new_n7111_);
  not g_10177 (not_pi207, pi207);
  or g_10178 (new_n6089_, not_new_n5862_, not_new_n6159_);
  or g_10179 (new_n2613_, not_new_n609__10, not_new_n4454_);
  not g_10180 (not_pi106, pi106);
  not g_10181 (not_new_n588__4, new_n588_);
  not g_10182 (not_new_n8825_, new_n8825_);
  and g_10183 (and_and_new_n6357__new_n6356__new_n6404_, and_new_n6357__new_n6356_, new_n6404_);
  or g_10184 (new_n1035_, not_new_n3407_, not_new_n3408_);
  not g_10185 (new_n6517_, new_n1067_);
  not g_10186 (not_new_n8470_, new_n8470_);
  or g_10187 (new_n4066_, not_pi033_5, not_new_n3993_);
  not g_10188 (not_new_n4438__0, new_n4438_);
  not g_10189 (not_new_n5714_, new_n5714_);
  or g_10190 (new_n5836_, not_new_n6221_, not_new_n6222_);
  or g_10191 (new_n2729_, not_new_n1616_, not_new_n2719_);
  not g_10192 (not_new_n5843_, new_n5843_);
  not g_10193 (not_new_n5522_, new_n5522_);
  not g_10194 (not_new_n7524_, new_n7524_);
  and g_10195 (and_new_n1934__new_n1937_, new_n1937_, new_n1934_);
  or g_10196 (new_n2824_, not_pi256_0, not_po296_125892552985318850263419623839875454447587430);
  or g_10197 (new_n6757_, not_new_n6507__0, not_new_n625__19773267430);
  not g_10198 (new_n9617_, new_n9497_);
  not g_10199 (not_new_n6333_, new_n6333_);
  not g_10200 (not_new_n639__490, new_n639_);
  not g_10201 (not_new_n639__2824752490, new_n639_);
  not g_10202 (not_new_n1598__1176490, new_n1598_);
  not g_10203 (not_new_n1971_, new_n1971_);
  and g_10204 (new_n5889_, new_n6144_, new_n6143_);
  not g_10205 (new_n4734_, new_n1045_);
  and g_10206 (new_n7079_, new_n7205_, new_n6966_);
  not g_10207 (not_new_n3864_, new_n3864_);
  not g_10208 (not_new_n1035__9, new_n1035_);
  not g_10209 (not_new_n6509_, new_n6509_);
  not g_10210 (not_new_n1011__0, new_n1011_);
  or g_10211 (new_n3191_, not_new_n634__7, not_new_n589__1);
  or g_10212 (new_n8387_, not_new_n8134__1, not_new_n1601__332329305696010);
  not g_10213 (not_new_n3846_, new_n3846_);
  not g_10214 (not_pi012_0, pi012);
  not g_10215 (new_n4165_, new_n4092_);
  not g_10216 (not_new_n7206_, new_n7206_);
  not g_10217 (not_new_n8707_, new_n8707_);
  not g_10218 (not_new_n928__797922662976120010, new_n928_);
  and g_10219 (new_n9993_, new_n10144_, new_n9862_);
  not g_10220 (not_new_n4614_, new_n4614_);
  not g_10221 (not_new_n9521_, new_n9521_);
  or g_10222 (new_n4209_, not_new_n4092_, not_pi249_2);
  and g_10223 (new_n8091_, new_n8371_, new_n8090_);
  or g_10224 (new_n2044_, not_new_n6568_, not_new_n1580__24010);
  not g_10225 (not_new_n1599__138412872010, new_n1599_);
  or g_10226 (new_n2969_, not_new_n621__3, not_new_n604__47475615099430);
  not g_10227 (not_new_n9388_, new_n9388_);
  not g_10228 (not_new_n595__1, new_n595_);
  not g_10229 (not_pi270_2, pi270);
  not g_10230 (new_n2509_, new_n988_);
  not g_10231 (not_new_n2896_, new_n2896_);
  not g_10232 (not_new_n4916_, new_n4916_);
  not g_10233 (not_new_n4263_, new_n4263_);
  not g_10234 (not_pi247_1, pi247);
  not g_10235 (not_new_n4101_, new_n4101_);
  not g_10236 (not_new_n9879_, new_n9879_);
  or g_10237 (new_n2958_, not_new_n595__6782230728490, not_new_n7058_);
  or g_10238 (new_n8492_, not_new_n8251_, not_new_n1607__24010);
  or g_10239 (new_n7671_, not_new_n7658_, not_new_n7886_);
  or g_10240 (new_n8519_, not_new_n8225_, not_new_n8257_);
  not g_10241 (not_new_n3991_, new_n3991_);
  not g_10242 (not_new_n5156__0, new_n5156_);
  or g_10243 (new_n3333_, not_new_n1534__8, not_pi038_0);
  not g_10244 (new_n1943_, new_n626_);
  not g_10245 (not_pi130, pi130);
  or g_10246 (new_n2235_, not_new_n1591__968890104070, not_new_n8912_);
  not g_10247 (not_new_n7858_, new_n7858_);
  or g_10248 (new_n8312_, not_new_n8280_, not_new_n648__47475615099430);
  not g_10249 (not_pi042, pi042);
  or g_10250 (new_n9436_, not_new_n9756_, not_new_n9757_);
  or g_10251 (or_not_new_n2881__not_new_n2880_, not_new_n2880_, not_new_n2881_);
  and g_10252 (new_n3982_, new_n4055_, new_n4056_);
  not g_10253 (not_new_n9948_, new_n9948_);
  not g_10254 (new_n4842_, new_n4763_);
  or g_10255 (new_n3900_, not_new_n9923_, not_new_n1057__7);
  not g_10256 (not_new_n1584__1, new_n1584_);
  and g_10257 (new_n6580_, new_n6654_, new_n6856_);
  and g_10258 (new_n9496_, new_n9792_, new_n9791_);
  and g_10259 (and_new_n2181__new_n2184_, new_n2181_, new_n2184_);
  or g_10260 (new_n9660_, new_n637_, new_n1065_);
  not g_10261 (not_new_n8318_, new_n8318_);
  and g_10262 (and_and_and_new_n1053__new_n6232__new_n6395__new_n6317_, and_and_new_n1053__new_n6232__new_n6395_, new_n6317_);
  or g_10263 (new_n7976_, not_new_n7975_, not_new_n7974_);
  or g_10264 (new_n6043_, not_new_n5803_, not_new_n646__168070);
  or g_10265 (new_n3500_, not_pi116_0, not_new_n1537__57648010);
  not g_10266 (not_new_n10261_, new_n10261_);
  or g_10267 (new_n2014_, not_new_n1276_, not_new_n2009_);
  not g_10268 (not_new_n7681_, new_n7681_);
  not g_10269 (not_new_n5489__0, new_n5489_);
  not g_10270 (not_new_n3023_, new_n3023_);
  or g_10271 (new_n2814_, not_new_n7047_, not_new_n595__8);
  not g_10272 (not_new_n8112__0, new_n8112_);
  or g_10273 (new_n3690_, not_pi231, not_new_n989__8235430);
  or g_10274 (new_n2148_, not_new_n586__2824752490, not_pi182);
  not g_10275 (not_new_n1626__0, new_n1626_);
  and g_10276 (new_n6358_, and_and_new_n6357__new_n6356__new_n6404_, new_n6367_);
  not g_10277 (new_n6801_, new_n6632_);
  not g_10278 (not_new_n1061__968890104070, new_n1061_);
  or g_10279 (new_n5642_, not_new_n1010__5, not_new_n5431__0);
  and g_10280 (new_n8688_, and_new_n8750__new_n8736_, new_n8718_);
  or g_10281 (new_n1714_, not_new_n596__332329305696010, key_gate_89);
  not g_10282 (new_n6267_, new_n645_);
  xnor g_10283 (key_gate_59, not_new_n1642_, key_59);
  not g_10284 (not_new_n9860_, new_n9860_);
  and g_10285 (new_n4919_, new_n5131_, new_n5134_);
  not g_10286 (not_new_n1037_, new_n1037_);
  and g_10287 (and_new_n8997__new_n8998_, new_n8998_, new_n8997_);
  or g_10288 (new_n3588_, not_new_n1538__797922662976120010, not_pi160_0);
  not g_10289 (not_new_n8153__0, new_n8153_);
  not g_10290 (not_new_n6512__0, new_n6512_);
  not g_10291 (not_new_n9110_, new_n9110_);
  or g_10292 (new_n1049_, not_new_n3442_, not_new_n3443_);
  not g_10293 (not_new_n589__11044276742439206463052992010, new_n589_);
  and g_10294 (new_n5883_, new_n6120_, new_n6121_);
  not g_10295 (not_new_n7773__0, new_n7773_);
  not g_10296 (not_new_n4236_, new_n4236_);
  not g_10297 (not_new_n6088_, new_n6088_);
  not g_10298 (new_n5456_, new_n1018_);
  or g_10299 (or_not_new_n3173__not_new_n3172_, not_new_n3172_, not_new_n3173_);
  or g_10300 (new_n2624_, not_new_n607__9, not_new_n1004_);
  not g_10301 (not_new_n2633_, new_n2633_);
  not g_10302 (new_n7427_, new_n7029_);
  or g_10303 (new_n9191_, not_new_n8850_, not_new_n8984__2);
  not g_10304 (not_pi197, pi197);
  or g_10305 (new_n763_, not_new_n3237_, not_new_n3236_);
  or g_10306 (new_n9583_, not_new_n9581_, not_new_n9466_);
  or g_10307 (new_n8523_, not_new_n8522_, not_new_n8436_);
  or g_10308 (new_n3301_, not_new_n1031__8, not_new_n589__7490483309651862334944941026945644936490);
  not g_10309 (not_new_n9534_, new_n9534_);
  or g_10310 (new_n996_, not_new_n1474_, not_new_n2725_);
  or g_10311 (new_n1722_, not_pi002_0, not_po296_113988951853731430);
  or g_10312 (new_n8481_, not_new_n8331_, not_new_n8248__2);
  or g_10313 (new_n8712_, not_new_n1599__57648010, not_new_n8779_);
  or g_10314 (new_n8747_, not_new_n8604_, not_new_n1152__0);
  and g_10315 (new_n3926_, new_n4027_, new_n3984_);
  or g_10316 (new_n8529_, not_new_n8092_, not_new_n8289__0);
  not g_10317 (not_new_n2654_, new_n2654_);
  not g_10318 (not_pi056_1, pi056);
  not g_10319 (not_new_n3266_, new_n3266_);
  not g_10320 (not_new_n648__968890104070, new_n648_);
  not g_10321 (not_new_n5515_, new_n5515_);
  not g_10322 (not_new_n642__490, new_n642_);
  not g_10323 (not_pi134_2, pi134);
  and g_10324 (po116, pi095, key_gate_101);
  not g_10325 (new_n9425_, new_n640_);
  not g_10326 (not_pi040_1, pi040);
  not g_10327 (not_new_n9012_, new_n9012_);
  not g_10328 (not_new_n2509__5, new_n2509_);
  not g_10329 (not_new_n8350__0, new_n8350_);
  not g_10330 (not_new_n9346_, new_n9346_);
  or g_10331 (new_n1682_, not_pi049, not_new_n1631__168070);
  or g_10332 (new_n9080_, not_new_n9079_, not_new_n8897_);
  and g_10333 (new_n1450_, and_new_n2672__new_n2671_, new_n2670_);
  not g_10334 (not_new_n585__6782230728490, new_n585_);
  not g_10335 (not_new_n10155_, new_n10155_);
  not g_10336 (not_pi033, pi033);
  or g_10337 (or_not_new_n1271__not_new_n1269_, not_new_n1269_, not_new_n1271_);
  not g_10338 (not_new_n9268_, new_n9268_);
  not g_10339 (not_new_n672_, new_n672_);
  not g_10340 (not_pi266_0, pi266);
  not g_10341 (not_new_n5451_, new_n5451_);
  and g_10342 (new_n4480_, new_n4615_, new_n4616_);
  or g_10343 (new_n5422_, not_new_n626__1176490, not_new_n4960_);
  not g_10344 (not_new_n1828_, new_n1828_);
  not g_10345 (not_new_n8851__0, new_n8851_);
  not g_10346 (not_new_n9793_, new_n9793_);
  not g_10347 (new_n8608_, new_n1179_);
  not g_10348 (not_new_n1869_, new_n1869_);
  not g_10349 (new_n8380_, new_n8253_);
  not g_10350 (not_new_n8405_, new_n8405_);
  not g_10351 (not_pi043_1, pi043);
  not g_10352 (not_new_n3251_, new_n3251_);
  not g_10353 (new_n4448_, new_n1012_);
  not g_10354 (not_new_n4909_, new_n4909_);
  not g_10355 (not_po296_797922662976120010, po296);
  or g_10356 (new_n9823_, not_new_n9821_, not_new_n9594__0);
  or g_10357 (new_n4621_, not_new_n4619_, not_new_n4525_);
  or g_10358 (new_n10033_, not_new_n1057__47475615099430, not_new_n636__113988951853731430);
  or g_10359 (new_n10103_, not_new_n10099_, not_new_n10101_);
  or g_10360 (new_n8983_, not_new_n636__47475615099430, not_new_n1057__19773267430);
  not g_10361 (not_new_n5384_, new_n5384_);
  not g_10362 (not_new_n5811__0, new_n5811_);
  or g_10363 (new_n4991_, or_not_new_n5291__not_new_n5290_, not_new_n5200_);
  or g_10364 (new_n7018_, not_new_n7332_, not_new_n7333_);
  not g_10365 (not_new_n596__113988951853731430, key_gate_88);
  or g_10366 (new_n2372_, not_new_n631__1, not_new_n603__3);
  and g_10367 (and_new_n1230__new_n1799_, new_n1230_, new_n1799_);
  not g_10368 (new_n4286_, new_n681_);
  not g_10369 (not_new_n2898_, new_n2898_);
  and g_10370 (new_n1404_, new_n2496_, new_n2495_);
  not g_10371 (not_new_n9659_, new_n9659_);
  not g_10372 (not_new_n10151_, new_n10151_);
  not g_10373 (not_new_n4178_, new_n4178_);
  and g_10374 (and_and_new_n2517__new_n2518__new_n2516_, new_n2516_, and_new_n2517__new_n2518_);
  not g_10375 (not_new_n10210_, new_n10210_);
  not g_10376 (new_n3464_, new_n1057_);
  not g_10377 (not_new_n639__10, new_n639_);
  not g_10378 (not_new_n5536_, new_n5536_);
  not g_10379 (not_new_n1612__138412872010, new_n1612_);
  or g_10380 (new_n5667_, not_pi145_2, not_new_n5469_);
  not g_10381 (not_new_n5079__0, new_n5079_);
  not g_10382 (not_new_n6933_, new_n6933_);
  not g_10383 (not_new_n1600__490, new_n1600_);
  not g_10384 (not_new_n1045__10, new_n1045_);
  or g_10385 (new_n7761_, not_new_n7935_, not_new_n7827_);
  or g_10386 (new_n5662_, not_pi146_3, not_new_n5471__0);
  or g_10387 (new_n1888_, not_new_n7593_, not_new_n1583__5);
  not g_10388 (not_new_n5038_, new_n5038_);
  not g_10389 (not_new_n7596__0, new_n7596_);
  or g_10390 (new_n1958_, not_pi172, not_new_n586__10);
  not g_10391 (new_n8706_, new_n1180_);
  not g_10392 (not_new_n1424_, new_n1424_);
  not g_10393 (new_n10156_, new_n9947_);
  not g_10394 (not_new_n3185__24010, new_n3185_);
  or g_10395 (new_n9701_, not_new_n9337_, not_new_n9506__1);
  or g_10396 (new_n1899_, not_new_n1045_, not_new_n1588__6);
  not g_10397 (not_new_n4782_, new_n4782_);
  or g_10398 (new_n6174_, not_new_n5866_, not_new_n5897_);
  or g_10399 (new_n4215_, not_new_n4150_, not_pi246_1);
  or g_10400 (new_n1662_, not_po296_9, not_pi022);
  not g_10401 (not_new_n4487_, new_n4487_);
  not g_10402 (not_new_n6970_, new_n6970_);
  or g_10403 (new_n8101_, not_new_n8319_, not_new_n8317_);
  not g_10404 (not_pi107, pi107);
  not g_10405 (not_new_n1167_, new_n1167_);
  or g_10406 (new_n9738_, not_new_n9355_, not_new_n1043__47475615099430);
  not g_10407 (not_new_n622__3430, new_n622_);
  or g_10408 (new_n2492_, not_new_n603__2326305139872070, not_new_n619__0);
  not g_10409 (not_new_n1478_, new_n1478_);
  or g_10410 (new_n6843_, not_new_n6841_, not_new_n6842_);
  not g_10411 (new_n9523_, new_n9361_);
  not g_10412 (new_n1971_, new_n953_);
  not g_10413 (not_new_n1576__403536070, new_n1576_);
  not g_10414 (not_new_n6582_, new_n6582_);
  not g_10415 (not_new_n7496_, new_n7496_);
  not g_10416 (not_new_n9796_, new_n9796_);
  not g_10417 (not_new_n5544_, new_n5544_);
  not g_10418 (not_new_n6547_, new_n6547_);
  not g_10419 (not_new_n1183_, key_gate_48);
  not g_10420 (not_new_n10013__1, new_n10013_);
  and g_10421 (and_new_n1820__new_n1823_, new_n1820_, new_n1823_);
  not g_10422 (not_new_n5182__0, new_n5182_);
  or g_10423 (new_n2600_, not_new_n1019__0, not_new_n608__8);
  or g_10424 (new_n8055_, not_new_n1061__57648010, not_new_n7657__0);
  or g_10425 (new_n3629_, not_new_n1611__57648010, not_new_n962_);
  not g_10426 (not_new_n1063__70, new_n1063_);
  not g_10427 (not_new_n7016__1, new_n7016_);
  not g_10428 (not_new_n4251_, new_n4251_);
  not g_10429 (not_new_n7130_, new_n7130_);
  not g_10430 (not_new_n1313_, new_n1313_);
  not g_10431 (not_new_n637__168070, new_n637_);
  or g_10432 (new_n6546_, not_new_n6534_, not_new_n6760_);
  or g_10433 (new_n6864_, not_new_n6619__0, not_new_n619__24010);
  not g_10434 (not_new_n2775_, new_n2775_);
  or g_10435 (new_n2069_, not_new_n4798_, not_new_n591__168070);
  not g_10436 (not_new_n7004__2, new_n7004_);
  not g_10437 (not_new_n1631__332329305696010, key_gate_76);
  or g_10438 (or_not_new_n6042__not_new_n5927_, not_new_n5927_, not_new_n6042_);
  or g_10439 (new_n7754_, not_new_n7946_, not_new_n7907_);
  or g_10440 (new_n7900_, not_new_n7768_, not_new_n7672_);
  not g_10441 (not_new_n9910_, new_n9910_);
  or g_10442 (new_n9011_, new_n1049_, new_n648_);
  not g_10443 (not_new_n6803_, new_n6803_);
  not g_10444 (not_new_n1811_, new_n1811_);
  and g_10445 (new_n3916_, new_n3955_, new_n4046_);
  or g_10446 (new_n7901_, not_new_n7648__1, not_new_n1055__138412872010);
  or g_10447 (new_n7138_, not_new_n7267_, not_new_n7012_);
  or g_10448 (new_n7380_, not_new_n7379_, not_new_n7378_);
  not g_10449 (not_new_n8399_, new_n8399_);
  or g_10450 (new_n6385_, not_new_n640__8235430, not_new_n6292_);
  not g_10451 (not_new_n9963_, new_n9963_);
  or g_10452 (new_n5390_, not_new_n4983_, not_new_n1067__10);
  or g_10453 (new_n4226_, not_new_n4157__1, not_new_n4082_);
  not g_10454 (new_n5437_, pi132);
  buf g_10455 (po034, pi230);
  not g_10456 (not_new_n8627_, new_n8627_);
  or g_10457 (new_n5632_, not_new_n5631_, not_new_n5630__0);
  not g_10458 (not_new_n1604__0, new_n1604_);
  not g_10459 (not_new_n5917_, new_n5917_);
  not g_10460 (not_new_n4685_, new_n4685_);
  or g_10461 (new_n3761_, not_new_n977_, not_new_n2266_);
  and g_10462 (new_n1377_, new_n2427_, new_n2428_);
  or g_10463 (new_n2951_, not_new_n625__3, not_new_n604__968890104070);
  not g_10464 (not_new_n1003__0, new_n1003_);
  not g_10465 (not_new_n4124__1, new_n4124_);
  not g_10466 (not_new_n7386_, new_n7386_);
  or g_10467 (new_n4133_, not_new_n4217_, not_new_n4218_);
  not g_10468 (not_new_n10343_, new_n10343_);
  xnor g_10469 (key_gate_43, new_n3930_, key_43);
  or g_10470 (new_n4214_, not_new_n4163__1, not_new_n4091_);
  not g_10471 (not_new_n1600__168070, new_n1600_);
  not g_10472 (not_new_n5007_, new_n5007_);
  or g_10473 (new_n6622_, not_new_n6587_, not_new_n6745_);
  not g_10474 (not_new_n2313_, new_n2313_);
  not g_10475 (not_new_n595__7, new_n595_);
  or g_10476 (new_n2024_, not_new_n1581__490, not_new_n8188_);
  not g_10477 (not_new_n3694_, new_n3694_);
  or g_10478 (or_not_new_n1560__not_new_n2459_, not_new_n2459_, not_new_n1560_);
  or g_10479 (new_n4195_, not_pi262_1, not_new_n4106_);
  not g_10480 (not_pi131_3, pi131);
  or g_10481 (new_n5006_, not_new_n5314_, not_new_n5315_);
  not g_10482 (not_new_n1597__490, new_n1597_);
  and g_10483 (and_new_n9168__new_n9167_, new_n9167_, new_n9168_);
  not g_10484 (not_new_n9520_, new_n9520_);
  or g_10485 (new_n6371_, not_new_n623__6, not_new_n6305_);
  not g_10486 (new_n7623_, new_n622_);
  not g_10487 (new_n8124_, new_n647_);
  or g_10488 (new_n4222_, not_new_n4085_, not_new_n4159__1);
  not g_10489 (not_new_n2989_, new_n2989_);
  not g_10490 (not_new_n6869_, new_n6869_);
  not g_10491 (not_new_n609__2, new_n609_);
  not g_10492 (not_new_n599__332329305696010, new_n599_);
  not g_10493 (not_new_n8892__0, new_n8892_);
  not g_10494 (not_new_n629__10, new_n629_);
  not g_10495 (not_new_n7658_, new_n7658_);
  not g_10496 (not_new_n628__797922662976120010, new_n628_);
  not g_10497 (not_new_n1576__2824752490, new_n1576_);
  not g_10498 (new_n8610_, new_n1035_);
  not g_10499 (not_new_n9132_, new_n9132_);
  or g_10500 (new_n5612_, not_new_n5444__0, not_pi135_3);
  not g_10501 (not_new_n9218_, new_n9218_);
  not g_10502 (not_pi209, pi209);
  or g_10503 (new_n2214_, not_new_n1581__138412872010, not_new_n8096_);
  or g_10504 (new_n1852_, not_new_n9434_, not_new_n1584__3);
  not g_10505 (not_new_n5503_, new_n5503_);
  or g_10506 (or_or_not_new_n2110__not_new_n2111__not_new_n2113_, not_new_n2113_, or_not_new_n2110__not_new_n2111_);
  not g_10507 (not_new_n5095_, new_n5095_);
  or g_10508 (new_n9507_, not_new_n9713_, not_new_n9712_);
  not g_10509 (new_n4232_, new_n709_);
  not g_10510 (not_new_n6480_, new_n6480_);
  not g_10511 (not_new_n8115_, new_n8115_);
  or g_10512 (new_n4559_, not_new_n4558_, not_new_n4502_);
  not g_10513 (new_n9405_, new_n646_);
  not g_10514 (not_new_n8159__0, new_n8159_);
  not g_10515 (not_new_n2954_, new_n2954_);
  not g_10516 (not_new_n638__24010, new_n638_);
  not g_10517 (not_new_n4044_, new_n4044_);
  not g_10518 (not_new_n593__2326305139872070, new_n593_);
  or g_10519 (new_n6776_, not_new_n6610_, not_new_n6774_);
  not g_10520 (not_new_n696_, new_n696_);
  not g_10521 (not_new_n9907_, new_n9907_);
  or g_10522 (new_n9662_, not_new_n9661_, not_new_n9478_);
  not g_10523 (not_new_n612__1, new_n612_);
  or g_10524 (new_n2678_, not_new_n610__1176490, not_new_n4460__0);
  not g_10525 (not_new_n3319_, new_n3319_);
  not g_10526 (not_new_n3161_, new_n3161_);
  or g_10527 (new_n6059_, not_new_n5900__0, not_new_n5727_);
  not g_10528 (not_new_n1324_, new_n1324_);
  not g_10529 (not_new_n5082_, new_n5082_);
  or g_10530 (new_n5267_, or_not_new_n4899__0_not_new_n5096__0, not_new_n4898__1);
  not g_10531 (not_new_n4576_, new_n4576_);
  or g_10532 (new_n4057_, not_pi060_2, not_new_n3984_);
  or g_10533 (new_n5198_, not_new_n5079_, not_new_n5087_);
  not g_10534 (new_n5438_, pi133);
  not g_10535 (not_new_n644__24010, new_n644_);
  or g_10536 (or_not_new_n1259__not_new_n1257_, not_new_n1257_, not_new_n1259_);
  not g_10537 (not_po296_6782230728490, po296);
  not g_10538 (not_new_n4120__2, new_n4120_);
  not g_10539 (not_new_n1051__8235430, new_n1051_);
  or g_10540 (new_n3445_, not_pi105_0, not_new_n1537__7);
  not g_10541 (not_new_n1053__2824752490, new_n1053_);
  not g_10542 (not_new_n8938_, new_n8938_);
  not g_10543 (not_new_n7576_, new_n7576_);
  not g_10544 (not_new_n1041__3, new_n1041_);
  not g_10545 (not_new_n3957__0, new_n3957_);
  or g_10546 (new_n8582_, not_new_n8445_, not_new_n8581_);
  not g_10547 (not_new_n2199_, new_n2199_);
  not g_10548 (not_new_n2695_, new_n2695_);
  or g_10549 (new_n4400_, not_new_n651_, not_new_n4282_);
  or g_10550 (new_n3874_, not_new_n1576__138412872010, not_new_n637__490);
  not g_10551 (new_n9181_, new_n8891_);
  not g_10552 (not_new_n990_, new_n990_);
  not g_10553 (not_new_n8106__1, new_n8106_);
  not g_10554 (not_new_n1164__0, new_n1164_);
  or g_10555 (new_n2254_, not_new_n8911_, not_new_n1591__6782230728490);
  not g_10556 (not_new_n1599__57648010, new_n1599_);
  not g_10557 (not_new_n646__2, new_n646_);
  or g_10558 (new_n10339_, not_new_n10337_, not_new_n10110__0);
  or g_10559 (new_n8336_, not_new_n626__797922662976120010, not_new_n8158_);
  or g_10560 (new_n6920_, not_new_n6825_, not_new_n6919_);
  or g_10561 (new_n10292_, not_new_n10291_, not_new_n10290_);
  not g_10562 (not_new_n9365__1, new_n9365_);
  not g_10563 (not_new_n604__168070, new_n604_);
  not g_10564 (not_new_n1588__0, new_n1588_);
  not g_10565 (not_pi053_1, pi053);
  not g_10566 (not_new_n964_, new_n964_);
  not g_10567 (not_new_n1063__7, new_n1063_);
  not g_10568 (not_new_n5747_, new_n5747_);
  not g_10569 (not_new_n4574_, new_n4574_);
  not g_10570 (new_n1584_, new_n931_);
  or g_10571 (new_n5622_, not_new_n1007__6, not_new_n5438_);
  not g_10572 (not_new_n9321_, new_n9321_);
  not g_10573 (not_new_n2838_, new_n2838_);
  or g_10574 (new_n4861_, not_new_n4841__1, not_new_n4765__1);
  or g_10575 (new_n10323_, not_new_n9903_, not_new_n645__113988951853731430);
  not g_10576 (not_new_n7809_, new_n7809_);
  not g_10577 (new_n1616_, new_n995_);
  not g_10578 (not_new_n2150_, new_n2150_);
  or g_10579 (new_n1698_, not_po296_19773267430, not_pi010_0);
  not g_10580 (not_new_n1061__2326305139872070, new_n1061_);
  or g_10581 (new_n2200_, not_new_n594__19773267430, not_new_n9966_);
  or g_10582 (new_n9687_, not_new_n9644_, not_new_n9512__0);
  or g_10583 (new_n7217_, not_new_n731_, not_new_n7034_);
  or g_10584 (new_n8788_, not_new_n1161__0, not_new_n8649_);
  and g_10585 (new_n9474_, new_n9642_, new_n9507_);
  not g_10586 (not_pi007, pi007);
  or g_10587 (new_n6481_, not_new_n632__403536070, not_new_n6483_);
  or g_10588 (new_n6737_, not_new_n6505_, not_new_n1603__24010);
  not g_10589 (not_new_n8696_, new_n8696_);
  not g_10590 (not_new_n4486_, new_n4486_);
  not g_10591 (not_new_n1008__6, new_n1008_);
  and g_10592 (new_n1416_, new_n1011_, new_n607_);
  and g_10593 (new_n1274_, new_n2005_, new_n2006_);
  or g_10594 (new_n8346_, not_new_n8149_, not_new_n637__138412872010);
  not g_10595 (not_new_n5047_, new_n5047_);
  not g_10596 (not_new_n2129_, new_n2129_);
  not g_10597 (new_n4834_, new_n4783_);
  or g_10598 (new_n10249_, not_new_n9877_, not_new_n1045__273687473400809163430);
  or g_10599 (new_n9746_, not_new_n9744_, not_new_n9745_);
  not g_10600 (not_new_n619__7, new_n619_);
  not g_10601 (not_new_n5179_, new_n5179_);
  not g_10602 (not_new_n7942_, new_n7942_);
  not g_10603 (new_n8115_, new_n1031_);
  or g_10604 (new_n1760_, not_new_n1728__16284135979104490, not_pi074);
  not g_10605 (not_new_n6305_, new_n6305_);
  not g_10606 (new_n8627_, new_n1071_);
  or g_10607 (po060, key_gate_109, not_new_n1187_);
  not g_10608 (not_new_n1536__57648010, new_n1536_);
  not g_10609 (not_new_n4758_, new_n4758_);
  not g_10610 (not_new_n5260_, new_n5260_);
  or g_10611 (new_n8989_, new_n631_, new_n1043_);
  and g_10612 (new_n8798_, new_n8990_, new_n8989_);
  not g_10613 (new_n6248_, new_n1605_);
  not g_10614 (not_new_n581__1070069044235980333563563003849377848070, new_n581_);
  or g_10615 (or_not_new_n2110__not_new_n2111_, not_new_n2110_, not_new_n2111_);
  or g_10616 (new_n6036_, not_new_n5814_, not_new_n5915_);
  not g_10617 (not_new_n1580__138412872010, new_n1580_);
  or g_10618 (new_n8334_, not_new_n1055__6782230728490, not_new_n8155_);
  not g_10619 (not_new_n3135_, new_n3135_);
  not g_10620 (not_new_n7630_, new_n7630_);
  not g_10621 (not_new_n5087_, new_n5087_);
  or g_10622 (new_n2836_, not_new_n994__3430, not_new_n4123__1);
  or g_10623 (new_n10129_, new_n1603_, new_n639_);
  or g_10624 (new_n3872_, not_new_n633__490, not_new_n1576__19773267430);
  not g_10625 (not_new_n3133_, new_n3133_);
  not g_10626 (not_new_n1071__24010, new_n1071_);
  or g_10627 (new_n4130_, not_new_n4211_, not_new_n4212_);
  not g_10628 (not_new_n2961_, new_n2961_);
  or g_10629 (new_n2569_, not_pi253, not_po296_657123623635342801395430);
  not g_10630 (not_new_n8454_, new_n8454_);
  not g_10631 (not_new_n3951_, new_n3951_);
  not g_10632 (not_new_n589__138412872010, new_n589_);
  not g_10633 (not_new_n6816_, new_n6816_);
  and g_10634 (and_new_n2667__new_n2668_, new_n2668_, new_n2667_);
  not g_10635 (not_pi190_0, pi190);
  not g_10636 (not_new_n3311__1, new_n3311_);
  or g_10637 (or_or_not_new_n1307__not_new_n1305__not_new_n2154_, not_new_n2154_, or_not_new_n1307__not_new_n1305_);
  not g_10638 (not_new_n10029__3, new_n10029_);
  not g_10639 (not_new_n599__10, new_n599_);
  not g_10640 (not_new_n7587_, new_n7587_);
  not g_10641 (not_new_n589__1577753820348458066150427430, new_n589_);
  or g_10642 (or_or_not_new_n1996__not_new_n1997__not_new_n1999_, or_not_new_n1996__not_new_n1997_, not_new_n1999_);
  not g_10643 (not_new_n4105_, new_n4105_);
  or g_10644 (or_not_new_n2874__not_new_n2877_, not_new_n2877_, not_new_n2874_);
  or g_10645 (or_or_not_new_n2567__not_new_n2571__not_new_n1429_, or_not_new_n2567__not_new_n2571_, not_new_n1429_);
  and g_10646 (and_new_n2257__new_n2260_, new_n2257_, new_n2260_);
  or g_10647 (new_n3033_, not_new_n1600__2, not_new_n581__24010);
  not g_10648 (not_new_n5054_, new_n5054_);
  not g_10649 (not_new_n6648_, new_n6648_);
  not g_10650 (not_new_n697_, new_n697_);
  not g_10651 (not_new_n5781__0, new_n5781_);
  or g_10652 (new_n957_, not_new_n2039_, or_or_not_new_n1283__not_new_n1281__not_new_n2040_);
  not g_10653 (not_new_n7672_, new_n7672_);
  or g_10654 (or_or_not_new_n1339__not_new_n1337__not_new_n2306_, or_not_new_n1339__not_new_n1337_, not_new_n2306_);
  not g_10655 (not_new_n7599__0, new_n7599_);
  not g_10656 (not_new_n3315__8235430, new_n3315_);
  or g_10657 (new_n2408_, not_new_n600__10, not_new_n4136__0);
  not g_10658 (not_new_n625__1176490, new_n625_);
  not g_10659 (not_new_n1452_, new_n1452_);
  not g_10660 (not_new_n635__70, new_n635_);
  or g_10661 (new_n9294_, not_new_n9163_, not_new_n8899__3);
  or g_10662 (or_not_new_n2939__not_new_n1485_, not_new_n1485_, not_new_n2939_);
  not g_10663 (not_pi020, pi020);
  not g_10664 (not_new_n7899_, new_n7899_);
  and g_10665 (new_n8948_, new_n9275_, and_new_n8874__new_n9276_);
  not g_10666 (not_new_n5832_, new_n5832_);
  not g_10667 (not_new_n7205_, new_n7205_);
  not g_10668 (not_new_n1051__19773267430, new_n1051_);
  or g_10669 (new_n8175_, not_new_n8362_, not_new_n8422_);
  not g_10670 (not_new_n581__225393402906922580878632490, new_n581_);
  not g_10671 (not_new_n8368__0, new_n8368_);
  not g_10672 (not_new_n1002__4, new_n1002_);
  or g_10673 (new_n3867_, not_new_n645__70, not_new_n6443__403536070);
  not g_10674 (not_new_n4837__1, new_n4837_);
  not g_10675 (not_new_n1279_, new_n1279_);
  xnor g_10676 (key_gate_73, key_73, new_n1672_);
  or g_10677 (new_n9154_, not_new_n8982__0, not_new_n9014_);
  or g_10678 (or_or_not_new_n1563__not_new_n2474__not_new_n1395_, not_new_n1395_, or_not_new_n1563__not_new_n2474_);
  or g_10679 (new_n3258_, not_new_n3184__5, not_new_n628__8);
  not g_10680 (not_new_n4321__0, new_n4321_);
  not g_10681 (not_new_n3554_, new_n3554_);
  not g_10682 (not_pi258_0, pi258);
  or g_10683 (new_n8846_, not_new_n9026_, not_new_n8930_);
  or g_10684 (or_or_not_new_n2892__not_new_n2895__not_new_n2894_, or_not_new_n2892__not_new_n2895_, not_new_n2894_);
  or g_10685 (new_n6808_, not_new_n6635__3, not_new_n6599_);
  or g_10686 (or_not_new_n7939__not_new_n7913_, not_new_n7913_, not_new_n7939_);
  or g_10687 (new_n3582_, not_pi157_0, not_new_n1538__2326305139872070);
  or g_10688 (po121, not_new_n3421_, not_new_n3420_);
  and g_10689 (new_n1421_, new_n2530_, new_n2532_);
  not g_10690 (not_new_n3440_, new_n3440_);
  or g_10691 (new_n2248_, not_new_n601__968890104070, not_new_n629__0);
  or g_10692 (new_n4895_, not_new_n4807__1, not_new_n4825__1);
  not g_10693 (not_pi027_0, pi027);
  or g_10694 (new_n2165_, not_new_n1604_, not_new_n1588__2824752490);
  or g_10695 (new_n8351_, not_new_n1065__968890104070, not_new_n8162__0);
  or g_10696 (new_n8384_, not_new_n8169__0, not_new_n8284_);
  buf g_10697 (po041, pi223);
  not g_10698 (not_new_n9186__0, new_n9186_);
  not g_10699 (not_new_n3499_, new_n3499_);
  or g_10700 (new_n1751_, not_pi067, not_new_n1728__403536070);
  not g_10701 (not_new_n5172_, new_n5172_);
  not g_10702 (not_new_n1039__273687473400809163430, new_n1039_);
  not g_10703 (not_new_n2712_, new_n2712_);
  not g_10704 (not_new_n1570_, new_n1570_);
  not g_10705 (not_new_n9828_, new_n9828_);
  not g_10706 (not_new_n1037__19773267430, new_n1037_);
  or g_10707 (new_n9120_, not_new_n9119_, not_new_n8947_);
  or g_10708 (new_n2404_, not_new_n9867__0, not_new_n599__9);
  and g_10709 (new_n596_, pi275, key_gate_77);
  or g_10710 (new_n9743_, not_new_n9556__0, not_new_n9741_);
  not g_10711 (new_n8357_, new_n8267_);
  not g_10712 (not_new_n1035__8, new_n1035_);
  not g_10713 (not_new_n9422__0, new_n9422_);
  not g_10714 (not_new_n7275_, new_n7275_);
  not g_10715 (not_new_n1602__168070, new_n1602_);
  or g_10716 (new_n3706_, not_pi239, not_new_n989__47475615099430);
  not g_10717 (not_pi038, pi038);
  and g_10718 (and_new_n2637__new_n2638_, new_n2638_, new_n2637_);
  not g_10719 (not_new_n3310__1176490, new_n3310_);
  not g_10720 (not_new_n3699_, new_n3699_);
  not g_10721 (not_new_n4137_, new_n4137_);
  or g_10722 (new_n4363_, not_new_n4304_, not_new_n4360_);
  not g_10723 (not_new_n3185__138412872010, new_n3185_);
  not g_10724 (not_new_n4206_, new_n4206_);
  not g_10725 (not_new_n1538__6782230728490, new_n1538_);
  or g_10726 (new_n6716_, not_new_n638__19773267430, not_new_n6519_);
  or g_10727 (new_n3452_, not_new_n1536__968890104070, not_pi022_0);
  not g_10728 (not_new_n1027__332329305696010, new_n1027_);
  or g_10729 (or_or_not_new_n1566__not_new_n2489__not_new_n1401_, or_not_new_n1566__not_new_n2489_, not_new_n1401_);
  and g_10730 (new_n5509_, new_n5652_, new_n5653_);
  not g_10731 (not_new_n2894_, new_n2894_);
  not g_10732 (not_new_n3420_, new_n3420_);
  not g_10733 (not_new_n8943_, new_n8943_);
  or g_10734 (new_n7951_, not_new_n7800_, not_new_n7734_);
  or g_10735 (new_n6108_, not_new_n631__403536070, not_new_n5742__2);
  not g_10736 (not_new_n4543_, new_n4543_);
  not g_10737 (not_new_n5180_, new_n5180_);
  not g_10738 (not_pi002_0, pi002);
  not g_10739 (not_new_n5106_, new_n5106_);
  not g_10740 (not_new_n1008_, new_n1008_);
  and g_10741 (and_new_n9696__new_n9695_, new_n9696_, new_n9695_);
  or g_10742 (new_n5268_, or_not_new_n5095__1_not_new_n4899__1, not_new_n4898__2);
  and g_10743 (new_n4143_, pi273, pi267);
  not g_10744 (new_n10231_, new_n10024_);
  not g_10745 (new_n4929_, new_n1043_);
  or g_10746 (or_not_new_n3136__not_new_n3137_, not_new_n3137_, not_new_n3136_);
  or g_10747 (new_n5950_, not_new_n5740__0, not_new_n5942_);
  not g_10748 (not_new_n5611_, new_n5611_);
  or g_10749 (new_n10086_, not_new_n1037__16284135979104490, not_new_n632__39098210485829880490);
  or g_10750 (new_n3405_, not_pi097_0, not_new_n1537_);
  not g_10751 (new_n10148_, new_n10015_);
  not g_10752 (not_new_n2874_, new_n2874_);
  not g_10753 (not_new_n1538__3430, new_n1538_);
  or g_10754 (new_n5336_, not_new_n5205_, not_new_n5334_);
  not g_10755 (not_new_n9909__0, new_n9909_);
  or g_10756 (new_n6212_, not_new_n636__8235430, not_new_n5790__0);
  or g_10757 (new_n7385_, not_new_n7360__1, not_new_n740__1);
  not g_10758 (not_new_n1364_, new_n1364_);
  not g_10759 (not_new_n1844_, new_n1844_);
  not g_10760 (not_new_n1600__9, new_n1600_);
  not g_10761 (not_new_n1014__3, new_n1014_);
  not g_10762 (not_new_n601__0, new_n601_);
  or g_10763 (new_n3090_, not_new_n581__273687473400809163430, not_new_n648__6);
  or g_10764 (new_n8782_, not_new_n1598__2824752490, not_new_n8657_);
  or g_10765 (or_or_not_new_n6340__not_new_n6341__not_new_n6342_, or_not_new_n6340__not_new_n6341_, not_new_n6342_);
  or g_10766 (new_n2239_, not_new_n622_, not_new_n593__968890104070);
  not g_10767 (not_new_n1017__2, new_n1017_);
  and g_10768 (new_n9344_, new_n9650_, new_n9648_);
  not g_10769 (not_new_n4127__1, new_n4127_);
  not g_10770 (not_new_n1583__138412872010, new_n1583_);
  or g_10771 (new_n8015_, not_new_n7628__0, not_new_n1602__8235430);
  or g_10772 (new_n3702_, not_new_n989__968890104070, not_pi237);
  not g_10773 (not_new_n7415__1, new_n7415_);
  or g_10774 (new_n3216_, not_new_n1604__4, not_new_n3185__24010);
  or g_10775 (po182, not_new_n1347_, not_new_n1348_);
  not g_10776 (not_new_n5954_, new_n5954_);
  not g_10777 (not_new_n4258_, new_n4258_);
  not g_10778 (not_new_n605__8, new_n605_);
  or g_10779 (new_n6004_, not_new_n6001_, not_new_n6003_);
  not g_10780 (not_new_n2059_, new_n2059_);
  not g_10781 (not_new_n2509__57648010, new_n2509_);
  not g_10782 (not_new_n4520_, new_n4520_);
  not g_10783 (not_new_n4771__0, new_n4771_);
  not g_10784 (not_new_n5434__0, new_n5434_);
  or g_10785 (new_n8378_, not_new_n8377_, not_new_n8129_);
  or g_10786 (new_n1929_, not_new_n8101_, not_new_n1581__7);
  not g_10787 (not_new_n660_, new_n660_);
  and g_10788 (new_n8683_, new_n8719_, new_n8682_);
  not g_10789 (not_new_n5509_, new_n5509_);
  not g_10790 (not_new_n8105__0, new_n8105_);
  not g_10791 (not_new_n9692_, new_n9692_);
  not g_10792 (not_new_n1039__57648010, new_n1039_);
  or g_10793 (new_n4890_, not_new_n1059__8, not_new_n4739_);
  or g_10794 (new_n8003_, not_new_n7624__0, not_new_n622__19773267430);
  not g_10795 (not_new_n7472_, new_n7472_);
  or g_10796 (new_n5946_, not_new_n648__168070, not_new_n5914_);
  not g_10797 (not_new_n3184__10, new_n3184_);
  and g_10798 (new_n6356_, new_n6410_, new_n6416_);
  or g_10799 (new_n3564_, not_new_n1538__57648010, not_pi148_0);
  or g_10800 (new_n5905_, or_not_new_n6073__not_new_n6048_, not_new_n5978_);
  not g_10801 (not_new_n1603__0, new_n1603_);
  not g_10802 (not_new_n643__39098210485829880490, new_n643_);
  not g_10803 (not_new_n607__24010, new_n607_);
  not g_10804 (not_new_n1027__1176490, new_n1027_);
  and g_10805 (new_n1232_, and_and_new_n1801__new_n1804__new_n1802_, new_n1803_);
  xnor g_10806 (key_gate_46, not_new_n3996_, key_46);
  not g_10807 (not_pi004, pi004);
  not g_10808 (not_new_n9995_, new_n9995_);
  or g_10809 (new_n7338_, not_new_n7018__2, not_new_n6988__0);
  or g_10810 (new_n9706_, not_new_n9338_, not_new_n9427__1);
  or g_10811 (new_n1885_, not_new_n4115_, not_new_n585__6);
  not g_10812 (not_new_n7970_, new_n7970_);
  not g_10813 (not_new_n5433_, new_n5433_);
  not g_10814 (not_new_n8234_, new_n8234_);
  not g_10815 (not_new_n6500__0, new_n6500_);
  and g_10816 (new_n1352_, new_n2365_, and_new_n1541__new_n2366_);
  or g_10817 (new_n8919_, not_new_n9308_, not_new_n9309_);
  not g_10818 (not_new_n4973_, new_n4973_);
  not g_10819 (not_new_n5281_, new_n5281_);
  not g_10820 (not_new_n5604_, new_n5604_);
  or g_10821 (new_n10283_, not_new_n617__657123623635342801395430, not_new_n9943__0);
  not g_10822 (not_new_n9255_, new_n9255_);
  and g_10823 (new_n7154_, new_n7559_, new_n7558_);
  not g_10824 (not_new_n5126_, new_n5126_);
  or g_10825 (new_n2990_, not_new_n581__0, not_new_n1051__2);
  and g_10826 (and_new_n6373__new_n6398_, new_n6373_, new_n6398_);
  not g_10827 (new_n2000_, new_n644_);
  or g_10828 (or_not_new_n9704__not_new_n9705_, not_new_n9705_, not_new_n9704_);
  not g_10829 (not_new_n5831_, new_n5831_);
  not g_10830 (not_new_n1051__47475615099430, new_n1051_);
  not g_10831 (not_new_n1211_, new_n1211_);
  buf g_10832 (po037, pi227);
  or g_10833 (new_n7051_, not_new_n7388_, not_new_n7389_);
  not g_10834 (not_new_n9165_, new_n9165_);
  not g_10835 (not_new_n8361_, new_n8361_);
  not g_10836 (not_new_n3721_, new_n3721_);
  not g_10837 (not_new_n600__8235430, new_n600_);
  not g_10838 (not_new_n6677_, new_n6677_);
  not g_10839 (not_new_n3407_, new_n3407_);
  not g_10840 (not_pi198, pi198);
  not g_10841 (not_new_n590__4, new_n590_);
  or g_10842 (new_n2524_, not_new_n607_, not_new_n1012_);
  not g_10843 (not_new_n8152_, new_n8152_);
  or g_10844 (new_n7520_, not_new_n7433__1, not_new_n727__1);
  not g_10845 (not_new_n4984__0, new_n4984_);
  or g_10846 (new_n2436_, not_new_n4796__0, not_new_n597__168070);
  not g_10847 (not_new_n4123__0, new_n4123_);
  not g_10848 (not_new_n1584__24010, new_n1584_);
  and g_10849 (new_n6598_, new_n625_, new_n6507_);
  not g_10850 (not_new_n2922_, new_n2922_);
  not g_10851 (not_new_n628__2, new_n628_);
  or g_10852 (new_n6680_, not_new_n6479_, not_new_n6679_);
  not g_10853 (not_new_n7613__0, new_n7613_);
  not g_10854 (not_new_n7817_, new_n7817_);
  not g_10855 (not_new_n727_, new_n727_);
  not g_10856 (not_new_n1037__4, new_n1037_);
  not g_10857 (not_new_n1069__2, new_n1069_);
  not g_10858 (not_pi143, pi143);
  not g_10859 (not_new_n6802_, new_n6802_);
  not g_10860 (not_new_n7503_, new_n7503_);
  not g_10861 (not_new_n8845__1, new_n8845_);
  or g_10862 (new_n9103_, new_n617_, new_n1597_);
  not g_10863 (not_new_n9941_, new_n9941_);
  not g_10864 (not_new_n9797_, new_n9797_);
  not g_10865 (not_new_n8879__0, new_n8879_);
  or g_10866 (new_n3654_, not_pi213, not_new_n989_);
  or g_10867 (new_n2001_, not_new_n627__0, not_new_n601__10);
  not g_10868 (not_new_n8218_, new_n8218_);
  not g_10869 (not_new_n607__1176490, new_n607_);
  or g_10870 (new_n2564_, not_new_n607__3, not_new_n1016_);
  not g_10871 (not_new_n634__5585458640832840070, new_n634_);
  not g_10872 (not_new_n6834_, new_n6834_);
  or g_10873 (new_n9098_, not_new_n8987_, not_new_n8979_);
  not g_10874 (not_pi248_2, pi248);
  not g_10875 (not_new_n5259_, new_n5259_);
  not g_10876 (not_pi171_2, pi171);
  not g_10877 (not_new_n1343_, new_n1343_);
  or g_10878 (or_or_not_new_n2129__not_new_n2130__not_new_n2132_, not_new_n2132_, or_not_new_n2129__not_new_n2130_);
  or g_10879 (new_n5489_, not_new_n5689_, not_new_n5690_);
  or g_10880 (or_not_new_n1479__not_new_n1480_, not_new_n1479_, not_new_n1480_);
  not g_10881 (not_new_n612__6, new_n612_);
  not g_10882 (not_new_n4808__0, new_n4808_);
  or g_10883 (new_n2498_, not_new_n599__16284135979104490, not_new_n9960__0);
  or g_10884 (new_n3754_, not_new_n1601__6, not_new_n630__10);
  or g_10885 (new_n4452_, not_new_n4717_, not_new_n4716_);
  not g_10886 (not_new_n9488_, new_n9488_);
  or g_10887 (new_n5418_, not_new_n1055__10, not_new_n4965_);
  or g_10888 (new_n6372_, not_new_n6304_, not_new_n619__490);
  not g_10889 (not_new_n1049__24010, new_n1049_);
  or g_10890 (new_n3945_, not_new_n3970_, not_new_n4017_);
  not g_10891 (not_new_n9009_, new_n9009_);
  not g_10892 (not_pi159, pi159);
  not g_10893 (not_new_n645__113988951853731430, new_n645_);
  not g_10894 (not_new_n639__968890104070, new_n639_);
  not g_10895 (not_new_n601__2326305139872070, new_n601_);
  not g_10896 (not_new_n4843_, new_n4843_);
  not g_10897 (not_new_n6758_, new_n6758_);
  not g_10898 (not_po296_17984650426474121466202803405696493492512490, po296);
  not g_10899 (not_new_n6974__138412872010, new_n6974_);
  not g_10900 (not_new_n10006__0, new_n10006_);
  or g_10901 (new_n2870_, not_new_n629__2, not_new_n604__24010);
  not g_10902 (not_new_n7351__0, new_n7351_);
  not g_10903 (not_new_n6503__2, new_n6503_);
  xnor g_10904 (key_gate_89, key_89, not_new_n3985_);
  or g_10905 (new_n1780_, not_new_n1588__0, not_new_n1031__1);
  or g_10906 (new_n701_, not_new_n3075_, not_new_n1525_);
  and g_10907 (new_n1566_, new_n3645_, new_n3644_);
  or g_10908 (new_n8558_, not_new_n1067__57648010, not_new_n8147__0);
  and g_10909 (and_new_n5084__new_n5345_, new_n5345_, new_n5084_);
  not g_10910 (not_new_n3100_, new_n3100_);
  not g_10911 (not_new_n9826_, new_n9826_);
  or g_10912 (new_n6646_, not_new_n6634__0, not_new_n6633_);
  not g_10913 (not_new_n586__1176490, new_n586_);
  or g_10914 (new_n2378_, not_new_n4117__0, not_new_n600__4);
  not g_10915 (not_new_n3984_, new_n3984_);
  not g_10916 (not_new_n7561_, new_n7561_);
  and g_10917 (new_n4471_, new_n4584_, new_n4652_);
  or g_10918 (new_n6642_, not_new_n6813_, not_new_n6709_);
  not g_10919 (not_new_n4004_, new_n4004_);
  not g_10920 (not_new_n1763_, new_n1763_);
  or g_10921 (new_n4995_, not_new_n5279_, not_new_n5188_);
  not g_10922 (new_n5579_, new_n5474_);
  or g_10923 (new_n1803_, not_new_n4748_, not_new_n591__1);
  or g_10924 (new_n5569_, not_new_n5674_, not_new_n1014__5);
  not g_10925 (not_new_n6815_, new_n6815_);
  or g_10926 (new_n3892_, not_new_n3894_, not_new_n10228_);
  or g_10927 (new_n9132_, new_n637_, new_n1065_);
  or g_10928 (po216, not_new_n1420_, or_or_not_new_n2527__not_new_n2531__not_new_n1421_);
  not g_10929 (not_new_n7853_, new_n7853_);
  or g_10930 (new_n7931_, not_new_n7709_, not_new_n7754__3);
  and g_10931 (new_n1390_, new_n2461_, new_n2460_);
  not g_10932 (not_new_n7583_, new_n7583_);
  and g_10933 (new_n4911_, new_n5193_, new_n5199_);
  not g_10934 (not_new_n1631__70, key_gate_76);
  not g_10935 (not_new_n9179_, new_n9179_);
  not g_10936 (not_new_n641__5, new_n641_);
  or g_10937 (new_n3255_, not_new_n1041__5, not_new_n589__273687473400809163430);
  not g_10938 (not_new_n4829_, new_n4829_);
  not g_10939 (not_new_n7549_, new_n7549_);
  not g_10940 (not_new_n10049_, new_n10049_);
  not g_10941 (not_new_n7135_, new_n7135_);
  not g_10942 (not_new_n10011_, new_n10011_);
  not g_10943 (not_new_n3184__6782230728490, new_n3184_);
  not g_10944 (not_new_n6443__332329305696010, new_n6443_);
  not g_10945 (not_new_n637__490, new_n637_);
  or g_10946 (new_n3871_, not_new_n633__70, not_new_n6443__19773267430);
  or g_10947 (new_n7115_, not_new_n7176_, not_new_n7071_);
  not g_10948 (not_new_n1071__1176490, new_n1071_);
  or g_10949 (new_n6931_, not_new_n6637_, not_new_n6605_);
  or g_10950 (new_n2499_, not_new_n1607__0, not_new_n598__16284135979104490);
  not g_10951 (not_new_n619_, new_n619_);
  not g_10952 (not_new_n3697_, new_n3697_);
  or g_10953 (new_n7724_, not_new_n8029_, not_new_n8028_);
  or g_10954 (new_n5603_, not_new_n5446_, not_pi136_2);
  not g_10955 (not_new_n5905__1, new_n5905_);
  not g_10956 (not_new_n6027_, new_n6027_);
  not g_10957 (not_new_n1612__0, new_n1612_);
  not g_10958 (new_n6979_, new_n740_);
  not g_10959 (not_new_n745_, new_n745_);
  or g_10960 (new_n10058_, not_new_n1047__332329305696010, not_new_n10055_);
  not g_10961 (not_pi123_0, pi123);
  not g_10962 (not_new_n928__113988951853731430, new_n928_);
  not g_10963 (not_new_n6913_, new_n6913_);
  not g_10964 (not_new_n3875_, new_n3875_);
  not g_10965 (not_new_n4128_, new_n4128_);
  not g_10966 (not_new_n6183_, new_n6183_);
  not g_10967 (not_pi271_0, pi271);
  not g_10968 (not_new_n4733_, new_n4733_);
  not g_10969 (not_new_n640__57648010, new_n640_);
  or g_10970 (new_n5158_, not_new_n5078_, not_new_n4907_);
  not g_10971 (not_new_n9486_, new_n9486_);
  not g_10972 (not_new_n8342_, new_n8342_);
  or g_10973 (po125, not_new_n3440_, not_new_n3441_);
  or g_10974 (new_n766_, not_new_n3189_, not_new_n3188_);
  not g_10975 (not_new_n7619_, new_n7619_);
  not g_10976 (not_new_n638__16284135979104490, new_n638_);
  or g_10977 (new_n4593_, not_new_n4591_, not_new_n4541_);
  not g_10978 (not_new_n9938_, new_n9938_);
  or g_10979 (new_n5696_, not_new_n5514_, not_new_n5515__0);
  or g_10980 (or_not_new_n7463__not_new_n7312_, not_new_n7312_, not_new_n7463_);
  not g_10981 (new_n7168_, new_n7145_);
  not g_10982 (new_n5750_, new_n1037_);
  not g_10983 (not_new_n2912_, new_n2912_);
  or g_10984 (new_n2904_, not_new_n595__57648010, not_new_n7061_);
  not g_10985 (not_new_n6579_, new_n6579_);
  not g_10986 (not_new_n638__113988951853731430, new_n638_);
  or g_10987 (new_n10202_, not_new_n10083_, not_new_n10041__0);
  or g_10988 (new_n2803_, not_new_n1604__1, not_new_n613__1);
  not g_10989 (not_new_n6992_, new_n6992_);
  not g_10990 (not_new_n1196_, new_n1196_);
  or g_10991 (new_n9008_, not_new_n9005_, not_new_n1047__2824752490);
  not g_10992 (not_new_n8273_, new_n8273_);
  not g_10993 (not_new_n1069__19773267430, new_n1069_);
  not g_10994 (not_new_n1598__19773267430, new_n1598_);
  or g_10995 (new_n8064_, not_new_n1057__57648010, not_new_n7653__0);
  not g_10996 (not_new_n1616__2824752490, new_n1616_);
  not g_10997 (not_new_n9119_, new_n9119_);
  not g_10998 (not_new_n627__138412872010, new_n627_);
  or g_10999 (new_n5250_, not_new_n5054_, not_new_n5249_);
  and g_11000 (new_n615_, new_n1227_, new_n584_);
  or g_11001 (new_n3838_, not_new_n624__490, not_new_n1576__4);
  or g_11002 (or_or_not_new_n1763__not_new_n1764__not_new_n1766_, or_not_new_n1763__not_new_n1764_, not_new_n1766_);
  not g_11003 (not_new_n5506_, new_n5506_);
  not g_11004 (not_new_n6781_, new_n6781_);
  not g_11005 (not_new_n8641_, new_n8641_);
  or g_11006 (new_n9796_, not_new_n9496_, not_new_n9497_);
  not g_11007 (not_new_n4770__0, new_n4770_);
  not g_11008 (not_new_n2173_, new_n2173_);
  or g_11009 (new_n5393_, not_new_n5391_, not_new_n5392_);
  not g_11010 (not_new_n4790_, new_n4790_);
  not g_11011 (not_new_n8438_, new_n8438_);
  not g_11012 (not_new_n1534__6782230728490, key_gate_5);
  and g_11013 (new_n1417_, new_n2515_, and_and_new_n2517__new_n2518__new_n2516_);
  or g_11014 (new_n767_, not_new_n3190_, not_new_n3191_);
  not g_11015 (not_new_n5195_, new_n5195_);
  or g_11016 (or_not_new_n1027__not_new_n1028__0, not_new_n1027_, not_new_n1028__0);
  not g_11017 (new_n1583_, new_n929_);
  not g_11018 (not_pi138_3, pi138);
  not g_11019 (new_n7643_, new_n1063_);
  or g_11020 (new_n2674_, not_new_n607__24010, not_new_n1009_);
  not g_11021 (not_new_n628__2824752490, new_n628_);
  or g_11022 (or_not_new_n3161__not_new_n3160_, not_new_n3160_, not_new_n3161_);
  not g_11023 (not_new_n1019__3, new_n1019_);
  not g_11024 (not_new_n7292_, new_n7292_);
  or g_11025 (po143, not_new_n3512_, not_new_n3513_);
  and g_11026 (new_n7734_, new_n7949_, new_n7948_);
  or g_11027 (new_n4336_, not_new_n4238_, not_new_n706_);
  or g_11028 (new_n7886_, not_new_n7759__0, not_new_n7837_);
  not g_11029 (not_new_n4577__0, new_n4577_);
  or g_11030 (new_n9901_, not_new_n9982_, not_new_n10071_);
  or g_11031 (new_n10093_, new_n626_, new_n1053_);
  or g_11032 (new_n6545_, not_new_n1602__24010, not_new_n6504_);
  or g_11033 (new_n4124_, not_new_n4199_, not_new_n4200_);
  and g_11034 (new_n1445_, new_n2650_, and_new_n2652__new_n2651_);
  not g_11035 (not_new_n2001_, new_n2001_);
  or g_11036 (new_n9575_, not_new_n9462_, not_new_n9573_);
  or g_11037 (new_n1948_, not_new_n8190_, not_new_n1581__8);
  not g_11038 (new_n2266_, new_n617_);
  not g_11039 (not_new_n6511__0, new_n6511_);
  or g_11040 (new_n4455_, not_new_n4606_, not_new_n4607_);
  or g_11041 (new_n1643_, not_pi036, not_new_n1631__2);
  not g_11042 (not_new_n7510_, new_n7510_);
  or g_11043 (new_n3554_, not_new_n1538__3430, not_pi143_0);
  not g_11044 (not_new_n5194_, new_n5194_);
  buf g_11045 (po027, pi237);
  or g_11046 (or_not_new_n1825__not_new_n1826_, not_new_n1825_, not_new_n1826_);
  or g_11047 (new_n3776_, not_new_n1059__6, not_new_n644__10);
  not g_11048 (not_new_n3311__2, new_n3311_);
  not g_11049 (not_new_n6974__2, new_n6974_);
  or g_11050 (new_n8234_, not_new_n8548_, not_new_n8549_);
  or g_11051 (new_n3066_, not_new_n1174_, not_new_n1027__16284135979104490);
  not g_11052 (not_new_n624__1176490, new_n624_);
  or g_11053 (new_n953_, not_new_n1963_, or_or_not_new_n1267__not_new_n1265__not_new_n1964_);
  or g_11054 (new_n8733_, not_new_n8725_, not_new_n8658_);
  not g_11055 (not_new_n9973__0, new_n9973_);
  not g_11056 (not_new_n8697_, new_n8697_);
  not g_11057 (not_new_n9960_, new_n9960_);
  or g_11058 (new_n8200_, not_new_n8590_, not_new_n8589_);
  not g_11059 (not_new_n10022_, new_n10022_);
  not g_11060 (not_new_n6978__0, new_n6978_);
  not g_11061 (not_new_n2960_, new_n2960_);
  not g_11062 (not_new_n9070_, new_n9070_);
  or g_11063 (new_n6789_, not_new_n6640__1, not_new_n6582_);
  not g_11064 (not_new_n3688_, new_n3688_);
  not g_11065 (not_new_n8967_, new_n8967_);
  or g_11066 (new_n9568_, not_new_n9358__1, not_new_n9361__0);
  or g_11067 (new_n663_, or_not_new_n3152__not_new_n3151_, not_new_n3150_);
  not g_11068 (new_n7293_, new_n7017_);
  not g_11069 (not_new_n634__6782230728490, new_n634_);
  or g_11070 (or_not_new_n6354__not_new_n6373__8, not_new_n6354_, not_new_n6373__8);
  not g_11071 (not_po296_57648010, po296);
  not g_11072 (not_new_n6901_, new_n6901_);
  or g_11073 (new_n10244_, not_new_n10006__0, not_new_n10199_);
  not g_11074 (not_new_n6581_, new_n6581_);
  not g_11075 (not_new_n2908_, new_n2908_);
  not g_11076 (not_new_n9915_, new_n9915_);
  not g_11077 (new_n5457_, pi141);
  not g_11078 (not_new_n1016__1, new_n1016_);
  and g_11079 (new_n8808_, new_n9086_, new_n8805_);
  not g_11080 (not_new_n994__0, new_n994_);
  not g_11081 (not_new_n7992_, new_n7992_);
  or g_11082 (new_n9142_, not_new_n8900_, not_new_n9141_);
  not g_11083 (not_new_n633__10, new_n633_);
  or g_11084 (new_n7975_, not_new_n7610__1, not_new_n628__47475615099430);
  not g_11085 (not_new_n4117__2, new_n4117_);
  not g_11086 (not_new_n3564_, new_n3564_);
  and g_11087 (new_n4300_, new_n4349_, and_new_n4348__new_n4301_);
  and g_11088 (new_n6446_, new_n6650_, new_n6703_);
  not g_11089 (not_new_n6259_, new_n6259_);
  not g_11090 (not_pi046, pi046);
  and g_11091 (new_n1254_, new_n1911_, new_n1910_);
  not g_11092 (not_new_n4133__0, new_n4133_);
  not g_11093 (not_new_n4120__1, new_n4120_);
  not g_11094 (not_pi098_0, pi098);
  or g_11095 (new_n2716_, not_new_n604_, not_new_n643__2);
  and g_11096 (new_n9998_, new_n10319_, and_new_n9905__new_n10320_);
  not g_11097 (not_new_n9568_, new_n9568_);
  not g_11098 (not_new_n3913_, new_n3913_);
  not g_11099 (new_n4079_, pi256);
  not g_11100 (not_new_n599__19773267430, new_n599_);
  and g_11101 (new_n1518_, new_n3053_, and_new_n3055__new_n998_);
  and g_11102 (new_n1187_, new_n1652_, new_n1650_);
  not g_11103 (not_new_n6294_, new_n6294_);
  or g_11104 (new_n5819_, not_new_n6173_, not_new_n6174_);
  or g_11105 (new_n7251_, not_new_n722_, not_new_n7041_);
  not g_11106 (not_new_n6317__0, new_n6317_);
  not g_11107 (not_new_n602__1176490, new_n602_);
  not g_11108 (not_new_n643__5585458640832840070, new_n643_);
  not g_11109 (new_n8993_, new_n8971_);
  not g_11110 (not_new_n1580__57648010, new_n1580_);
  not g_11111 (not_new_n7023_, new_n7023_);
  not g_11112 (not_new_n10163_, new_n10163_);
  not g_11113 (not_new_n9505_, new_n9505_);
  not g_11114 (new_n3993_, pi034);
  or g_11115 (new_n7559_, not_new_n6999__0, not_new_n7033__0);
  not g_11116 (not_new_n8384_, new_n8384_);
  not g_11117 (not_new_n1613__0, new_n1613_);
  not g_11118 (not_new_n646__403536070, new_n646_);
  or g_11119 (new_n3263_, not_new_n589__657123623635342801395430, not_new_n1598__5);
  not g_11120 (not_new_n8975_, new_n8975_);
  not g_11121 (not_new_n595__0, new_n595_);
  or g_11122 (new_n5310_, not_new_n1043__10, not_new_n4927_);
  or g_11123 (new_n3581_, not_new_n1612__332329305696010, not_new_n2299__0);
  not g_11124 (not_new_n8284_, new_n8284_);
  not g_11125 (not_new_n608_, new_n608_);
  not g_11126 (not_new_n635__168070, new_n635_);
  or g_11127 (new_n3361_, not_pi033_1, not_new_n1534__138412872010);
  or g_11128 (new_n6430_, not_new_n6347_, not_new_n6346_);
  or g_11129 (new_n5130_, not_new_n4946_, not_new_n5129_);
  or g_11130 (new_n3753_, not_new_n3752_, not_new_n3751_);
  not g_11131 (not_new_n9951__1, new_n9951_);
  not g_11132 (not_new_n3831_, new_n3831_);
  not g_11133 (not_new_n4134__1, new_n4134_);
  not g_11134 (not_new_n621__39098210485829880490, new_n621_);
  and g_11135 (new_n1521_, and_new_n3064__new_n998_, new_n3062_);
  not g_11136 (not_new_n6312_, new_n6312_);
  or g_11137 (new_n4146_, or_not_pi257_3_not_pi260_3, not_pi269_3);
  not g_11138 (not_new_n638__3, new_n638_);
  not g_11139 (not_new_n1067__47475615099430, new_n1067_);
  and g_11140 (new_n8090_, new_n8089_, new_n8087_);
  and g_11141 (new_n9452_, new_n628_, new_n1039_);
  not g_11142 (not_new_n6443__8, new_n6443_);
  or g_11143 (new_n2487_, not_new_n618__1, not_new_n603__332329305696010);
  not g_11144 (not_new_n9813_, new_n9813_);
  not g_11145 (not_new_n7772_, new_n7772_);
  not g_11146 (not_new_n1069__168070, new_n1069_);
  or g_11147 (new_n8016_, not_new_n625__332329305696010, not_new_n7631__2);
  not g_11148 (new_n5544_, new_n5447_);
  or g_11149 (po059, key_gate_54, not_new_n1186_);
  or g_11150 (new_n9399_, not_new_n9589_, not_new_n9702_);
  not g_11151 (not_new_n3182_, new_n3182_);
  not g_11152 (not_new_n1645_, key_gate_67);
  or g_11153 (new_n924_, key_gate_112, key_gate_38);
  not g_11154 (not_new_n644__10, new_n644_);
  not g_11155 (new_n7252_, new_n7139_);
  or g_11156 (new_n10330_, not_new_n10329_, not_new_n10328_);
  and g_11157 (new_n9480_, and_new_n9511__new_n9839_, new_n9838_);
  not g_11158 (not_new_n6888_, new_n6888_);
  or g_11159 (new_n10262_, not_new_n10260_, not_new_n10261_);
  and g_11160 (new_n4299_, new_n4247_, new_n668_);
  not g_11161 (not_new_n2166_, new_n2166_);
  not g_11162 (not_new_n1043__332329305696010, new_n1043_);
  not g_11163 (not_new_n8049_, new_n8049_);
  and g_11164 (new_n5047_, new_n5182_, new_n5070_);
  or g_11165 (new_n5763_, not_new_n5911_, or_not_new_n6042__not_new_n5927_);
  not g_11166 (not_new_n940_, new_n940_);
  not g_11167 (not_new_n7159_, new_n7159_);
  not g_11168 (not_new_n6498__1, new_n6498_);
  not g_11169 (not_new_n636__19773267430, new_n636_);
  or g_11170 (new_n7489_, not_new_n7487_, not_new_n7488_);
  not g_11171 (not_new_n589__968890104070, new_n589_);
  not g_11172 (not_new_n6443__4, new_n6443_);
  and g_11173 (new_n1479_, new_n2811_, new_n2812_);
  not g_11174 (not_new_n610__4, new_n610_);
  or g_11175 (new_n9535_, not_new_n634__16284135979104490, not_new_n9534_);
  not g_11176 (not_new_n6647__0, new_n6647_);
  not g_11177 (not_new_n5779_, new_n5779_);
  not g_11178 (not_new_n10150_, new_n10150_);
  and g_11179 (new_n5715_, new_n5970_, new_n5969_);
  or g_11180 (new_n3367_, not_pi060_0, not_new_n1534__6782230728490);
  not g_11181 (not_new_n8275__0, new_n8275_);
  or g_11182 (new_n9750_, not_new_n9350_, not_new_n1037__332329305696010);
  or g_11183 (new_n8904_, not_new_n9200_, not_new_n9201_);
  and g_11184 (new_n1399_, new_n2483_, new_n2482_);
  not g_11185 (not_new_n1585__7, new_n1585_);
  or g_11186 (new_n9016_, not_new_n9015_, not_new_n8845__0);
  not g_11187 (not_new_n6917_, new_n6917_);
  not g_11188 (not_new_n1604__168070, new_n1604_);
  or g_11189 (new_n6882_, not_new_n6753_, not_new_n6625__1);
  not g_11190 (not_new_n598__57648010, new_n598_);
  or g_11191 (new_n9194_, not_new_n9193_, not_new_n9192_);
  or g_11192 (new_n8260_, not_new_n8139_, not_new_n8385_);
  not g_11193 (not_new_n7022__1, new_n7022_);
  not g_11194 (not_new_n8021_, new_n8021_);
  not g_11195 (not_new_n3315_, new_n3315_);
  not g_11196 (not_new_n1601__10, new_n1601_);
  not g_11197 (not_new_n624__168070, new_n624_);
  not g_11198 (not_new_n6609_, new_n6609_);
  or g_11199 (new_n620_, not_new_n2341_, or_not_new_n2339__not_new_n2340_);
  or g_11200 (new_n2080_, not_new_n1584__168070, not_new_n9445_);
  not g_11201 (not_pi158_0, pi158);
  and g_11202 (new_n8672_, new_n8607_, new_n1157_);
  not g_11203 (not_new_n3384__2, new_n3384_);
  or g_11204 (new_n1794_, not_new_n5820_, not_new_n1585__0);
  not g_11205 (not_new_n1039__70, new_n1039_);
  or g_11206 (new_n6983_, not_new_n7024_, not_new_n743_);
  or g_11207 (or_or_not_new_n1311__not_new_n1309__not_new_n2173_, or_not_new_n1311__not_new_n1309_, not_new_n2173_);
  and g_11208 (new_n6327_, new_n6232_, new_n6277_);
  or g_11209 (or_not_new_n2635__not_new_n2634_, not_new_n2634_, not_new_n2635_);
  not g_11210 (new_n5565_, new_n5462_);
  not g_11211 (not_new_n641__6, new_n641_);
  not g_11212 (not_new_n10207_, new_n10207_);
  not g_11213 (not_new_n3990__0, new_n3990_);
  not g_11214 (not_pi265, pi265);
  not g_11215 (not_new_n2878_, new_n2878_);
  not g_11216 (not_pi153, pi153);
  buf g_11217 (po022, pi242);
  or g_11218 (new_n5101_, not_new_n5081_, not_new_n1043__8);
  not g_11219 (not_new_n1047__2326305139872070, new_n1047_);
  or g_11220 (new_n1696_, key_gate_45, not_new_n596__2824752490);
  or g_11221 (new_n9634_, not_new_n9491__0, not_new_n1596__16284135979104490);
  not g_11222 (not_new_n1591__2824752490, new_n1591_);
  not g_11223 (not_new_n4791__0, new_n4791_);
  not g_11224 (not_new_n4969__0, new_n4969_);
  or g_11225 (new_n5261_, not_new_n4974__1, not_new_n5231_);
  not g_11226 (not_new_n1534__8235430, key_gate_5);
  not g_11227 (not_pi161_0, pi161);
  not g_11228 (not_new_n6706_, new_n6706_);
  or g_11229 (new_n2333_, not_new_n5008_, not_new_n1589__16284135979104490);
  not g_11230 (not_new_n6215_, new_n6215_);
  not g_11231 (not_new_n1055__138412872010, new_n1055_);
  not g_11232 (not_new_n2891_, new_n2891_);
  not g_11233 (not_new_n3586_, new_n3586_);
  or g_11234 (new_n3546_, not_pi139_0, not_new_n1538__9);
  not g_11235 (not_new_n7344_, new_n7344_);
  or g_11236 (new_n5477_, not_new_n5601_, not_new_n5600_);
  or g_11237 (po202, or_or_not_new_n1559__not_new_n2454__not_new_n1387_, not_new_n1388_);
  not g_11238 (not_new_n3994_, new_n3994_);
  or g_11239 (new_n5077_, not_new_n5158_, not_new_n5159_);
  not g_11240 (not_new_n5453_, new_n5453_);
  or g_11241 (new_n7950_, not_new_n7802_, not_new_n7735__3);
  or g_11242 (new_n753_, not_new_n3214_, not_new_n3215_);
  not g_11243 (not_new_n7483_, new_n7483_);
  not g_11244 (not_new_n1045__2824752490, new_n1045_);
  not g_11245 (not_new_n634__113988951853731430, new_n634_);
  not g_11246 (new_n3439_, new_n1047_);
  not g_11247 (not_new_n8443_, new_n8443_);
  or g_11248 (new_n9196_, not_new_n9194_, not_new_n9013__0);
  not g_11249 (not_new_n6585_, new_n6585_);
  not g_11250 (not_new_n621__10, new_n621_);
  not g_11251 (not_new_n5726_, new_n5726_);
  not g_11252 (not_new_n9899__0, new_n9899_);
  not g_11253 (not_new_n928__57648010, new_n928_);
  not g_11254 (not_new_n7144_, new_n7144_);
  or g_11255 (new_n3781_, not_new_n3409_, not_new_n1767_);
  or g_11256 (new_n10131_, new_n625_, new_n1602_);
  not g_11257 (not_new_n4490_, new_n4490_);
  or g_11258 (po201, not_new_n1386_, or_or_not_new_n1558__not_new_n2449__not_new_n1385_);
  not g_11259 (not_new_n593__168070, new_n593_);
  not g_11260 (not_new_n589__6, new_n589_);
  or g_11261 (new_n1801_, not_new_n594__0, not_new_n9953_);
  not g_11262 (not_new_n3310_, new_n3310_);
  and g_11263 (new_n9867_, new_n10197_, new_n10194_);
  or g_11264 (new_n5706_, not_new_n5454_, not_new_n5551_);
  not g_11265 (new_n4167_, new_n4096_);
  or g_11266 (new_n2132_, not_new_n585__403536070, not_new_n4127_);
  or g_11267 (new_n1833_, not_new_n1584__2, not_new_n9435_);
  and g_11268 (new_n8663_, new_n8767_, new_n8769_);
  not g_11269 (not_new_n3188_, new_n3188_);
  and g_11270 (new_n5062_, new_n5330_, new_n5331_);
  and g_11271 (and_new_n1953__new_n1956_, new_n1956_, new_n1953_);
  or g_11272 (new_n9747_, not_new_n9686_, not_new_n9485_);
  not g_11273 (not_new_n1588__2824752490, new_n1588_);
  not g_11274 (not_new_n3108_, new_n3108_);
  not g_11275 (not_new_n1035__70, new_n1035_);
  not g_11276 (not_new_n6348_, new_n6348_);
  not g_11277 (not_new_n5369_, new_n5369_);
  or g_11278 (new_n3295_, not_new_n589__21838143759917965991093122527538323430, not_new_n1055__5);
  not g_11279 (not_new_n8874_, new_n8874_);
  not g_11280 (not_new_n4170_, new_n4170_);
  or g_11281 (new_n1666_, not_new_n596__10, key_gate_16);
  not g_11282 (not_new_n9951_, new_n9951_);
  and g_11283 (and_new_n8983__new_n9311_, new_n9311_, new_n8983_);
  or g_11284 (new_n9213_, not_new_n9211_, not_new_n9212_);
  not g_11285 (not_new_n9096_, new_n9096_);
  or g_11286 (new_n2883_, not_new_n1057__1, not_new_n3311__70);
  not g_11287 (not_new_n4919_, new_n4919_);
  not g_11288 (not_new_n587__1176490, new_n587_);
  not g_11289 (not_new_n7002__1, new_n7002_);
  or g_11290 (new_n5707_, not_pi139_3, not_new_n5452__1);
  not g_11291 (not_new_n5930_, new_n5930_);
  not g_11292 (not_new_n1588__138412872010, new_n1588_);
  not g_11293 (not_new_n5713_, new_n5713_);
  not g_11294 (new_n8120_, new_n624_);
  or g_11295 (new_n3113_, not_new_n618__4, not_new_n3315__9);
  not g_11296 (not_new_n8238_, new_n8238_);
  or g_11297 (new_n9167_, not_new_n8798__1, or_not_new_n8799__0_not_new_n8996__0);
  not g_11298 (not_new_n1611__1176490, new_n1611_);
  or g_11299 (new_n1162_, not_new_n3854_, not_new_n3853_);
  not g_11300 (not_new_n6673__0, new_n6673_);
  not g_11301 (not_new_n1599__0, new_n1599_);
  not g_11302 (new_n7177_, new_n7115_);
  or g_11303 (new_n6782_, or_not_new_n6590__not_new_n6589_, not_new_n6745__0);
  or g_11304 (new_n6707_, not_new_n6447_, not_new_n6706_);
  not g_11305 (not_new_n1583__2326305139872070, new_n1583_);
  not g_11306 (not_new_n590__3, new_n590_);
  or g_11307 (new_n5951_, not_new_n5843_, not_new_n5950_);
  not g_11308 (not_new_n2057_, new_n2057_);
  not g_11309 (not_new_n3387__2, new_n3387_);
  or g_11310 (new_n2703_, or_not_new_n1470__not_new_n3824_, not_new_n3823_);
  not g_11311 (not_new_n1061__2824752490, new_n1061_);
  or g_11312 (new_n3435_, not_pi103_0, not_new_n1537__5);
  not g_11313 (not_new_n8323_, new_n8323_);
  not g_11314 (not_new_n2951_, new_n2951_);
  not g_11315 (not_new_n8388_, new_n8388_);
  or g_11316 (new_n9786_, not_new_n630__113988951853731430, not_new_n9414__0);
  not g_11317 (not_new_n604__8, new_n604_);
  not g_11318 (not_new_n8253__0, new_n8253_);
  not g_11319 (new_n8649_, new_n1598_);
  or g_11320 (new_n6860_, not_new_n6618_, not_new_n6663__0);
  or g_11321 (new_n2373_, not_new_n600__3, not_new_n4118__0);
  not g_11322 (not_new_n637__332329305696010, new_n637_);
  and g_11323 (new_n5054_, and_new_n5082__new_n5423_, new_n5422_);
  not g_11324 (not_new_n3174_, new_n3174_);
  not g_11325 (not_new_n5638_, new_n5638_);
  and g_11326 (new_n8085_, new_n8314_, new_n8077_);
  and g_11327 (new_n1308_, and_and_new_n2162__new_n2165__new_n2163_, new_n2164_);
  not g_11328 (not_new_n9556__0, new_n9556_);
  not g_11329 (not_new_n8010_, new_n8010_);
  not g_11330 (not_new_n7231_, new_n7231_);
  not g_11331 (new_n5768_, new_n629_);
  not g_11332 (not_new_n581__152867006319425761937651857692768264010, new_n581_);
  or g_11333 (new_n7111_, not_new_n7317_, not_new_n7322_);
  not g_11334 (not_new_n7006__0, new_n7006_);
  not g_11335 (not_new_n645__2824752490, new_n645_);
  not g_11336 (not_new_n925__0, new_n925_);
  or g_11337 (new_n4145_, or_or_not_pi269_2_not_pi248_2_not_pi257_2, not_pi260_2);
  and g_11338 (new_n6237_, new_n6372_, and_and_new_n6251__new_n6371__new_n1597_);
  not g_11339 (not_new_n5440__0, new_n5440_);
  not g_11340 (not_new_n9889__0, new_n9889_);
  not g_11341 (not_new_n3997_, new_n3997_);
  or g_11342 (or_not_new_n7047__0_not_new_n3369__0, not_new_n7047__0, not_new_n3369__0);
  not g_11343 (not_new_n5487__0, new_n5487_);
  not g_11344 (new_n4233_, new_n708_);
  or g_11345 (new_n6123_, not_new_n5883_, not_new_n5928__0);
  not g_11346 (not_new_n6688_, new_n6688_);
  not g_11347 (not_new_n1923_, new_n1923_);
  not g_11348 (not_new_n1825_, new_n1825_);
  not g_11349 (not_new_n4132_, new_n4132_);
  not g_11350 (not_new_n598__2824752490, new_n598_);
  or g_11351 (new_n7276_, not_new_n7240_, not_new_n7146__0);
  not g_11352 (not_new_n6026_, new_n6026_);
  not g_11353 (not_new_n5983_, new_n5983_);
  not g_11354 (new_n3321_, new_n999_);
  and g_11355 (new_n1464_, new_n3756_, and_and_new_n3750__new_n3753__new_n3759_);
  or g_11356 (new_n5591_, not_new_n1002__7, not_new_n5451__0);
  not g_11357 (not_new_n5110_, new_n5110_);
  not g_11358 (not_pi042_2, pi042);
  or g_11359 (new_n7227_, not_new_n7029_, not_new_n7226_);
  or g_11360 (new_n8497_, not_new_n8093_, or_not_new_n8172__0_not_new_n1596__138412872010);
  or g_11361 (new_n7260_, not_new_n7084_, not_new_n7139_);
  not g_11362 (not_new_n8889_, new_n8889_);
  or g_11363 (or_not_new_n4319__0_not_new_n713_, not_new_n4319__0, not_new_n713_);
  not g_11364 (not_pi044_3, pi044);
  not g_11365 (new_n4990_, new_n622_);
  or g_11366 (new_n685_, not_new_n1500_, not_new_n3023_);
  and g_11367 (new_n1524_, new_n3071_, and_new_n3073__new_n998_);
  not g_11368 (not_new_n7310_, new_n7310_);
  or g_11369 (new_n2710_, or_not_new_n1572__0_not_new_n1028__6, not_new_n581_);
  not g_11370 (not_new_n8156_, new_n8156_);
  or g_11371 (new_n3735_, not_new_n3734_, not_new_n3733_);
  not g_11372 (not_new_n5086_, new_n5086_);
  not g_11373 (not_new_n8036_, new_n8036_);
  or g_11374 (new_n1675_, key_gate_55, not_new_n596__3430);
  not g_11375 (not_new_n6474__2, new_n6474_);
  and g_11376 (new_n605_, new_n3369_, new_n2505_);
  not g_11377 (not_new_n4729_, new_n4729_);
  not g_11378 (not_pi099_0, pi099);
  not g_11379 (not_new_n1589_, new_n1589_);
  not g_11380 (not_new_n9008_, new_n9008_);
  or g_11381 (new_n4020_, pi033, pi034);
  or g_11382 (new_n6420_, not_new_n6242__0, or_or_not_new_n6328__not_new_n6373__3_not_new_n6329_);
  not g_11383 (not_new_n645__8235430, new_n645_);
  not g_11384 (not_new_n1613__1, new_n1613_);
  and g_11385 (new_n1330_, new_n2271_, new_n2272_);
  not g_11386 (not_new_n3347_, new_n3347_);
  or g_11387 (new_n7922_, not_new_n7860_, not_new_n7667_);
  not g_11388 (not_pi191_0, pi191);
  or g_11389 (new_n2421_, not_new_n597__490, not_new_n4803__0);
  not g_11390 (not_new_n1596__0, new_n1596_);
  or g_11391 (new_n2305_, not_new_n601__332329305696010, not_new_n617__0);
  or g_11392 (new_n3667_, not_po298_6, not_new_n635__9);
  not g_11393 (not_new_n1490_, new_n1490_);
  not g_11394 (new_n5464_, pi143);
  not g_11395 (not_new_n985__0, new_n985_);
  and g_11396 (and_new_n6473__new_n6833_, new_n6833_, new_n6473_);
  not g_11397 (new_n4241_, new_n671_);
  not g_11398 (not_pi271, pi271);
  not g_11399 (not_new_n1609_, new_n1609_);
  or g_11400 (new_n7266_, not_new_n7406__0, not_new_n7014__0);
  or g_11401 (new_n5382_, not_new_n5261_, not_new_n4998__1);
  or g_11402 (new_n7039_, not_new_n7437_, not_new_n7438_);
  not g_11403 (not_new_n1339_, new_n1339_);
  not g_11404 (not_new_n1585__8235430, new_n1585_);
  not g_11405 (not_new_n5707_, new_n5707_);
  or g_11406 (new_n8478_, not_new_n8322__0, not_new_n8246_);
  not g_11407 (not_new_n9151_, new_n9151_);
  not g_11408 (not_new_n6988_, new_n6988_);
  not g_11409 (not_new_n6974__5, new_n6974_);
  not g_11410 (not_new_n1601__9, new_n1601_);
  and g_11411 (new_n1552_, new_n3616_, new_n3617_);
  not g_11412 (not_new_n8099_, new_n8099_);
  not g_11413 (not_new_n9265_, new_n9265_);
  or g_11414 (new_n5631_, not_new_n5435__1, not_pi132_3);
  or g_11415 (new_n4125_, not_new_n4201_, not_new_n4202_);
  and g_11416 (new_n9466_, new_n9511_, new_n9582_);
  not g_11417 (not_new_n5128__0, new_n5128_);
  not g_11418 (not_new_n643__57648010, new_n643_);
  not g_11419 (not_new_n7622__0, new_n7622_);
  not g_11420 (not_new_n763_, new_n763_);
  or g_11421 (new_n5232_, new_n637_, new_n1065_);
  not g_11422 (not_new_n6470_, new_n6470_);
  or g_11423 (new_n9684_, not_new_n9549_, not_new_n9365__1);
  not g_11424 (not_new_n10056_, new_n10056_);
  or g_11425 (new_n8257_, not_new_n8427_, not_new_n8437_);
  and g_11426 (new_n1248_, and_and_new_n1877__new_n1880__new_n1878_, new_n1879_);
  or g_11427 (or_or_not_new_n2982__not_new_n2985__not_new_n2984_, or_not_new_n2982__not_new_n2985_, not_new_n2984_);
  not g_11428 (not_new_n6205_, new_n6205_);
  or g_11429 (new_n8741_, not_new_n1149__0, not_new_n8601_);
  not g_11430 (not_new_n5765__0, new_n5765_);
  not g_11431 (new_n4970_, new_n643_);
  not g_11432 (not_new_n7762_, new_n7762_);
  not g_11433 (not_new_n8062_, new_n8062_);
  not g_11434 (not_new_n9971__0, new_n9971_);
  and g_11435 (new_n6352_, new_n6373_, new_n6436_);
  not g_11436 (not_new_n1538__2326305139872070, new_n1538_);
  not g_11437 (not_new_n6974__490, new_n6974_);
  not g_11438 (not_new_n1603__57648010, new_n1603_);
  not g_11439 (not_new_n9458_, new_n9458_);
  not g_11440 (not_new_n599__2326305139872070, new_n599_);
  not g_11441 (not_new_n2991_, new_n2991_);
  not g_11442 (not_pi235, pi235);
  not g_11443 (not_new_n6623_, new_n6623_);
  or g_11444 (new_n1005_, not_new_n3332_, not_new_n3331_);
  and g_11445 (new_n4495_, new_n4667_, new_n4668_);
  not g_11446 (not_new_n1518_, new_n1518_);
  not g_11447 (not_new_n5062_, new_n5062_);
  not g_11448 (not_new_n4318_, new_n4318_);
  not g_11449 (not_new_n2071_, new_n2071_);
  not g_11450 (not_new_n6443__6782230728490, new_n6443_);
  not g_11451 (not_new_n1613__16284135979104490, new_n1613_);
  and g_11452 (new_n8943_, new_n8979_, new_n8811_);
  not g_11453 (not_new_n8855__0, new_n8855_);
  or g_11454 (or_not_new_n2685__not_new_n2684_, not_new_n2684_, not_new_n2685_);
  not g_11455 (not_new_n4797__0, new_n4797_);
  not g_11456 (not_new_n1027__5585458640832840070, new_n1027_);
  and g_11457 (new_n8950_, and_new_n8884__new_n9290_, new_n9289_);
  not g_11458 (not_new_n609__8, new_n609_);
  not g_11459 (new_n5752_, new_n642_);
  or g_11460 (new_n2965_, not_new_n4133__2, not_new_n3310__1176490);
  and g_11461 (po107, pi086, key_gate_101);
  not g_11462 (not_new_n6443__490, new_n6443_);
  or g_11463 (new_n7312_, not_new_n7086_, not_new_n7260__0);
  not g_11464 (not_new_n1611__1, new_n1611_);
  or g_11465 (new_n2451_, not_new_n597__57648010, not_new_n4788__0);
  or g_11466 (new_n2431_, not_new_n4798__0, not_new_n597__24010);
  not g_11467 (not_new_n1616__10, new_n1616_);
  or g_11468 (new_n9292_, not_new_n8882_, not_new_n1065__16284135979104490);
  or g_11469 (new_n2717_, not_new_n602_, not_new_n637__2);
  not g_11470 (not_new_n8675_, new_n8675_);
  or g_11471 (new_n4821_, not_new_n4730_, not_new_n1043__7);
  or g_11472 (new_n3551_, not_new_n1612__70, not_new_n2014__0);
  and g_11473 (and_new_n1258__new_n1932_, new_n1932_, new_n1258_);
  or g_11474 (new_n961_, not_new_n2115_, or_or_not_new_n1299__not_new_n1297__not_new_n2116_);
  not g_11475 (not_new_n9324_, new_n9324_);
  not g_11476 (not_new_n3671_, new_n3671_);
  not g_11477 (not_new_n2724_, new_n2724_);
  not g_11478 (not_new_n6640__1, new_n6640_);
  not g_11479 (not_new_n4799__0, new_n4799_);
  or g_11480 (or_or_not_new_n2727__not_new_n2730__not_new_n2729_, not_new_n2729_, or_not_new_n2727__not_new_n2730_);
  not g_11481 (not_new_n1055__1, new_n1055_);
  not g_11482 (not_new_n1593_, new_n1593_);
  not g_11483 (not_new_n9040_, new_n9040_);
  not g_11484 (not_new_n9903_, new_n9903_);
  not g_11485 (not_new_n5808__0, new_n5808_);
  not g_11486 (not_new_n6754_, new_n6754_);
  not g_11487 (not_new_n775__47475615099430, new_n775_);
  or g_11488 (new_n768_, not_new_n3193_, not_new_n3192_);
  not g_11489 (new_n9384_, new_n625_);
  not g_11490 (not_new_n3315__6782230728490, new_n3315_);
  not g_11491 (not_new_n3490_, new_n3490_);
  not g_11492 (new_n5568_, new_n5465_);
  not g_11493 (not_new_n1410_, new_n1410_);
  not g_11494 (not_new_n2110_, new_n2110_);
  not g_11495 (not_new_n1957__0, new_n1957_);
  not g_11496 (not_new_n1059__168070, new_n1059_);
  or g_11497 (new_n7173_, not_new_n6983_, not_new_n6984__0);
  not g_11498 (not_new_n8554_, new_n8554_);
  not g_11499 (not_pi145_2, pi145);
  not g_11500 (not_new_n1037__1176490, new_n1037_);
  not g_11501 (not_new_n7240__0, new_n7240_);
  not g_11502 (not_pi050_1, pi050);
  or g_11503 (po196, or_not_new_n1553__not_new_n1376_, not_new_n1375_);
  or g_11504 (new_n4664_, not_new_n4662_, not_new_n4663_);
  not g_11505 (not_new_n633__6782230728490, new_n633_);
  not g_11506 (not_new_n588__403536070, new_n588_);
  not g_11507 (not_new_n1386_, new_n1386_);
  not g_11508 (not_new_n3184__3, new_n3184_);
  not g_11509 (not_new_n10052_, new_n10052_);
  not g_11510 (not_new_n3920_, new_n3920_);
  or g_11511 (po277, or_or_or_not_new_n2820__not_new_n2823__not_new_n2822__not_new_n2824_, not_new_n2821_);
  not g_11512 (not_pi155_0, pi155);
  not g_11513 (not_new_n4439_, new_n4439_);
  not g_11514 (not_new_n1194_, new_n1194_);
  or g_11515 (new_n3349_, not_new_n1534__1176490, not_pi048_0);
  not g_11516 (not_new_n1611__138412872010, new_n1611_);
  not g_11517 (not_new_n645__332329305696010, new_n645_);
  or g_11518 (new_n7143_, not_new_n7243_, not_new_n7242_);
  or g_11519 (new_n5012_, not_new_n5354_, not_new_n5355_);
  not g_11520 (not_new_n1616__7, new_n1616_);
  not g_11521 (not_new_n8138_, new_n8138_);
  not g_11522 (not_new_n595__19773267430, new_n595_);
  not g_11523 (not_pi048, pi048);
  not g_11524 (not_new_n1605__6, new_n1605_);
  or g_11525 (new_n7006_, not_new_n7037_, not_new_n726_);
  not g_11526 (not_new_n1846_, new_n1846_);
  or g_11527 (new_n9113_, not_new_n8984_, not_new_n9109_);
  not g_11528 (not_new_n1604__3430, new_n1604_);
  not g_11529 (not_new_n9092_, new_n9092_);
  or g_11530 (new_n3855_, not_new_n6443__3430, not_new_n629__70);
  not g_11531 (not_new_n5859_, new_n5859_);
  not g_11532 (not_new_n8158_, new_n8158_);
  or g_11533 (new_n9753_, not_new_n619__138412872010, not_new_n9487__0);
  not g_11534 (not_new_n581__2326305139872070, new_n581_);
  not g_11535 (not_new_n5767__0, new_n5767_);
  and g_11536 (new_n7733_, new_n7768_, new_n8071_);
  not g_11537 (new_n1786_, new_n632_);
  not g_11538 (not_new_n7178_, new_n7178_);
  or g_11539 (new_n4686_, not_new_n4499_, not_new_n4500__0);
  not g_11540 (not_new_n4727__0, new_n4727_);
  not g_11541 (not_new_n7926_, new_n7926_);
  not g_11542 (not_new_n4778_, new_n4778_);
  not g_11543 (not_pi030_0, pi030);
  or g_11544 (new_n5920_, not_new_n5755_, not_new_n1043__70);
  not g_11545 (not_new_n9908_, new_n9908_);
  not g_11546 (not_new_n7465_, new_n7465_);
  not g_11547 (not_new_n5294_, new_n5294_);
  and g_11548 (new_n8659_, new_n8615_, new_n1057_);
  or g_11549 (new_n2771_, not_pi250_4, not_po296_1070069044235980333563563003849377848070);
  not g_11550 (not_new_n9897_, new_n9897_);
  not g_11551 (not_new_n1611__332329305696010, new_n1611_);
  not g_11552 (not_new_n6296_, new_n6296_);
  not g_11553 (not_new_n1705_, key_gate_18);
  not g_11554 (new_n6489_, new_n624_);
  not g_11555 (not_new_n7617__0, new_n7617_);
  not g_11556 (new_n6279_, new_n622_);
  not g_11557 (not_new_n1023__4, new_n1023_);
  not g_11558 (not_new_n1576__16284135979104490, new_n1576_);
  not g_11559 (new_n5755_, new_n631_);
  not g_11560 (not_new_n4532_, new_n4532_);
  not g_11561 (not_new_n2509__490, new_n2509_);
  not g_11562 (not_new_n6973_, new_n6973_);
  or g_11563 (new_n9593_, not_new_n1063__968890104070, not_new_n638__93874803376477543056490);
  not g_11564 (not_new_n1069__490, new_n1069_);
  or g_11565 (new_n8319_, not_new_n8206_, not_new_n8318_);
  or g_11566 (new_n3537_, not_new_n1612__4, not_new_n1881__0);
  not g_11567 (not_new_n1980_, new_n1980_);
  not g_11568 (not_new_n636__57648010, new_n636_);
  not g_11569 (not_new_n4419__0, new_n4419_);
  not g_11570 (not_new_n625__168070, new_n625_);
  or g_11571 (new_n4498_, not_new_n4563_, not_new_n4564_);
  or g_11572 (or_not_new_n4833__not_new_n4782_, not_new_n4833_, not_new_n4782_);
  not g_11573 (not_new_n5386_, new_n5386_);
  not g_11574 (not_pi180_1, pi180);
  not g_11575 (not_pi009, pi009);
  not g_11576 (not_new_n10164_, new_n10164_);
  or g_11577 (new_n6786_, not_new_n6711_, not_new_n6709__0);
  not g_11578 (not_new_n6819_, new_n6819_);
  not g_11579 (not_new_n5435_, new_n5435_);
  or g_11580 (new_n5762_, not_new_n5955_, not_new_n5757_);
  or g_11581 (new_n2337_, not_new_n1588__113988951853731430, not_new_n1607_);
  or g_11582 (po200, or_or_not_new_n1557__not_new_n2444__not_new_n1383_, not_new_n1384_);
  or g_11583 (new_n5122_, not_new_n5092_, not_new_n5096_);
  or g_11584 (new_n4383_, not_new_n656_, not_new_n4273_);
  and g_11585 (new_n5859_, new_n5809_, new_n5918_);
  and g_11586 (new_n1336_, and_and_new_n2295__new_n2298__new_n2296_, new_n2297_);
  or g_11587 (new_n8316_, not_new_n8104__0, not_new_n8308_);
  not g_11588 (not_new_n643__273687473400809163430, new_n643_);
  not g_11589 (not_new_n7096_, new_n7096_);
  not g_11590 (not_new_n2094_, new_n2094_);
  and g_11591 (new_n8687_, new_n1166_, new_n8620_);
  or g_11592 (new_n2393_, not_new_n4114__0, not_new_n600__7);
  or g_11593 (or_not_new_n3164__not_new_n3163_, not_new_n3163_, not_new_n3164_);
  not g_11594 (not_new_n8110_, new_n8110_);
  not g_11595 (not_new_n2565_, new_n2565_);
  not g_11596 (not_new_n1611__168070, new_n1611_);
  not g_11597 (not_new_n5778_, new_n5778_);
  not g_11598 (not_new_n3748_, new_n3748_);
  buf g_11599 (po018, pi211);
  or g_11600 (new_n10007_, not_new_n10081_, not_new_n10069_);
  not g_11601 (not_new_n1191_, new_n1191_);
  not g_11602 (new_n8392_, new_n8177_);
  not g_11603 (not_new_n9117_, new_n9117_);
  not g_11604 (not_new_n589_, new_n589_);
  not g_11605 (not_new_n5706__0, new_n5706_);
  not g_11606 (new_n8288_, new_n8165_);
  not g_11607 (not_new_n3094_, new_n3094_);
  not g_11608 (not_new_n7072_, new_n7072_);
  or g_11609 (new_n8044_, not_new_n633__19773267430, not_new_n7641__0);
  not g_11610 (not_new_n9480_, new_n9480_);
  not g_11611 (not_new_n7013__0, new_n7013_);
  or g_11612 (new_n4563_, not_new_n4500_, not_new_n4562_);
  not g_11613 (new_n8599_, new_n1163_);
  not g_11614 (not_new_n3794_, new_n3794_);
  not g_11615 (new_n4230_, new_n676_);
  or g_11616 (po252, not_new_n3691_, not_new_n3690_);
  not g_11617 (not_new_n2895_, new_n2895_);
  not g_11618 (not_new_n4161__0, new_n4161_);
  or g_11619 (new_n3634_, not_new_n984__19773267430, not_pi183_0);
  not g_11620 (not_new_n604__9, new_n604_);
  and g_11621 (new_n1466_, new_n3765_, new_n3762_);
  not g_11622 (not_new_n603__168070, new_n603_);
  not g_11623 (not_new_n6996_, new_n6996_);
  or g_11624 (new_n3671_, not_new_n648__9, not_po298_8);
  not g_11625 (not_new_n9884_, new_n9884_);
  not g_11626 (not_new_n1010__2, new_n1010_);
  or g_11627 (po233, not_new_n1457_, not_new_n1456_);
  or g_11628 (new_n7831_, not_new_n644__138412872010, not_new_n7646_);
  not g_11629 (new_n5798_, new_n637_);
  or g_11630 (new_n10083_, not_new_n628__93874803376477543056490, not_new_n1039__39098210485829880490);
  or g_11631 (new_n2185_, not_new_n2180_, not_new_n1312_);
  not g_11632 (not_new_n958_, new_n958_);
  not g_11633 (not_new_n4344_, new_n4344_);
  not g_11634 (not_new_n1027__57648010, new_n1027_);
  not g_11635 (not_new_n1606__6, new_n1606_);
  or g_11636 (new_n2826_, not_new_n602__10, not_new_n631__3);
  not g_11637 (new_n10213_, new_n9894_);
  not g_11638 (not_new_n7406__1, new_n7406_);
  or g_11639 (new_n5152_, new_n1057_, new_n636_);
  or g_11640 (new_n5730_, not_new_n6038_, not_new_n6035_);
  or g_11641 (new_n3774_, not_new_n3773_, not_new_n3772_);
  not g_11642 (not_new_n2892_, new_n2892_);
  and g_11643 (new_n4918_, new_n5139_, new_n5142_);
  not g_11644 (not_new_n8268_, new_n8268_);
  not g_11645 (not_new_n7019__0, new_n7019_);
  not g_11646 (not_new_n9395_, new_n9395_);
  or g_11647 (new_n8761_, not_new_n8681_, not_new_n8596_);
  or g_11648 (or_not_new_n1787__not_new_n1788_, not_new_n1788_, not_new_n1787_);
  not g_11649 (not_new_n4076_, new_n4076_);
  or g_11650 (new_n3552_, not_pi142_0, not_new_n1538__490);
  not g_11651 (not_new_n945_, new_n945_);
  or g_11652 (new_n2416_, not_new_n4806__0, not_new_n597__70);
  not g_11653 (new_n4943_, new_n1051_);
  not g_11654 (not_new_n6247_, new_n6247_);
  or g_11655 (new_n6056_, not_new_n6002__0, not_new_n5812__0);
  not g_11656 (not_new_n6214_, new_n6214_);
  or g_11657 (new_n7397_, not_new_n7351__0, not_new_n742__1);
  and g_11658 (new_n4470_, new_n4648_, and_new_n4580__new_n4649_);
  or g_11659 (new_n3203_, not_new_n589__7, not_new_n617__7);
  not g_11660 (not_new_n1534__332329305696010, key_gate_5);
  not g_11661 (not_new_n6522__0, new_n6522_);
  not g_11662 (not_new_n6915_, new_n6915_);
  or g_11663 (new_n3370_, not_pi055_0, not_new_n1534__47475615099430);
  or g_11664 (new_n9267_, not_new_n9265_, not_new_n9266_);
  not g_11665 (not_new_n10068_, new_n10068_);
  and g_11666 (new_n9335_, new_n9330_, new_n9584_);
  or g_11667 (new_n1870_, not_new_n5828_, not_new_n1585__4);
  and g_11668 (new_n1483_, new_n1484_, new_n2901_);
  not g_11669 (not_new_n1831_, new_n1831_);
  not g_11670 (not_new_n5084_, new_n5084_);
  or g_11671 (new_n7141_, not_new_n7246_, not_new_n7247_);
  not g_11672 (not_new_n594__168070, new_n594_);
  not g_11673 (not_new_n1071__168070, new_n1071_);
  not g_11674 (not_new_n1057__57648010, new_n1057_);
  not g_11675 (not_new_n1611__10, new_n1611_);
  or g_11676 (new_n5389_, not_new_n633__168070, not_new_n4985__0);
  or g_11677 (new_n3465_, not_pi109_0, not_new_n1537__70);
  not g_11678 (not_new_n1061__332329305696010, new_n1061_);
  or g_11679 (or_not_new_n1572__0_not_new_n1028__6, not_new_n1028__6, not_new_n1572__0);
  or g_11680 (new_n5496_, not_new_n5546_, not_new_n5545_);
  not g_11681 (not_new_n8906_, new_n8906_);
  or g_11682 (new_n9555_, not_new_n1039__16284135979104490, not_new_n628__39098210485829880490);
  not g_11683 (not_new_n9327__1, new_n9327_);
  or g_11684 (new_n6061_, not_new_n5728_, not_new_n5900__1);
  not g_11685 (new_n8451_, new_n8248_);
  not g_11686 (new_n7415_, new_n7030_);
  or g_11687 (or_not_new_n8172__0_not_new_n1596__138412872010, not_new_n1596__138412872010, not_new_n8172__0);
  not g_11688 (not_new_n9037_, new_n9037_);
  or g_11689 (new_n9270_, not_new_n639__332329305696010, not_new_n8879_);
  not g_11690 (not_new_n9259_, new_n9259_);
  not g_11691 (not_new_n9063_, new_n9063_);
  not g_11692 (not_new_n4901_, new_n4901_);
  not g_11693 (not_new_n605_, new_n605_);
  not g_11694 (not_new_n6979_, new_n6979_);
  not g_11695 (not_new_n2863_, new_n2863_);
  or g_11696 (new_n2153_, not_new_n601__57648010, not_new_n645__0);
  not g_11697 (not_new_n7530_, new_n7530_);
  not g_11698 (not_new_n6729_, new_n6729_);
  not g_11699 (not_new_n1591__968890104070, new_n1591_);
  not g_11700 (not_new_n2071__0, new_n2071_);
  not g_11701 (not_new_n3993_, new_n3993_);
  not g_11702 (not_new_n1603__6782230728490, new_n1603_);
  not g_11703 (not_new_n1006__2, new_n1006_);
  or g_11704 (new_n7178_, not_new_n7342_, not_new_n6981_);
  not g_11705 (not_new_n3379_, new_n3379_);
  not g_11706 (not_new_n1359_, new_n1359_);
  not g_11707 (not_new_n1603__8235430, new_n1603_);
  or g_11708 (new_n5835_, not_new_n6205_, not_new_n6204_);
  not g_11709 (not_new_n1149_, new_n1149_);
  not g_11710 (not_new_n1536__168070, new_n1536_);
  not g_11711 (not_new_n4986__0, new_n4986_);
  or g_11712 (new_n4693_, not_new_n4501_, not_new_n4502__0);
  or g_11713 (new_n6831_, not_new_n6682_, not_new_n6612_);
  not g_11714 (not_new_n1600__1176490, new_n1600_);
  or g_11715 (new_n9519_, new_n628_, new_n1039_);
  not g_11716 (not_new_n1606_, new_n1606_);
  not g_11717 (not_new_n1045__3430, new_n1045_);
  or g_11718 (new_n9815_, not_new_n9501__0, not_new_n9690_);
  not g_11719 (not_new_n7209_, new_n7209_);
  not g_11720 (not_new_n9501_, new_n9501_);
  and g_11721 (new_n1205_, new_n1704_, new_n1706_);
  not g_11722 (not_new_n5064_, new_n5064_);
  or g_11723 (new_n2605_, not_new_n605__9, not_new_n5476_);
  not g_11724 (not_new_n3521_, new_n3521_);
  or g_11725 (new_n2204_, not_new_n1316_, not_new_n2199_);
  or g_11726 (new_n7306_, not_new_n7006__0, not_new_n7240__0);
  or g_11727 (new_n5147_, not_new_n5145_, not_new_n5034_);
  and g_11728 (new_n8093_, new_n8493_, new_n8492_);
  not g_11729 (not_new_n601__968890104070, new_n601_);
  or g_11730 (new_n10211_, not_new_n9854__1, or_not_new_n9855__0_not_new_n10046__0);
  or g_11731 (po232, not_new_n1454_, not_new_n1455_);
  not g_11732 (not_pi130_2, pi130);
  not g_11733 (not_new_n2503_, new_n2503_);
  not g_11734 (not_pi066, pi066);
  not g_11735 (not_new_n724__1, new_n724_);
  not g_11736 (not_new_n3540_, new_n3540_);
  not g_11737 (not_new_n5091__0, new_n5091_);
  not g_11738 (not_new_n928__8, new_n928_);
  not g_11739 (not_new_n7025__1, new_n7025_);
  not g_11740 (not_new_n4278_, new_n4278_);
  not g_11741 (not_new_n1002__5, new_n1002_);
  or g_11742 (new_n8405_, not_new_n8178_, not_new_n8281_);
  or g_11743 (new_n9433_, not_new_n9736_, not_new_n9735_);
  not g_11744 (not_new_n5882_, new_n5882_);
  not g_11745 (not_new_n6629_, new_n6629_);
  not g_11746 (not_new_n1045__490, new_n1045_);
  or g_11747 (new_n2423_, not_new_n4133__0, not_new_n600__3430);
  and g_11748 (new_n6227_, new_n6315_, new_n6226_);
  not g_11749 (not_new_n3896_, new_n3896_);
  not g_11750 (not_new_n735__1, new_n735_);
  not g_11751 (not_new_n1611__2, new_n1611_);
  not g_11752 (not_new_n6812_, new_n6812_);
  or g_11753 (po228, not_new_n1445_, not_new_n1444_);
  not g_11754 (not_new_n1601__19773267430, new_n1601_);
  and g_11755 (and_and_and_new_n2325__new_n2332__new_n2333__new_n2329_, and_and_new_n2325__new_n2332__new_n2333_, new_n2329_);
  not g_11756 (not_new_n767_, new_n767_);
  or g_11757 (new_n3397_, not_new_n3375__5, not_new_n1023__3);
  not g_11758 (not_new_n7036__0, new_n7036_);
  not g_11759 (new_n4428_, new_n1004_);
  not g_11760 (not_new_n1580__7, new_n1580_);
  not g_11761 (new_n8848_, new_n1597_);
  not g_11762 (not_new_n6920_, new_n6920_);
  or g_11763 (po172, not_new_n3571_, not_new_n3570_);
  not g_11764 (not_new_n1583__3, new_n1583_);
  not g_11765 (not_new_n3770_, new_n3770_);
  not g_11766 (not_new_n5617__1, new_n5617_);
  or g_11767 (new_n8096_, not_new_n8529_, or_or_or_not_new_n8528__not_new_n8429__not_new_n8457__not_new_n8458_);
  and g_11768 (and_new_n3082__new_n998_, new_n998_, new_n3082_);
  or g_11769 (or_not_new_n7313__not_new_n7314_, not_new_n7314_, not_new_n7313_);
  or g_11770 (or_or_or_not_new_n2883__not_new_n2886__not_new_n2885__not_new_n2887_, not_new_n2887_, or_or_not_new_n2883__not_new_n2886__not_new_n2885_);
  or g_11771 (new_n4717_, not_new_n4413_, not_pi161_3);
  not g_11772 (not_new_n1041__10, new_n1041_);
  or g_11773 (or_not_new_n7908__not_new_n7743_, not_new_n7908_, not_new_n7743_);
  or g_11774 (new_n6987_, not_new_n775_, not_new_n745_);
  not g_11775 (not_new_n7419_, new_n7419_);
  xnor g_11776 (key_gate_58, new_n1684_, key_58);
  not g_11777 (not_new_n1581__138412872010, new_n1581_);
  or g_11778 (new_n3093_, not_new_n581__1915812313805664144010, not_new_n634__6);
  not g_11779 (not_new_n3486_, new_n3486_);
  or g_11780 (new_n4590_, not_pi170_3, not_new_n4431__0);
  not g_11781 (not_new_n7448_, new_n7448_);
  not g_11782 (not_new_n3220_, new_n3220_);
  not g_11783 (not_new_n4160_, new_n4160_);
  not g_11784 (not_new_n7187_, new_n7187_);
  not g_11785 (not_new_n5488_, new_n5488_);
  not g_11786 (not_new_n8148_, new_n8148_);
  not g_11787 (not_new_n4592_, new_n4592_);
  not g_11788 (new_n5756_, new_n624_);
  not g_11789 (new_n7121_, new_n760_);
  not g_11790 (not_new_n632__968890104070, new_n632_);
  and g_11791 (new_n1262_, new_n1948_, new_n1949_);
  not g_11792 (not_new_n9944__0, new_n9944_);
  and g_11793 (and_and_new_n2219__new_n2222__new_n2220_, new_n2220_, and_new_n2219__new_n2222_);
  not g_11794 (not_new_n1039__8, new_n1039_);
  not g_11795 (new_n8959_, new_n1607_);
  or g_11796 (new_n4203_, not_pi264_1, not_new_n4098_);
  not g_11797 (not_new_n3682_, new_n3682_);
  or g_11798 (new_n5621_, not_new_n5619_, not_new_n1006__6);
  and g_11799 (new_n1211_, new_n1722_, new_n1724_);
  or g_11800 (new_n974_, not_new_n2248_, or_or_not_new_n1327__not_new_n1325__not_new_n2249_);
  and g_11801 (new_n4315_, new_n4395_, new_n4394_);
  and g_11802 (new_n1292_, and_and_new_n2086__new_n2089__new_n2087_, new_n2088_);
  not g_11803 (not_new_n597__3, new_n597_);
  not g_11804 (not_new_n8716__0, new_n8716_);
  not g_11805 (not_new_n8083_, new_n8083_);
  not g_11806 (not_new_n8117__0, new_n8117_);
  or g_11807 (new_n6002_, not_new_n5772_, not_new_n1603__70);
  not g_11808 (not_new_n6209_, new_n6209_);
  not g_11809 (not_new_n622__1176490, new_n622_);
  not g_11810 (not_new_n3170_, new_n3170_);
  or g_11811 (new_n2656_, or_not_new_n2655__not_new_n2654_, not_new_n2653_);
  not g_11812 (not_new_n6353_, new_n6353_);
  not g_11813 (not_new_n1537__6782230728490, new_n1537_);
  not g_11814 (not_new_n627__403536070, new_n627_);
  not g_11815 (not_new_n7802_, new_n7802_);
  not g_11816 (not_new_n4307_, new_n4307_);
  buf g_11817 (po023, pi241);
  or g_11818 (new_n7860_, not_new_n7623_, not_new_n1599__24010);
  not g_11819 (not_new_n3366__0, new_n3366_);
  xor g_11820 (key_gate_120, new_n1723_, key_120);
  or g_11821 (new_n5387_, not_new_n5262_, not_new_n5073__0);
  not g_11822 (not_new_n581__5585458640832840070, new_n581_);
  not g_11823 (not_new_n1538__2, new_n1538_);
  or g_11824 (new_n1032_, not_new_n3402_, not_new_n3403_);
  not g_11825 (not_new_n4003__0, new_n4003_);
  or g_11826 (new_n5999_, not_new_n625__1176490, not_new_n5774_);
  or g_11827 (new_n3259_, not_new_n589__13410686196639649008070, not_new_n1596__5);
  not g_11828 (not_new_n1063__2, new_n1063_);
  and g_11829 (new_n7075_, new_n6961_, new_n7193_);
  not g_11830 (not_new_n7873_, new_n7873_);
  not g_11831 (not_new_n2743_, new_n2743_);
  not g_11832 (not_new_n617__113988951853731430, new_n617_);
  or g_11833 (or_not_new_n2845__not_new_n2844_, not_new_n2845_, not_new_n2844_);
  not g_11834 (new_n7936_, new_n7761_);
  or g_11835 (new_n7897_, not_new_n7651__0, not_new_n626__2326305139872070);
  not g_11836 (not_new_n618__5, new_n618_);
  or g_11837 (new_n5664_, not_new_n5510_, not_new_n5511__0);
  not g_11838 (not_new_n607__9, new_n607_);
  or g_11839 (new_n8183_, not_new_n8542_, not_new_n8541_);
  not g_11840 (new_n4510_, new_n4415_);
  not g_11841 (not_new_n8987_, new_n8987_);
  or g_11842 (new_n5861_, not_new_n6152_, not_new_n6153_);
  or g_11843 (new_n4136_, not_new_n4223_, not_new_n4224_);
  not g_11844 (not_new_n6180_, new_n6180_);
  not g_11845 (not_new_n9416__0, new_n9416_);
  or g_11846 (new_n2311_, not_new_n1591__2326305139872070, not_new_n8909_);
  not g_11847 (not_new_n4937_, new_n4937_);
  not g_11848 (new_n9565_, new_n9485_);
  not g_11849 (not_new_n1598__70, new_n1598_);
  not g_11850 (not_new_n10280_, new_n10280_);
  not g_11851 (not_new_n1536__0, new_n1536_);
  not g_11852 (not_new_n7085_, new_n7085_);
  and g_11853 (new_n8681_, and_and_new_n8723__new_n1174__new_n8719_, new_n8619_);
  not g_11854 (not_new_n1016__6, new_n1016_);
  not g_11855 (new_n8862_, new_n1057_);
  or g_11856 (or_not_new_n2557__not_new_n2561_, not_new_n2561_, not_new_n2557_);
  not g_11857 (not_new_n9713_, new_n9713_);
  not g_11858 (not_new_n588__2326305139872070, new_n588_);
  and g_11859 (new_n1440_, and_new_n2627__new_n2628_, new_n2629_);
  or g_11860 (new_n10095_, new_n644_, new_n1059_);
  and g_11861 (new_n1320_, and_and_new_n2219__new_n2222__new_n2220_, new_n2221_);
  not g_11862 (not_pi189, pi189);
  not g_11863 (not_new_n1027__2824752490, new_n1027_);
  not g_11864 (not_new_n4618_, new_n4618_);
  or g_11865 (or_not_new_n1552__not_new_n2419_, not_new_n1552_, not_new_n2419_);
  not g_11866 (not_new_n640__10, new_n640_);
  not g_11867 (not_new_n3344_, new_n3344_);
  not g_11868 (not_new_n1045__8235430, new_n1045_);
  not g_11869 (not_new_n8609_, new_n8609_);
  not g_11870 (not_new_n1069__3430, new_n1069_);
  or g_11871 (new_n3167_, not_new_n3315__2326305139872070, not_new_n627__5);
  or g_11872 (new_n3245_, not_new_n1051__5, not_new_n589__16284135979104490);
  not g_11873 (not_new_n1001__0, new_n1001_);
  not g_11874 (new_n5806_, new_n1598_);
  or g_11875 (new_n9153_, not_new_n8955_, not_new_n9151_);
  or g_11876 (new_n7832_, not_new_n1065__57648010, not_new_n7655_);
  not g_11877 (not_new_n588__168070, new_n588_);
  not g_11878 (not_new_n7584_, new_n7584_);
  not g_11879 (not_new_n7065_, new_n7065_);
  not g_11880 (not_pi027, pi027);
  not g_11881 (not_new_n6497_, new_n6497_);
  not g_11882 (new_n1952_, new_n952_);
  not g_11883 (not_new_n602__6782230728490, new_n602_);
  not g_11884 (not_new_n2281_, new_n2281_);
  or g_11885 (new_n2243_, not_pi187, not_new_n586__47475615099430);
  not g_11886 (not_new_n636__168070, new_n636_);
  not g_11887 (not_po298_7, po298);
  not g_11888 (not_new_n5153_, new_n5153_);
  not g_11889 (not_new_n4224_, new_n4224_);
  not g_11890 (not_new_n6591_, new_n6591_);
  not g_11891 (not_new_n4472_, new_n4472_);
  or g_11892 (new_n4538_, pi169, new_n1003_);
  and g_11893 (new_n1287_, and_new_n1286__new_n2065_, new_n2064_);
  not g_11894 (not_new_n4246_, new_n4246_);
  not g_11895 (not_pi005, pi005);
  not g_11896 (not_new_n639__403536070, new_n639_);
  not g_11897 (not_pi030, pi030);
  not g_11898 (not_new_n600__19773267430, new_n600_);
  or g_11899 (new_n2806_, not_new_n595__7, not_new_n7060_);
  or g_11900 (new_n6469_, not_new_n6697_, not_new_n6694_);
  or g_11901 (new_n4631_, not_new_n4419__0, not_new_n1008__4);
  not g_11902 (not_new_n1012__6, new_n1012_);
  not g_11903 (not_new_n7685_, new_n7685_);
  not g_11904 (not_new_n6924_, new_n6924_);
  or g_11905 (new_n8043_, not_new_n7640__0, not_new_n1067__1176490);
  not g_11906 (new_n4986_, new_n1601_);
  not g_11907 (not_new_n1016__5, new_n1016_);
  or g_11908 (new_n3277_, not_new_n589__541169560379521116689596608490, not_new_n1037__5);
  not g_11909 (not_new_n7793_, new_n7793_);
  not g_11910 (not_new_n1043__6782230728490, new_n1043_);
  or g_11911 (new_n8263_, not_new_n8431_, not_new_n8144_);
  not g_11912 (not_new_n9439_, new_n9439_);
  not g_11913 (not_new_n1557_, new_n1557_);
  not g_11914 (not_new_n9710_, new_n9710_);
  not g_11915 (new_n4529_, new_n4479_);
  or g_11916 (new_n2435_, not_new_n1065__0, not_new_n598__168070);
  or g_11917 (new_n3758_, not_new_n971_, not_new_n2209_);
  not g_11918 (not_new_n4952_, new_n4952_);
  not g_11919 (not_new_n594__3430, new_n594_);
  not g_11920 (not_new_n7752__0, new_n7752_);
  not g_11921 (not_pi248_1, pi248);
  or g_11922 (new_n1884_, not_new_n588__6, not_pi104);
  not g_11923 (not_new_n7690_, new_n7690_);
  or g_11924 (or_not_new_n1251__not_new_n1249_, not_new_n1249_, not_new_n1251_);
  not g_11925 (not_pi064_2, pi064);
  or g_11926 (new_n9940_, not_new_n629__16284135979104490, not_new_n1600__47475615099430);
  not g_11927 (not_new_n5538_, new_n5538_);
  or g_11928 (new_n3403_, not_new_n1728__797922662976120010, not_pi065_0);
  not g_11929 (not_new_n5521_, new_n5521_);
  or g_11930 (new_n2550_, not_new_n608__3, not_new_n1014__0);
  or g_11931 (new_n9009_, not_new_n8845_, not_new_n8800_);
  not g_11932 (not_new_n1039__3, new_n1039_);
  not g_11933 (not_new_n7415__2, new_n7415_);
  not g_11934 (not_new_n9484__0, new_n9484_);
  or g_11935 (new_n8537_, not_new_n8261_, not_new_n8434_);
  not g_11936 (not_new_n3384_, new_n3384_);
  not g_11937 (not_new_n7277__0, new_n7277_);
  or g_11938 (new_n9036_, not_new_n8992__0, not_new_n8995__0);
  not g_11939 (not_new_n5321_, new_n5321_);
  not g_11940 (not_new_n8649_, new_n8649_);
  or g_11941 (new_n7455_, not_new_n775__2326305139872070, not_new_n7133_);
  or g_11942 (new_n3877_, not_new_n6443__6782230728490, not_new_n643__70);
  not g_11943 (not_new_n7348_, new_n7348_);
  not g_11944 (not_pi084, pi084);
  not g_11945 (not_new_n1061__2, new_n1061_);
  not g_11946 (not_new_n1583__968890104070, new_n1583_);
  or g_11947 (new_n3856_, not_new_n1576__3430, not_new_n629__490);
  not g_11948 (new_n8279_, new_n8112_);
  or g_11949 (new_n4595_, not_pi169_2, not_new_n4430_);
  and g_11950 (new_n4507_, new_n4710_, new_n4709_);
  or g_11951 (new_n10124_, not_new_n10123_, not_new_n10122_);
  not g_11952 (not_new_n2058_, new_n2058_);
  not g_11953 (not_new_n1663_, key_gate_61);
  not g_11954 (not_new_n8138__0, new_n8138_);
  not g_11955 (not_new_n1576__19773267430, new_n1576_);
  not g_11956 (not_new_n622__19773267430, new_n622_);
  or g_11957 (or_not_new_n1158__1_not_new_n8715__0, not_new_n8715__0, not_new_n1158__1);
  and g_11958 (new_n5904_, new_n6202_, new_n6203_);
  not g_11959 (not_new_n7557_, new_n7557_);
  not g_11960 (not_new_n1583__2824752490, new_n1583_);
  or g_11961 (new_n4978_, not_new_n1069__8, not_new_n646__3430);
  not g_11962 (not_new_n581__57648010, new_n581_);
  or g_11963 (new_n6696_, not_new_n6487__1, not_new_n1045__8235430);
  or g_11964 (new_n9430_, not_new_n9852_, not_new_n9853_);
  not g_11965 (not_new_n1071__968890104070, new_n1071_);
  or g_11966 (new_n9967_, not_new_n10326_, not_new_n10327_);
  not g_11967 (not_new_n7751_, new_n7751_);
  or g_11968 (new_n4339_, not_new_n4243_, not_new_n672_);
  not g_11969 (not_new_n1612__1176490, new_n1612_);
  not g_11970 (not_new_n10322_, new_n10322_);
  not g_11971 (not_new_n1031__4, new_n1031_);
  not g_11972 (not_new_n8439_, new_n8439_);
  not g_11973 (not_new_n1051__9, new_n1051_);
  or g_11974 (new_n6884_, not_new_n6499__0, not_new_n1599__3430);
  not g_11975 (not_new_n1612__490, new_n1612_);
  or g_11976 (new_n3692_, not_new_n989__57648010, not_pi232);
  not g_11977 (not_new_n606__490, new_n606_);
  not g_11978 (not_new_n1631__2824752490, key_gate_76);
  not g_11979 (not_new_n628__6782230728490, new_n628_);
  not g_11980 (new_n7123_, new_n757_);
  not g_11981 (new_n6540_, new_n1596_);
  and g_11982 (new_n6572_, new_n6453_, new_n6452_);
  not g_11983 (not_new_n3311__70, new_n3311_);
  not g_11984 (not_new_n1179__0, new_n1179_);
  not g_11985 (not_new_n8090_, new_n8090_);
  not g_11986 (not_new_n5314_, new_n5314_);
  or g_11987 (or_not_new_n6541__0_not_new_n1596__1176490, not_new_n6541__0, not_new_n1596__1176490);
  not g_11988 (new_n9884_, new_n628_);
  not g_11989 (new_n4985_, new_n1067_);
  not g_11990 (not_new_n3881_, new_n3881_);
  not g_11991 (not_new_n5606_, new_n5606_);
  or g_11992 (new_n7957_, not_new_n1047__1176490, not_new_n7596__0);
  not g_11993 (not_pi164_1, pi164);
  not g_11994 (not_new_n5753__1, new_n5753_);
  not g_11995 (not_new_n581__1577753820348458066150427430, new_n581_);
  or g_11996 (new_n6678_, not_new_n6474_, not_new_n1049__24010);
  not g_11997 (not_new_n5973_, new_n5973_);
  not g_11998 (not_new_n587__47475615099430, new_n587_);
  or g_11999 (new_n8494_, not_new_n8251__0, not_new_n1607__168070);
  not g_12000 (not_pi169_0, pi169);
  not g_12001 (not_new_n4751_, new_n4751_);
  or g_12002 (new_n2948_, not_new_n2945_, not_new_n1616__138412872010);
  not g_12003 (not_new_n6081_, new_n6081_);
  or g_12004 (or_not_new_n6352__not_new_n6242__5, not_new_n6352_, not_new_n6242__5);
  or g_12005 (new_n8894_, not_new_n9108_, not_new_n8854_);
  or g_12006 (new_n3011_, not_new_n1156_, not_new_n1027__10);
  not g_12007 (not_new_n6662_, new_n6662_);
  not g_12008 (not_new_n579_, new_n579_);
  or g_12009 (new_n10081_, not_new_n10042__0, not_new_n10045__0);
  or g_12010 (new_n5977_, not_new_n1059__490, not_new_n5788_);
  not g_12011 (not_new_n8061_, new_n8061_);
  not g_12012 (not_new_n639__4, new_n639_);
  or g_12013 (new_n5674_, not_new_n5467_, not_new_n5568_);
  not g_12014 (not_new_n633__8, new_n633_);
  and g_12015 (new_n1508_, new_n1509_, new_n3037_);
  not g_12016 (not_new_n1336_, new_n1336_);
  not g_12017 (not_new_n9701_, new_n9701_);
  or g_12018 (new_n2514_, not_pi193, not_new_n2509_);
  or g_12019 (new_n7339_, not_new_n7338_, not_new_n7337_);
  not g_12020 (not_new_n7442__0, new_n7442_);
  and g_12021 (new_n616_, and_and_and_new_n2325__new_n2332__new_n2333__new_n2329_, new_n2326_);
  not g_12022 (new_n8620_, new_n1603_);
  not g_12023 (not_new_n8190_, new_n8190_);
  not g_12024 (not_new_n6635__1, new_n6635_);
  and g_12025 (new_n8083_, and_new_n8304__new_n8299_, new_n8286_);
  or g_12026 (new_n5604_, not_new_n1004__7, not_new_n5445__0);
  not g_12027 (not_new_n1244_, new_n1244_);
  or g_12028 (new_n7410_, not_new_n7118_, not_new_n775__490);
  not g_12029 (new_n1614_, key_gate_101);
  and g_12030 (new_n8593_, new_n8732_, new_n8592_);
  not g_12031 (new_n9118_, new_n8898_);
  not g_12032 (not_new_n9965_, new_n9965_);
  not g_12033 (not_new_n6506_, new_n6506_);
  or g_12034 (new_n10094_, not_new_n10093_, not_new_n10092_);
  or g_12035 (new_n4329_, not_new_n677_, not_new_n4232_);
  not g_12036 (not_new_n6654_, new_n6654_);
  not g_12037 (not_new_n1631__403536070, key_gate_76);
  or g_12038 (new_n2917_, not_new_n4119__1, not_new_n994__138412872010);
  not g_12039 (not_new_n7704_, new_n7704_);
  not g_12040 (not_new_n947_, new_n947_);
  or g_12041 (new_n5645_, or_not_new_n5430__0_not_pi130_2, not_new_n5431__1);
  not g_12042 (not_new_n7076_, new_n7076_);
  or g_12043 (new_n3777_, not_new_n3775_, not_new_n3776_);
  or g_12044 (new_n9643_, not_new_n9474_, not_new_n9641_);
  not g_12045 (new_n3950_, pi055);
  not g_12046 (not_new_n5432_, new_n5432_);
  not g_12047 (not_new_n1166_, new_n1166_);
  not g_12048 (not_new_n7772__0, new_n7772_);
  not g_12049 (not_new_n775__9, new_n775_);
  not g_12050 (not_new_n4671_, new_n4671_);
  not g_12051 (not_new_n629__57648010, new_n629_);
  or g_12052 (new_n3440_, not_new_n1537__6, not_pi104_0);
  not g_12053 (new_n9703_, new_n9399_);
  not g_12054 (not_new_n1598__490, new_n1598_);
  not g_12055 (not_new_n644__39098210485829880490, new_n644_);
  or g_12056 (new_n9818_, not_new_n9411_, not_new_n1067__6782230728490);
  and g_12057 (and_new_n6433__new_n6432_, new_n6433_, new_n6432_);
  not g_12058 (not_new_n3549_, new_n3549_);
  not g_12059 (not_new_n3843_, new_n3843_);
  and g_12060 (new_n9990_, new_n10033_, new_n10098_);
  or g_12061 (new_n2414_, not_new_n9972__0, not_new_n599__70);
  or g_12062 (new_n1957_, not_new_n1952_, not_new_n1264_);
  not g_12063 (not_new_n1603__70, new_n1603_);
  not g_12064 (not_new_n6223_, new_n6223_);
  or g_12065 (new_n1168_, not_new_n3865_, not_new_n3866_);
  not g_12066 (not_new_n1885_, new_n1885_);
  not g_12067 (not_new_n4259_, new_n4259_);
  or g_12068 (new_n7685_, not_new_n7959_, not_new_n7960_);
  or g_12069 (new_n5321_, not_new_n4921_, not_new_n632__168070);
  not g_12070 (not_new_n7424_, new_n7424_);
  not g_12071 (not_new_n1041__968890104070, new_n1041_);
  or g_12072 (or_not_new_n8169__1_not_new_n8508_, not_new_n8169__1, not_new_n8508_);
  or g_12073 (new_n4644_, not_new_n4414_, not_new_n4510__0);
  not g_12074 (not_new_n7141__0, new_n7141_);
  not g_12075 (not_new_n5524_, new_n5524_);
  not g_12076 (not_new_n9781_, new_n9781_);
  or g_12077 (new_n9112_, not_new_n8945_, not_new_n9111_);
  not g_12078 (not_new_n1613__8235430, new_n1613_);
  and g_12079 (new_n1491_, and_new_n3004__new_n998_, new_n3002_);
  and g_12080 (new_n4289_, and_new_n4405__new_n4330_, new_n4329_);
  not g_12081 (not_new_n7014__0, new_n7014_);
  or g_12082 (new_n3607_, not_new_n1611__7, not_new_n951_);
  not g_12083 (not_new_n1583__6782230728490, new_n1583_);
  not g_12084 (not_new_n3898_, new_n3898_);
  xor g_12085 (key_gate_117, not_new_n3925_, key_117);
  or g_12086 (new_n2880_, not_new_n602__1176490, not_new_n644__2);
  not g_12087 (not_new_n6596_, new_n6596_);
  not g_12088 (not_new_n4134_, new_n4134_);
  not g_12089 (new_n4173_, new_n4108_);
  and g_12090 (and_new_n6373__new_n6386_, new_n6373_, new_n6386_);
  and g_12091 (new_n5032_, new_n5133_, new_n4898_);
  not g_12092 (new_n4792_, new_n1067_);
  not g_12093 (not_new_n3372__968890104070, new_n3372_);
  or g_12094 (new_n5386_, not_new_n5385_, not_new_n5384_);
  or g_12095 (new_n3840_, not_new_n620__4, not_new_n1576__5);
  not g_12096 (not_new_n1311_, new_n1311_);
  not g_12097 (not_po296_10, po296);
  not g_12098 (not_new_n1045__1176490, new_n1045_);
  not g_12099 (not_new_n4100_, new_n4100_);
  not g_12100 (not_new_n5740__0, new_n5740_);
  or g_12101 (new_n1939_, not_pi171, not_new_n586__9);
  or g_12102 (new_n3725_, not_new_n2322_, not_new_n982_);
  and g_12103 (new_n1188_, new_n1653_, new_n1655_);
  not g_12104 (not_new_n5069_, new_n5069_);
  not g_12105 (not_new_n634__2, new_n634_);
  not g_12106 (not_new_n2868_, new_n2868_);
  not g_12107 (new_n8111_, new_n632_);
  or g_12108 (new_n10241_, not_new_n648__273687473400809163430, not_new_n9895_);
  not g_12109 (not_new_n9873__0, new_n9873_);
  not g_12110 (not_new_n4573_, new_n4573_);
  and g_12111 (new_n1332_, new_n2278_, and_and_new_n2276__new_n2279__new_n2277_);
  not g_12112 (new_n3396_, new_n1031_);
  not g_12113 (not_new_n6153_, new_n6153_);
  not g_12114 (not_new_n8972_, new_n8972_);
  or g_12115 (new_n6438_, not_new_n6233__1, or_or_not_new_n6353__not_new_n6232__5_not_new_n1069__3430);
  not g_12116 (not_new_n1000_, new_n1000_);
  not g_12117 (not_new_n621__113988951853731430, new_n621_);
  not g_12118 (new_n5466_, new_n1014_);
  not g_12119 (new_n8856_, new_n625_);
  not g_12120 (not_new_n5763_, new_n5763_);
  not g_12121 (not_new_n9949_, new_n9949_);
  not g_12122 (not_new_n7816_, new_n7816_);
  not g_12123 (not_new_n10339_, new_n10339_);
  and g_12124 (new_n4312_, new_n4385_, new_n4386_);
  not g_12125 (not_new_n581__26517308458596534717790233816010, new_n581_);
  or g_12126 (new_n6114_, not_new_n5881_, not_new_n6076_);
  not g_12127 (not_new_n1537__8235430, new_n1537_);
  not g_12128 (not_new_n7770_, new_n7770_);
  and g_12129 (new_n9341_, new_n9674_, new_n9671_);
  not g_12130 (not_new_n6443__2326305139872070, new_n6443_);
  not g_12131 (not_new_n1976_, new_n1976_);
  not g_12132 (not_new_n7368_, new_n7368_);
  not g_12133 (new_n4736_, new_n1041_);
  not g_12134 (not_new_n1067__57648010, new_n1067_);
  not g_12135 (not_new_n3310__4, new_n3310_);
  or g_12136 (new_n5117_, not_new_n5028_, not_new_n5116_);
  not g_12137 (not_new_n8524_, new_n8524_);
  or g_12138 (new_n10102_, not_new_n9864_, not_new_n10029__0);
  not g_12139 (new_n8172_, new_n618_);
  not g_12140 (not_pi165, pi165);
  or g_12141 (new_n8526_, not_new_n630__968890104070, not_new_n8137__0);
  not g_12142 (not_new_n1597__5, new_n1597_);
  not g_12143 (not_new_n1027__490, new_n1027_);
  or g_12144 (new_n2168_, not_new_n587__19773267430, not_pi151);
  not g_12145 (not_new_n8964_, new_n8964_);
  not g_12146 (not_new_n10023_, new_n10023_);
  or g_12147 (new_n5335_, not_new_n5063__1, not_new_n5062_);
  not g_12148 (not_new_n9109__0, new_n9109_);
  not g_12149 (not_new_n2280_, new_n2280_);
  not g_12150 (not_new_n8544_, new_n8544_);
  or g_12151 (new_n9900_, not_new_n9979_, not_new_n9978_);
  or g_12152 (new_n6102_, not_new_n5761__0, not_new_n5954_);
  or g_12153 (new_n3177_, not_new_n1031__6, not_new_n928__797922662976120010);
  not g_12154 (not_new_n9382_, new_n9382_);
  not g_12155 (not_new_n3492_, new_n3492_);
  not g_12156 (not_new_n3580_, new_n3580_);
  or g_12157 (new_n3044_, not_new_n1027__19773267430, not_new_n1167_);
  not g_12158 (not_new_n1613__70, new_n1613_);
  or g_12159 (new_n1724_, not_pi063, not_new_n1631__113988951853731430);
  not g_12160 (not_new_n4430_, new_n4430_);
  or g_12161 (new_n5020_, not_new_n5416_, not_new_n5415_);
  not g_12162 (not_new_n628__47475615099430, new_n628_);
  or g_12163 (new_n721_, not_new_n3268_, not_new_n3267_);
  not g_12164 (new_n8171_, new_n1596_);
  and g_12165 (new_n4301_, new_n4353_, new_n4352_);
  or g_12166 (or_or_or_not_new_n2794__not_new_n2797__not_new_n2796__not_new_n2798_, not_new_n2798_, or_or_not_new_n2794__not_new_n2797__not_new_n2796_);
  not g_12167 (not_new_n631__5, new_n631_);
  not g_12168 (not_new_n636__1176490, new_n636_);
  or g_12169 (new_n7850_, not_new_n7627_, not_new_n1601__2824752490);
  not g_12170 (new_n5767_, new_n617_);
  or g_12171 (new_n2677_, not_new_n2676_, not_new_n611__2824752490);
  or g_12172 (new_n6857_, not_new_n6480__0, not_new_n1037__168070);
  not g_12173 (not_new_n1039__403536070, new_n1039_);
  and g_12174 (new_n8809_, new_n8807_, new_n9061_);
  not g_12175 (new_n4825_, new_n4738_);
  not g_12176 (not_new_n646__8235430, new_n646_);
  not g_12177 (not_new_n621_, new_n621_);
  or g_12178 (new_n1785_, not_new_n585__0, not_pi250);
  or g_12179 (or_not_new_n9176__not_new_n9177_, not_new_n9177_, not_new_n9176_);
  not g_12180 (not_new_n4521_, new_n4521_);
  not g_12181 (not_new_n3728_, new_n3728_);
  or g_12182 (new_n3497_, not_new_n1536__39098210485829880490, not_pi013_0);
  not g_12183 (not_new_n5468_, new_n5468_);
  not g_12184 (not_new_n618__403536070, new_n618_);
  not g_12185 (not_new_n581__10, new_n581_);
  and g_12186 (and_new_n3052__new_n998_, new_n998_, new_n3052_);
  or g_12187 (new_n951_, not_new_n1925_, or_or_not_new_n1259__not_new_n1257__not_new_n1926_);
  not g_12188 (not_new_n4477_, new_n4477_);
  not g_12189 (not_new_n6058_, new_n6058_);
  or g_12190 (or_or_not_new_n6897__not_new_n6798__not_new_n6826_, or_not_new_n6897__not_new_n6798_, not_new_n6826_);
  not g_12191 (not_pi002, pi002);
  or g_12192 (new_n2983_, not_new_n4115__2, not_new_n3310__8235430);
  not g_12193 (new_n8447_, new_n8272_);
  not g_12194 (not_new_n593__490, new_n593_);
  not g_12195 (not_new_n642__138412872010, new_n642_);
  or g_12196 (new_n3703_, not_new_n629__9, not_po298_6782230728490);
  or g_12197 (new_n8725_, not_new_n8610_, not_new_n1179__0);
  not g_12198 (not_new_n4804_, new_n4804_);
  not g_12199 (not_new_n626__490, new_n626_);
  not g_12200 (not_new_n2053_, new_n2053_);
  or g_12201 (new_n10268_, not_new_n1607__2824752490, not_new_n10008_);
  or g_12202 (po161, not_new_n3549_, not_new_n3548_);
  not g_12203 (not_pi061, pi061);
  not g_12204 (not_new_n7623__0, new_n7623_);
  not g_12205 (new_n9578_, new_n9506_);
  or g_12206 (new_n7675_, not_new_n8006_, not_new_n8005_);
  not g_12207 (not_new_n1010__4, new_n1010_);
  not g_12208 (not_new_n1533_, new_n1533_);
  not g_12209 (new_n4174_, new_n4110_);
  or g_12210 (new_n967_, not_new_n1536__1, not_pi010);
  and g_12211 (and_new_n3070__new_n998_, new_n998_, new_n3070_);
  not g_12212 (not_new_n1020__5, new_n1020_);
  or g_12213 (new_n4619_, not_new_n4617_, not_new_n4618_);
  not g_12214 (new_n8995_, new_n8833_);
  not g_12215 (new_n6512_, new_n1604_);
  not g_12216 (not_new_n991__0, new_n991_);
  not g_12217 (not_new_n8602_, new_n8602_);
  and g_12218 (new_n6324_, new_n6232_, new_n6383_);
  or g_12219 (new_n10317_, not_new_n1603__113988951853731430, not_new_n9911__0);
  not g_12220 (not_new_n601__5, new_n601_);
  or g_12221 (new_n2705_, not_new_n2704_, not_new_n1622__0);
  not g_12222 (new_n2304_, new_n619_);
  not g_12223 (not_new_n3824_, new_n3824_);
  not g_12224 (not_new_n627__16284135979104490, new_n627_);
  not g_12225 (not_new_n8845__2, new_n8845_);
  or g_12226 (new_n1664_, not_pi043, not_new_n1631__9);
  not g_12227 (not_new_n7601_, new_n7601_);
  not g_12228 (not_new_n4772__0, new_n4772_);
  not g_12229 (not_new_n598__3430, new_n598_);
  not g_12230 (not_new_n587__797922662976120010, new_n587_);
  not g_12231 (not_new_n7445_, new_n7445_);
  not g_12232 (not_new_n8504_, new_n8504_);
  or g_12233 (new_n5381_, not_new_n5379_, not_new_n5380_);
  not g_12234 (not_new_n7670__0, new_n7670_);
  not g_12235 (not_new_n4748__0, new_n4748_);
  or g_12236 (po191, not_new_n1365_, or_not_new_n1548__not_new_n1366_);
  or g_12237 (new_n1637_, not_new_n1631__0, not_pi034);
  not g_12238 (not_new_n10146_, new_n10146_);
  or g_12239 (new_n9126_, not_new_n9118_, not_new_n8874__0);
  not g_12240 (not_new_n3375__1, new_n3375_);
  or g_12241 (new_n7188_, not_new_n737_, not_new_n7019_);
  not g_12242 (not_new_n6717_, new_n6717_);
  or g_12243 (new_n8363_, not_new_n1601__6782230728490, not_new_n8134_);
  not g_12244 (not_new_n5433__0, new_n5433_);
  not g_12245 (not_new_n5470__0, new_n5470_);
  not g_12246 (new_n8135_, new_n625_);
  not g_12247 (not_new_n609__9, new_n609_);
  not g_12248 (not_new_n589__185621159210175743024531636712070, new_n589_);
  not g_12249 (not_new_n5572_, new_n5572_);
  not g_12250 (not_new_n4107_, new_n4107_);
  not g_12251 (new_n4837_, new_n4744_);
  or g_12252 (new_n2197_, not_new_n8914_, not_new_n1591__19773267430);
  not g_12253 (not_new_n1534__6, key_gate_5);
  or g_12254 (po242, not_new_n3670_, not_new_n3671_);
  not g_12255 (not_new_n6868_, new_n6868_);
  or g_12256 (new_n9006_, not_new_n8838_, not_new_n8837_);
  not g_12257 (not_new_n4948_, new_n4948_);
  or g_12258 (new_n2829_, not_new_n1041__1, not_new_n3311__7);
  not g_12259 (not_new_n1963_, new_n1963_);
  not g_12260 (not_new_n7006_, new_n7006_);
  or g_12261 (or_not_new_n1406__not_new_n1407_, not_new_n1407_, not_new_n1406_);
  not g_12262 (not_new_n3569_, new_n3569_);
  not g_12263 (new_n1829_, new_n624_);
  not g_12264 (not_new_n768_, new_n768_);
  or g_12265 (new_n3652_, not_pi192_0, not_new_n984__797922662976120010);
  and g_12266 (new_n1242_, new_n1853_, new_n1854_);
  or g_12267 (new_n2778_, not_new_n1616__4, not_new_n2775_);
  not g_12268 (not_new_n3923_, new_n3923_);
  not g_12269 (not_new_n9967__0, new_n9967_);
  not g_12270 (not_new_n8285__0, new_n8285_);
  or g_12271 (po289, not_new_n2929_, or_or_or_not_new_n2928__not_new_n2931__not_new_n2930__not_new_n2932_);
  or g_12272 (new_n8042_, not_new_n7726_, not_new_n7755__0);
  not g_12273 (not_pi179_4, pi179);
  not g_12274 (not_new_n3315__2824752490, new_n3315_);
  not g_12275 (new_n9420_, new_n618_);
  not g_12276 (not_new_n6538__1, new_n6538_);
  not g_12277 (new_n3956_, pi043);
  not g_12278 (new_n8025_, new_n7723_);
  or g_12279 (new_n3261_, not_new_n589__93874803376477543056490, not_new_n1597__5);
  not g_12280 (not_new_n9684_, new_n9684_);
  or g_12281 (new_n6715_, not_new_n6518_, not_new_n637__57648010);
  or g_12282 (new_n10115_, not_new_n633__797922662976120010, not_new_n10114_);
  not g_12283 (not_new_n9819_, new_n9819_);
  not g_12284 (not_new_n6502__0, new_n6502_);
  or g_12285 (new_n2636_, or_not_new_n2635__not_new_n2634_, not_new_n2633_);
  not g_12286 (not_po296_367033682172941254412302110320336601888010, po296);
  not g_12287 (new_n9552_, new_n9375_);
  not g_12288 (not_new_n595__57648010, new_n595_);
  or g_12289 (new_n4596_, not_new_n1003__4, not_new_n4429__0);
  or g_12290 (new_n2048_, not_new_n594__3430, not_new_n9971_);
  not g_12291 (not_new_n4792__0, new_n4792_);
  not g_12292 (not_new_n638__5585458640832840070, new_n638_);
  not g_12293 (not_pi009_0, pi009);
  or g_12294 (new_n1807_, not_pi132, not_new_n587__2);
  or g_12295 (new_n7726_, not_new_n8038_, not_new_n8039_);
  not g_12296 (not_new_n5135_, new_n5135_);
  not g_12297 (not_new_n626__1, new_n626_);
  not g_12298 (not_new_n1159__0, new_n1159_);
  or g_12299 (new_n7444_, not_new_n752_, not_new_n6974__138412872010);
  not g_12300 (not_new_n9159_, new_n9159_);
  not g_12301 (not_new_n6413_, new_n6413_);
  or g_12302 (new_n4688_, not_new_n1016__3, not_new_n4439_);
  not g_12303 (not_new_n5147_, new_n5147_);
  not g_12304 (not_new_n4797_, new_n4797_);
  not g_12305 (not_new_n647__138412872010, new_n647_);
  xor g_12306 (key_gate_110, not_new_n1705_, key_110);
  or g_12307 (new_n4928_, not_new_n624__3430, not_new_n1041__8);
  not g_12308 (not_pi056_2, pi056);
  or g_12309 (new_n6097_, not_new_n5741__2, not_new_n1049__490);
  not g_12310 (not_pi033_5, pi033);
  not g_12311 (not_new_n3115_, new_n3115_);
  not g_12312 (not_new_n3274_, new_n3274_);
  not g_12313 (not_new_n1061__1, new_n1061_);
  or g_12314 (new_n6751_, not_new_n618__2824752490, not_new_n6540_);
  or g_12315 (new_n4696_, not_pi173_2, not_new_n4438_);
  not g_12316 (not_pi259, pi259);
  not g_12317 (new_n7130_, new_n751_);
  not g_12318 (not_new_n644__4, new_n644_);
  or g_12319 (new_n5459_, not_new_n5560_, not_new_n5561_);
  and g_12320 (new_n1244_, and_and_new_n1858__new_n1861__new_n1859_, new_n1860_);
  not g_12321 (not_new_n1904_, new_n1904_);
  or g_12322 (new_n1632_, key_gate_4, key_gate_90);
  or g_12323 (new_n7490_, not_new_n7141__0, not_new_n7140_);
  or g_12324 (new_n3476_, not_new_n1613__3430, not_new_n2052_);
  not g_12325 (not_pi257_2, pi257);
  or g_12326 (new_n10101_, new_n644_, new_n1059_);
  or g_12327 (new_n6012_, not_new_n5767__0, not_new_n5766_);
  not g_12328 (not_new_n9741_, new_n9741_);
  not g_12329 (not_new_n9576_, new_n9576_);
  or g_12330 (new_n2529_, not_pi259, not_po296_273687473400809163430);
  or g_12331 (new_n10085_, not_new_n9890__1, not_new_n9893__0);
  and g_12332 (new_n1304_, and_and_new_n2143__new_n2146__new_n2144_, new_n2145_);
  not g_12333 (not_new_n7197_, new_n7197_);
  or g_12334 (new_n7491_, not_new_n7248_, not_new_n7489_);
  or g_12335 (new_n9715_, or_not_new_n9631__not_new_n9515__0, not_new_n9507__0);
  or g_12336 (new_n9696_, not_new_n9326__2, or_not_new_n9523__1_not_new_n9327__1);
  not g_12337 (not_new_n1212_, new_n1212_);
  and g_12338 (new_n7586_, new_n7981_, new_n7982_);
  or g_12339 (new_n9721_, not_new_n1051__968890104070, not_new_n9370_);
  or g_12340 (new_n2993_, not_new_n1049__2, not_new_n581__1);
  or g_12341 (or_not_new_n2964__not_new_n2967_, not_new_n2964_, not_new_n2967_);
  not g_12342 (not_new_n584__0, new_n584_);
  not g_12343 (not_new_n1168__0, new_n1168_);
  not g_12344 (not_new_n2959_, new_n2959_);
  not g_12345 (not_new_n589__332329305696010, new_n589_);
  or g_12346 (new_n8584_, not_new_n8155__2, not_new_n1055__2326305139872070);
  not g_12347 (not_new_n4015_, new_n4015_);
  not g_12348 (not_new_n687_, new_n687_);
  not g_12349 (not_new_n586__968890104070, new_n586_);
  not g_12350 (not_new_n10042__0, new_n10042_);
  or g_12351 (new_n2278_, not_new_n4769_, not_new_n591__332329305696010);
  not g_12352 (not_pi055_1, pi055);
  not g_12353 (not_new_n4999__0, new_n4999_);
  and g_12354 (new_n6351_, new_n6434_, new_n6435_);
  not g_12355 (not_new_n599__138412872010, new_n599_);
  not g_12356 (not_new_n3690_, new_n3690_);
  or g_12357 (new_n3149_, not_new_n633__5, not_new_n3315__19773267430);
  or g_12358 (new_n6034_, not_new_n6033_, not_new_n6068_);
  or g_12359 (new_n9713_, not_new_n1598__47475615099430, not_new_n9625__0);
  not g_12360 (not_new_n1583__8, new_n1583_);
  or g_12361 (new_n3039_, not_new_n1602__2, not_new_n581__1176490);
  not g_12362 (not_new_n3683_, new_n3683_);
  not g_12363 (not_new_n1037__70, new_n1037_);
  not g_12364 (not_new_n1440_, new_n1440_);
  or g_12365 (or_or_not_new_n2189__not_new_n2186__not_new_n2187_, not_new_n2187_, or_not_new_n2189__not_new_n2186_);
  not g_12366 (not_new_n9108_, new_n9108_);
  or g_12367 (new_n7280_, not_new_n7279_, not_new_n7091_);
  not g_12368 (not_new_n8800_, new_n8800_);
  not g_12369 (not_new_n5084__2, new_n5084_);
  not g_12370 (not_new_n6504__0, new_n6504_);
  or g_12371 (new_n9528_, not_new_n631__13410686196639649008070, not_new_n9527_);
  and g_12372 (new_n6322_, and_and_and_new_n6227__new_n6232__new_n6229__new_n6317_, new_n6231_);
  not g_12373 (not_new_n8065_, new_n8065_);
  not g_12374 (not_new_n646__2326305139872070, new_n646_);
  not g_12375 (not_new_n7396_, new_n7396_);
  not g_12376 (not_new_n1041__5, new_n1041_);
  or g_12377 (new_n636_, or_or_not_new_n1977__not_new_n1978__not_new_n1980_, not_new_n1979_);
  not g_12378 (not_new_n8471_, new_n8471_);
  not g_12379 (not_new_n1213_, new_n1213_);
  not g_12380 (not_new_n1065__39098210485829880490, new_n1065_);
  not g_12381 (not_new_n3235_, new_n3235_);
  not g_12382 (not_new_n642__5, new_n642_);
  and g_12383 (and_new_n1217__new_n1218_, new_n1218_, new_n1217_);
  or g_12384 (new_n6065_, not_new_n5900__3, not_new_n5851_);
  not g_12385 (not_new_n4807__0, new_n4807_);
  and g_12386 (and_new_n2992__new_n998_, new_n998_, new_n2992_);
  or g_12387 (new_n9435_, not_new_n9748_, not_new_n9747_);
  not g_12388 (not_new_n2611_, new_n2611_);
  and g_12389 (new_n7702_, new_n7570_, new_n7814_);
  not g_12390 (not_new_n8191_, new_n8191_);
  not g_12391 (not_new_n3785_, new_n3785_);
  not g_12392 (not_new_n4424_, new_n4424_);
  not g_12393 (not_new_n4596_, new_n4596_);
  or g_12394 (new_n6936_, not_new_n638__6782230728490, not_new_n6519__2);
  not g_12395 (not_new_n2091_, new_n2091_);
  not g_12396 (not_new_n1041__6, new_n1041_);
  or g_12397 (new_n6389_, not_new_n6289_, not_new_n645__8235430);
  not g_12398 (not_new_n5341_, new_n5341_);
  or g_12399 (new_n8896_, not_new_n9072_, not_new_n9071_);
  not g_12400 (not_new_n1597__968890104070, new_n1597_);
  not g_12401 (not_new_n1035__24010, new_n1035_);
  or g_12402 (new_n10321_, not_new_n10043_, not_new_n10023_);
  not g_12403 (new_n9109_, new_n8894_);
  not g_12404 (not_new_n7303_, new_n7303_);
  not g_12405 (not_new_n1049__0, new_n1049_);
  not g_12406 (not_new_n10218_, new_n10218_);
  and g_12407 (new_n6365_, and_new_n6440__new_n6441_, new_n6442_);
  not g_12408 (not_new_n1613__113988951853731430, new_n1613_);
  not g_12409 (new_n4767_, new_n1598_);
  not g_12410 (not_new_n7642__0, new_n7642_);
  not g_12411 (not_new_n4715_, new_n4715_);
  or g_12412 (new_n2270_, not_new_n9345_, not_new_n1584__47475615099430);
  or g_12413 (new_n1179_, not_new_n3887_, not_new_n3888_);
  not g_12414 (not_pi059_2, pi059);
  or g_12415 (new_n7554_, not_new_n7032__0, not_new_n6996__0);
  not g_12416 (not_new_n9889_, new_n9889_);
  not g_12417 (not_new_n1413_, new_n1413_);
  not g_12418 (not_new_n3148_, new_n3148_);
  and g_12419 (and_not_pi040_3_not_pi041_2, not_pi041_2, not_pi040_3);
  or g_12420 (new_n6769_, not_new_n6768_, not_new_n6651__0);
  not g_12421 (not_new_n607__4, new_n607_);
  not g_12422 (not_new_n8294_, new_n8294_);
  not g_12423 (not_new_n1588__6782230728490, new_n1588_);
  and g_12424 (new_n4313_, new_n4388_, new_n4389_);
  not g_12425 (not_new_n639__39098210485829880490, new_n639_);
  or g_12426 (new_n3727_, not_new_n640__10, not_new_n1604__6);
  or g_12427 (new_n3086_, not_new_n1051__3, not_new_n928_);
  not g_12428 (new_n9903_, new_n1071_);
  and g_12429 (new_n1487_, new_n2990_, and_new_n2992__new_n998_);
  not g_12430 (not_new_n7146_, new_n7146_);
  and g_12431 (new_n8230_, new_n8368_, new_n8089_);
  not g_12432 (not_new_n950_, new_n950_);
  not g_12433 (not_new_n610__24010, new_n610_);
  not g_12434 (not_new_n626__47475615099430, new_n626_);
  not g_12435 (not_new_n3368_, new_n3368_);
  not g_12436 (not_new_n633__968890104070, new_n633_);
  not g_12437 (not_new_n9636_, new_n9636_);
  or g_12438 (new_n6827_, not_new_n6598_, not_new_n6896_);
  not g_12439 (not_new_n5116_, new_n5116_);
  not g_12440 (not_new_n647__332329305696010, new_n647_);
  not g_12441 (not_new_n8992_, new_n8992_);
  not g_12442 (not_new_n4451_, new_n4451_);
  not g_12443 (not_new_n8225_, new_n8225_);
  not g_12444 (not_new_n7759_, new_n7759_);
  not g_12445 (not_new_n1830_, new_n1830_);
  not g_12446 (new_n2104_, new_n960_);
  or g_12447 (or_not_new_n10219__not_new_n10220_, not_new_n10220_, not_new_n10219_);
  or g_12448 (new_n6850_, not_new_n6617__2, not_new_n6700_);
  not g_12449 (not_new_n1031__70, new_n1031_);
  not g_12450 (not_new_n9934_, new_n9934_);
  not g_12451 (not_new_n1591__7, new_n1591_);
  not g_12452 (not_new_n6457_, new_n6457_);
  not g_12453 (not_new_n2653_, new_n2653_);
  or g_12454 (or_not_new_n2980__not_new_n2979_, not_new_n2980_, not_new_n2979_);
  not g_12455 (not_new_n599__16284135979104490, new_n599_);
  or g_12456 (new_n5337_, not_new_n4948_, not_new_n617__24010);
  or g_12457 (new_n4731_, not_new_n4735_, or_not_new_n4814__not_new_n4734_);
  not g_12458 (not_new_n1603__403536070, new_n1603_);
  or g_12459 (new_n7053_, not_new_n7402_, not_new_n7403_);
  not g_12460 (not_new_n1604__6782230728490, new_n1604_);
  not g_12461 (new_n4780_, new_n1603_);
  not g_12462 (new_n8106_, new_n1043_);
  or g_12463 (new_n8911_, not_new_n9249_, not_new_n9250_);
  not g_12464 (not_new_n7124_, new_n7124_);
  not g_12465 (not_new_n648__7, new_n648_);
  not g_12466 (not_new_n1027__39098210485829880490, new_n1027_);
  not g_12467 (not_new_n5183_, new_n5183_);
  not g_12468 (not_new_n628__8, new_n628_);
  or g_12469 (new_n5273_, not_new_n5078__1, not_new_n4909_);
  not g_12470 (not_new_n5452_, new_n5452_);
  not g_12471 (not_pi176_3, pi176);
  not g_12472 (not_new_n3387_, new_n3387_);
  or g_12473 (new_n7985_, not_new_n7984_, not_new_n7983_);
  not g_12474 (not_new_n1599__19773267430, new_n1599_);
  not g_12475 (not_new_n3661_, new_n3661_);
  not g_12476 (not_pi154, pi154);
  not g_12477 (new_n5917_, new_n5893_);
  not g_12478 (not_new_n1611__2824752490, new_n1611_);
  and g_12479 (new_n8922_, new_n8923_, new_n8991_);
  not g_12480 (not_new_n629__70, new_n629_);
  not g_12481 (not_new_n2757_, new_n2757_);
  not g_12482 (not_new_n8333_, new_n8333_);
  not g_12483 (not_new_n1377_, new_n1377_);
  not g_12484 (not_new_n6663_, new_n6663_);
  not g_12485 (not_new_n5066__0, new_n5066_);
  not g_12486 (not_new_n7020__0, new_n7020_);
  or g_12487 (new_n4453_, not_new_n4593_, not_new_n4592_);
  not g_12488 (not_new_n9972__0, new_n9972_);
  not g_12489 (not_new_n7721_, new_n7721_);
  not g_12490 (not_new_n1067__19773267430, new_n1067_);
  or g_12491 (new_n8724_, not_new_n8637_, not_new_n1053__2824752490);
  or g_12492 (new_n4880_, not_new_n4790_, not_new_n1069__7);
  not g_12493 (new_n5508_, pi148);
  not g_12494 (not_new_n1604_, new_n1604_);
  or g_12495 (new_n2647_, not_new_n611__8235430, not_new_n2646_);
  not g_12496 (not_new_n9816_, new_n9816_);
  not g_12497 (not_new_n5741__2, new_n5741_);
  not g_12498 (not_new_n7004__0, new_n7004_);
  not g_12499 (not_new_n699_, new_n699_);
  not g_12500 (not_new_n928__2824752490, new_n928_);
  or g_12501 (or_not_new_n2747__not_new_n2746_, not_new_n2746_, not_new_n2747_);
  not g_12502 (not_new_n4983_, new_n4983_);
  or g_12503 (new_n5695_, not_new_n5694_, not_new_n5693_);
  or g_12504 (new_n1002_, not_new_n3325_, not_new_n3326_);
  or g_12505 (new_n6711_, not_new_n6523_, not_new_n636__403536070);
  or g_12506 (new_n7159_, not_new_n733_, not_new_n7030_);
  not g_12507 (new_n9354_, new_n624_);
  and g_12508 (new_n4291_, and_new_n4327__new_n4331_, new_n4328_);
  or g_12509 (new_n3133_, not_new_n625__6, not_new_n581__1299348114471230201171721456984490);
  not g_12510 (not_new_n2586_, new_n2586_);
  and g_12511 (and_and_new_n2707__new_n2708__new_n3822_, new_n3822_, and_new_n2707__new_n2708_);
  or g_12512 (new_n7594_, not_new_n7804_, not_new_n7806_);
  not g_12513 (not_new_n6075_, new_n6075_);
  not g_12514 (not_new_n1631_, key_gate_76);
  not g_12515 (not_new_n6068__0, new_n6068_);
  or g_12516 (new_n3446_, not_new_n1613__7, not_new_n1938_);
  or g_12517 (new_n6980_, not_new_n740_, not_new_n7022_);
  not g_12518 (not_new_n4124__2, new_n4124_);
  or g_12519 (new_n1782_, not_pi163, not_new_n586__0);
  and g_12520 (new_n6630_, new_n6904_, new_n6903_);
  and g_12521 (new_n6363_, and_new_n6362__new_n6430_, new_n6429_);
  not g_12522 (not_new_n1175_, new_n1175_);
  not g_12523 (not_new_n3488_, new_n3488_);
  not g_12524 (not_new_n7907_, new_n7907_);
  or g_12525 (new_n3767_, not_new_n1049__6, not_new_n648__10);
  not g_12526 (not_new_n3105_, new_n3105_);
  not g_12527 (not_new_n3928__0, new_n3928_);
  not g_12528 (not_pi059_1, pi059);
  or g_12529 (new_n8543_, not_new_n1035__490, not_new_n8116_);
  not g_12530 (not_new_n7620__1, new_n7620_);
  not g_12531 (not_new_n9225_, new_n9225_);
  not g_12532 (not_new_n8119_, new_n8119_);
  not g_12533 (not_new_n3816_, new_n3816_);
  and g_12534 (new_n1378_, new_n2431_, new_n2430_);
  not g_12535 (not_new_n2563_, new_n2563_);
  not g_12536 (not_new_n5597__1, new_n5597_);
  not g_12537 (not_new_n591__7, new_n591_);
  or g_12538 (new_n3111_, not_new_n928__8, not_new_n1607__2);
  not g_12539 (not_new_n1055__490, new_n1055_);
  or g_12540 (po237, not_new_n3660_, not_new_n3661_);
  not g_12541 (not_new_n625__657123623635342801395430, new_n625_);
  or g_12542 (new_n5190_, new_n625_, new_n1602_);
  not g_12543 (new_n9403_, new_n1604_);
  or g_12544 (new_n6115_, not_new_n5749__1, not_new_n1039__490);
  or g_12545 (new_n10122_, not_new_n10121_, not_new_n9949_);
  not g_12546 (new_n8825_, new_n1041_);
  not g_12547 (not_new_n7594_, new_n7594_);
  not g_12548 (new_n5439_, new_n1007_);
  or g_12549 (new_n3796_, not_new_n1867_, not_new_n3434_);
  or g_12550 (new_n954_, or_or_not_new_n1271__not_new_n1269__not_new_n1983_, not_new_n1982_);
  not g_12551 (not_pi221, pi221);
  not g_12552 (not_new_n8048_, new_n8048_);
  not g_12553 (not_new_n1584__2824752490, new_n1584_);
  or g_12554 (new_n5245_, not_new_n1059__10, not_new_n644__168070);
  not g_12555 (not_new_n992_, new_n992_);
  not g_12556 (not_new_n5706_, new_n5706_);
  or g_12557 (new_n3117_, not_new_n928__10, not_new_n1597__3);
  not g_12558 (new_n9910_, new_n1603_);
  not g_12559 (not_new_n7912_, new_n7912_);
  not g_12560 (not_new_n5093_, new_n5093_);
  not g_12561 (not_po296_9095436801298611408202050198891430, po296);
  not g_12562 (not_new_n4946__0, new_n4946_);
  or g_12563 (new_n5940_, not_new_n5721_, not_new_n5882_);
  and g_12564 (new_n8805_, new_n9077_, new_n8804_);
  or g_12565 (new_n9969_, not_new_n10339_, not_new_n10338_);
  not g_12566 (not_new_n2920_, new_n2920_);
  not g_12567 (not_new_n8650_, new_n8650_);
  or g_12568 (or_not_new_n7906__not_new_n7780_, not_new_n7906_, not_new_n7780_);
  or g_12569 (po188, not_new_n1359_, or_not_new_n1545__not_new_n1360_);
  or g_12570 (or_not_new_n8448__not_new_n8419_, not_new_n8419_, not_new_n8448_);
  and g_12571 (new_n7093_, and_new_n6993__new_n7526_, new_n7525_);
  or g_12572 (new_n3343_, not_new_n1534__3430, not_pi051_0);
  and g_12573 (new_n7090_, new_n6965_, new_n7273_);
  not g_12574 (not_new_n598__113988951853731430, new_n598_);
  and g_12575 (new_n1561_, new_n3635_, new_n3634_);
  not g_12576 (not_new_n6245_, new_n6245_);
  not g_12577 (not_new_n1069__10, new_n1069_);
  or g_12578 (new_n2663_, not_new_n609__168070, not_new_n4459_);
  and g_12579 (new_n604_, new_n1595_, new_n1021_);
  or g_12580 (new_n1642_, key_gate_31, not_new_n596__2);
  not g_12581 (not_new_n5412_, new_n5412_);
  and g_12582 (and_new_n2276__new_n2279_, new_n2276_, new_n2279_);
  or g_12583 (new_n7543_, not_new_n7542_, not_new_n7541_);
  not g_12584 (not_new_n8854_, new_n8854_);
  not g_12585 (not_new_n7162_, new_n7162_);
  or g_12586 (new_n6045_, not_new_n5941_, not_new_n5722_);
  or g_12587 (new_n4758_, not_new_n4760__0, not_new_n4843__0);
  or g_12588 (new_n10326_, not_new_n10205_, not_new_n9950__1);
  or g_12589 (new_n5255_, not_new_n5111__0, not_new_n4959__0);
  and g_12590 (new_n5028_, new_n5302_, and_new_n4937__new_n5303_);
  or g_12591 (new_n1681_, key_gate_46, not_new_n596__168070);
  not g_12592 (not_new_n8368_, new_n8368_);
  not g_12593 (not_new_n4089_, new_n4089_);
  and g_12594 (new_n7078_, new_n7159_, new_n7210_);
  not g_12595 (not_new_n8082_, new_n8082_);
  not g_12596 (not_new_n4926_, new_n4926_);
  or g_12597 (new_n6687_, not_new_n6656_, not_new_n6494_);
  not g_12598 (not_new_n7432_, new_n7432_);
  not g_12599 (not_new_n5800_, new_n5800_);
  not g_12600 (not_new_n5975_, new_n5975_);
  or g_12601 (new_n6468_, not_new_n6701_, not_new_n6822_);
  or g_12602 (new_n8900_, not_new_n8866_, not_new_n9139_);
  not g_12603 (not_new_n7244_, new_n7244_);
  not g_12604 (not_new_n8351_, new_n8351_);
  not g_12605 (not_new_n4232_, new_n4232_);
  and g_12606 (new_n1475_, new_n590_, new_n2724_);
  not g_12607 (not_new_n4802__0, new_n4802_);
  not g_12608 (new_n2294_, new_n978_);
  and g_12609 (new_n7757_, new_n8052_, new_n8051_);
  not g_12610 (not_new_n6671_, new_n6671_);
  not g_12611 (not_pi136_3, pi136);
  not g_12612 (not_new_n9645_, new_n9645_);
  or g_12613 (new_n2469_, not_new_n599__138412872010, not_new_n9965__0);
  and g_12614 (new_n1249_, new_n1889_, new_n1890_);
  not g_12615 (not_new_n9854__2, new_n9854_);
  not g_12616 (not_new_n8201_, new_n8201_);
  not g_12617 (not_new_n8426_, new_n8426_);
  not g_12618 (not_new_n3185__7, new_n3185_);
  or g_12619 (new_n1973_, not_new_n593__9, not_new_n627_);
  not g_12620 (not_new_n1041__3430, new_n1041_);
  or g_12621 (new_n3040_, not_new_n3372__2824752490, not_new_n625__4);
  not g_12622 (new_n9920_, new_n1053_);
  or g_12623 (new_n9214_, not_new_n8846__0, not_new_n9157_);
  or g_12624 (or_or_not_new_n2946__not_new_n2949__not_new_n2948_, not_new_n2948_, or_not_new_n2946__not_new_n2949_);
  not g_12625 (not_new_n644__332329305696010, new_n644_);
  or g_12626 (new_n5825_, not_new_n6214_, not_new_n6215_);
  or g_12627 (new_n8548_, not_new_n8142__0, not_new_n1071__57648010);
  not g_12628 (not_new_n9725_, new_n9725_);
  not g_12629 (not_new_n631__2824752490, new_n631_);
  not g_12630 (not_new_n1441_, new_n1441_);
  not g_12631 (not_new_n1015__2, new_n1015_);
  not g_12632 (not_new_n5380_, new_n5380_);
  or g_12633 (new_n4473_, not_new_n4540_, not_new_n4539_);
  not g_12634 (not_new_n640__113988951853731430, new_n640_);
  not g_12635 (not_pi261_1, pi261);
  not g_12636 (not_new_n3919__0, new_n3919_);
  not g_12637 (not_new_n4663_, new_n4663_);
  or g_12638 (new_n3211_, not_new_n589__70, not_new_n630__7);
  or g_12639 (po079, not_new_n1206_, key_gate_96);
  not g_12640 (not_new_n9537_, new_n9537_);
  or g_12641 (new_n8731_, not_new_n1041__403536070, not_new_n8631_);
  and g_12642 (and_new_n2200__new_n2203_, new_n2203_, new_n2200_);
  or g_12643 (new_n5559_, pi141, new_n1017_);
  not g_12644 (not_new_n7049_, new_n7049_);
  not g_12645 (not_new_n2074_, new_n2074_);
  not g_12646 (not_new_n2553_, new_n2553_);
  or g_12647 (new_n8309_, not_new_n8105_, not_new_n1049__2824752490);
  not g_12648 (not_new_n647__70, new_n647_);
  or g_12649 (new_n8355_, not_new_n8147_, not_new_n1067__8235430);
  or g_12650 (or_not_new_n6373__not_new_n6413_, not_new_n6373_, not_new_n6413_);
  not g_12651 (not_new_n8883_, new_n8883_);
  not g_12652 (not_new_n4934_, new_n4934_);
  not g_12653 (not_new_n7607_, new_n7607_);
  and g_12654 (and_new_n1858__new_n1861_, new_n1858_, new_n1861_);
  or g_12655 (new_n3447_, not_pi023_0, not_new_n1536__138412872010);
  or g_12656 (new_n8507_, not_new_n8170__2, not_new_n1597__138412872010);
  not g_12657 (not_new_n8271_, new_n8271_);
  or g_12658 (new_n4646_, or_not_new_n4414__0_not_new_n1010__3, not_new_n4415__1);
  not g_12659 (not_pi224, pi224);
  not g_12660 (not_new_n7329_, new_n7329_);
  not g_12661 (not_new_n1053__47475615099430, new_n1053_);
  not g_12662 (not_new_n8139__0, new_n8139_);
  not g_12663 (not_new_n1596__16284135979104490, new_n1596_);
  not g_12664 (not_new_n4031_, new_n4031_);
  not g_12665 (not_new_n628__657123623635342801395430, new_n628_);
  not g_12666 (not_new_n1602__2, new_n1602_);
  or g_12667 (new_n4620_, not_new_n4480_, not_new_n4481__0);
  not g_12668 (not_new_n3372__5, new_n3372_);
  not g_12669 (not_new_n3162_, new_n3162_);
  not g_12670 (not_new_n4619_, new_n4619_);
  not g_12671 (not_new_n1247_, new_n1247_);
  not g_12672 (not_pi095, pi095);
  or g_12673 (new_n6374_, not_new_n6302_, not_new_n617__403536070);
  not g_12674 (not_new_n1437_, new_n1437_);
  or g_12675 (or_not_new_n2497__not_new_n1568_, not_new_n2497_, not_new_n1568_);
  not g_12676 (not_new_n4123_, new_n4123_);
  or g_12677 (new_n3640_, not_new_n984__6782230728490, not_pi186_0);
  not g_12678 (not_new_n1248_, new_n1248_);
  not g_12679 (not_new_n7644__0, new_n7644_);
  and g_12680 (new_n1391_, new_n2462_, new_n2463_);
  and g_12681 (and_new_n1801__new_n1804_, new_n1804_, new_n1801_);
  not g_12682 (not_new_n1576__9, new_n1576_);
  or g_12683 (new_n7502_, not_new_n7004__2, not_new_n7039__0);
  not g_12684 (not_new_n6373__4, new_n6373_);
  not g_12685 (not_new_n1037__6782230728490, new_n1037_);
  or g_12686 (new_n3007_, not_new_n3372__9, not_new_n624__4);
  or g_12687 (new_n4571_, not_new_n4570_, not_new_n4496_);
  or g_12688 (new_n6178_, not_new_n6177_, not_new_n5926_);
  not g_12689 (not_new_n2676_, new_n2676_);
  not g_12690 (new_n8981_, new_n8828_);
  not g_12691 (not_new_n7470_, new_n7470_);
  not g_12692 (not_new_n5460_, new_n5460_);
  not g_12693 (not_new_n3667_, new_n3667_);
  not g_12694 (not_new_n585__490, new_n585_);
  not g_12695 (not_new_n4168_, new_n4168_);
  not g_12696 (not_new_n1601__24010, new_n1601_);
  not g_12697 (not_new_n1538__3, new_n1538_);
  or g_12698 (or_or_not_new_n1331__not_new_n1329__not_new_n2268_, or_not_new_n1331__not_new_n1329_, not_new_n2268_);
  not g_12699 (not_new_n9318_, new_n9318_);
  not g_12700 (not_new_n8177_, new_n8177_);
  not g_12701 (not_new_n600__1, new_n600_);
  not g_12702 (new_n8605_, new_n1043_);
  not g_12703 (not_new_n643__70, new_n643_);
  not g_12704 (not_new_n5425_, new_n5425_);
  not g_12705 (not_new_n7007__0, new_n7007_);
  not g_12706 (not_new_n6918_, new_n6918_);
  not g_12707 (not_new_n2887_, new_n2887_);
  or g_12708 (new_n8473_, not_new_n8107__0, not_new_n635__968890104070);
  not g_12709 (not_new_n1611__0, new_n1611_);
  not g_12710 (not_new_n9540_, new_n9540_);
  or g_12711 (new_n8895_, not_new_n9179_, not_new_n9088_);
  not g_12712 (not_new_n7367_, new_n7367_);
  or g_12713 (new_n4730_, or_not_new_n4812__not_new_n4736_, not_new_n4737_);
  not g_12714 (not_new_n1531_, new_n1531_);
  or g_12715 (or_not_new_n4835__not_new_n4777_, not_new_n4835_, not_new_n4777_);
  not g_12716 (not_new_n4780__0, new_n4780_);
  not g_12717 (not_new_n2605_, new_n2605_);
  not g_12718 (not_new_n7906_, new_n7906_);
  or g_12719 (new_n3890_, not_new_n1576__797922662976120010, not_new_n641__10);
  not g_12720 (new_n5742_, new_n1043_);
  not g_12721 (not_new_n3976__0, new_n3976_);
  not g_12722 (not_new_n6577_, new_n6577_);
  or g_12723 (new_n5975_, not_new_n5796_, not_new_n1057__70);
  not g_12724 (not_new_n1613__2326305139872070, new_n1613_);
  or g_12725 (new_n2640_, not_new_n1005__0, not_new_n608__490);
  or g_12726 (new_n8052_, not_new_n7643__2, not_new_n638__16284135979104490);
  not g_12727 (not_new_n9403_, new_n9403_);
  not g_12728 (not_new_n6737__1, new_n6737_);
  or g_12729 (new_n5965_, not_new_n5938__0, not_new_n5757__0);
  or g_12730 (new_n2129_, not_new_n586__403536070, not_pi181);
  not g_12731 (not_new_n7651__2, new_n7651_);
  not g_12732 (not_new_n10041__0, new_n10041_);
  not g_12733 (new_n2076_, new_n633_);
  or g_12734 (new_n10248_, not_new_n9876_, not_new_n635__113988951853731430);
  not g_12735 (new_n6256_, new_n631_);
  not g_12736 (not_new_n630__8235430, new_n630_);
  or g_12737 (new_n3374_, not_pi064_332329305696010, not_new_n3923__0);
  or g_12738 (new_n6159_, not_new_n6157_, not_new_n6158_);
  not g_12739 (new_n6986_, new_n745_);
  not g_12740 (not_new_n4930_, new_n4930_);
  not g_12741 (not_new_n1598__3, new_n1598_);
  or g_12742 (new_n8757_, not_new_n8659_, not_new_n8756_);
  not g_12743 (new_n5554_, new_n5517_);
  not g_12744 (not_new_n594__1, new_n594_);
  or g_12745 (new_n4049_, not_new_n3936_, not_pi041_3);
  not g_12746 (not_new_n4802_, new_n4802_);
  not g_12747 (not_new_n5210_, new_n5210_);
  or g_12748 (new_n4201_, not_pi252_1, not_new_n4100_);
  or g_12749 (new_n2364_, not_new_n599__1, not_new_n9873__0);
  not g_12750 (not_new_n1921_, new_n1921_);
  not g_12751 (not_new_n618__19773267430, new_n618_);
  or g_12752 (new_n5392_, not_new_n1065__9, not_new_n4982_);
  not g_12753 (new_n4078_, pi266);
  or g_12754 (new_n3547_, not_new_n1976__0, not_new_n1612__9);
  or g_12755 (new_n2366_, not_new_n4723__0, not_new_n597__1);
  not g_12756 (not_new_n3216_, new_n3216_);
  or g_12757 (new_n1686_, not_pi014, not_po296_8235430);
  not g_12758 (not_new_n581__0, new_n581_);
  not g_12759 (not_pi268, pi268);
  not g_12760 (new_n4034_, new_n3989_);
  not g_12761 (not_new_n3035_, new_n3035_);
  not g_12762 (not_new_n9351_, new_n9351_);
  not g_12763 (not_new_n8897__0, new_n8897_);
  not g_12764 (not_new_n5196_, new_n5196_);
  not g_12765 (not_new_n640__5, new_n640_);
  or g_12766 (new_n5168_, new_n637_, new_n1065_);
  or g_12767 (po152, not_new_n3531_, not_new_n3530_);
  not g_12768 (new_n6010_, new_n5890_);
  not g_12769 (new_n6304_, new_n1607_);
  or g_12770 (po124, not_new_n3435_, not_new_n3436_);
  not g_12771 (not_new_n1041__0, new_n1041_);
  not g_12772 (not_new_n607__0, new_n607_);
  not g_12773 (not_new_n1416_, new_n1416_);
  not g_12774 (not_new_n4115_, new_n4115_);
  not g_12775 (not_new_n9523_, new_n9523_);
  or g_12776 (new_n5692_, not_pi141_2, not_new_n5458_);
  not g_12777 (not_new_n1055__57648010, new_n1055_);
  not g_12778 (not_new_n8064_, new_n8064_);
  not g_12779 (not_new_n5199_, new_n5199_);
  or g_12780 (new_n1880_, not_new_n1588__5, not_new_n1043_);
  not g_12781 (not_new_n6452_, new_n6452_);
  not g_12782 (not_new_n5889_, new_n5889_);
  not g_12783 (not_new_n3677_, new_n3677_);
  and g_12784 (po108, key_gate_101, pi087);
  not g_12785 (not_new_n6146_, new_n6146_);
  or g_12786 (new_n9842_, not_new_n9840_, not_new_n9841_);
  or g_12787 (or_not_new_n9612__not_new_n9611_, not_new_n9612_, not_new_n9611_);
  not g_12788 (not_new_n9987_, new_n9987_);
  or g_12789 (new_n3302_, not_new_n3184__2326305139872070, not_new_n641__6);
  not g_12790 (not_pi109, pi109);
  not g_12791 (new_n5446_, new_n1004_);
  not g_12792 (not_new_n999__1, new_n999_);
  not g_12793 (not_new_n1065_, new_n1065_);
  not g_12794 (not_pi250_2, pi250);
  not g_12795 (not_new_n5108_, new_n5108_);
  not g_12796 (not_new_n1598__7, new_n1598_);
  or g_12797 (new_n4598_, not_new_n4596_, not_new_n4597_);
  or g_12798 (or_not_new_n2695__not_new_n2694_, not_new_n2694_, not_new_n2695_);
  not g_12799 (new_n3988_, pi056);
  not g_12800 (not_new_n7996_, new_n7996_);
  not g_12801 (not_new_n7890_, new_n7890_);
  or g_12802 (new_n2287_, not_new_n7590_, not_new_n1583__332329305696010);
  or g_12803 (or_not_new_n3091__not_new_n3090_, not_new_n3090_, not_new_n3091_);
  or g_12804 (po218, not_new_n1424_, or_or_not_new_n2547__not_new_n2551__not_new_n1425_);
  not g_12805 (not_new_n9894_, new_n9894_);
  or g_12806 (new_n2036_, not_pi112, not_new_n588__24010);
  not g_12807 (not_new_n6544_, new_n6544_);
  and g_12808 (new_n8684_, new_n1172_, new_n8611_);
  or g_12809 (new_n9048_, new_n626_, new_n1053_);
  not g_12810 (not_pi031_0, pi031);
  not g_12811 (not_new_n1764_, new_n1764_);
  or g_12812 (new_n2318_, not_new_n2313_, not_new_n1340_);
  not g_12813 (not_new_n4484_, new_n4484_);
  and g_12814 (new_n4720_, new_n4722_, new_n4721_);
  not g_12815 (not_new_n8963__1, new_n8963_);
  and g_12816 (new_n4771_, new_n4864_, new_n4865_);
  not g_12817 (not_new_n645__19773267430, new_n645_);
  not g_12818 (not_new_n2931_, new_n2931_);
  not g_12819 (not_new_n5527_, new_n5527_);
  or g_12820 (new_n2623_, not_new_n4455_, not_new_n609__70);
  not g_12821 (not_new_n6051_, new_n6051_);
  not g_12822 (not_new_n3374_, new_n3374_);
  or g_12823 (new_n7753_, not_new_n7673_, not_new_n1031__1176490);
  or g_12824 (new_n1864_, not_new_n587__5, not_pi135);
  not g_12825 (not_new_n622__2326305139872070, new_n622_);
  or g_12826 (new_n8749_, not_new_n8675_, not_new_n8746_);
  and g_12827 (new_n6338_, new_n6228_, new_n1047_);
  or g_12828 (or_not_new_n3110__not_new_n3109_, not_new_n3110_, not_new_n3109_);
  not g_12829 (not_new_n1187_, new_n1187_);
  not g_12830 (not_pi215, pi215);
  not g_12831 (not_pi016, pi016);
  or g_12832 (new_n923_, not_new_n1626_, not_new_n3315__0);
  not g_12833 (not_new_n758_, new_n758_);
  xnor g_12834 (key_gate_76, new_n1631_, key_76);
  or g_12835 (new_n3156_, not_new_n1063__3, not_new_n928__968890104070);
  or g_12836 (new_n8075_, not_new_n7762_, not_new_n7934__0);
  or g_12837 (new_n2295_, not_new_n594__332329305696010, not_new_n9962_);
  not g_12838 (not_new_n9635_, new_n9635_);
  not g_12839 (not_new_n1445_, new_n1445_);
  or g_12840 (new_n9674_, not_new_n9481_, not_new_n9672_);
  or g_12841 (new_n2615_, not_new_n605__10, not_new_n5477_);
  or g_12842 (new_n6613_, not_new_n6784_, not_new_n6574_);
  not g_12843 (not_new_n1605__1, new_n1605_);
  not g_12844 (not_new_n4683_, new_n4683_);
  and g_12845 (new_n1497_, new_n998_, new_n3018_);
  or g_12846 (po142, not_new_n3511_, not_new_n3510_);
  and g_12847 (and_new_n1238__new_n1837_, new_n1837_, new_n1238_);
  or g_12848 (new_n5816_, not_new_n6134_, not_new_n6135_);
  not g_12849 (new_n6492_, new_n1051_);
  or g_12850 (new_n3841_, not_new_n6443__6, not_new_n4718_);
  not g_12851 (not_new_n4431__0, new_n4431_);
  or g_12852 (new_n8549_, not_new_n645__968890104070, not_new_n8145__0);
  not g_12853 (not_new_n9550_, new_n9550_);
  not g_12854 (not_new_n611__5, new_n611_);
  not g_12855 (not_new_n602__19773267430, new_n602_);
  not g_12856 (new_n5924_, new_n5757_);
  not g_12857 (not_pi123, pi123);
  not g_12858 (not_new_n3282_, new_n3282_);
  or g_12859 (new_n6189_, not_new_n5869_, not_new_n5901__0);
  not g_12860 (not_new_n7328_, new_n7328_);
  and g_12861 (and_new_n2105__new_n2108_, new_n2105_, new_n2108_);
  not g_12862 (not_new_n622__168070, new_n622_);
  not g_12863 (not_new_n1601__3, new_n1601_);
  not g_12864 (not_new_n8596__3, new_n8596_);
  or g_12865 (new_n1017_, not_new_n3356_, not_new_n3355_);
  or g_12866 (new_n7864_, not_new_n7662_, not_new_n7663__0);
  and g_12867 (new_n8212_, new_n8343_, new_n8088_);
  not g_12868 (not_new_n4975__0, new_n4975_);
  not g_12869 (not_new_n6541_, new_n6541_);
  not g_12870 (not_new_n1819_, new_n1819_);
  or g_12871 (new_n7403_, not_new_n7401_, not_new_n7170__0);
  or g_12872 (po178, not_new_n3583_, not_new_n3582_);
  not g_12873 (not_new_n1045__47475615099430, new_n1045_);
  not g_12874 (not_new_n1611__24010, new_n1611_);
  or g_12875 (new_n9117_, not_new_n8973_, not_new_n9086_);
  not g_12876 (not_new_n1403_, new_n1403_);
  not g_12877 (new_n9350_, new_n632_);
  not g_12878 (not_new_n5039_, new_n5039_);
  or g_12879 (new_n8372_, not_new_n629__138412872010, not_new_n8133_);
  not g_12880 (new_n4158_, new_n4152_);
  and g_12881 (new_n3971_, and_and_not_pi048_2_not_pi047_2_not_pi050_2, not_pi049_2);
  not g_12882 (not_new_n8278__0, new_n8278_);
  not g_12883 (not_new_n5482__0, new_n5482_);
  not g_12884 (not_pi171_1, pi171);
  or g_12885 (new_n2745_, not_new_n631__2, not_new_n604__1);
  not g_12886 (not_new_n1919__0, new_n1919_);
  not g_12887 (not_new_n5427__0, new_n5427_);
  not g_12888 (not_pi169_3, pi169);
  not g_12889 (new_n9363_, new_n635_);
  not g_12890 (not_new_n6537_, new_n6537_);
  or g_12891 (new_n3768_, not_new_n3766_, not_new_n3767_);
  not g_12892 (not_new_n7443_, new_n7443_);
  not g_12893 (not_new_n1069__4, new_n1069_);
  not g_12894 (not_new_n4776__0, new_n4776_);
  not g_12895 (not_new_n9362_, new_n9362_);
  or g_12896 (new_n5403_, not_new_n4969_, not_new_n643__1176490);
  not g_12897 (not_new_n1576__8235430, new_n1576_);
  not g_12898 (new_n6792_, new_n6544_);
  not g_12899 (new_n1578_, new_n937_);
  or g_12900 (new_n6190_, not_new_n1067__490, not_new_n5783__0);
  not g_12901 (not_po296_21838143759917965991093122527538323430, po296);
  or g_12902 (new_n5410_, not_new_n4967_, not_new_n644__1176490);
  not g_12903 (not_new_n6634_, new_n6634_);
  and g_12904 (new_n1201_, new_n1694_, new_n1692_);
  and g_12905 (and_new_n1242__new_n1856_, new_n1242_, new_n1856_);
  not g_12906 (not_new_n5924_, new_n5924_);
  not g_12907 (not_new_n621__332329305696010, new_n621_);
  not g_12908 (not_new_n3510_, new_n3510_);
  not g_12909 (not_new_n1055_, new_n1055_);
  not g_12910 (not_new_n5111__0, new_n5111_);
  not g_12911 (not_new_n581__1176490, new_n581_);
  not g_12912 (not_new_n8446_, new_n8446_);
  or g_12913 (new_n8777_, not_new_n8718_, not_new_n8697_);
  not g_12914 (not_new_n5841_, new_n5841_);
  not g_12915 (not_new_n5479_, new_n5479_);
  or g_12916 (new_n9648_, not_new_n9475_, not_new_n9647_);
  not g_12917 (not_new_n3331_, new_n3331_);
  and g_12918 (new_n9502_, new_n9824_, new_n9825_);
  not g_12919 (not_new_n2946_, new_n2946_);
  not g_12920 (not_new_n5463_, new_n5463_);
  not g_12921 (new_n8618_, new_n1059_);
  not g_12922 (not_new_n6761__0, new_n6761_);
  or g_12923 (new_n6791_, not_new_n6729_, not_new_n6730_);
  or g_12924 (new_n8102_, not_new_n8265_, not_new_n8410_);
  not g_12925 (not_new_n4188_, new_n4188_);
  not g_12926 (not_new_n7110_, new_n7110_);
  and g_12927 (and_new_n933__new_n935_, new_n935_, new_n933_);
  not g_12928 (not_new_n617__3430, new_n617_);
  not g_12929 (not_new_n9616_, new_n9616_);
  not g_12930 (new_n8865_, new_n627_);
  not g_12931 (not_new_n3315__2326305139872070, new_n3315_);
  or g_12932 (new_n6437_, not_new_n6232__4, or_not_new_n6352__not_new_n6242__5);
  not g_12933 (not_new_n7703_, new_n7703_);
  or g_12934 (new_n2472_, not_new_n603__968890104070, not_new_n622__1);
  and g_12935 (new_n7077_, new_n6960_, new_n7200_);
  not g_12936 (not_new_n4898__1, new_n4898_);
  not g_12937 (not_new_n4468__0, new_n4468_);
  not g_12938 (not_new_n1253_, new_n1253_);
  not g_12939 (not_new_n4843__1, new_n4843_);
  not g_12940 (not_new_n1205_, new_n1205_);
  or g_12941 (new_n10150_, not_new_n10015_, not_new_n10149_);
  and g_12942 (new_n1256_, and_and_new_n1915__new_n1918__new_n1916_, new_n1917_);
  or g_12943 (or_not_new_n2727__not_new_n2730_, not_new_n2730_, not_new_n2727_);
  not g_12944 (not_new_n8801_, new_n8801_);
  not g_12945 (not_new_n7304_, new_n7304_);
  or g_12946 (new_n6135_, not_new_n5858_, not_new_n5887__0);
  not g_12947 (not_new_n10127_, new_n10127_);
  and g_12948 (new_n5871_, new_n6028_, new_n5717_);
  not g_12949 (not_pi162_0, pi162);
  not g_12950 (not_po296_332329305696010, po296);
  or g_12951 (new_n9609_, not_new_n9403_, not_new_n9402_);
  or g_12952 (new_n10233_, not_new_n10232_, not_new_n10000_);
  or g_12953 (new_n1739_, not_new_n1728__7, not_pi083);
  not g_12954 (new_n4093_, pi249);
  not g_12955 (not_pi167_1, pi167);
  or g_12956 (new_n4335_, not_new_n4337__0, not_new_n4293_);
  not g_12957 (new_n7604_, new_n632_);
  not g_12958 (new_n7647_, new_n1057_);
  not g_12959 (new_n8615_, new_n1176_);
  not g_12960 (not_new_n2885_, new_n2885_);
  not g_12961 (not_new_n5354_, new_n5354_);
  not g_12962 (not_new_n7628__0, new_n7628_);
  not g_12963 (not_new_n4739_, new_n4739_);
  or g_12964 (new_n1953_, not_new_n9955_, not_new_n594__8);
  or g_12965 (or_not_new_n2776__not_new_n2779_, not_new_n2779_, not_new_n2776_);
  not g_12966 (new_n4754_, new_n1605_);
  not g_12967 (new_n4934_, new_n1045_);
  not g_12968 (not_new_n1041__1176490, new_n1041_);
  not g_12969 (not_new_n7261_, new_n7261_);
  or g_12970 (new_n6768_, not_new_n638__968890104070, not_new_n6519__1);
  or g_12971 (new_n5976_, not_new_n5790_, not_new_n636__1176490);
  not g_12972 (not_new_n10006_, new_n10006_);
  and g_12973 (new_n1310_, new_n2177_, new_n2176_);
  not g_12974 (not_new_n2033__0, new_n2033_);
  not g_12975 (not_new_n4582_, new_n4582_);
  not g_12976 (not_new_n9852_, new_n9852_);
  not g_12977 (not_new_n6595_, new_n6595_);
  not g_12978 (new_n4802_, new_n1059_);
  not g_12979 (not_new_n8127_, new_n8127_);
  not g_12980 (not_new_n588__0, new_n588_);
  not g_12981 (not_new_n740__1, new_n740_);
  not g_12982 (not_new_n4393_, new_n4393_);
  xor g_12983 (key_gate_105, key_105, not_new_n1675_);
  xor g_12984 (key_gate_20, not_new_n3924_, key_20);
  and g_12985 (and_and_not_pi060_1_not_pi059_1_not_pi058_1, not_pi058_1, and_not_pi060_1_not_pi059_1);
  not g_12986 (not_new_n589__445676403263631959001900459745680070, new_n589_);
  not g_12987 (not_new_n589__490, new_n589_);
  and g_12988 (new_n4503_, new_n4695_, new_n4696_);
  not g_12989 (not_new_n7818_, new_n7818_);
  not g_12990 (not_new_n9944_, new_n9944_);
  not g_12991 (not_new_n3867_, new_n3867_);
  or g_12992 (new_n7037_, not_new_n7440_, not_new_n7441_);
  not g_12993 (not_new_n3190_, new_n3190_);
  not g_12994 (not_new_n6691__0, new_n6691_);
  not g_12995 (not_new_n5381_, new_n5381_);
  or g_12996 (or_or_not_new_n6239__not_new_n6350__not_new_n6232__3, not_new_n6232__3, or_not_new_n6239__not_new_n6350_);
  or g_12997 (new_n8918_, not_new_n9302_, not_new_n9301_);
  or g_12998 (new_n9058_, not_new_n8807_, not_new_n8978_);
  not g_12999 (not_new_n1043__19773267430, new_n1043_);
  not g_13000 (not_new_n3577_, new_n3577_);
  or g_13001 (or_or_not_new_n2865__not_new_n2868__not_new_n2867_, or_not_new_n2865__not_new_n2868_, not_new_n2867_);
  not g_13002 (not_new_n3934__0, new_n3934_);
  not g_13003 (not_new_n7420_, new_n7420_);
  not g_13004 (not_new_n8549_, new_n8549_);
  and g_13005 (po089, key_gate_101, pi068);
  not g_13006 (not_new_n6160_, new_n6160_);
  not g_13007 (not_new_n3372__7, new_n3372_);
  not g_13008 (not_new_n9215_, new_n9215_);
  not g_13009 (not_new_n600__168070, new_n600_);
  not g_13010 (not_new_n9788_, new_n9788_);
  not g_13011 (not_new_n1027__1, new_n1027_);
  not g_13012 (not_new_n1600__8, new_n1600_);
  not g_13013 (not_new_n9926_, new_n9926_);
  not g_13014 (not_new_n4829__1, new_n4829_);
  and g_13015 (new_n1443_, and_new_n2642__new_n2641_, new_n2640_);
  or g_13016 (new_n3124_, not_new_n581__3788186922656647816827176259430, not_new_n622__6);
  or g_13017 (new_n6797_, not_new_n6542_, not_new_n6742_);
  not g_13018 (not_new_n8579_, new_n8579_);
  not g_13019 (not_new_n596__5, key_gate_88);
  or g_13020 (new_n8444_, not_new_n8085_, not_new_n8244__0);
  and g_13021 (new_n6348_, and_new_n6373__new_n6398_, new_n6276_);
  and g_13022 (new_n1212_, new_n1725_, new_n1727_);
  not g_13023 (not_new_n587__490, new_n587_);
  not g_13024 (not_new_n1603__1, new_n1603_);
  or g_13025 (new_n6001_, not_new_n6000_, not_new_n5719_);
  and g_13026 (new_n6962_, new_n7208_, new_n7207_);
  not g_13027 (not_new_n642__24010, new_n642_);
  or g_13028 (new_n3413_, not_new_n1009__1, not_new_n1594__1);
  or g_13029 (new_n3864_, not_new_n640__490, not_new_n1576__8235430);
  not g_13030 (not_new_n621__797922662976120010, new_n621_);
  or g_13031 (new_n3525_, not_new_n1613__797922662976120010, not_new_n2348_);
  not g_13032 (not_new_n1055__19773267430, new_n1055_);
  not g_13033 (not_new_n7031__1, new_n7031_);
  and g_13034 (and_new_n1298__new_n2122_, new_n1298_, new_n2122_);
  not g_13035 (not_new_n7267_, new_n7267_);
  not g_13036 (not_new_n4432_, new_n4432_);
  not g_13037 (not_new_n6414_, new_n6414_);
  not g_13038 (new_n8423_, new_n8175_);
  not g_13039 (not_new_n626__4, new_n626_);
  or g_13040 (new_n4354_, not_new_n4300_, not_new_n4347_);
  not g_13041 (not_new_n3315__138412872010, new_n3315_);
  not g_13042 (not_new_n8936_, new_n8936_);
  not g_13043 (not_new_n1611_, new_n1611_);
  and g_13044 (new_n9974_, new_n10041_, new_n9975_);
  or g_13045 (new_n2818_, not_new_n4113__1, not_new_n994__70);
  or g_13046 (or_not_new_n1024__2_not_new_n1028__3, not_new_n1028__3, not_new_n1024__2);
  or g_13047 (new_n7882_, not_new_n7721_, not_new_n7880_);
  not g_13048 (not_new_n9403__0, new_n9403_);
  not g_13049 (new_n4843_, new_n4747_);
  not g_13050 (not_new_n749_, new_n749_);
  and g_13051 (new_n9345_, new_n9640_, new_n9643_);
  or g_13052 (new_n4694_, not_new_n4692_, not_new_n4557_);
  not g_13053 (not_new_n7872_, new_n7872_);
  or g_13054 (new_n7054_, not_new_n7465_, not_new_n7464_);
  not g_13055 (not_new_n6839_, new_n6839_);
  or g_13056 (new_n5896_, not_new_n6059_, not_new_n6052_);
  or g_13057 (new_n8462_, not_new_n8313_, not_new_n8243_);
  not g_13058 (not_new_n9800_, new_n9800_);
  not g_13059 (not_new_n6181_, new_n6181_);
  or g_13060 (new_n3799_, not_new_n1886_, not_new_n3439_);
  or g_13061 (new_n10289_, not_new_n9942_, not_new_n1598__113988951853731430);
  not g_13062 (not_new_n5820_, new_n5820_);
  not g_13063 (not_new_n6982__2, new_n6982_);
  or g_13064 (new_n10227_, not_new_n9987_, not_new_n9900__1);
  not g_13065 (not_new_n4203_, new_n4203_);
  or g_13066 (new_n6955_, not_new_n6953_, not_new_n6954_);
  not g_13067 (not_new_n6020_, new_n6020_);
  not g_13068 (not_new_n1027__403536070, new_n1027_);
  not g_13069 (not_new_n2982_, new_n2982_);
  not g_13070 (not_new_n2593_, new_n2593_);
  not g_13071 (not_new_n9198_, new_n9198_);
  not g_13072 (not_new_n10200_, new_n10200_);
  not g_13073 (not_new_n2858_, new_n2858_);
  not g_13074 (not_new_n6588_, new_n6588_);
  not g_13075 (not_new_n7234_, new_n7234_);
  not g_13076 (not_new_n623__4, new_n623_);
  not g_13077 (not_new_n1009__2, new_n1009_);
  not g_13078 (not_new_n619__490, new_n619_);
  not g_13079 (not_new_n6373__2, new_n6373_);
  or g_13080 (new_n6050_, not_new_n5987_, not_new_n5989_);
  not g_13081 (not_new_n586__24010, new_n586_);
  not g_13082 (not_po296_3430, po296);
  not g_13083 (new_n4765_, new_n1597_);
  not g_13084 (not_new_n6974__968890104070, new_n6974_);
  and g_13085 (new_n1285_, new_n2060_, new_n2061_);
  not g_13086 (not_new_n605__168070, new_n605_);
  not g_13087 (not_new_n617__93874803376477543056490, new_n617_);
  or g_13088 (po193, or_not_new_n1550__not_new_n1370_, not_new_n1369_);
  not g_13089 (not_new_n8281_, new_n8281_);
  not g_13090 (not_new_n591__9, new_n591_);
  not g_13091 (not_new_n3706_, new_n3706_);
  not g_13092 (not_new_n6636__0, new_n6636_);
  or g_13093 (new_n3026_, not_new_n1027__168070, not_new_n1161_);
  or g_13094 (new_n10311_, not_new_n10310_, not_new_n10309_);
  not g_13095 (not_new_n4620_, new_n4620_);
  not g_13096 (not_new_n1005_, new_n1005_);
  or g_13097 (new_n2959_, not_pi271, not_po296_597682638941559493067901192655856192170251494124306816490);
  or g_13098 (new_n4202_, not_new_n4169__0, not_new_n4101_);
  not g_13099 (not_new_n1520_, new_n1520_);
  and g_13100 (new_n5048_, new_n5375_, and_new_n4974__new_n5376_);
  or g_13101 (new_n9705_, not_new_n9703_, not_new_n9592_);
  or g_13102 (new_n2727_, not_new_n3311_, not_new_n1063__1);
  not g_13103 (not_new_n9875_, new_n9875_);
  not g_13104 (not_new_n10193_, new_n10193_);
  or g_13105 (new_n7245_, not_new_n7445_, not_new_n7008_);
  or g_13106 (new_n3641_, not_new_n974_, not_new_n1611__6782230728490);
  not g_13107 (not_new_n1589__8, new_n1589_);
  not g_13108 (not_new_n645__4, new_n645_);
  or g_13109 (new_n2298_, not_new_n1597_, not_new_n1588__2326305139872070);
  not g_13110 (not_new_n9685_, new_n9685_);
  not g_13111 (not_new_n619__24010, new_n619_);
  or g_13112 (new_n5007_, not_new_n5320_, not_new_n5319_);
  and g_13113 (new_n5514_, new_n5691_, new_n5692_);
  and g_13114 (new_n8227_, new_n8368_, new_n8092_);
  not g_13115 (not_new_n6508__0, new_n6508_);
  and g_13116 (new_n9457_, new_n9328_, new_n9547_);
  or g_13117 (new_n5324_, not_new_n5058_, not_new_n1607__5);
  not g_13118 (new_n1602_, new_n967_);
  not g_13119 (not_new_n647__1176490, new_n647_);
  not g_13120 (not_new_n6150_, new_n6150_);
  or g_13121 (new_n4946_, not_new_n5126_, not_new_n5030_);
  not g_13122 (not_new_n3535_, new_n3535_);
  not g_13123 (not_new_n1581__403536070, new_n1581_);
  not g_13124 (new_n5085_, new_n4966_);
  not g_13125 (not_pi035_1, pi035);
  not g_13126 (new_n7777_, new_n7614_);
  or g_13127 (new_n9810_, not_new_n9426__1, not_new_n9689_);
  not g_13128 (new_n9362_, new_n1045_);
  or g_13129 (new_n3222_, not_new_n1069__4, not_new_n3185__8235430);
  not g_13130 (not_new_n3860_, new_n3860_);
  not g_13131 (not_new_n2801_, new_n2801_);
  not g_13132 (not_new_n4416__0, new_n4416_);
  not g_13133 (not_new_n1596__57648010, new_n1596_);
  not g_13134 (not_new_n634__5, new_n634_);
  not g_13135 (not_new_n4092_, new_n4092_);
  not g_13136 (not_new_n8507_, new_n8507_);
  not g_13137 (new_n9921_, new_n626_);
  not g_13138 (not_new_n8455_, new_n8455_);
  not g_13139 (not_pi160_0, pi160);
  or g_13140 (new_n9442_, not_new_n9797_, not_new_n9796_);
  not g_13141 (not_new_n4528_, new_n4528_);
  not g_13142 (not_new_n618__16284135979104490, new_n618_);
  not g_13143 (not_new_n10062_, new_n10062_);
  or g_13144 (new_n6695_, not_new_n6655__0, not_new_n6495_);
  not g_13145 (not_new_n6035_, new_n6035_);
  not g_13146 (not_new_n6946_, new_n6946_);
  not g_13147 (not_new_n5774__0, new_n5774_);
  not g_13148 (not_new_n3955_, new_n3955_);
  or g_13149 (new_n8535_, not_new_n639__6782230728490, not_new_n8140__0);
  xnor g_13150 (key_gate_18, new_n1705_, key_18);
  or g_13151 (new_n3585_, not_new_n1612__16284135979104490, not_new_n2338__0);
  not g_13152 (not_new_n635__4, new_n635_);
  or g_13153 (new_n2525_, not_new_n5485_, not_new_n605__1);
  not g_13154 (not_new_n742__1, new_n742_);
  not g_13155 (not_new_n1580__490, new_n1580_);
  not g_13156 (not_new_n6140_, new_n6140_);
  not g_13157 (new_n7008_, new_n723_);
  not g_13158 (not_new_n647__47475615099430, new_n647_);
  not g_13159 (not_new_n4753_, new_n4753_);
  or g_13160 (new_n2887_, not_po296_103677930763188441902487387275962551382129494864490, not_pi263_0);
  not g_13161 (not_new_n4716_, new_n4716_);
  not g_13162 (not_pi119_0, pi119);
  not g_13163 (not_new_n7363_, new_n7363_);
  not g_13164 (new_n6258_, new_n1600_);
  or g_13165 (new_n7155_, or_not_new_n7311__not_new_n7203_, not_new_n7157_);
  not g_13166 (new_n6478_, new_n1047_);
  not g_13167 (not_new_n5478_, new_n5478_);
  not g_13168 (not_new_n8047_, new_n8047_);
  not g_13169 (not_new_n9242_, new_n9242_);
  not g_13170 (not_new_n644_, new_n644_);
  not g_13171 (not_new_n8256__0, new_n8256_);
  and g_13172 (new_n3977_, new_n4050_, new_n4049_);
  not g_13173 (not_new_n7718_, new_n7718_);
  not g_13174 (not_pi108, pi108);
  or g_13175 (new_n2543_, not_new_n4464_, not_new_n609__3);
  or g_13176 (new_n4878_, not_new_n4742_, not_new_n1071__7);
  or g_13177 (new_n9081_, not_new_n8874_, not_new_n8875_);
  or g_13178 (or_not_new_n1958__not_new_n1959_, not_new_n1958_, not_new_n1959_);
  or g_13179 (new_n1649_, not_new_n1631__4, not_pi038);
  not g_13180 (not_new_n2171_, new_n2171_);
  or g_13181 (new_n667_, not_new_n3162_, or_not_new_n3164__not_new_n3163_);
  not g_13182 (not_new_n634__2824752490, new_n634_);
  not g_13183 (not_new_n7435_, new_n7435_);
  or g_13184 (new_n1617_, not_pi275_2, not_new_n996_);
  not g_13185 (new_n1895_, new_n949_);
  not g_13186 (not_new_n8787_, new_n8787_);
  not g_13187 (new_n4569_, new_n4496_);
  not g_13188 (new_n4537_, new_n4475_);
  or g_13189 (new_n5075_, not_new_n4971_, not_new_n5273_);
  or g_13190 (or_not_new_n1570__not_new_n2502_, not_new_n2502_, not_new_n1570_);
  or g_13191 (new_n4865_, not_new_n4770__1, not_new_n4839__1);
  or g_13192 (new_n8320_, not_new_n8287__0, not_new_n8104__1);
  not g_13193 (not_new_n9600_, new_n9600_);
  or g_13194 (new_n1897_, not_new_n593__5, not_new_n634_);
  not g_13195 (not_new_n4135__1, new_n4135_);
  and g_13196 (new_n7758_, new_n8056_, new_n8055_);
  not g_13197 (new_n3424_, new_n1041_);
  not g_13198 (not_new_n4771_, new_n4771_);
  not g_13199 (not_new_n9401_, new_n9401_);
  and g_13200 (new_n1363_, and_new_n2394__new_n2393_, new_n2392_);
  or g_13201 (new_n9141_, new_n1057_, new_n636_);
  or g_13202 (new_n7241_, not_new_n7436__0, not_new_n7007__0);
  not g_13203 (not_new_n1583__0, new_n1583_);
  not g_13204 (not_new_n3315__5, new_n3315_);
  not g_13205 (not_new_n5186__0, new_n5186_);
  or g_13206 (new_n3050_, not_new_n1071__2, not_new_n581__2824752490);
  not g_13207 (not_new_n7658__0, new_n7658_);
  not g_13208 (not_new_n5686__1, new_n5686_);
  not g_13209 (new_n5533_, new_n5440_);
  or g_13210 (new_n6654_, not_new_n1037__24010, not_new_n6480_);
  or g_13211 (new_n10333_, not_new_n9916__0, not_new_n633__39098210485829880490);
  not g_13212 (not_new_n8994_, new_n8994_);
  or g_13213 (new_n2903_, not_new_n1616__8235430, not_new_n2900_);
  not g_13214 (not_new_n6373__7, new_n6373_);
  not g_13215 (not_new_n4161_, new_n4161_);
  not g_13216 (not_new_n8976_, new_n8976_);
  not g_13217 (new_n7651_, new_n1053_);
  not g_13218 (not_new_n9147_, new_n9147_);
  not g_13219 (not_new_n2911_, new_n2911_);
  not g_13220 (not_new_n3829_, new_n3829_);
  not g_13221 (not_new_n5295_, new_n5295_);
  not g_13222 (not_new_n4988__0, new_n4988_);
  or g_13223 (new_n9076_, new_n645_, new_n1071_);
  not g_13224 (not_new_n4444__0, new_n4444_);
  and g_13225 (new_n6618_, new_n6858_, new_n6857_);
  not g_13226 (not_new_n622__5, new_n622_);
  not g_13227 (not_new_n595__968890104070, new_n595_);
  not g_13228 (not_new_n638__332329305696010, new_n638_);
  not g_13229 (not_new_n626__797922662976120010, new_n626_);
  not g_13230 (new_n4490_, new_n1028_);
  not g_13231 (not_new_n630__10, new_n630_);
  not g_13232 (not_new_n3184__24010, new_n3184_);
  or g_13233 (new_n6830_, not_new_n6613__3, not_new_n6684_);
  not g_13234 (not_pi142_2, pi142);
  not g_13235 (not_new_n5188_, new_n5188_);
  not g_13236 (not_new_n4757_, new_n4757_);
  not g_13237 (not_new_n620__4, new_n620_);
  or g_13238 (new_n2189_, not_new_n4124_, not_new_n585__138412872010);
  and g_13239 (new_n4909_, new_n5161_, new_n4907_);
  or g_13240 (new_n1818_, not_new_n4918_, not_new_n1589__1);
  not g_13241 (not_new_n633__113988951853731430, new_n633_);
  or g_13242 (new_n2134_, not_new_n601__8235430, not_new_n646__0);
  or g_13243 (new_n10164_, not_new_n10024_, not_new_n10128_);
  or g_13244 (or_not_new_n3170__not_new_n3169_, not_new_n3170_, not_new_n3169_);
  not g_13245 (not_new_n9361__0, new_n9361_);
  not g_13246 (not_new_n9951__0, new_n9951_);
  not g_13247 (not_new_n1728__332329305696010, new_n1728_);
  not g_13248 (not_new_n7069_, new_n7069_);
  not g_13249 (not_new_n8147_, new_n8147_);
  not g_13250 (not_new_n1595_, new_n1595_);
  not g_13251 (not_new_n2624_, new_n2624_);
  not g_13252 (new_n6985_, new_n744_);
  or g_13253 (new_n5318_, not_new_n5317_, not_new_n5316_);
  not g_13254 (not_po296_7, po296);
  not g_13255 (not_new_n7204_, new_n7204_);
  not g_13256 (not_new_n1583__168070, new_n1583_);
  and g_13257 (new_n8970_, new_n9271_, new_n9270_);
  not g_13258 (not_new_n7653_, new_n7653_);
  and g_13259 (and_and_new_n2143__new_n2146__new_n2144_, new_n2144_, and_new_n2143__new_n2146_);
  or g_13260 (new_n2265_, not_new_n585__332329305696010, not_new_n4120_);
  not g_13261 (not_new_n8702_, new_n8702_);
  or g_13262 (new_n5397_, not_new_n1063__9, not_new_n4958_);
  not g_13263 (not_new_n775__490, new_n775_);
  or g_13264 (new_n9625_, new_n1599_, new_n622_);
  or g_13265 (new_n10318_, not_new_n10316_, not_new_n10317_);
  or g_13266 (new_n2115_, not_new_n601__1176490, not_new_n633__0);
  not g_13267 (not_new_n7153__0, new_n7153_);
  not g_13268 (not_new_n3973_, new_n3973_);
  not g_13269 (not_new_n989_, new_n989_);
  not g_13270 (not_new_n1580__9, new_n1580_);
  not g_13271 (not_new_n593__3430, new_n593_);
  not g_13272 (not_new_n6373__0, new_n6373_);
  not g_13273 (not_new_n618__273687473400809163430, new_n618_);
  not g_13274 (new_n5759_, new_n1051_);
  not g_13275 (not_new_n2034_, new_n2034_);
  or g_13276 (new_n7739_, not_new_n7941_, not_new_n7696_);
  not g_13277 (not_new_n5441_, new_n5441_);
  or g_13278 (new_n2353_, not_pi255_0, not_new_n600_);
  not g_13279 (not_new_n960_, new_n960_);
  not g_13280 (not_new_n4451__0, new_n4451_);
  not g_13281 (not_new_n3315__10, new_n3315_);
  or g_13282 (new_n3018_, not_new_n1607__1, not_new_n581__9);
  not g_13283 (not_new_n603__2, new_n603_);
  not g_13284 (not_new_n2306_, new_n2306_);
  or g_13285 (new_n2942_, not_new_n647__3, not_new_n604__138412872010);
  and g_13286 (new_n3917_, new_n4045_, new_n3941_);
  not g_13287 (new_n9896_, new_n648_);
  not g_13288 (not_new_n5956__0, new_n5956_);
  not g_13289 (not_new_n9716_, new_n9716_);
  or g_13290 (new_n8496_, not_new_n8494_, not_new_n8495_);
  or g_13291 (new_n4328_, not_new_n4290_, not_new_n4330__0);
  not g_13292 (new_n6254_, new_n632_);
  and g_13293 (new_n6590_, new_n6462_, new_n6751_);
  not g_13294 (not_new_n8506_, new_n8506_);
  or g_13295 (new_n2592_, not_pi201, not_new_n2509__7);
  not g_13296 (not_new_n1588__3, new_n1588_);
  xor g_13297 (key_gate_83, new_n1720_, key_83);
  not g_13298 (not_new_n2344_, new_n2344_);
  or g_13299 (new_n6528_, not_new_n6492_, not_new_n647__57648010);
  not g_13300 (not_new_n8172_, new_n8172_);
  or g_13301 (new_n3364_, not_new_n1534__968890104070, not_pi061_0);
  and g_13302 (and_new_n1839__new_n1842_, new_n1839_, new_n1842_);
  not g_13303 (not_pi037_3, pi037);
  and g_13304 (new_n1544_, new_n3601_, new_n3600_);
  or g_13305 (new_n8442_, not_new_n8244_, not_new_n8314__0);
  not g_13306 (new_n7809_, new_n7619_);
  not g_13307 (not_new_n6611_, new_n6611_);
  not g_13308 (not_new_n4818__1, new_n4818_);
  not g_13309 (not_new_n7809__0, new_n7809_);
  or g_13310 (new_n9243_, not_new_n9102_, not_new_n9241_);
  not g_13311 (not_new_n637__70, new_n637_);
  not g_13312 (new_n8621_, new_n1602_);
  not g_13313 (not_new_n6499_, new_n6499_);
  not g_13314 (not_pi017_0, pi017);
  not g_13315 (not_new_n1063__47475615099430, new_n1063_);
  not g_13316 (not_new_n617__3, new_n617_);
  not g_13317 (not_pi255, pi255);
  not g_13318 (not_new_n3450_, new_n3450_);
  not g_13319 (not_new_n642__8235430, new_n642_);
  not g_13320 (not_new_n2958_, new_n2958_);
  not g_13321 (not_new_n9284_, new_n9284_);
  not g_13322 (not_new_n6475__1, new_n6475_);
  not g_13323 (not_new_n6685_, new_n6685_);
  not g_13324 (not_new_n6474_, new_n6474_);
  not g_13325 (not_new_n7321__0, new_n7321_);
  or g_13326 (new_n706_, not_new_n1490_, not_new_n3000_);
  not g_13327 (new_n5994_, new_n5780_);
  not g_13328 (not_new_n4718__0, new_n4718_);
  not g_13329 (not_new_n3215_, new_n3215_);
  or g_13330 (new_n8177_, not_new_n8165_, not_new_n8391_);
  not g_13331 (not_new_n1597__8, new_n1597_);
  not g_13332 (not_new_n6053_, new_n6053_);
  not g_13333 (not_new_n1962_, new_n1962_);
  not g_13334 (not_new_n7528_, new_n7528_);
  not g_13335 (new_n9028_, new_n8846_);
  not g_13336 (not_new_n7692_, new_n7692_);
  not g_13337 (not_new_n7900_, new_n7900_);
  or g_13338 (new_n8469_, not_new_n8109__0, not_new_n634__6782230728490);
  not g_13339 (not_new_n5005_, new_n5005_);
  not g_13340 (not_new_n5137_, new_n5137_);
  or g_13341 (new_n2432_, not_new_n603__168070, not_new_n633__1);
  not g_13342 (not_new_n7010_, new_n7010_);
  not g_13343 (not_new_n9226_, new_n9226_);
  not g_13344 (not_pi153_0, pi153);
  not g_13345 (not_new_n646__0, new_n646_);
  not g_13346 (not_new_n4264_, new_n4264_);
  not g_13347 (not_new_n6546__0, new_n6546_);
  not g_13348 (not_new_n7667_, new_n7667_);
  or g_13349 (new_n9957_, not_new_n10252_, not_new_n10251_);
  not g_13350 (not_new_n5050_, new_n5050_);
  or g_13351 (new_n8375_, not_new_n8170_, not_new_n1597__2824752490);
  or g_13352 (new_n5478_, not_new_n5607_, not_new_n5608_);
  not g_13353 (not_new_n632__5585458640832840070, new_n632_);
  not g_13354 (not_new_n1585__3, new_n1585_);
  not g_13355 (not_new_n9062_, new_n9062_);
  and g_13356 (new_n1215_, new_n1777_, new_n1779_);
  not g_13357 (not_new_n2799_, new_n2799_);
  or g_13358 (new_n5681_, not_pi143_3, not_new_n5462__1);
  not g_13359 (not_new_n7439__2, new_n7439_);
  or g_13360 (new_n7943_, not_new_n7772__0, not_new_n7620__0);
  or g_13361 (new_n8828_, not_new_n624__6782230728490, not_new_n1041__2824752490);
  not g_13362 (not_new_n1051__2824752490, new_n1051_);
  not g_13363 (not_new_n1611__8235430, new_n1611_);
  or g_13364 (new_n3709_, not_new_n617__9, not_po298_2326305139872070);
  not g_13365 (not_new_n5674__0, new_n5674_);
  not g_13366 (not_new_n1597__47475615099430, new_n1597_);
  or g_13367 (new_n7303_, not_new_n7275_, not_new_n7161_);
  not g_13368 (not_new_n4535_, new_n4535_);
  or g_13369 (new_n1936_, not_new_n591__8, not_new_n4753_);
  not g_13370 (not_new_n635__24010, new_n635_);
  or g_13371 (new_n7042_, not_new_n7455_, not_new_n7456_);
  or g_13372 (new_n723_, not_new_n3271_, not_new_n3272_);
  or g_13373 (new_n4866_, not_new_n4773_, not_new_n1600__7);
  not g_13374 (not_new_n1035__168070, new_n1035_);
  or g_13375 (new_n4984_, not_new_n637__3430, not_new_n1065__8);
  not g_13376 (not_new_n8745_, new_n8745_);
  not g_13377 (not_pi053_3, pi053);
  not g_13378 (not_new_n1584__403536070, new_n1584_);
  not g_13379 (not_new_n7269_, new_n7269_);
  not g_13380 (not_pi129_2, pi129);
  not g_13381 (not_new_n9508_, new_n9508_);
  or g_13382 (new_n4225_, not_pi270_2, not_new_n4080_);
  not g_13383 (not_new_n10224_, new_n10224_);
  not g_13384 (not_new_n7556_, new_n7556_);
  or g_13385 (new_n6780_, not_new_n642__57648010, not_new_n6633__0);
  or g_13386 (new_n2031_, not_new_n591__3430, not_new_n4803_);
  and g_13387 (new_n9865_, new_n10128_, new_n9861_);
  not g_13388 (not_new_n1583__1176490, new_n1583_);
  not g_13389 (not_new_n5476_, new_n5476_);
  not g_13390 (not_new_n7607__0, new_n7607_);
  not g_13391 (not_new_n4475_, new_n4475_);
  and g_13392 (and_and_and_new_n1463__new_n1465__new_n1464__new_n3720_, and_and_new_n1463__new_n1465__new_n1464_, new_n3720_);
  or g_13393 (po297, not_pi275, not_new_n1629_);
  or g_13394 (new_n9657_, new_n642_, new_n1035_);
  or g_13395 (new_n3560_, not_pi146_0, not_new_n1538__1176490);
  not g_13396 (new_n9360_, new_n641_);
  or g_13397 (new_n7863_, not_new_n7711_, not_new_n7666_);
  not g_13398 (not_new_n747_, new_n747_);
  not g_13399 (not_new_n603__5, new_n603_);
  not g_13400 (not_new_n775__968890104070, new_n775_);
  not g_13401 (not_new_n723__1, new_n723_);
  not g_13402 (not_new_n2783_, new_n2783_);
  not g_13403 (not_new_n1053__1, new_n1053_);
  not g_13404 (not_new_n7101_, new_n7101_);
  not g_13405 (not_new_n9298_, new_n9298_);
  not g_13406 (not_new_n4569_, new_n4569_);
  not g_13407 (not_new_n643__3430, new_n643_);
  not g_13408 (not_new_n1149__0, new_n1149_);
  not g_13409 (new_n7007_, new_n724_);
  not g_13410 (not_new_n8963_, new_n8963_);
  and g_13411 (and_and_new_n1972__new_n1975__new_n1973_, and_new_n1972__new_n1975_, new_n1973_);
  or g_13412 (new_n7195_, not_new_n6976__1, not_new_n7366__1);
  and g_13413 (new_n1408_, new_n930_, new_n931_);
  or g_13414 (new_n10108_, new_n1063_, new_n638_);
  not g_13415 (not_new_n4922_, new_n4922_);
  not g_13416 (not_new_n4132__0, new_n4132_);
  and g_13417 (new_n8261_, new_n8535_, new_n8534_);
  not g_13418 (not_new_n1601__2, new_n1601_);
  not g_13419 (not_new_n6159_, new_n6159_);
  not g_13420 (not_new_n621__1176490, new_n621_);
  not g_13421 (not_new_n9394_, new_n9394_);
  not g_13422 (not_new_n10041_, new_n10041_);
  not g_13423 (new_n8128_, new_n1598_);
  or g_13424 (new_n5417_, not_new_n627__168070, not_new_n4964_);
  or g_13425 (or_not_new_n3097__not_new_n3096_, not_new_n3097_, not_new_n3096_);
  not g_13426 (not_new_n1585__9, new_n1585_);
  or g_13427 (new_n10070_, not_new_n10045_, not_new_n9855_);
  or g_13428 (new_n9828_, not_new_n9826_, not_new_n9827_);
  not g_13429 (not_pi140_1, pi140);
  not g_13430 (not_new_n8595__6, new_n8595_);
  not g_13431 (not_pi174_1, pi174);
  not g_13432 (not_new_n610__2, new_n610_);
  not g_13433 (not_new_n1011__5, new_n1011_);
  not g_13434 (not_new_n4526_, new_n4526_);
  not g_13435 (new_n4980_, new_n639_);
  not g_13436 (not_new_n8822_, new_n8822_);
  or g_13437 (new_n4481_, not_new_n4524_, not_new_n4523_);
  and g_13438 (new_n1348_, and_new_n1539__new_n2356_, new_n2355_);
  not g_13439 (not_new_n7436__1, new_n7436_);
  or g_13440 (or_not_new_n929__not_new_n931_, not_new_n931_, not_new_n929_);
  or g_13441 (new_n10116_, not_new_n10113_, not_new_n1067__47475615099430);
  not g_13442 (not_new_n5601_, new_n5601_);
  or g_13443 (new_n643_, or_or_not_new_n2015__not_new_n2016__not_new_n2018_, not_new_n2017_);
  not g_13444 (not_new_n8946_, new_n8946_);
  not g_13445 (not_new_n7330_, new_n7330_);
  not g_13446 (not_new_n8963__0, new_n8963_);
  not g_13447 (not_new_n5465__0, new_n5465_);
  not g_13448 (not_new_n1031__7, new_n1031_);
  or g_13449 (or_not_new_n6363__not_new_n6358_, not_new_n6363_, not_new_n6358_);
  not g_13450 (not_new_n7034__1, new_n7034_);
  and g_13451 (new_n8241_, new_n8078_, new_n8406_);
  or g_13452 (new_n9449_, not_new_n9848_, not_new_n9849_);
  or g_13453 (new_n4189_, not_new_n4148_, not_pi267_0);
  or g_13454 (new_n5699_, not_pi140_2, not_new_n5456_);
  and g_13455 (po115, key_gate_101, pi094);
  not g_13456 (not_new_n615_, new_n615_);
  not g_13457 (not_new_n3551_, new_n3551_);
  not g_13458 (new_n6676_, new_n6491_);
  and g_13459 (new_n1339_, new_n2311_, and_new_n1338__new_n2312_);
  not g_13460 (not_new_n5074_, new_n5074_);
  not g_13461 (not_new_n4496_, new_n4496_);
  or g_13462 (new_n2087_, not_new_n633_, not_new_n593__168070);
  not g_13463 (new_n8864_, new_n1055_);
  not g_13464 (new_n8647_, new_n1601_);
  not g_13465 (not_new_n1312_, new_n1312_);
  not g_13466 (not_new_n6772_, new_n6772_);
  or g_13467 (new_n3716_, not_new_n989__797922662976120010, not_pi244);
  not g_13468 (not_pi061_0, pi061);
  not g_13469 (not_new_n1581__24010, new_n1581_);
  and g_13470 (and_new_n7597__new_n7953_, new_n7597_, new_n7953_);
  not g_13471 (not_new_n581__47475615099430, new_n581_);
  not g_13472 (not_new_n740__0, new_n740_);
  not g_13473 (not_new_n2187_, new_n2187_);
  not g_13474 (not_pi169_1, pi169);
  not g_13475 (not_new_n8713_, new_n8713_);
  or g_13476 (new_n6161_, not_new_n6018_, or_not_new_n5917__not_new_n5719__0);
  xnor g_13477 (key_gate_115, key_115, new_n1666_);
  or g_13478 (new_n9129_, new_n642_, new_n1035_);
  or g_13479 (new_n5120_, not_new_n5029_, not_new_n5118_);
  or g_13480 (or_not_new_n2034__not_new_n2035_, not_new_n2035_, not_new_n2034_);
  not g_13481 (not_new_n1027__3430, new_n1027_);
  not g_13482 (not_new_n618__0, new_n618_);
  not g_13483 (not_new_n3184__3430, new_n3184_);
  and g_13484 (new_n6224_, new_n6389_, new_n6390_);
  or g_13485 (new_n9845_, not_new_n9392_, not_new_n627__2326305139872070);
  or g_13486 (new_n9302_, not_new_n9063_, not_new_n9300_);
  not g_13487 (not_new_n3883_, new_n3883_);
  not g_13488 (not_new_n6165_, new_n6165_);
  and g_13489 (new_n8954_, new_n9322_, and_new_n8982__new_n9323_);
  or g_13490 (new_n6160_, not_new_n5811_, or_not_new_n5893__0_not_new_n6159__0);
  not g_13491 (new_n8322_, new_n8126_);
  and g_13492 (and_new_n1754__new_n1755_, new_n1755_, new_n1754_);
  not g_13493 (not_new_n5427_, new_n5427_);
  not g_13494 (not_po296_4, po296);
  or g_13495 (new_n3823_, not_new_n990_, not_new_n3315__5585458640832840070);
  not g_13496 (not_new_n1534__7, key_gate_5);
  not g_13497 (not_new_n1051__10, new_n1051_);
  or g_13498 (new_n5084_, not_new_n622__3430, not_new_n1599__8);
  or g_13499 (new_n5625_, not_pi133_3, not_new_n5439__0);
  or g_13500 (new_n5619_, not_new_n5618_, not_new_n5617__0);
  not g_13501 (not_new_n9414__0, new_n9414_);
  not g_13502 (not_new_n598__70, new_n598_);
  and g_13503 (new_n6317_, new_n6241_, new_n6375_);
  not g_13504 (new_n5451_, pi138);
  or g_13505 (new_n10271_, not_new_n10270_, not_new_n10269_);
  not g_13506 (not_new_n591__968890104070, new_n591_);
  or g_13507 (new_n7747_, not_new_n7927_, not_new_n7919_);
  not g_13508 (not_new_n8798__2, new_n8798_);
  and g_13509 (new_n5039_, new_n4910_, new_n5190_);
  not g_13510 (not_new_n4218_, new_n4218_);
  or g_13511 (or_not_new_n2545__not_new_n2544_, not_new_n2545_, not_new_n2544_);
  not g_13512 (not_new_n6242__3, new_n6242_);
  or g_13513 (new_n4662_, not_new_n4447__0, not_new_n1012__4);
  not g_13514 (not_new_n1728__0, new_n1728_);
  or g_13515 (or_not_new_n2547__not_new_n2551_, not_new_n2547_, not_new_n2551_);
  not g_13516 (not_new_n6640__2, new_n6640_);
  not g_13517 (new_n8832_, new_n641_);
  not g_13518 (not_new_n9217_, new_n9217_);
  and g_13519 (and_new_n8753__new_n8754_, new_n8753_, new_n8754_);
  not g_13520 (not_new_n628__968890104070, new_n628_);
  not g_13521 (not_new_n9900_, new_n9900_);
  not g_13522 (not_new_n638__47475615099430, new_n638_);
  not g_13523 (not_new_n3977_, key_gate_37);
  not g_13524 (not_new_n8320_, new_n8320_);
  not g_13525 (not_new_n5442_, new_n5442_);
  or g_13526 (new_n6436_, not_new_n6223__0, not_new_n6351_);
  not g_13527 (not_new_n1165_, new_n1165_);
  not g_13528 (not_new_n2800_, new_n2800_);
  and g_13529 (new_n581_, new_n998_, new_n1768_);
  not g_13530 (not_new_n4600_, new_n4600_);
  not g_13531 (not_new_n596__8, key_gate_88);
  or g_13532 (new_n1750_, not_pi094, not_new_n1728__57648010);
  not g_13533 (not_new_n5742_, new_n5742_);
  not g_13534 (not_new_n1047__490, new_n1047_);
  not g_13535 (new_n9538_, new_n9484_);
  not g_13536 (not_new_n9598_, new_n9598_);
  or g_13537 (new_n3701_, not_po298_968890104070, not_new_n630__9);
  or g_13538 (new_n9766_, not_new_n9377_, not_new_n1597__16284135979104490);
  not g_13539 (not_new_n9721_, new_n9721_);
  not g_13540 (not_new_n5658_, new_n5658_);
  not g_13541 (not_new_n7555_, new_n7555_);
  not g_13542 (not_new_n1506_, new_n1506_);
  not g_13543 (not_pi273_1, pi273);
  or g_13544 (new_n4479_, not_new_n4528_, not_new_n4527_);
  or g_13545 (new_n6035_, not_new_n5876_, not_new_n6034_);
  or g_13546 (new_n9253_, not_new_n9251_, not_new_n9252_);
  not g_13547 (not_new_n7632__0, new_n7632_);
  or g_13548 (new_n7501_, not_new_n725__0, not_new_n7439__2);
  or g_13549 (new_n6210_, not_new_n5906_, not_new_n5873_);
  or g_13550 (or_or_not_new_n3944__not_new_n3914__1_not_new_n4014__4, or_not_new_n3944__not_new_n3914__1, not_new_n4014__4);
  not g_13551 (not_new_n3209_, new_n3209_);
  not g_13552 (not_new_n7094_, new_n7094_);
  or g_13553 (new_n9423_, not_new_n9616_, not_new_n9707_);
  not g_13554 (not_new_n1510_, new_n1510_);
  not g_13555 (not_new_n9855__0, new_n9855_);
  not g_13556 (not_new_n9880__0, new_n9880_);
  not g_13557 (not_new_n6676_, new_n6676_);
  not g_13558 (not_new_n5481__0, new_n5481_);
  not g_13559 (not_new_n609__490, new_n609_);
  and g_13560 (new_n5033_, new_n5092_, new_n5141_);
  not g_13561 (not_new_n3695_, new_n3695_);
  or g_13562 (or_or_or_not_new_n2847__not_new_n2850__not_new_n2849__not_new_n2851_, not_new_n2851_, or_or_not_new_n2847__not_new_n2850__not_new_n2849_);
  not g_13563 (not_new_n628__39098210485829880490, new_n628_);
  and g_13564 (new_n5895_, new_n6167_, new_n6166_);
  or g_13565 (new_n2250_, not_new_n5817_, not_new_n1585__6782230728490);
  not g_13566 (not_new_n9966__0, new_n9966_);
  or g_13567 (new_n8770_, not_new_n1604__2824752490, not_new_n8643_);
  or g_13568 (or_not_new_n1319__not_new_n1317_, not_new_n1319_, not_new_n1317_);
  or g_13569 (new_n5626_, not_new_n5624_, not_new_n5625_);
  not g_13570 (not_new_n4511_, new_n4511_);
  not g_13571 (not_new_n8686_, new_n8686_);
  not g_13572 (not_new_n6958_, new_n6958_);
  or g_13573 (new_n3338_, not_new_n3930__0, not_pi064_10);
  or g_13574 (new_n2579_, not_pi263, not_po296_4599865365447399609768010);
  not g_13575 (not_new_n7598__1, new_n7598_);
  not g_13576 (not_new_n10260_, new_n10260_);
  not g_13577 (not_new_n5643_, new_n5643_);
  not g_13578 (not_new_n1535_, key_gate_101);
  not g_13579 (not_new_n633__5, new_n633_);
  or g_13580 (new_n3213_, not_new_n589__490, not_new_n625__7);
  or g_13581 (new_n5972_, not_new_n5971_, not_new_n5715_);
  not g_13582 (not_new_n2764_, new_n2764_);
  not g_13583 (new_n4417_, pi163);
  and g_13584 (and_and_new_n2010__new_n2013__new_n2011_, and_new_n2010__new_n2013_, new_n2011_);
  and g_13585 (new_n6312_, new_n6301_, new_n633_);
  or g_13586 (new_n8458_, not_new_n8527_, not_new_n8229_);
  not g_13587 (not_new_n4284_, new_n4284_);
  not g_13588 (not_new_n1597__4, new_n1597_);
  or g_13589 (new_n1648_, key_gate_19, not_new_n596__4);
  not g_13590 (not_new_n8590_, new_n8590_);
  not g_13591 (not_new_n3129_, new_n3129_);
  or g_13592 (new_n9111_, not_new_n9110_, not_new_n8894_);
  or g_13593 (new_n7152_, not_new_n7080_, not_new_n7330_);
  not g_13594 (not_new_n1580__24010, new_n1580_);
  not g_13595 (not_new_n1061__0, new_n1061_);
  not g_13596 (not_new_n7516_, new_n7516_);
  or g_13597 (new_n3148_, not_new_n646__6, not_new_n581__21838143759917965991093122527538323430);
  not g_13598 (not_new_n594__47475615099430, new_n594_);
  or g_13599 (new_n5650_, not_new_n5507__0, not_pi148_2);
  not g_13600 (not_new_n4130__1, new_n4130_);
  not g_13601 (not_pi253_0, pi253);
  not g_13602 (not_new_n6808_, new_n6808_);
  not g_13603 (not_new_n8541_, new_n8541_);
  not g_13604 (not_new_n625__4, new_n625_);
  or g_13605 (new_n10204_, not_new_n10144__0, not_new_n9940__0);
  or g_13606 (new_n4583_, not_new_n4577_, not_new_n4582_);
  or g_13607 (new_n3660_, not_new_n989__2, not_pi216);
  not g_13608 (not_new_n9663_, new_n9663_);
  or g_13609 (new_n10088_, new_n1051_, new_n647_);
  not g_13610 (new_n7673_, new_n641_);
  not g_13611 (new_n9410_, new_n637_);
  not g_13612 (not_new_n4635_, new_n4635_);
  not g_13613 (not_new_n6978__1, new_n6978_);
  not g_13614 (not_new_n6630_, new_n6630_);
  not g_13615 (not_new_n1351_, new_n1351_);
  or g_13616 (new_n759_, not_new_n3228_, not_new_n3229_);
  or g_13617 (new_n6125_, not_new_n619__10, not_new_n5884_);
  or g_13618 (or_or_not_new_n1863__not_new_n1864__not_new_n1866_, not_new_n1866_, or_not_new_n1863__not_new_n1864_);
  or g_13619 (new_n3221_, not_new_n645__7, not_new_n589__1176490);
  not g_13620 (not_new_n1049__2326305139872070, new_n1049_);
  not g_13621 (not_new_n4471_, new_n4471_);
  not g_13622 (not_new_n7580_, new_n7580_);
  not g_13623 (not_new_n9161_, new_n9161_);
  not g_13624 (not_new_n9899_, new_n9899_);
  or g_13625 (new_n6694_, not_new_n6693_, not_new_n6578_);
  not g_13626 (new_n10036_, new_n9909_);
  not g_13627 (not_new_n628__138412872010, new_n628_);
  or g_13628 (new_n6087_, not_new_n5992_, not_new_n5901_);
  or g_13629 (new_n5018_, not_new_n5402_, not_new_n5401_);
  not g_13630 (not_new_n600__70, new_n600_);
  not g_13631 (not_new_n3364_, new_n3364_);
  not g_13632 (not_new_n633__47475615099430, new_n633_);
  or g_13633 (new_n1628_, not_new_n1627_, not_new_n3315__1);
  not g_13634 (new_n4992_, new_n618_);
  not g_13635 (not_new_n7663__2, new_n7663_);
  not g_13636 (not_new_n630__2326305139872070, new_n630_);
  or g_13637 (new_n6243_, not_new_n6364_, or_or_or_not_new_n6363__not_new_n6358__not_new_n6361__not_new_n6366_);
  not g_13638 (not_new_n595__3430, new_n595_);
  or g_13639 (new_n7296_, not_new_n7295_, not_new_n7095_);
  or g_13640 (or_not_new_n2265__not_new_n2262_, not_new_n2265_, not_new_n2262_);
  not g_13641 (not_new_n2346_, new_n2346_);
  not g_13642 (not_new_n6394_, new_n6394_);
  and g_13643 (new_n4499_, new_n4681_, new_n4682_);
  not g_13644 (not_new_n9418_, new_n9418_);
  not g_13645 (new_n9396_, new_n644_);
  not g_13646 (new_n8617_, new_n1055_);
  or g_13647 (new_n2943_, not_new_n627__3, not_new_n602__968890104070);
  not g_13648 (not_new_n587__19773267430, new_n587_);
  and g_13649 (new_n6965_, new_n7253_, new_n7254_);
  not g_13650 (not_new_n8901_, new_n8901_);
  or g_13651 (new_n4467_, not_new_n4701_, not_new_n4700_);
  or g_13652 (or_or_or_not_new_n2946__not_new_n2949__not_new_n2948__not_new_n2950_, not_new_n2950_, or_or_not_new_n2946__not_new_n2949__not_new_n2948_);
  or g_13653 (po081, key_gate_106, not_new_n1208_);
  not g_13654 (not_pi026_0, pi026);
  and g_13655 (new_n7136_, new_n7466_, new_n7467_);
  not g_13656 (not_new_n7768_, new_n7768_);
  and g_13657 (and_new_n1326__new_n2255_, new_n2255_, new_n1326_);
  or g_13658 (new_n5289_, not_new_n5203__0, not_new_n5281_);
  not g_13659 (not_new_n9842_, new_n9842_);
  or g_13660 (new_n1654_, not_new_n596__6, key_gate_121);
  or g_13661 (new_n5546_, not_pi137_1, not_new_n5447_);
  not g_13662 (not_new_n6242_, new_n6242_);
  not g_13663 (not_new_n3185__19773267430, new_n3185_);
  not g_13664 (not_new_n4122__2, new_n4122_);
  not g_13665 (not_new_n6475_, new_n6475_);
  not g_13666 (not_pi258_1, pi258);
  not g_13667 (not_new_n4000__0, new_n4000_);
  not g_13668 (not_new_n745__0, new_n745_);
  or g_13669 (new_n9664_, not_new_n633__16284135979104490, not_new_n1067__968890104070);
  or g_13670 (or_or_not_new_n2547__not_new_n2551__not_new_n1425_, not_new_n1425_, or_not_new_n2547__not_new_n2551_);
  not g_13671 (new_n5450_, new_n1002_);
  not g_13672 (not_po296_1742514982336908143055105517947102601079450420187483430, po296);
  not g_13673 (not_new_n1576__3, new_n1576_);
  not g_13674 (not_new_n8181_, new_n8181_);
  not g_13675 (not_new_n1602__2824752490, new_n1602_);
  not g_13676 (not_new_n621__968890104070, new_n621_);
  or g_13677 (new_n7459_, not_new_n6974__2326305139872070, not_new_n717_);
  not g_13678 (not_new_n4425__0, new_n4425_);
  xnor g_13679 (key_gate_54, key_54, not_new_n1648_);
  or g_13680 (new_n970_, not_new_n2210_, or_or_not_new_n1319__not_new_n1317__not_new_n2211_);
  or g_13681 (new_n10279_, not_new_n10012_, not_new_n10013__1);
  or g_13682 (new_n3049_, not_new_n3372__968890104070, not_new_n632__4);
  not g_13683 (not_new_n989__70, new_n989_);
  not g_13684 (not_new_n4156_, new_n4156_);
  or g_13685 (po245, not_new_n3677_, not_new_n3676_);
  or g_13686 (new_n2335_, not_new_n594__16284135979104490, not_new_n9960_);
  or g_13687 (new_n4887_, not_new_n4797__1, not_new_n4829__1);
  or g_13688 (new_n2207_, not_pi121, not_new_n588__968890104070);
  not g_13689 (not_new_n9815_, new_n9815_);
  not g_13690 (new_n4553_, new_n4504_);
  not g_13691 (not_new_n3998_, key_gate_114);
  not g_13692 (not_new_n1018__7, new_n1018_);
  or g_13693 (or_not_new_n2655__not_new_n2654_, not_new_n2655_, not_new_n2654_);
  not g_13694 (not_new_n3107_, new_n3107_);
  or g_13695 (new_n7320_, not_new_n7179_, not_new_n7113_);
  or g_13696 (or_or_not_new_n1977__not_new_n1978__not_new_n1980_, not_new_n1980_, or_not_new_n1977__not_new_n1978_);
  not g_13697 (not_new_n4209_, new_n4209_);
  not g_13698 (not_new_n611__9, new_n611_);
  not g_13699 (not_pi262, pi262);
  or g_13700 (new_n2238_, not_new_n9964_, not_new_n594__968890104070);
  not g_13701 (new_n8308_, new_n8125_);
  and g_13702 (new_n5837_, new_n5929_, new_n5919_);
  not g_13703 (not_new_n7629_, new_n7629_);
  not g_13704 (not_new_n7515_, new_n7515_);
  not g_13705 (not_new_n1585__490, new_n1585_);
  not g_13706 (not_new_n3482_, new_n3482_);
  not g_13707 (not_new_n2693_, new_n2693_);
  or g_13708 (new_n6031_, not_new_n6030_, not_new_n5916__0);
  not g_13709 (not_new_n3144_, new_n3144_);
  not g_13710 (not_new_n4500__0, new_n4500_);
  not g_13711 (not_new_n1028__10, new_n1028_);
  not g_13712 (new_n4237_, new_n675_);
  and g_13713 (new_n8946_, new_n9114_, new_n8979_);
  not g_13714 (not_pi193, pi193);
  or g_13715 (new_n5325_, not_new_n619__9, not_new_n5059__0);
  not g_13716 (not_new_n586__6, new_n586_);
  or g_13717 (new_n9284_, not_new_n8876_, not_new_n646__47475615099430);
  or g_13718 (new_n9531_, new_n1047_, new_n634_);
  not g_13719 (new_n4071_, pi269);
  or g_13720 (new_n7539_, not_new_n731__0, not_new_n7421__0);
  not g_13721 (not_new_n4686_, new_n4686_);
  or g_13722 (new_n7196_, not_new_n6982__0, not_new_n7354__0);
  not g_13723 (not_new_n8913_, new_n8913_);
  or g_13724 (new_n5395_, not_new_n5393_, not_new_n5166__0);
  not g_13725 (not_new_n775__1, new_n775_);
  and g_13726 (and_new_n1338__new_n2312_, new_n1338_, new_n2312_);
  or g_13727 (new_n1620_, not_po298, not_new_n776_);
  or g_13728 (new_n6199_, not_new_n5786__2, not_new_n638__403536070);
  or g_13729 (or_or_or_not_new_n2776__not_new_n2779__not_new_n2778__not_new_n2780_, or_or_not_new_n2776__not_new_n2779__not_new_n2778_, not_new_n2780_);
  not g_13730 (not_new_n600__5, new_n600_);
  or g_13731 (new_n5440_, not_new_n5532_, not_new_n5531_);
  and g_13732 (new_n1265_, new_n1965_, new_n1966_);
  not g_13733 (not_new_n4137__1, new_n4137_);
  not g_13734 (not_new_n1534__797922662976120010, key_gate_5);
  not g_13735 (not_new_n647__5, new_n647_);
  and g_13736 (and_and_new_n1053__new_n6232__new_n6395_, and_new_n1053__new_n6232_, new_n6395_);
  not g_13737 (not_new_n6631__1, new_n6631_);
  not g_13738 (not_new_n1045__2, new_n1045_);
  or g_13739 (new_n3681_, not_po298_3430, not_new_n644__9);
  not g_13740 (not_new_n1061__3, new_n1061_);
  xor g_13741 (key_gate_86, not_new_n3932_, key_86);
  and g_13742 (new_n1498_, new_n3022_, new_n1499_);
  not g_13743 (not_new_n4257_, new_n4257_);
  not g_13744 (not_new_n7380_, new_n7380_);
  not g_13745 (not_new_n1028__4, new_n1028_);
  not g_13746 (not_new_n4285_, new_n4285_);
  or g_13747 (new_n10114_, not_new_n9915_, not_new_n9916_);
  not g_13748 (not_new_n7554_, new_n7554_);
  not g_13749 (not_new_n2975_, new_n2975_);
  not g_13750 (not_new_n581__445676403263631959001900459745680070, new_n581_);
  not g_13751 (not_new_n1006__4, new_n1006_);
  not g_13752 (not_new_n984__490, new_n984_);
  not g_13753 (not_new_n6093_, new_n6093_);
  or g_13754 (new_n9757_, not_new_n9635_, not_new_n9755_);
  or g_13755 (new_n10332_, not_new_n10330_, not_new_n10231_);
  or g_13756 (new_n3625_, not_new_n960_, not_new_n1611__1176490);
  not g_13757 (new_n4829_, new_n4740_);
  not g_13758 (not_new_n9929__0, new_n9929_);
  or g_13759 (new_n5375_, not_new_n4975__0, not_new_n640__24010);
  not g_13760 (new_n7317_, new_n6989_);
  or g_13761 (new_n8400_, not_new_n8282__0, not_new_n8399_);
  or g_13762 (new_n6878_, not_new_n6876_, or_not_new_n6538__1_not_new_n6877_);
  not g_13763 (not_new_n10005_, new_n10005_);
  not g_13764 (new_n6988_, new_n736_);
  not g_13765 (not_new_n9934__0, new_n9934_);
  not g_13766 (not_new_n1537__1176490, new_n1537_);
  or g_13767 (new_n8847_, not_new_n9023_, not_new_n9022_);
  or g_13768 (or_not_new_n2615__not_new_n2614_, not_new_n2615_, not_new_n2614_);
  not g_13769 (not_new_n600__3430, new_n600_);
  and g_13770 (new_n9978_, and_new_n10047__new_n10048_, new_n10050_);
  and g_13771 (new_n6453_, new_n6678_, new_n6656_);
  not g_13772 (not_new_n598__138412872010, new_n598_);
  or g_13773 (new_n9189_, not_new_n9103__0, not_new_n9181_);
  not g_13774 (not_new_n8875_, new_n8875_);
  or g_13775 (new_n2879_, not_new_n627__2, not_new_n604__168070);
  or g_13776 (new_n3132_, not_new_n1602__3, not_new_n928__168070);
  or g_13777 (new_n3618_, not_pi175_0, not_new_n984__3430);
  not g_13778 (not_new_n7739__2, new_n7739_);
  buf g_13779 (po045, pi219);
  not g_13780 (not_new_n4084_, new_n4084_);
  or g_13781 (new_n1937_, not_new_n1049_, not_new_n1588__8);
  not g_13782 (not_new_n7115__0, new_n7115_);
  not g_13783 (not_po296, po296);
  not g_13784 (not_new_n9552_, new_n9552_);
  or g_13785 (new_n3062_, not_new_n581__6782230728490, not_new_n1063__2);
  not g_13786 (not_new_n8357_, new_n8357_);
  not g_13787 (not_new_n6242__1, new_n6242_);
  and g_13788 (new_n6366_, and_and_new_n6365__new_n6439__new_n6438_, new_n6437_);
  not g_13789 (not_new_n765_, new_n765_);
  or g_13790 (new_n625_, or_or_not_new_n2170__not_new_n2167__not_new_n2168_, not_new_n2169_);
  not g_13791 (not_new_n591__8235430, new_n591_);
  not g_13792 (not_new_n6354_, new_n6354_);
  or g_13793 (new_n8465_, not_new_n1049__138412872010, not_new_n8105__2);
  and g_13794 (and_new_n2314__new_n2317_, new_n2314_, new_n2317_);
  not g_13795 (not_new_n1027__13410686196639649008070, new_n1027_);
  not g_13796 (not_po296_5585458640832840070, po296);
  not g_13797 (not_new_n3462_, new_n3462_);
  not g_13798 (not_new_n1018__6, new_n1018_);
  not g_13799 (not_new_n3399_, new_n3399_);
  not g_13800 (not_new_n645__1, new_n645_);
  or g_13801 (new_n7984_, not_new_n7741__0, not_new_n619__1176490);
  or g_13802 (new_n10023_, not_new_n9890_, not_new_n10176_);
  or g_13803 (new_n7398_, not_new_n7025__1, not_new_n6984__1);
  or g_13804 (new_n4514_, pi163, new_n1009_);
  not g_13805 (not_new_n677_, new_n677_);
  not g_13806 (not_new_n605__24010, new_n605_);
  not g_13807 (not_new_n581__9, new_n581_);
  xor g_13808 (key_gate_102, key_102, not_new_n1699_);
  not g_13809 (not_new_n1479_, new_n1479_);
  or g_13810 (new_n7620_, or_not_new_n7906__not_new_n7780_, not_new_n7764_);
  not g_13811 (not_new_n1601__93874803376477543056490, new_n1601_);
  not g_13812 (not_new_n638__2824752490, new_n638_);
  or g_13813 (new_n3356_, not_pi064_403536070, not_new_n3998__0);
  not g_13814 (not_new_n9935_, new_n9935_);
  not g_13815 (not_new_n1537__797922662976120010, new_n1537_);
  or g_13816 (new_n5511_, not_new_n5574_, not_new_n5573_);
  not g_13817 (not_new_n4946_, new_n4946_);
  not g_13818 (not_new_n1581__168070, new_n1581_);
  not g_13819 (not_new_n8167_, new_n8167_);
  or g_13820 (new_n5379_, not_new_n4972_, not_new_n645__24010);
  or g_13821 (new_n9007_, not_new_n9006_, not_new_n634__47475615099430);
  or g_13822 (new_n3515_, not_new_n1613__47475615099430, not_new_n2280_);
  and g_13823 (new_n602_, new_n1595_, new_n3366_);
  or g_13824 (new_n3458_, not_new_n1018__1, not_new_n1594__10);
  and g_13825 (new_n4306_, new_n4367_, new_n4368_);
  or g_13826 (new_n1763_, not_pi162, not_new_n586_);
  not g_13827 (new_n8607_, new_n1039_);
  not g_13828 (not_new_n3530_, new_n3530_);
  not g_13829 (not_new_n6963_, new_n6963_);
  or g_13830 (new_n1956_, not_new_n1051_, not_new_n1588__9);
  not g_13831 (not_pi260_3, pi260);
  or g_13832 (po256, not_new_n3698_, not_new_n3699_);
  or g_13833 (new_n7475_, not_new_n7454__2, not_new_n720__0);
  not g_13834 (not_new_n7143__0, new_n7143_);
  not g_13835 (not_new_n4223_, new_n4223_);
  not g_13836 (not_new_n10122_, new_n10122_);
  not g_13837 (not_new_n989__24010, new_n989_);
  buf g_13838 (po043, pi221);
  not g_13839 (not_new_n9038_, new_n9038_);
  not g_13840 (not_new_n6233_, new_n6233_);
  or g_13841 (or_or_not_new_n2577__not_new_n2581__not_new_n1431_, or_not_new_n2577__not_new_n2581_, not_new_n1431_);
  or g_13842 (or_not_new_n1553__not_new_n1376_, not_new_n1553_, not_new_n1376_);
  not g_13843 (not_new_n4098_, new_n4098_);
  not g_13844 (not_new_n6090_, new_n6090_);
  or g_13845 (new_n7458_, not_new_n7134_, not_new_n775__16284135979104490);
  not g_13846 (not_new_n775__2824752490, new_n775_);
  or g_13847 (new_n6564_, not_new_n6883_, not_new_n6882_);
  or g_13848 (new_n5082_, not_new_n647__3430, not_new_n1051__8);
  not g_13849 (not_new_n3272_, new_n3272_);
  not g_13850 (new_n8853_, new_n629_);
  not g_13851 (not_new_n7610_, new_n7610_);
  not g_13852 (not_new_n3210_, new_n3210_);
  or g_13853 (new_n5997_, not_new_n1601__70, not_new_n5770_);
  not g_13854 (new_n8134_, new_n630_);
  or g_13855 (new_n4011_, not_new_n3938_, not_pi036_3);
  not g_13856 (not_new_n2916_, new_n2916_);
  not g_13857 (not_pi021, pi021);
  not g_13858 (not_pi139_1, pi139);
  not g_13859 (not_new_n5096_, new_n5096_);
  or g_13860 (new_n6113_, not_new_n5882__2, not_new_n5965_);
  not g_13861 (not_po296_3788186922656647816827176259430, po296);
  not g_13862 (not_pi064_0, pi064);
  not g_13863 (not_new_n4965_, new_n4965_);
  or g_13864 (new_n10226_, not_new_n9980_, not_new_n10225_);
  not g_13865 (not_new_n9382__0, new_n9382_);
  not g_13866 (not_new_n1597__10, new_n1597_);
  or g_13867 (new_n2405_, not_new_n1053__1, not_new_n598__9);
  or g_13868 (new_n3328_, not_pi064_5, not_new_n3977__0);
  not g_13869 (not_new_n1614_, new_n1614_);
  not g_13870 (not_new_n2734_, new_n2734_);
  or g_13871 (new_n2696_, or_not_new_n2695__not_new_n2694_, not_new_n2693_);
  not g_13872 (not_new_n9118__0, new_n9118_);
  and g_13873 (new_n5722_, new_n5921_, new_n5943_);
  or g_13874 (new_n4883_, not_new_n4831__1, not_new_n4792__1);
  not g_13875 (not_new_n1881__0, new_n1881_);
  and g_13876 (new_n8247_, new_n8479_, new_n8480_);
  not g_13877 (not_new_n645__2, new_n645_);
  or g_13878 (new_n7678_, not_new_n8031_, not_new_n8032_);
  or g_13879 (po253, not_new_n3693_, not_new_n3692_);
  or g_13880 (or_or_or_not_new_n6226__0_not_new_n6336__not_new_n6373__5_not_new_n6242__2, not_new_n6242__2, or_or_not_new_n6226__0_not_new_n6336__not_new_n6373__5);
  not g_13881 (not_new_n594__0, new_n594_);
  not g_13882 (not_new_n3901_, new_n3901_);
  not g_13883 (new_n9401_, new_n645_);
  not g_13884 (not_new_n9406_, new_n9406_);
  not g_13885 (not_new_n10029__0, new_n10029_);
  not g_13886 (not_new_n8966_, new_n8966_);
  not g_13887 (not_new_n6979__0, new_n6979_);
  not g_13888 (not_new_n3497_, new_n3497_);
  and g_13889 (new_n1328_, new_n2259_, and_and_new_n2257__new_n2260__new_n2258_);
  and g_13890 (new_n1321_, new_n2231_, new_n2232_);
  or g_13891 (new_n9299_, not_new_n1063__138412872010, not_new_n8858__0);
  and g_13892 (new_n8699_, new_n8708_, new_n8717_);
  not g_13893 (not_new_n6443__6, new_n6443_);
  or g_13894 (new_n7256_, not_new_n719_, not_new_n7043_);
  not g_13895 (new_n5529_, new_n5502_);
  not g_13896 (not_new_n7627__2, new_n7627_);
  not g_13897 (new_n8887_, new_n630_);
  not g_13898 (not_new_n724__0, new_n724_);
  or g_13899 (po086, not_new_n3378_, not_new_n3379_);
  not g_13900 (not_new_n586__490, new_n586_);
  not g_13901 (not_new_n1602__19773267430, new_n1602_);
  or g_13902 (new_n7044_, not_new_n7453_, not_new_n7452_);
  or g_13903 (new_n2527_, not_new_n2526_, not_new_n611__5);
  not g_13904 (not_new_n5916__0, new_n5916_);
  not g_13905 (not_new_n1013__3, new_n1013_);
  not g_13906 (not_new_n2502_, new_n2502_);
  and g_13907 (new_n7585_, new_n7858_, new_n7584_);
  not g_13908 (not_new_n3481_, new_n3481_);
  or g_13909 (new_n3642_, not_new_n984__47475615099430, not_pi187_0);
  not g_13910 (not_new_n5322_, new_n5322_);
  not g_13911 (not_new_n1585__138412872010, new_n1585_);
  not g_13912 (not_new_n4179_, new_n4179_);
  not g_13913 (not_new_n1232_, new_n1232_);
  or g_13914 (new_n4705_, not_pi172_3, not_new_n4436__0);
  or g_13915 (new_n3745_, not_new_n1598__6, not_new_n621__10);
  or g_13916 (new_n3675_, not_new_n626__9, not_po298_10);
  and g_13917 (new_n1342_, and_and_new_n2327__new_n2328__new_n2331_, new_n2330_);
  and g_13918 (new_n4316_, new_n4398_, new_n4397_);
  not g_13919 (not_pi263_1, pi263);
  not g_13920 (not_new_n5752_, new_n5752_);
  not g_13921 (not_new_n1039__113988951853731430, new_n1039_);
  not g_13922 (not_new_n5408_, new_n5408_);
  not g_13923 (not_new_n2591_, new_n2591_);
  not g_13924 (not_new_n5782_, new_n5782_);
  not g_13925 (not_new_n9667_, new_n9667_);
  not g_13926 (not_new_n9914_, new_n9914_);
  not g_13927 (not_new_n7091_, new_n7091_);
  not g_13928 (not_new_n8216_, new_n8216_);
  not g_13929 (not_new_n7611_, new_n7611_);
  not g_13930 (not_new_n3130_, new_n3130_);
  or g_13931 (new_n5346_, not_new_n622__24010, not_new_n4989_);
  not g_13932 (not_new_n9854__1, new_n9854_);
  not g_13933 (not_new_n688_, new_n688_);
  or g_13934 (new_n4768_, not_new_n4770__0, not_new_n4839__0);
  not g_13935 (not_new_n4110_, new_n4110_);
  not g_13936 (not_new_n1589__403536070, new_n1589_);
  not g_13937 (not_new_n4996_, new_n4996_);
  and g_13938 (new_n1331_, and_new_n1330__new_n2274_, new_n2273_);
  or g_13939 (new_n9158_, not_new_n9038_, not_new_n8991__0);
  or g_13940 (new_n10068_, not_new_n632__5585458640832840070, not_new_n1037__2326305139872070);
  not g_13941 (new_n4103_, pi271);
  not g_13942 (new_n10052_, new_n9900_);
  not g_13943 (not_new_n5443_, new_n5443_);
  or g_13944 (new_n8302_, not_new_n8290_, not_new_n8286_);
  or g_13945 (new_n10111_, new_n1067_, new_n633_);
  not g_13946 (not_new_n8898_, new_n8898_);
  not g_13947 (not_new_n589__4, new_n589_);
  or g_13948 (new_n2580_, not_new_n1017__0, not_new_n608__6);
  or g_13949 (new_n6567_, not_new_n6938_, not_new_n6937_);
  or g_13950 (new_n8794_, not_new_n8796_, not_new_n8714_);
  not g_13951 (not_po296_8235430, po296);
  not g_13952 (not_new_n4316_, new_n4316_);
  and g_13953 (new_n4898_, new_n5090_, new_n5089_);
  not g_13954 (new_n4957_, new_n1063_);
  not g_13955 (not_new_n7664__0, new_n7664_);
  or g_13956 (new_n4528_, not_pi166_1, not_new_n1006__2);
  not g_13957 (not_new_n3781_, new_n3781_);
  or g_13958 (new_n10143_, not_new_n10141_, not_new_n9994_);
  not g_13959 (not_new_n1024__0, new_n1024_);
  or g_13960 (new_n679_, or_not_new_n3176__not_new_n3175_, not_new_n3174_);
  not g_13961 (not_new_n7904_, new_n7904_);
  or g_13962 (new_n6725_, not_new_n6517_, not_new_n633__57648010);
  or g_13963 (new_n6896_, not_new_n6894_, not_new_n6895_);
  not g_13964 (new_n4444_, new_n1014_);
  or g_13965 (or_not_new_n1323__not_new_n1321_, not_new_n1323_, not_new_n1321_);
  not g_13966 (not_new_n4676_, new_n4676_);
  or g_13967 (new_n8787_, not_new_n8650_, not_new_n1160__0);
  not g_13968 (not_new_n1596__19773267430, new_n1596_);
  not g_13969 (not_new_n6332_, new_n6332_);
  not g_13970 (not_new_n610__5, new_n610_);
  not g_13971 (new_n6301_, new_n1067_);
  not g_13972 (not_new_n2342_, new_n2342_);
  not g_13973 (not_new_n1055__1176490, new_n1055_);
  or g_13974 (new_n3020_, not_new_n1159_, not_new_n1027__3430);
  not g_13975 (not_new_n606__70, new_n606_);
  not g_13976 (not_new_n2167_, new_n2167_);
  not g_13977 (not_new_n4135__0, new_n4135_);
  not g_13978 (new_n9516_, new_n9387_);
  not g_13979 (not_new_n6303_, new_n6303_);
  not g_13980 (not_new_n611__8, new_n611_);
  not g_13981 (not_new_n588__9, new_n588_);
  not g_13982 (not_new_n8515_, new_n8515_);
  and g_13983 (new_n6346_, new_n6373_, new_n6274_);
  not g_13984 (not_new_n1580__332329305696010, new_n1580_);
  not g_13985 (not_new_n5894_, new_n5894_);
  not g_13986 (not_new_n8275_, new_n8275_);
  or g_13987 (new_n3262_, not_new_n617__8, not_new_n3184__7);
  or g_13988 (new_n4044_, not_new_n3997_, not_new_n4013_);
  not g_13989 (not_new_n8658_, new_n8658_);
  not g_13990 (not_new_n5193_, new_n5193_);
  or g_13991 (new_n7212_, not_new_n6996_, not_new_n7409_);
  not g_13992 (not_new_n9339_, new_n9339_);
  or g_13993 (new_n9286_, not_new_n9285_, not_new_n9284_);
  or g_13994 (new_n2399_, not_new_n599__8, not_new_n9955__0);
  not g_13995 (not_new_n1199_, new_n1199_);
  not g_13996 (not_new_n6777_, new_n6777_);
  or g_13997 (new_n8063_, not_new_n7730_, not_new_n7760_);
  and g_13998 (new_n1298_, new_n2119_, new_n2120_);
  not g_13999 (not_new_n2247_, new_n2247_);
  or g_14000 (new_n9444_, not_new_n9816_, not_new_n9815_);
  or g_14001 (new_n7692_, not_new_n8053_, not_new_n8054_);
  not g_14002 (not_new_n1045__1, new_n1045_);
  not g_14003 (not_new_n4170__0, new_n4170_);
  not g_14004 (new_n5796_, new_n636_);
  not g_14005 (not_new_n2795_, new_n2795_);
  or g_14006 (new_n6822_, not_new_n6579_, not_new_n6821_);
  or g_14007 (new_n1772_, not_new_n8102_, not_new_n1581_);
  not g_14008 (not_new_n1576__3430, new_n1576_);
  or g_14009 (new_n9261_, not_new_n8967_, not_new_n8888__0);
  not g_14010 (not_new_n2634_, new_n2634_);
  or g_14011 (new_n3619_, not_new_n957_, not_new_n1611__3430);
  not g_14012 (not_new_n8884_, new_n8884_);
  not g_14013 (not_pi097_0, pi097);
  not g_14014 (not_new_n631__2, new_n631_);
  or g_14015 (new_n6306_, not_new_n6415_, not_new_n6414_);
  not g_14016 (not_new_n5377_, new_n5377_);
  or g_14017 (new_n1980_, not_new_n4135_, not_new_n585__70);
  not g_14018 (not_new_n3940_, new_n3940_);
  or g_14019 (new_n9779_, not_new_n629__2326305139872070, not_new_n9380_);
  or g_14020 (new_n2861_, not_new_n604__3430, not_new_n638__2);
  not g_14021 (not_new_n1585__0, new_n1585_);
  not g_14022 (not_new_n4445__0, new_n4445_);
  not g_14023 (new_n9169_, new_n8839_);
  not g_14024 (new_n7926_, new_n7750_);
  not g_14025 (not_new_n5581_, new_n5581_);
  not g_14026 (not_new_n629__0, new_n629_);
  not g_14027 (not_new_n8870_, new_n8870_);
  not g_14028 (not_new_n9015_, new_n9015_);
  not g_14029 (not_new_n4122_, new_n4122_);
  or g_14030 (new_n1701_, not_po296_138412872010, not_pi009_0);
  or g_14031 (new_n3406_, not_new_n1613_, not_new_n1781_);
  or g_14032 (new_n3519_, not_new_n2318_, not_new_n1613__2326305139872070);
  or g_14033 (new_n7359_, not_new_n769_, not_new_n6974__6);
  or g_14034 (new_n3097_, not_new_n3315__5, not_new_n631__5);
  not g_14035 (not_pi176_1, pi176);
  or g_14036 (new_n9716_, not_new_n9714__0, or_not_new_n9469__not_new_n9339_);
  and g_14037 (and_new_n3804__new_n3807_, new_n3804_, new_n3807_);
  not g_14038 (not_new_n10248_, new_n10248_);
  not g_14039 (not_new_n1323_, new_n1323_);
  not g_14040 (not_new_n1621_, new_n1621_);
  not g_14041 (not_new_n637_, new_n637_);
  not g_14042 (new_n5470_, pi146);
  not g_14043 (new_n6296_, new_n1049_);
  and g_14044 (and_new_n2517__new_n2518_, new_n2517_, new_n2518_);
  not g_14045 (not_new_n1576__57648010, new_n1576_);
  not g_14046 (new_n6891_, new_n6595_);
  not g_14047 (not_new_n4713_, new_n4713_);
  or g_14048 (new_n4655_, not_new_n1011__4, not_new_n4449__0);
  not g_14049 (not_new_n4993__0, new_n4993_);
  or g_14050 (new_n8448_, not_new_n8212_, not_new_n8244__2);
  or g_14051 (or_not_new_n1158__0_not_new_n8713__1, not_new_n8713__1, not_new_n1158__0);
  not g_14052 (not_new_n4842_, new_n4842_);
  not g_14053 (not_new_n1583__70, new_n1583_);
  or g_14054 (new_n659_, not_new_n3135_, or_not_new_n3136__not_new_n3137_);
  not g_14055 (not_new_n1341_, new_n1341_);
  not g_14056 (not_new_n4245_, new_n4245_);
  not g_14057 (not_new_n1071__138412872010, new_n1071_);
  or g_14058 (new_n3534_, not_pi133_0, not_new_n1538__3);
  not g_14059 (not_new_n3959_, new_n3959_);
  or g_14060 (new_n6136_, not_new_n1597__490, not_new_n5767__1);
  not g_14061 (not_new_n9079_, new_n9079_);
  not g_14062 (not_new_n626__332329305696010, new_n626_);
  not g_14063 (not_new_n764_, new_n764_);
  or g_14064 (new_n7171_, not_new_n6984_, not_new_n7351_);
  and g_14065 (new_n7583_, new_n7846_, new_n7848_);
  not g_14066 (new_n5925_, new_n5795_);
  not g_14067 (new_n4440_, new_n1016_);
  not g_14068 (not_new_n8849_, new_n8849_);
  not g_14069 (not_new_n6126_, new_n6126_);
  not g_14070 (not_new_n7620__0, new_n7620_);
  or g_14071 (or_not_new_n10045__1_not_new_n9855__1, not_new_n9855__1, not_new_n10045__1);
  or g_14072 (new_n3083_, not_new_n1031__5, not_new_n581__5585458640832840070);
  not g_14073 (not_new_n628__3430, new_n628_);
  not g_14074 (new_n8143_, new_n1604_);
  or g_14075 (new_n2277_, not_new_n593__47475615099430, not_new_n617_);
  or g_14076 (new_n7402_, not_new_n7302_, not_new_n6991__1);
  not g_14077 (not_new_n1535__0, key_gate_101);
  or g_14078 (new_n3509_, not_new_n1613__138412872010, not_new_n2223_);
  not g_14079 (new_n4431_, new_n1002_);
  not g_14080 (not_new_n2134_, new_n2134_);
  not g_14081 (not_new_n7448__0, new_n7448_);
  not g_14082 (not_new_n5769_, new_n5769_);
  not g_14083 (not_new_n1020__7, new_n1020_);
  not g_14084 (not_new_n643__6782230728490, new_n643_);
  or g_14085 (new_n7763_, not_new_n7713_, not_new_n7744_);
  not g_14086 (not_new_n10083_, new_n10083_);
  not g_14087 (not_new_n1491_, new_n1491_);
  not g_14088 (not_new_n622__7, new_n622_);
  not g_14089 (not_new_n647__0, new_n647_);
  or g_14090 (new_n6424_, not_new_n6233_, or_or_not_new_n6335__not_new_n6373__4_not_new_n1071__490);
  xor g_14091 (key_gate_38, not_pi275_0, key_38);
  not g_14092 (not_new_n3925_, key_gate_85);
  or g_14093 (new_n9722_, not_new_n9721_, not_new_n9720_);
  not g_14094 (not_new_n1730__0, new_n1730_);
  not g_14095 (not_new_n7019_, new_n7019_);
  not g_14096 (not_new_n10329_, new_n10329_);
  or g_14097 (po280, not_new_n2848_, or_or_or_not_new_n2847__not_new_n2850__not_new_n2849__not_new_n2851_);
  not g_14098 (not_new_n4779__0, new_n4779_);
  or g_14099 (new_n1945_, not_new_n1583__8, not_new_n7684_);
  not g_14100 (not_new_n9866_, new_n9866_);
  or g_14101 (new_n7725_, not_new_n8034_, not_new_n8033_);
  or g_14102 (new_n3430_, not_new_n1537__4, not_pi102_0);
  not g_14103 (not_new_n4226_, new_n4226_);
  not g_14104 (not_new_n4835_, new_n4835_);
  not g_14105 (not_new_n8235_, new_n8235_);
  not g_14106 (not_new_n5681_, new_n5681_);
  not g_14107 (not_new_n1043__8235430, new_n1043_);
  or g_14108 (po266, not_new_n2714_, not_new_n1471_);
  not g_14109 (not_new_n1059__4, new_n1059_);
  not g_14110 (not_new_n3372__39098210485829880490, new_n3372_);
  not g_14111 (not_new_n3185__3, new_n3185_);
  or g_14112 (new_n5698_, not_new_n1018__6, not_new_n5455_);
  or g_14113 (new_n7298_, not_new_n7031__0, not_new_n732__0);
  not g_14114 (not_pi165_0, pi165);
  or g_14115 (or_not_new_n6897__not_new_n6798_, not_new_n6798_, not_new_n6897_);
  or g_14116 (new_n2795_, not_new_n3310__4, not_new_n4134__2);
  not g_14117 (not_new_n7427__0, new_n7427_);
  and g_14118 (new_n1337_, new_n2307_, new_n2308_);
  and g_14119 (and_new_n1043__new_n6232_, new_n6232_, new_n1043_);
  or g_14120 (new_n3813_, not_new_n3811_, not_new_n3812_);
  not g_14121 (not_new_n1591__3, new_n1591_);
  not g_14122 (not_new_n5920__0, new_n5920_);
  or g_14123 (new_n5372_, not_new_n639__168070, not_new_n4979__0);
  not g_14124 (not_new_n644__2824752490, new_n644_);
  or g_14125 (or_or_or_not_new_n2874__not_new_n2877__not_new_n2876__not_new_n2878_, not_new_n2878_, or_or_not_new_n2874__not_new_n2877__not_new_n2876_);
  not g_14126 (not_new_n5078_, new_n5078_);
  not g_14127 (not_new_n7781__0, new_n7781_);
  or g_14128 (new_n8406_, not_new_n1055__332329305696010, not_new_n8155__1);
  not g_14129 (not_new_n634__0, new_n634_);
  not g_14130 (not_new_n4200_, new_n4200_);
  not g_14131 (not_new_n664_, new_n664_);
  not g_14132 (not_new_n1069__968890104070, new_n1069_);
  not g_14133 (not_new_n6709_, new_n6709_);
  or g_14134 (new_n2143_, not_new_n9967_, not_new_n594__57648010);
  not g_14135 (new_n4175_, new_n4148_);
  or g_14136 (new_n7358_, not_new_n775__7, not_new_n7106_);
  not g_14137 (not_new_n9248_, new_n9248_);
  or g_14138 (new_n9309_, not_new_n9060_, not_new_n9307_);
  not g_14139 (new_n7665_, new_n618_);
  or g_14140 (new_n6977_, not_new_n7020_, not_new_n739_);
  not g_14141 (not_new_n6000_, new_n6000_);
  not g_14142 (not_new_n6607_, new_n6607_);
  not g_14143 (new_n10031_, new_n9888_);
  or g_14144 (new_n2899_, not_pi265_2, not_new_n994__2824752490);
  not g_14145 (not_new_n595__5, new_n595_);
  not g_14146 (not_new_n1159_, new_n1159_);
  not g_14147 (not_new_n10198_, new_n10198_);
  not g_14148 (not_new_n4265_, new_n4265_);
  not g_14149 (not_new_n922__1, new_n922_);
  or g_14150 (new_n2517_, not_new_n611__4, or_not_new_n5484__not_new_n605__0);
  not g_14151 (not_new_n9761_, new_n9761_);
  not g_14152 (new_n9908_, new_n646_);
  not g_14153 (not_new_n7773_, new_n7773_);
  or g_14154 (new_n2991_, not_new_n1027__3, not_new_n1149_);
  and g_14155 (and_new_n2697__new_n2698_, new_n2697_, new_n2698_);
  or g_14156 (new_n9729_, not_new_n9727_, not_new_n9538_);
  not g_14157 (not_new_n606__5, new_n606_);
  or g_14158 (new_n6105_, not_new_n635__1176490, not_new_n5743__0);
  or g_14159 (new_n2659_, not_pi257, not_po296_26517308458596534717790233816010);
  not g_14160 (not_new_n585__2326305139872070, new_n585_);
  not g_14161 (new_n4281_, new_n684_);
  not g_14162 (new_n4565_, new_n4498_);
  not g_14163 (not_new_n5704_, new_n5704_);
  not g_14164 (not_new_n2888_, new_n2888_);
  or g_14165 (new_n7474_, not_new_n7043__1, not_new_n7013__1);
  or g_14166 (new_n8491_, not_new_n8249_, not_new_n8294__0);
  not g_14167 (not_new_n928__7, new_n928_);
  and g_14168 (new_n3987_, new_n4059_, new_n4060_);
  not g_14169 (not_new_n7152__0, new_n7152_);
  or g_14170 (or_not_new_n5203__not_new_n5087__0, not_new_n5087__0, not_new_n5203_);
  or g_14171 (new_n8057_, not_new_n7896_, not_new_n7759__2);
  or g_14172 (new_n3571_, not_new_n2204__0, not_new_n1612__19773267430);
  or g_14173 (new_n4607_, not_new_n4605_, not_new_n4533_);
  not g_14174 (not_new_n3397_, new_n3397_);
  or g_14175 (new_n6151_, not_new_n5860_, not_new_n5891__0);
  not g_14176 (not_pi144_2, pi144);
  or g_14177 (new_n3329_, not_new_n1534__6, not_pi040_0);
  not g_14178 (not_new_n6479_, new_n6479_);
  not g_14179 (not_new_n610__70, new_n610_);
  not g_14180 (not_new_n5200_, new_n5200_);
  not g_14181 (not_new_n610__8235430, new_n610_);
  not g_14182 (not_new_n989__19773267430, new_n989_);
  not g_14183 (not_new_n8660_, new_n8660_);
  not g_14184 (not_new_n4158_, new_n4158_);
  not g_14185 (not_new_n5595_, new_n5595_);
  not g_14186 (new_n4033_, new_n3949_);
  not g_14187 (not_new_n3214_, new_n3214_);
  not g_14188 (not_new_n10177_, new_n10177_);
  not g_14189 (new_n7001_, new_n731_);
  or g_14190 (new_n5647_, not_new_n5508_, not_new_n1028__70);
  or g_14191 (new_n4585_, not_new_n4471_, not_new_n4583_);
  not g_14192 (not_new_n9381_, new_n9381_);
  not g_14193 (not_new_n7167_, new_n7167_);
  or g_14194 (new_n2747_, not_new_n4116__1, not_new_n994__3);
  not g_14195 (not_new_n644__16284135979104490, new_n644_);
  not g_14196 (not_new_n4113_, new_n4113_);
  not g_14197 (not_new_n597__8, new_n597_);
  or g_14198 (new_n9244_, not_new_n621__2326305139872070, not_new_n8851__0);
  not g_14199 (not_new_n734__0, new_n734_);
  or g_14200 (new_n1979_, not_pi109, not_new_n588__70);
  not g_14201 (not_new_n3011_, new_n3011_);
  not g_14202 (not_new_n618__10, new_n618_);
  not g_14203 (not_new_n617__138412872010, new_n617_);
  and g_14204 (and_and_not_pi048_2_not_pi047_2_not_pi050_2, not_pi050_2, and_not_pi048_2_not_pi047_2);
  not g_14205 (new_n5803_, new_n1069_);
  or g_14206 (new_n2535_, not_new_n605__2, not_new_n5486_);
  not g_14207 (not_new_n9013__0, new_n9013_);
  or g_14208 (new_n5911_, not_new_n5899__0, not_new_n5898_);
  or g_14209 (new_n4466_, not_new_n4693_, not_new_n4694_);
  not g_14210 (not_new_n7445__1, new_n7445_);
  or g_14211 (new_n2753_, not_pi248_0, not_po296_21838143759917965991093122527538323430);
  not g_14212 (not_new_n1368_, new_n1368_);
  not g_14213 (not_new_n3474_, new_n3474_);
  and g_14214 (new_n7080_, new_n7214_, new_n7319_);
  or g_14215 (new_n3852_, not_new_n621__490, not_new_n1576__70);
  not g_14216 (not_new_n775__332329305696010, new_n775_);
  or g_14217 (new_n8502_, not_new_n8380_, not_new_n8501_);
  or g_14218 (or_not_new_n1307__not_new_n1305_, not_new_n1305_, not_new_n1307_);
  not g_14219 (not_new_n3737_, new_n3737_);
  not g_14220 (not_new_n8246_, new_n8246_);
  or g_14221 (new_n10161_, not_new_n621__39098210485829880490, not_new_n1598__16284135979104490);
  or g_14222 (new_n3718_, not_new_n1607__3, not_new_n619__5);
  not g_14223 (not_new_n6299_, new_n6299_);
  or g_14224 (new_n5365_, not_new_n4955__0, not_new_n625__168070);
  or g_14225 (new_n6009_, not_new_n5804_, not_new_n622__168070);
  not g_14226 (not_new_n1537__19773267430, new_n1537_);
  not g_14227 (new_n9876_, new_n1045_);
  not g_14228 (not_new_n1296_, new_n1296_);
  not g_14229 (not_new_n2643_, new_n2643_);
  or g_14230 (new_n10174_, not_new_n1604__16284135979104490, not_new_n640__16284135979104490);
  not g_14231 (not_new_n4999__1, new_n4999_);
  xnor g_14232 (key_gate_107, not_new_n1660_, key_107);
  not g_14233 (not_new_n1031__8, new_n1031_);
  not g_14234 (not_new_n1782_, new_n1782_);
  not g_14235 (not_new_n5663_, new_n5663_);
  not g_14236 (not_new_n629__47475615099430, new_n629_);
  not g_14237 (not_new_n1616__968890104070, new_n1616_);
  not g_14238 (not_new_n8043_, new_n8043_);
  or g_14239 (new_n9164_, not_new_n9147_, not_new_n8983__0);
  or g_14240 (new_n10090_, not_new_n10038_, not_new_n9857_);
  not g_14241 (not_new_n6238_, new_n6238_);
  or g_14242 (po206, or_or_not_new_n1563__not_new_n2474__not_new_n1395_, not_new_n1396_);
  xor g_14243 (key_gate_44, key_44, new_n1634_);
  not g_14244 (not_new_n1512_, new_n1512_);
  not g_14245 (not_new_n6443__3430, new_n6443_);
  or g_14246 (new_n6790_, not_new_n6724_, not_new_n6722_);
  or g_14247 (new_n2463_, not_new_n600__19773267430, not_new_n4125__0);
  not g_14248 (new_n3404_, new_n1032_);
  and g_14249 (and_and_new_n2086__new_n2089__new_n2087_, new_n2087_, and_new_n2086__new_n2089_);
  not g_14250 (not_new_n9478_, new_n9478_);
  not g_14251 (not_new_n7778_, new_n7778_);
  not g_14252 (not_new_n3123_, new_n3123_);
  or g_14253 (new_n6542_, not_new_n6741_, not_new_n6795_);
  not g_14254 (not_new_n2644_, new_n2644_);
  not g_14255 (not_new_n4240_, new_n4240_);
  and g_14256 (new_n1562_, new_n3636_, new_n3637_);
  not g_14257 (new_n5209_, new_n4994_);
  or g_14258 (new_n3306_, not_new_n1583__113988951853731430, not_new_n7591__0);
  and g_14259 (new_n5845_, new_n5920_, new_n6106_);
  not g_14260 (not_new_n631__13410686196639649008070, new_n631_);
  not g_14261 (not_new_n9900__0, new_n9900_);
  not g_14262 (not_new_n1039__8235430, new_n1039_);
  not g_14263 (not_new_n9005_, new_n9005_);
  not g_14264 (not_new_n2810_, new_n2810_);
  not g_14265 (not_new_n3290_, new_n3290_);
  not g_14266 (new_n7776_, new_n7632_);
  not g_14267 (not_pi078, pi078);
  or g_14268 (or_pi033_pi035, pi035, pi033);
  or g_14269 (new_n696_, not_new_n1520_, not_new_n3060_);
  not g_14270 (not_new_n1581__5, new_n1581_);
  not g_14271 (not_new_n9436_, new_n9436_);
  not g_14272 (not_new_n4913_, new_n4913_);
  or g_14273 (new_n4671_, not_new_n4670_, not_new_n4669_);
  not g_14274 (not_new_n4155_, new_n4155_);
  or g_14275 (new_n7376_, not_new_n7363__0, not_new_n738__1);
  not g_14276 (not_new_n994__138412872010, new_n994_);
  not g_14277 (not_new_n10148_, new_n10148_);
  not g_14278 (not_new_n7018__1, new_n7018_);
  not g_14279 (not_new_n1049__3, new_n1049_);
  not g_14280 (not_new_n6621_, new_n6621_);
  not g_14281 (not_new_n5114_, new_n5114_);
  or g_14282 (new_n9650_, not_new_n9649_, not_new_n9802_);
  not g_14283 (not_new_n3556_, new_n3556_);
  or g_14284 (new_n9834_, not_new_n9398__0, not_new_n1061__2326305139872070);
  or g_14285 (or_not_new_n1596__403536070_not_new_n7586_, not_new_n7586_, not_new_n1596__403536070);
  not g_14286 (not_new_n7749_, new_n7749_);
  not g_14287 (not_new_n5057_, new_n5057_);
  or g_14288 (or_or_not_new_n6226__0_not_new_n6336__not_new_n6373__5, or_not_new_n6226__0_not_new_n6336_, not_new_n6373__5);
  not g_14289 (not_new_n1591__47475615099430, new_n1591_);
  not g_14290 (not_new_n5791__1, new_n5791_);
  not g_14291 (not_new_n602__138412872010, new_n602_);
  not g_14292 (not_new_n642__19773267430, new_n642_);
  not g_14293 (not_new_n1409_, new_n1409_);
  or g_14294 (new_n3436_, not_new_n1613__5, not_new_n1900_);
  not g_14295 (not_new_n5656_, new_n5656_);
  not g_14296 (not_new_n6661_, new_n6661_);
  not g_14297 (not_new_n594__8235430, new_n594_);
  not g_14298 (not_new_n621__5585458640832840070, new_n621_);
  not g_14299 (new_n7602_, new_n1047_);
  and g_14300 (new_n1214_, new_n1771_, new_n1772_);
  not g_14301 (not_new_n3300_, new_n3300_);
  not g_14302 (not_new_n6593_, new_n6593_);
  or g_14303 (new_n3485_, not_new_n1537__168070, not_pi113_0);
  or g_14304 (new_n6398_, not_new_n647__8235430, not_new_n6285_);
  not g_14305 (not_new_n628__4, new_n628_);
  not g_14306 (not_new_n8420_, new_n8420_);
  or g_14307 (new_n8785_, not_new_n8653__0, not_new_n1606__7);
  not g_14308 (new_n6974_, new_n775_);
  or g_14309 (new_n6138_, not_new_n6136_, not_new_n6137_);
  not g_14310 (not_new_n9670_, new_n9670_);
  not g_14311 (not_new_n4761__0, new_n4761_);
  and g_14312 (new_n1268_, new_n1974_, and_and_new_n1972__new_n1975__new_n1973_);
  not g_14313 (new_n4960_, new_n1053_);
  or g_14314 (new_n2341_, not_pi128, not_new_n588__797922662976120010);
  not g_14315 (new_n8881_, new_n1065_);
  not g_14316 (not_new_n1594__0, new_n1594_);
  or g_14317 (new_n8122_, not_new_n8305_, not_new_n8303_);
  not g_14318 (not_new_n9871_, new_n9871_);
  not g_14319 (not_new_n1611__6, new_n1611_);
  not g_14320 (not_new_n6272_, new_n6272_);
  not g_14321 (not_new_n2076_, new_n2076_);
  or g_14322 (new_n6641_, not_new_n6530_, not_new_n6815_);
  or g_14323 (new_n10325_, not_new_n10323_, not_new_n10324_);
  or g_14324 (new_n5868_, not_new_n6180_, not_new_n6181_);
  or g_14325 (new_n7846_, not_new_n1071__168070, not_new_n7635_);
  or g_14326 (new_n5057_, not_new_n5136_, not_new_n5124_);
  and g_14327 (new_n5838_, new_n5931_, new_n5932_);
  or g_14328 (new_n8341_, not_new_n8160_, not_new_n1057__403536070);
  not g_14329 (not_new_n7142_, new_n7142_);
  or g_14330 (new_n8723_, not_new_n1063__403536070, not_new_n8640_);
  or g_14331 (new_n5409_, not_new_n5407_, not_new_n5160_);
  or g_14332 (new_n5665_, not_new_n5575_, not_new_n5663_);
  not g_14333 (not_new_n1027__9, new_n1027_);
  or g_14334 (new_n4121_, not_new_n4194_, not_new_n4193_);
  not g_14335 (not_new_n624__8, new_n624_);
  not g_14336 (not_new_n5750_, new_n5750_);
  not g_14337 (not_new_n7876_, new_n7876_);
  not g_14338 (not_new_n5037_, new_n5037_);
  or g_14339 (new_n8180_, not_new_n8502_, not_new_n8503_);
  not g_14340 (not_new_n5336_, new_n5336_);
  and g_14341 (new_n1419_, new_n1418_, and_new_n2521__new_n2520_);
  not g_14342 (new_n4245_, new_n702_);
  or g_14343 (or_not_new_n6780__not_new_n6662_, not_new_n6780_, not_new_n6662_);
  not g_14344 (not_new_n6046_, new_n6046_);
  or g_14345 (new_n5184_, not_new_n1603__8, not_new_n639__3430);
  not g_14346 (not_new_n1585__2824752490, new_n1585_);
  or g_14347 (or_not_new_n6073__not_new_n6048_, not_new_n6048_, not_new_n6073_);
  not g_14348 (not_new_n2967_, new_n2967_);
  or g_14349 (new_n10337_, not_new_n10335_, not_new_n10336_);
  or g_14350 (new_n6098_, not_new_n648__8235430, not_new_n5746__1);
  not g_14351 (not_new_n723__0, new_n723_);
  not g_14352 (not_new_n1014__6, new_n1014_);
  or g_14353 (new_n3010_, not_new_n620__0, not_new_n3372__10);
  not g_14354 (new_n7005_, new_n726_);
  not g_14355 (not_new_n3850_, new_n3850_);
  or g_14356 (new_n2162_, not_new_n9870_, not_new_n594__403536070);
  not g_14357 (new_n4434_, new_n1019_);
  or g_14358 (new_n5066_, not_new_n5194_, not_new_n5195_);
  not g_14359 (not_new_n6173_, new_n6173_);
  not g_14360 (new_n4433_, pi171);
  not g_14361 (new_n8840_, new_n1049_);
  or g_14362 (new_n2675_, not_new_n5483_, not_new_n605__1176490);
  not g_14363 (not_new_n3318__0, new_n3318_);
  not g_14364 (not_new_n4317_, new_n4317_);
  not g_14365 (not_new_n9138_, new_n9138_);
  not g_14366 (not_new_n6059_, new_n6059_);
  or g_14367 (new_n6150_, not_new_n6149_, not_new_n6066_);
  or g_14368 (po064, key_gate_98, not_new_n1191_);
  or g_14369 (new_n2900_, or_not_new_n2899__not_new_n2898_, not_new_n2897_);
  not g_14370 (new_n1933_, new_n951_);
  or g_14371 (new_n3037_, not_new_n630__4, not_new_n3372__403536070);
  not g_14372 (not_new_n1589__3430, new_n1589_);
  not g_14373 (not_new_n1580__47475615099430, new_n1580_);
  or g_14374 (new_n6053_, not_new_n5812_, not_new_n5725_);
  not g_14375 (not_new_n1150_, new_n1150_);
  not g_14376 (not_new_n6270_, new_n6270_);
  not g_14377 (not_new_n639__3430, new_n639_);
  or g_14378 (new_n3699_, not_po298_138412872010, not_new_n625__9);
  not g_14379 (not_new_n641__8, new_n641_);
  or g_14380 (new_n1629_, not_new_n1536__70, not_new_n1628_);
  not g_14381 (not_new_n6524__2, new_n6524_);
  not g_14382 (new_n8138_, new_n1602_);
  or g_14383 (new_n1707_, not_pi007_0, not_po296_6782230728490);
  or g_14384 (new_n3738_, not_new_n3736_, not_new_n3737_);
  or g_14385 (new_n6605_, not_new_n6927_, not_new_n6928_);
  not g_14386 (not_new_n1182_, key_gate_122);
  not g_14387 (not_new_n7883_, new_n7883_);
  not g_14388 (not_new_n1037__47475615099430, new_n1037_);
  and g_14389 (new_n9863_, new_n9857_, new_n10059_);
  not g_14390 (not_new_n4512_, new_n4512_);
  not g_14391 (not_new_n1071__3, new_n1071_);
  and g_14392 (new_n4910_, new_n4908_, new_n4903_);
  or g_14393 (po219, or_or_not_new_n2557__not_new_n2561__not_new_n1427_, not_new_n1426_);
  not g_14394 (not_new_n608__8, new_n608_);
  or g_14395 (new_n2211_, not_new_n7589_, not_new_n1583__138412872010);
  or g_14396 (po263, not_new_n3713_, not_new_n3712_);
  not g_14397 (not_new_n3800_, new_n3800_);
  or g_14398 (new_n7929_, not_new_n7585_, not_new_n7754__2);
  not g_14399 (new_n7119_, new_n762_);
  not g_14400 (not_new_n7632_, new_n7632_);
  not g_14401 (not_new_n3531_, new_n3531_);
  not g_14402 (new_n6286_, new_n1063_);
  not g_14403 (not_new_n1631__168070, key_gate_76);
  not g_14404 (not_new_n5290_, new_n5290_);
  or g_14405 (new_n5887_, not_new_n6083_, not_new_n5853_);
  not g_14406 (not_po296_19773267430, po296);
  or g_14407 (new_n4847_, not_new_n1037__7, not_new_n4846_);
  not g_14408 (new_n8619_, new_n1061_);
  not g_14409 (not_new_n617__9, new_n617_);
  not g_14410 (not_new_n645__6782230728490, new_n645_);
  or g_14411 (new_n9150_, not_new_n8954_, not_new_n9149_);
  not g_14412 (not_new_n5825_, new_n5825_);
  not g_14413 (not_new_n8983_, new_n8983_);
  or g_14414 (new_n1835_, not_new_n6468_, not_new_n1580__3);
  not g_14415 (not_new_n586__0, new_n586_);
  not g_14416 (not_new_n3184__9, new_n3184_);
  or g_14417 (new_n8054_, not_new_n7757_, not_new_n7887__0);
  not g_14418 (not_new_n1631__2326305139872070, key_gate_76);
  or g_14419 (new_n9361_, not_new_n9453_, not_new_n9522_);
  or g_14420 (new_n3837_, not_new_n624__70, not_new_n6443__4);
  not g_14421 (not_new_n775__10, new_n775_);
  not g_14422 (not_new_n1251_, new_n1251_);
  not g_14423 (not_new_n1016__2, new_n1016_);
  or g_14424 (po068, key_gate_105, not_new_n1195_);
  or g_14425 (new_n7914_, not_new_n7759__1, not_new_n7707_);
  not g_14426 (not_new_n3241_, new_n3241_);
  or g_14427 (new_n8165_, not_new_n643__47475615099430, not_new_n8151_);
  not g_14428 (not_new_n8183_, new_n8183_);
  or g_14429 (or_not_new_n6337__not_new_n6373__6, not_new_n6373__6, not_new_n6337_);
  or g_14430 (new_n2708_, not_new_n1572_, not_new_n1579_);
  not g_14431 (not_new_n4458__0, new_n4458_);
  not g_14432 (not_new_n8897_, new_n8897_);
  not g_14433 (not_new_n2168_, new_n2168_);
  not g_14434 (not_new_n7808_, new_n7808_);
  not g_14435 (not_pi195, pi195);
  not g_14436 (not_new_n6765_, new_n6765_);
  not g_14437 (not_new_n5182_, new_n5182_);
  not g_14438 (not_new_n2348__0, new_n2348_);
  not g_14439 (not_new_n8261_, new_n8261_);
  not g_14440 (not_new_n1538__16284135979104490, new_n1538_);
  and g_14441 (new_n584_, new_n1221_, new_n1226_);
  not g_14442 (not_new_n9029_, new_n9029_);
  or g_14443 (new_n3691_, not_po298_57648010, not_new_n646__9);
  not g_14444 (not_new_n6443__1176490, new_n6443_);
  not g_14445 (not_new_n9082_, new_n9082_);
  not g_14446 (not_new_n8340_, new_n8340_);
  not g_14447 (not_new_n4613_, new_n4613_);
  not g_14448 (not_pi045_1, pi045);
  not g_14449 (not_new_n645_, new_n645_);
  or g_14450 (new_n2061_, not_new_n9446_, not_new_n1584__24010);
  or g_14451 (new_n6625_, not_new_n6809_, not_new_n6585_);
  not g_14452 (not_new_n1612__70, new_n1612_);
  or g_14453 (new_n10126_, not_new_n639__5585458640832840070, not_new_n1603__2326305139872070);
  not g_14454 (new_n6870_, new_n6591_);
  not g_14455 (not_new_n626__657123623635342801395430, new_n626_);
  not g_14456 (not_new_n8174_, new_n8174_);
  and g_14457 (new_n1203_, new_n1698_, new_n1700_);
  or g_14458 (new_n8921_, not_new_n9321_, not_new_n9320_);
  or g_14459 (new_n7356_, not_new_n6974__5, not_new_n766_);
  not g_14460 (not_new_n3309_, new_n3309_);
  not g_14461 (not_new_n6235_, new_n6235_);
  not g_14462 (not_new_n9028__0, new_n9028_);
  not g_14463 (not_new_n6339_, new_n6339_);
  not g_14464 (not_new_n10046__0, new_n10046_);
  not g_14465 (not_new_n593__968890104070, new_n593_);
  not g_14466 (not_pi274_2, pi274);
  not g_14467 (not_new_n1429_, new_n1429_);
  not g_14468 (not_new_n1069__2824752490, new_n1069_);
  or g_14469 (new_n1944_, not_new_n601__7, not_new_n648__0);
  not g_14470 (not_new_n3315__16284135979104490, new_n3315_);
  and g_14471 (new_n1553_, new_n3619_, new_n3618_);
  not g_14472 (not_new_n5890_, new_n5890_);
  or g_14473 (or_not_new_n3152__not_new_n3151_, not_new_n3152_, not_new_n3151_);
  or g_14474 (new_n6167_, not_new_n5776__0, not_new_n639__8235430);
  or g_14475 (new_n4051_, not_pi037_3, not_new_n3939_);
  not g_14476 (not_new_n2789_, new_n2789_);
  not g_14477 (not_new_n4764_, new_n4764_);
  not g_14478 (not_new_n1536__5, new_n1536_);
  not g_14479 (not_new_n1041__19773267430, new_n1041_);
  or g_14480 (new_n5253_, not_new_n5251_, not_new_n5055_);
  or g_14481 (new_n2242_, not_new_n2237_, not_new_n1324_);
  or g_14482 (new_n2973_, not_new_n613__7, not_new_n1597__1);
  and g_14483 (new_n1317_, new_n2212_, new_n2213_);
  not g_14484 (not_new_n4402_, new_n4402_);
  or g_14485 (po207, or_or_not_new_n1564__not_new_n2479__not_new_n1397_, not_new_n1398_);
  not g_14486 (new_n5163_, new_n5075_);
  or g_14487 (new_n8166_, not_new_n8349_, not_new_n8351_);
  not g_14488 (not_new_n6718_, new_n6718_);
  not g_14489 (not_pi140, pi140);
  and g_14490 (new_n5046_, new_n5214_, new_n5079_);
  not g_14491 (new_n4087_, pi246);
  or g_14492 (new_n3386_, not_pi064_16284135979104490, not_new_n3992__0);
  or g_14493 (new_n2329_, not_new_n1584__16284135979104490, not_new_n9436_);
  not g_14494 (not_new_n1631__16284135979104490, key_gate_76);
  not g_14495 (not_new_n9768_, new_n9768_);
  not g_14496 (not_pi272_2, pi272);
  not g_14497 (not_new_n1176__0, new_n1176_);
  not g_14498 (new_n6499_, new_n622_);
  or g_14499 (new_n3179_, not_new_n1593_, not_new_n1530_);
  or g_14500 (new_n10166_, not_new_n9860_, not_new_n9950_);
  not g_14501 (not_new_n8722_, new_n8722_);
  not g_14502 (not_new_n8135_, new_n8135_);
  or g_14503 (new_n10141_, not_new_n9862_, not_new_n10037_);
  not g_14504 (not_new_n612__0, new_n612_);
  not g_14505 (not_new_n5742__1, new_n5742_);
  not g_14506 (not_pi269_0, pi269);
  not g_14507 (not_new_n1982_, new_n1982_);
  not g_14508 (not_new_n9199_, new_n9199_);
  or g_14509 (new_n8467_, not_new_n8466_, not_new_n8465_);
  not g_14510 (not_new_n1057__70, new_n1057_);
  not g_14511 (not_new_n4801_, new_n4801_);
  not g_14512 (not_new_n984__2824752490, new_n984_);
  not g_14513 (new_n9107_, new_n8961_);
  and g_14514 (new_n4806_, new_n4893_, new_n4892_);
  not g_14515 (not_new_n8521_, new_n8521_);
  not g_14516 (not_new_n8123_, new_n8123_);
  and g_14517 (new_n6240_, and_and_new_n6395__new_n6396__new_n6228_, new_n6397_);
  not g_14518 (not_new_n1063__5, new_n1063_);
  not g_14519 (not_new_n3296_, new_n3296_);
  not g_14520 (not_new_n9387__0, new_n9387_);
  or g_14521 (new_n3559_, not_new_n1612__168070, not_new_n2090__0);
  or g_14522 (new_n1535_, not_new_n590__2, not_new_n927_);
  not g_14523 (not_new_n589__6782230728490, new_n589_);
  not g_14524 (not_new_n7028__0, new_n7028_);
  not g_14525 (not_new_n638__5, new_n638_);
  not g_14526 (not_new_n6498__0, new_n6498_);
  not g_14527 (not_new_n1024__1, new_n1024_);
  or g_14528 (new_n7263_, not_new_n7406_, not_new_n7014_);
  not g_14529 (not_pi064_2326305139872070, pi064);
  or g_14530 (new_n4527_, not_new_n4526_, not_new_n4481_);
  or g_14531 (new_n692_, not_new_n3044_, not_new_n1514_);
  not g_14532 (new_n7617_, new_n647_);
  and g_14533 (and_new_n2508__new_n2510_, new_n2510_, new_n2508_);
  not g_14534 (not_new_n8150_, new_n8150_);
  or g_14535 (new_n649_, not_new_n3104_, not_new_n3105_);
  not g_14536 (not_new_n1059__403536070, new_n1059_);
  or g_14537 (or_not_new_n1901__not_new_n1902_, not_new_n1902_, not_new_n1901_);
  not g_14538 (new_n3978_, pi037);
  or g_14539 (or_not_new_n2971__not_new_n2970_, not_new_n2970_, not_new_n2971_);
  not g_14540 (not_pi146_3, pi146);
  and g_14541 (new_n8223_, new_n8284_, new_n8506_);
  not g_14542 (not_new_n1537_, new_n1537_);
  not g_14543 (not_new_n3739_, new_n3739_);
  or g_14544 (new_n2731_, not_pi246_0, not_po296_445676403263631959001900459745680070);
  not g_14545 (not_new_n8419_, new_n8419_);
  not g_14546 (not_new_n6527_, new_n6527_);
  or g_14547 (new_n5217_, not_new_n5073_, not_new_n5186_);
  not g_14548 (new_n6919_, new_n6603_);
  not g_14549 (not_new_n8453_, new_n8453_);
  not g_14550 (not_new_n9101_, new_n9101_);
  and g_14551 (and_new_n3780__new_n3783_, new_n3780_, new_n3783_);
  or g_14552 (new_n1157_, not_new_n3843_, not_new_n3844_);
  not g_14553 (not_new_n5368_, new_n5368_);
  or g_14554 (new_n9448_, not_new_n9843_, not_new_n9844_);
  or g_14555 (new_n1883_, not_new_n587__6, not_pi136);
  or g_14556 (new_n3831_, not_new_n6443__1, not_new_n634__70);
  not g_14557 (not_new_n3930_, key_gate_43);
  not g_14558 (not_new_n9878_, new_n9878_);
  or g_14559 (new_n7830_, not_new_n1059__8235430, not_new_n7645_);
  not g_14560 (not_new_n3195_, new_n3195_);
  and g_14561 (new_n6587_, new_n6748_, new_n6747_);
  not g_14562 (not_new_n8189_, new_n8189_);
  not g_14563 (not_new_n603__0, new_n603_);
  not g_14564 (not_new_n5952_, new_n5952_);
  or g_14565 (new_n7192_, not_new_n7321_, not_new_n6977__0);
  not g_14566 (not_new_n5084__1, new_n5084_);
  not g_14567 (not_new_n589__152867006319425761937651857692768264010, new_n589_);
  not g_14568 (not_new_n8518_, new_n8518_);
  not g_14569 (not_new_n9614_, new_n9614_);
  and g_14570 (and_new_n1286__new_n2065_, new_n2065_, new_n1286_);
  not g_14571 (not_new_n732_, new_n732_);
  not g_14572 (not_new_n8155__2, new_n8155_);
  not g_14573 (not_new_n594__16284135979104490, new_n594_);
  or g_14574 (new_n3783_, not_new_n3782_, not_new_n3781_);
  not g_14575 (not_new_n7612_, new_n7612_);
  not g_14576 (not_new_n625__9, new_n625_);
  not g_14577 (not_new_n9769_, new_n9769_);
  or g_14578 (new_n4945_, not_new_n5027_, not_new_n5026_);
  not g_14579 (not_new_n4309_, new_n4309_);
  not g_14580 (not_new_n1565_, new_n1565_);
  not g_14581 (not_new_n7333_, new_n7333_);
  or g_14582 (new_n6388_, not_new_n6387_, not_new_n6312_);
  or g_14583 (new_n5219_, not_new_n4904_, not_new_n4998_);
  not g_14584 (not_new_n4845_, new_n4845_);
  not g_14585 (not_new_n6974__8, new_n6974_);
  not g_14586 (not_new_n624__0, new_n624_);
  not g_14587 (new_n3479_, new_n1063_);
  not g_14588 (not_new_n5906_, new_n5906_);
  not g_14589 (not_new_n8596_, new_n8596_);
  or g_14590 (new_n6117_, not_new_n5749__2, not_new_n1039__3430);
  or g_14591 (new_n3456_, not_new_n1613__9, not_new_n1976_);
  or g_14592 (new_n3327_, not_new_n1534__5, not_pi041_0);
  and g_14593 (new_n5725_, new_n6002_, new_n5718_);
  or g_14594 (new_n631_, or_or_not_new_n1844__not_new_n1845__not_new_n1847_, not_new_n1846_);
  or g_14595 (or_not_new_n7715__not_new_n7714_, not_new_n7715_, not_new_n7714_);
  not g_14596 (not_new_n1616__4, new_n1616_);
  not g_14597 (not_new_n5786__1, new_n5786_);
  not g_14598 (not_new_n5792__0, new_n5792_);
  or g_14599 (new_n984_, not_new_n2351_, not_new_n590_);
  not g_14600 (not_new_n7212__0, new_n7212_);
  not g_14601 (not_new_n6634__0, new_n6634_);
  not g_14602 (not_new_n6071_, new_n6071_);
  or g_14603 (new_n2465_, not_new_n598__19773267430, not_new_n1602__0);
  not g_14604 (not_new_n1631__3, key_gate_76);
  and g_14605 (and_new_n2513__new_n2512_, new_n2513_, new_n2512_);
  not g_14606 (not_new_n636__8, new_n636_);
  not g_14607 (not_new_n618__2824752490, new_n618_);
  or g_14608 (new_n8515_, not_new_n8130__0, not_new_n1599__8235430);
  or g_14609 (new_n4625_, not_pi165_3, not_new_n4422__0);
  not g_14610 (not_new_n6642_, new_n6642_);
  not g_14611 (not_new_n6145_, new_n6145_);
  not g_14612 (not_new_n2018_, new_n2018_);
  not g_14613 (not_new_n7131_, new_n7131_);
  not g_14614 (not_new_n6177_, new_n6177_);
  and g_14615 (and_and_new_n2200__new_n2203__new_n2201_, new_n2201_, and_new_n2200__new_n2203_);
  not g_14616 (not_new_n10249_, new_n10249_);
  and g_14617 (new_n1392_, new_n2465_, new_n2466_);
  or g_14618 (new_n7770_, not_new_n1602__1176490, not_new_n7628_);
  not g_14619 (not_new_n5640_, new_n5640_);
  not g_14620 (not_new_n4593_, new_n4593_);
  not g_14621 (not_new_n4237_, new_n4237_);
  or g_14622 (po278, not_new_n2829_, or_or_not_new_n2831__not_new_n1481__not_new_n2830_);
  and g_14623 (new_n1441_, and_new_n2632__new_n2631_, new_n2630_);
  not g_14624 (not_new_n595__2824752490, new_n595_);
  or g_14625 (new_n4971_, not_new_n5274_, not_new_n5161_);
  not g_14626 (not_new_n1598__2326305139872070, new_n1598_);
  not g_14627 (not_new_n10245_, new_n10245_);
  and g_14628 (and_new_n3306__new_n3305_, new_n3305_, new_n3306_);
  not g_14629 (not_new_n694_, new_n694_);
  not g_14630 (not_new_n619__1, new_n619_);
  not g_14631 (not_new_n5566_, new_n5566_);
  not g_14632 (not_new_n2749_, new_n2749_);
  or g_14633 (new_n5092_, new_n1037_, new_n632_);
  or g_14634 (new_n2067_, not_new_n9970_, not_new_n594__24010);
  not g_14635 (not_new_n3562_, new_n3562_);
  not g_14636 (not_new_n4939_, new_n4939_);
  and g_14637 (new_n1423_, new_n2542_, new_n2540_);
  or g_14638 (new_n2443_, not_new_n4129__0, not_new_n600__8235430);
  or g_14639 (new_n3084_, not_new_n1180_, not_new_n1027__1915812313805664144010);
  or g_14640 (new_n3425_, not_new_n1537__3, not_pi101_0);
  not g_14641 (not_new_n2794_, new_n2794_);
  not g_14642 (not_new_n4381_, new_n4381_);
  not g_14643 (not_pi260_2, pi260);
  not g_14644 (not_new_n636__5, new_n636_);
  or g_14645 (or_not_new_n1339__not_new_n1337_, not_new_n1337_, not_new_n1339_);
  not g_14646 (not_new_n581__6168735096280623662907561568153897267931784070, new_n581_);
  or g_14647 (new_n10119_, new_n1603_, new_n639_);
  or g_14648 (new_n7923_, not_new_n7846_, not_new_n7754_);
  or g_14649 (new_n6899_, not_new_n6504__0, not_new_n1602__168070);
  not g_14650 (not_pi179, pi179);
  not g_14651 (not_new_n5095__0, new_n5095_);
  or g_14652 (or_not_new_n4240__not_new_n4343_, not_new_n4240_, not_new_n4343_);
  not g_14653 (new_n7598_, new_n648_);
  or g_14654 (new_n6106_, not_new_n6104_, not_new_n6105_);
  not g_14655 (new_n4168_, new_n4098_);
  or g_14656 (new_n7189_, not_new_n7366__0, not_new_n6976__0);
  and g_14657 (new_n1361_, and_new_n2389__new_n2388_, new_n2387_);
  not g_14658 (not_new_n7896_, new_n7896_);
  not g_14659 (not_new_n7724_, new_n7724_);
  not g_14660 (not_new_n602__8235430, new_n602_);
  and g_14661 (new_n6347_, new_n6236_, and_and_and_new_n1053__new_n6232__new_n6395__new_n6317_);
  not g_14662 (not_new_n7670_, new_n7670_);
  or g_14663 (new_n743_, not_new_n3278_, not_new_n3277_);
  or g_14664 (new_n4540_, not_new_n1003__2, not_pi169_1);
  not g_14665 (not_new_n8850_, new_n8850_);
  not g_14666 (not_new_n7649__0, new_n7649_);
  not g_14667 (not_new_n9099__0, new_n9099_);
  or g_14668 (new_n9439_, not_new_n9778_, not_new_n9777_);
  not g_14669 (not_new_n4426_, new_n4426_);
  not g_14670 (not_new_n3245_, new_n3245_);
  not g_14671 (not_new_n8113_, new_n8113_);
  not g_14672 (not_new_n9956__0, new_n9956_);
  not g_14673 (not_new_n3101_, new_n3101_);
  or g_14674 (or_not_new_n6353__not_new_n6232__5, not_new_n6232__5, not_new_n6353_);
  not g_14675 (new_n6280_, new_n629_);
  not g_14676 (not_new_n9557_, new_n9557_);
  not g_14677 (not_new_n8106__0, new_n8106_);
  not g_14678 (not_new_n4612_, new_n4612_);
  or g_14679 (new_n4002_, not_new_n3937_, not_new_n4001__1);
  not g_14680 (not_new_n5884__0, new_n5884_);
  not g_14681 (not_po296_2, po296);
  not g_14682 (not_new_n6528_, new_n6528_);
  not g_14683 (not_new_n10171_, new_n10171_);
  not g_14684 (not_new_n2543_, new_n2543_);
  not g_14685 (not_new_n8348_, new_n8348_);
  not g_14686 (not_new_n10046_, new_n10046_);
  not g_14687 (not_new_n632__332329305696010, new_n632_);
  not g_14688 (new_n8624_, new_n1170_);
  not g_14689 (not_new_n4163__1, new_n4163_);
  not g_14690 (not_new_n1602__24010, new_n1602_);
  not g_14691 (not_new_n3471_, new_n3471_);
  not g_14692 (not_new_n595__2, new_n595_);
  or g_14693 (new_n8977_, not_new_n9059_, not_new_n9058_);
  not g_14694 (not_new_n5444__0, new_n5444_);
  or g_14695 (or_or_not_new_n1263__not_new_n1261__not_new_n1945_, or_not_new_n1263__not_new_n1261_, not_new_n1945_);
  or g_14696 (new_n3214_, not_new_n1603__4, not_new_n3185__3430);
  not g_14697 (not_new_n7138__0, new_n7138_);
  not g_14698 (not_new_n8265__2, new_n8265_);
  not g_14699 (not_new_n10154_, new_n10154_);
  not g_14700 (not_new_n6660_, new_n6660_);
  not g_14701 (not_new_n1381_, new_n1381_);
  not g_14702 (not_new_n633__3430, new_n633_);
  not g_14703 (not_new_n647__3, new_n647_);
  not g_14704 (not_new_n5959_, new_n5959_);
  not g_14705 (not_new_n1061__9, new_n1061_);
  not g_14706 (not_new_n8441_, new_n8441_);
  or g_14707 (new_n6003_, not_new_n5770__0, not_new_n1601__490);
  or g_14708 (new_n5740_, not_new_n5745_, not_new_n634__1176490);
  not g_14709 (not_new_n7044__0, new_n7044_);
  not g_14710 (not_new_n775__403536070, new_n775_);
  not g_14711 (not_new_n6030_, new_n6030_);
  not g_14712 (not_new_n604__6782230728490, new_n604_);
  not g_14713 (not_new_n7164_, new_n7164_);
  not g_14714 (not_new_n7856_, new_n7856_);
  not g_14715 (not_new_n4992__0, new_n4992_);
  not g_14716 (not_new_n7148_, new_n7148_);
  not g_14717 (not_new_n5393_, new_n5393_);
  or g_14718 (new_n3765_, not_new_n3764_, not_new_n3763_);
  not g_14719 (new_n4280_, new_n652_);
  not g_14720 (new_n9912_, new_n1065_);
  not g_14721 (not_new_n9584_, new_n9584_);
  not g_14722 (not_pi090, pi090);
  not g_14723 (not_pi175_3, pi175);
  not g_14724 (new_n10055_, new_n9879_);
  not g_14725 (new_n4975_, new_n1604_);
  or g_14726 (new_n1975_, not_new_n1588__10, not_new_n1053__0);
  or g_14727 (new_n9631_, new_n617_, new_n1597_);
  not g_14728 (not_new_n7132_, new_n7132_);
  and g_14729 (and_new_n8828__new_n9210_, new_n9210_, new_n8828_);
  not g_14730 (not_new_n8058_, new_n8058_);
  not g_14731 (new_n6536_, new_n1069_);
  or g_14732 (new_n9297_, not_new_n8858_, not_new_n1063__19773267430);
  not g_14733 (not_new_n1613__57648010, new_n1613_);
  not g_14734 (not_new_n647__2326305139872070, new_n647_);
  and g_14735 (new_n1428_, new_n2569_, new_n2568_);
  or g_14736 (new_n2330_, not_new_n1581__16284135979104490, not_new_n8098_);
  not g_14737 (not_new_n6350_, new_n6350_);
  not g_14738 (not_new_n1006__1, new_n1006_);
  not g_14739 (not_pi184, pi184);
  not g_14740 (not_new_n1007__6, new_n1007_);
  not g_14741 (not_new_n1063__16284135979104490, new_n1063_);
  not g_14742 (not_new_n6195_, new_n6195_);
  not g_14743 (not_new_n8344_, new_n8344_);
  not g_14744 (not_new_n3882_, new_n3882_);
  not g_14745 (new_n10184_, new_n9952_);
  not g_14746 (not_new_n9433_, new_n9433_);
  not g_14747 (not_new_n4677_, new_n4677_);
  or g_14748 (new_n3756_, not_new_n3754_, not_new_n3755_);
  or g_14749 (new_n4679_, not_new_n4497_, not_new_n4498__0);
  or g_14750 (new_n8726_, not_new_n8636_, not_new_n1051__403536070);
  or g_14751 (new_n9249_, not_new_n9159_, not_new_n8894__0);
  not g_14752 (new_n4513_, new_n4487_);
  or g_14753 (new_n3685_, not_po298_168070, not_new_n638__9);
  not g_14754 (not_pi223, pi223);
  not g_14755 (not_new_n940__0, new_n940_);
  or g_14756 (new_n6183_, not_new_n6182_, not_new_n6088_);
  or g_14757 (new_n4210_, not_new_n4093_, not_new_n4165__0);
  or g_14758 (new_n6166_, not_new_n5772__0, not_new_n1603__490);
  or g_14759 (new_n4068_, not_new_n4016__0, not_new_n3995__0);
  or g_14760 (new_n8366_, not_new_n8081_, not_new_n8289_);
  not g_14761 (not_new_n586__113988951853731430, new_n586_);
  not g_14762 (not_new_n4119__1, new_n4119_);
  not g_14763 (not_new_n4816__0, new_n4816_);
  not g_14764 (not_pi161, pi161);
  not g_14765 (not_new_n5599_, new_n5599_);
  or g_14766 (new_n640_, or_or_not_new_n2129__not_new_n2130__not_new_n2132_, not_new_n2131_);
  and g_14767 (new_n4761_, new_n4857_, new_n4856_);
  not g_14768 (not_new_n1061__138412872010, new_n1061_);
  not g_14769 (not_new_n1045__332329305696010, new_n1045_);
  or g_14770 (new_n6902_, not_new_n6755_, not_new_n6628_);
  not g_14771 (not_new_n3184__168070, new_n3184_);
  or g_14772 (or_not_new_n4816__not_new_n4751_, not_new_n4751_, not_new_n4816_);
  or g_14773 (new_n5811_, not_new_n5864_, not_new_n6063_);
  or g_14774 (new_n4988_, not_new_n5040_, not_new_n5282_);
  or g_14775 (new_n5265_, not_new_n5156__0, not_new_n4966__0);
  not g_14776 (not_new_n7578_, new_n7578_);
  or g_14777 (new_n3112_, not_new_n619__3, not_new_n581__1577753820348458066150427430);
  or g_14778 (new_n6667_, not_new_n628__2824752490, not_new_n6648_);
  not g_14779 (not_new_n4987_, new_n4987_);
  not g_14780 (not_new_n2526_, new_n2526_);
  not g_14781 (not_new_n2245_, new_n2245_);
  not g_14782 (not_new_n7479_, new_n7479_);
  and g_14783 (and_and_new_n2162__new_n2165__new_n2163_, and_new_n2162__new_n2165_, new_n2163_);
  not g_14784 (not_new_n6976_, new_n6976_);
  or g_14785 (new_n10284_, not_new_n1597__39098210485829880490, not_new_n9944__0);
  not g_14786 (not_new_n6446_, new_n6446_);
  or g_14787 (or_or_not_new_n2838__not_new_n2841__not_new_n2840_, not_new_n2840_, or_not_new_n2838__not_new_n2841_);
  not g_14788 (not_new_n1580__1, new_n1580_);
  not g_14789 (new_n6154_, new_n5861_);
  not g_14790 (not_new_n611__1176490, new_n611_);
  not g_14791 (not_new_n2741_, new_n2741_);
  or g_14792 (new_n6129_, or_not_new_n5764__0_not_new_n618__8235430, not_new_n6126_);
  or g_14793 (new_n7216_, not_new_n7152_, not_new_n7215_);
  not g_14794 (not_new_n1603__2824752490, new_n1603_);
  and g_14795 (new_n1245_, new_n1871_, new_n1870_);
  or g_14796 (new_n8059_, not_new_n7645__0, not_new_n1059__57648010);
  not g_14797 (not_new_n589__16284135979104490, new_n589_);
  not g_14798 (new_n6295_, new_n1053_);
  not g_14799 (not_new_n5621_, new_n5621_);
  not g_14800 (not_new_n2758_, new_n2758_);
  not g_14801 (not_new_n2161_, new_n2161_);
  or g_14802 (new_n4010_, not_new_n4009_, not_pi038_3);
  not g_14803 (new_n9923_, new_n636_);
  or g_14804 (or_or_not_new_n1473__not_new_n2722__not_new_n2723_, not_new_n2723_, or_not_new_n1473__not_new_n2722_);
  not g_14805 (new_n9380_, new_n1600_);
  and g_14806 (new_n3914_, new_n3964_, new_n3963_);
  or g_14807 (new_n1756_, not_pi070, not_new_n1728__6782230728490);
  not g_14808 (new_n1621_, new_n923_);
  not g_14809 (not_new_n607_, new_n607_);
  not g_14810 (not_new_n1065__57648010, new_n1065_);
  not g_14811 (not_new_n7645_, new_n7645_);
  not g_14812 (not_new_n8522_, new_n8522_);
  not g_14813 (not_new_n1063__19773267430, new_n1063_);
  not g_14814 (not_new_n3273_, new_n3273_);
  or g_14815 (po267, or_or_or_not_new_n2727__not_new_n2730__not_new_n2729__not_new_n2731_, not_new_n2728_);
  not g_14816 (not_new_n3767_, new_n3767_);
  not g_14817 (not_new_n617__2326305139872070, new_n617_);
  not g_14818 (not_new_n6010_, new_n6010_);
  not g_14819 (not_new_n5262_, new_n5262_);
  or g_14820 (new_n7793_, not_new_n7739_, not_new_n7577_);
  not g_14821 (not_new_n4340_, new_n4340_);
  or g_14822 (new_n4594_, not_new_n4429_, not_new_n1003__3);
  not g_14823 (not_pi073, pi073);
  or g_14824 (new_n7194_, not_new_n7192_, not_new_n7075_);
  not g_14825 (new_n6976_, new_n739_);
  not g_14826 (not_new_n594__1176490, new_n594_);
  and g_14827 (new_n1515_, new_n998_, new_n3045_);
  not g_14828 (not_new_n7662__0, new_n7662_);
  not g_14829 (new_n4423_, pi166);
  not g_14830 (not_new_n6761_, new_n6761_);
  not g_14831 (new_n7348_, new_n7027_);
  not g_14832 (not_new_n1581__8, new_n1581_);
  and g_14833 (new_n1525_, new_n3074_, and_new_n3076__new_n998_);
  not g_14834 (not_new_n6133_, new_n6133_);
  or g_14835 (new_n3795_, not_new_n3793_, not_new_n3794_);
  or g_14836 (new_n3291_, not_new_n589__445676403263631959001900459745680070, not_new_n1059__5);
  not g_14837 (not_new_n4118_, new_n4118_);
  not g_14838 (not_new_n8886_, new_n8886_);
  not g_14839 (not_new_n9554_, new_n9554_);
  not g_14840 (not_new_n10157_, new_n10157_);
  and g_14841 (new_n8092_, new_n8527_, new_n8176_);
  not g_14842 (not_new_n640__1176490, new_n640_);
  or g_14843 (new_n7405_, not_new_n6974__9, not_new_n747_);
  not g_14844 (not_new_n5056__0, new_n5056_);
  or g_14845 (new_n2949_, not_new_n595__968890104070, not_new_n7069_);
  not g_14846 (not_new_n3981_, new_n3981_);
  not g_14847 (not_new_n8595_, new_n8595_);
  not g_14848 (not_new_n7589_, new_n7589_);
  not g_14849 (not_new_n610__7, new_n610_);
  or g_14850 (new_n2992_, not_new_n3372__4, not_new_n647__4);
  or g_14851 (new_n1154_, not_new_n3838_, not_new_n3837_);
  and g_14852 (new_n8692_, new_n8764_, new_n8693_);
  not g_14853 (not_new_n6697_, new_n6697_);
  or g_14854 (new_n3648_, not_pi190_0, not_new_n984__16284135979104490);
  not g_14855 (not_new_n3982__0, new_n3982_);
  not g_14856 (not_new_n1067__7, new_n1067_);
  not g_14857 (not_new_n588__24010, new_n588_);
  not g_14858 (not_new_n1583__490, new_n1583_);
  not g_14859 (not_new_n1581__2824752490, new_n1581_);
  not g_14860 (new_n9359_, new_n1031_);
  not g_14861 (not_new_n7077_, new_n7077_);
  not g_14862 (not_new_n3340_, new_n3340_);
  not g_14863 (not_new_n3248_, new_n3248_);
  not g_14864 (not_new_n989__6, new_n989_);
  or g_14865 (new_n5488_, not_new_n5684_, not_new_n5683_);
  or g_14866 (new_n6855_, not_new_n6486__1, not_new_n628__138412872010);
  or g_14867 (new_n10341_, not_new_n1063__2326305139872070, not_new_n9918_);
  not g_14868 (not_new_n4072__0, new_n4072_);
  not g_14869 (not_new_n7481_, new_n7481_);
  not g_14870 (not_pi265_3, pi265);
  or g_14871 (new_n1805_, not_new_n1232_, not_new_n1800_);
  not g_14872 (not_new_n9585_, new_n9585_);
  or g_14873 (new_n1815_, not_new_n8194_, not_new_n1581__1);
  not g_14874 (not_new_n1977_, new_n1977_);
  or g_14875 (new_n2483_, not_new_n4121__0, not_new_n600__47475615099430);
  xnor g_14876 (key_gate_1, not_new_n1654_, key_1);
  not g_14877 (not_new_n8074_, new_n8074_);
  not g_14878 (new_n4242_, new_n670_);
  or g_14879 (new_n8457_, not_new_n8082__0, not_new_n8228_);
  not g_14880 (not_new_n589__225393402906922580878632490, new_n589_);
  or g_14881 (po241, not_new_n3668_, not_new_n3669_);
  not g_14882 (not_new_n586__9, new_n586_);
  not g_14883 (new_n8137_, new_n1601_);
  not g_14884 (not_new_n4669_, new_n4669_);
  and g_14885 (new_n4912_, new_n5253_, new_n5250_);
  and g_14886 (new_n1405_, and_new_n3306__new_n3305_, new_n3304_);
  or g_14887 (or_not_new_n1159__0_not_new_n8794__0, not_new_n8794__0, not_new_n1159__0);
  not g_14888 (not_new_n6613__3, new_n6613_);
  not g_14889 (new_n8251_, new_n619_);
  not g_14890 (not_new_n7489_, new_n7489_);
  not g_14891 (not_new_n6937_, new_n6937_);
  not g_14892 (not_new_n6540__1, new_n6540_);
  not g_14893 (not_new_n2348_, new_n2348_);
  or g_14894 (new_n7026_, not_new_n7343_, not_new_n7344_);
  not g_14895 (not_new_n10010_, new_n10010_);
  xor g_14896 (key_gate_84, key_84, not_new_n3917_);
  not g_14897 (not_pi034_2, pi034);
  or g_14898 (new_n9952_, not_new_n10183_, not_new_n9926_);
  or g_14899 (new_n5405_, not_new_n643__8235430, not_new_n4969__0);
  not g_14900 (not_new_n9477_, new_n9477_);
  or g_14901 (new_n7965_, not_new_n7599__2, not_new_n631__2326305139872070);
  not g_14902 (not_new_n4846_, new_n4846_);
  not g_14903 (not_new_n6906_, new_n6906_);
  or g_14904 (new_n4572_, not_new_n1013__2, not_pi177_1);
  not g_14905 (not_new_n731_, new_n731_);
  not g_14906 (not_new_n3929__0, key_gate_36);
  and g_14907 (and_new_n4405__new_n4330_, new_n4330_, new_n4405_);
  not g_14908 (new_n4004_, new_n3954_);
  or g_14909 (new_n2306_, not_new_n7674_, not_new_n1583__2326305139872070);
  not g_14910 (not_new_n10239_, new_n10239_);
  and g_14911 (new_n1184_, new_n1641_, new_n1643_);
  or g_14912 (new_n3949_, not_new_n3973_, not_new_n4032_);
  not g_14913 (not_new_n604__10, new_n604_);
  not g_14914 (not_new_n9606_, new_n9606_);
  or g_14915 (new_n7759_, or_not_new_n7939__not_new_n7913_, not_new_n7831_);
  or g_14916 (new_n3089_, not_new_n928__0, not_new_n1049__3);
  not g_14917 (not_new_n1398_, new_n1398_);
  not g_14918 (not_new_n4227_, new_n4227_);
  not g_14919 (not_new_n1208_, new_n1208_);
  not g_14920 (not_new_n4955_, new_n4955_);
  not g_14921 (not_new_n646__4, new_n646_);
  or g_14922 (new_n4100_, not_pi264_0, not_new_n4168_);
  or g_14923 (new_n3092_, not_new_n928__1, not_new_n1047__3);
  or g_14924 (new_n6415_, not_new_n1606__5, not_new_n6249_);
  or g_14925 (new_n5476_, not_new_n5595_, not_new_n5594_);
  or g_14926 (new_n6041_, not_new_n5751_, not_new_n641__3430);
  not g_14927 (not_new_n7648__2, new_n7648_);
  or g_14928 (new_n2871_, not_new_n602__168070, not_new_n621__2);
  not g_14929 (new_n6274_, new_n626_);
  or g_14930 (new_n952_, not_new_n1944_, or_or_not_new_n1263__not_new_n1261__not_new_n1945_);
  or g_14931 (new_n1755_, not_pi069, not_new_n1728__968890104070);
  not g_14932 (not_new_n6300_, new_n6300_);
  not g_14933 (new_n7013_, new_n719_);
  not g_14934 (not_new_n7930_, new_n7930_);
  not g_14935 (not_new_n3856_, new_n3856_);
  or g_14936 (po222, or_or_not_new_n2587__not_new_n2591__not_new_n1433_, not_new_n1432_);
  or g_14937 (new_n2246_, not_new_n4121_, not_new_n585__47475615099430);
  or g_14938 (new_n6872_, not_new_n6591_, not_new_n6622__0);
  not g_14939 (not_new_n622__70, new_n622_);
  or g_14940 (new_n8053_, not_new_n7671__0, not_new_n7895_);
  not g_14941 (new_n7622_, new_n1597_);
  not g_14942 (not_new_n4898__0, new_n4898_);
  not g_14943 (not_new_n8908_, new_n8908_);
  not g_14944 (not_new_n7113__2, new_n7113_);
  and g_14945 (new_n1346_, and_new_n1033__new_n3404_, new_n1592_);
  not g_14946 (not_new_n1027__968890104070, new_n1027_);
  or g_14947 (new_n9045_, not_new_n8801_, not_new_n8988_);
  not g_14948 (not_new_n6531__1, new_n6531_);
  not g_14949 (not_pi264_0, pi264);
  or g_14950 (new_n3005_, not_new_n581__5, not_new_n1041__2);
  and g_14951 (and_and_new_n2325__new_n2332__new_n2333_, new_n2333_, and_new_n2325__new_n2332_);
  not g_14952 (new_n7608_, new_n1031_);
  not g_14953 (not_new_n3383_, new_n3383_);
  not g_14954 (not_new_n8217_, new_n8217_);
  or g_14955 (new_n5210_, new_n1599_, new_n622_);
  or g_14956 (po295, or_or_or_not_new_n2982__not_new_n2985__not_new_n2984__not_new_n2986_, not_new_n2983_);
  not g_14957 (not_new_n7752_, new_n7752_);
  not g_14958 (new_n8501_, new_n8222_);
  or g_14959 (po056, key_gate_9, key_gate_21);
  not g_14960 (new_n4450_, new_n1011_);
  not g_14961 (not_new_n1601__797922662976120010, new_n1601_);
  and g_14962 (and_new_n2143__new_n2146_, new_n2146_, new_n2143_);
  or g_14963 (new_n3680_, not_new_n989__490, not_pi226);
  not g_14964 (not_new_n3776_, new_n3776_);
  not g_14965 (not_new_n599__8, new_n599_);
  or g_14966 (new_n6939_, not_new_n6533__0, not_new_n1061__1176490);
  not g_14967 (not_new_n1037__113988951853731430, new_n1037_);
  not g_14968 (not_new_n4452_, new_n4452_);
  not g_14969 (not_new_n8296_, new_n8296_);
  or g_14970 (new_n2447_, not_new_n603__57648010, not_new_n640__1);
  not g_14971 (not_new_n7830_, new_n7830_);
  not g_14972 (new_n5799_, new_n638_);
  or g_14973 (new_n6743_, not_new_n622__57648010, not_new_n6500_);
  or g_14974 (new_n8284_, not_new_n8168_, not_new_n1598__57648010);
  not g_14975 (not_new_n7230_, new_n7230_);
  not g_14976 (not_new_n7382_, new_n7382_);
  not g_14977 (new_n6052_, new_n5812_);
  or g_14978 (po122, not_new_n3425_, not_new_n3426_);
  not g_14979 (not_new_n1728__3, new_n1728_);
  or g_14980 (new_n5532_, not_pi133_1, not_new_n1007__5);
  not g_14981 (not_new_n1672_, key_gate_73);
  not g_14982 (not_new_n6248_, new_n6248_);
  not g_14983 (not_new_n1041__24010, new_n1041_);
  or g_14984 (new_n3078_, not_new_n1027__39098210485829880490, not_new_n1178_);
  not g_14985 (not_new_n5293_, new_n5293_);
  or g_14986 (new_n2673_, not_new_n609__1176490, not_new_n4460_);
  not g_14987 (not_new_n1617_, new_n1617_);
  not g_14988 (not_new_n1047__403536070, new_n1047_);
  and g_14989 (new_n6238_, and_and_new_n6244__new_n6372__new_n1596_, new_n6371_);
  not g_14990 (not_new_n5744_, new_n5744_);
  not g_14991 (not_pi166_1, pi166);
  not g_14992 (not_new_n989__8235430, new_n989_);
  not g_14993 (not_po298_10, po298);
  not g_14994 (not_new_n6443__1, new_n6443_);
  not g_14995 (not_new_n5559_, new_n5559_);
  or g_14996 (new_n2939_, not_new_n2936_, not_new_n1616__19773267430);
  or g_14997 (new_n8569_, not_new_n8269_, not_new_n8392__0);
  or g_14998 (new_n3819_, not_new_n3384__6, not_new_n2706_);
  not g_14999 (not_new_n7679_, new_n7679_);
  or g_15000 (or_not_new_n1055__168070_not_new_n6325_, not_new_n1055__168070, not_new_n6325_);
  not g_15001 (not_new_n3315__6, new_n3315_);
  not g_15002 (not_po298_9, po298);
  or g_15003 (or_or_or_not_pi269_1_not_pi260_1_not_pi257_1_not_pi248_1, or_or_not_pi269_1_not_pi260_1_not_pi257_1, not_pi248_1);
  or g_15004 (new_n4348_, or_or_not_new_n4246__not_new_n4350__not_new_n669_, not_new_n4351_);
  not g_15005 (not_new_n581__16284135979104490, new_n581_);
  not g_15006 (not_new_n607__5, new_n607_);
  not g_15007 (not_new_n3946_, new_n3946_);
  not g_15008 (not_new_n629__403536070, new_n629_);
  or g_15009 (new_n2072_, not_pi178, not_new_n586__1176490);
  or g_15010 (new_n9653_, not_new_n9652_, not_new_n9476_);
  or g_15011 (new_n3095_, not_new_n1045__3, not_new_n928__2);
  or g_15012 (or_or_not_new_n2284__not_new_n2281__not_new_n2282_, or_not_new_n2284__not_new_n2281_, not_new_n2282_);
  or g_15013 (new_n7690_, not_new_n8017_, not_new_n8018_);
  and g_15014 (new_n4904_, new_n5175_, new_n5176_);
  or g_15015 (new_n9257_, not_new_n8887_, not_new_n1601__113988951853731430);
  or g_15016 (new_n1859_, not_new_n593__3, not_new_n631_);
  or g_15017 (new_n2217_, not_new_n1589__138412872010, not_new_n5013_);
  not g_15018 (not_new_n5764__0, new_n5764_);
  not g_15019 (not_new_n3334_, new_n3334_);
  not g_15020 (not_new_n1554_, new_n1554_);
  not g_15021 (not_new_n1599__10, new_n1599_);
  not g_15022 (not_new_n1591_, new_n1591_);
  not g_15023 (not_new_n5662_, new_n5662_);
  and g_15024 (new_n7084_, new_n6965_, new_n7258_);
  not g_15025 (not_new_n5426_, new_n5426_);
  not g_15026 (not_new_n1616__9, new_n1616_);
  or g_15027 (new_n2108_, not_new_n1588__8235430, not_new_n1067_);
  not g_15028 (not_new_n2842_, new_n2842_);
  or g_15029 (new_n5601_, not_new_n5599_, not_new_n1003__6);
  not g_15030 (not_po296_43181145673964365640352930977077280875522488490, po296);
  or g_15031 (new_n2096_, not_new_n637__0, not_new_n601__168070);
  not g_15032 (not_new_n4838_, new_n4838_);
  not g_15033 (not_new_n7342_, new_n7342_);
  or g_15034 (new_n3510_, not_pi121_0, not_new_n1537__968890104070);
  or g_15035 (new_n6880_, not_new_n6537__0, not_new_n1598__168070);
  not g_15036 (not_new_n7005__0, new_n7005_);
  not g_15037 (not_new_n5000__0, new_n5000_);
  or g_15038 (new_n6774_, not_new_n6547_, not_new_n6650_);
  not g_15039 (not_new_n1598__10, new_n1598_);
  not g_15040 (not_new_n1067__24010, new_n1067_);
  not g_15041 (not_new_n9782_, new_n9782_);
  not g_15042 (new_n5956_, new_n5762_);
  not g_15043 (not_new_n8877_, new_n8877_);
  or g_15044 (or_not_new_n1555__not_new_n2434_, not_new_n1555_, not_new_n2434_);
  not g_15045 (not_new_n617__403536070, new_n617_);
  or g_15046 (new_n2039_, not_new_n644__0, not_new_n601__490);
  or g_15047 (new_n2398_, not_new_n4113__0, not_new_n600__8);
  or g_15048 (or_not_new_n6340__not_new_n6341_, not_new_n6340_, not_new_n6341_);
  and g_15049 (new_n6597_, new_n6756_, new_n6652_);
  or g_15050 (new_n1908_, not_new_n1585__6, not_new_n5827_);
  not g_15051 (not_new_n5446_, new_n5446_);
  not g_15052 (not_new_n8340__0, new_n8340_);
  or g_15053 (new_n2032_, not_new_n1588__3430, not_new_n1059_);
  not g_15054 (not_new_n1378_, new_n1378_);
  or g_15055 (new_n3817_, not_new_n3387__5, not_new_n3816_);
  or g_15056 (new_n947_, or_or_not_new_n1243__not_new_n1241__not_new_n1850_, not_new_n1849_);
  not g_15057 (not_new_n8826_, new_n8826_);
  or g_15058 (new_n3631_, not_new_n1611__403536070, not_new_n964_);
  xnor g_15059 (key_gate_98, not_new_n1663_, key_98);
  not g_15060 (not_new_n1551_, new_n1551_);
  and g_15061 (new_n6320_, new_n6406_, new_n6407_);
  not g_15062 (not_new_n4914_, new_n4914_);
  not g_15063 (not_new_n7013__1, new_n7013_);
  not g_15064 (not_new_n4426__0, new_n4426_);
  not g_15065 (new_n8858_, new_n638_);
  not g_15066 (not_new_n2072_, new_n2072_);
  not g_15067 (not_new_n8442_, new_n8442_);
  not g_15068 (new_n8354_, new_n8268_);
  not g_15069 (not_new_n5706__1, new_n5706_);
  not g_15070 (not_pi208, pi208);
  not g_15071 (new_n7132_, new_n749_);
  not g_15072 (not_new_n6193_, new_n6193_);
  or g_15073 (new_n6491_, not_new_n6674_, not_new_n6672_);
  not g_15074 (not_new_n1010__0, new_n1010_);
  or g_15075 (new_n5657_, not_new_n5474__0, not_new_n5509_);
  or g_15076 (new_n3623_, not_new_n1611__168070, not_new_n959_);
  not g_15077 (not_new_n1037__8235430, new_n1037_);
  or g_15078 (or_or_not_new_n1271__not_new_n1269__not_new_n1983_, not_new_n1983_, or_not_new_n1271__not_new_n1269_);
  or g_15079 (new_n10022_, not_new_n1031__138412872010, not_new_n641__138412872010);
  or g_15080 (new_n3102_, not_new_n581__657123623635342801395430, not_new_n624__6);
  or g_15081 (new_n2528_, not_new_n4462__0, not_new_n610__1);
  or g_15082 (new_n3620_, not_new_n984__24010, not_pi176_0);
  or g_15083 (new_n8978_, not_new_n9171_, not_new_n8936_);
  or g_15084 (or_or_not_new_n2091__not_new_n2092__not_new_n2094_, not_new_n2094_, or_not_new_n2091__not_new_n2092_);
  not g_15085 (not_new_n1767_, new_n1767_);
  not g_15086 (not_new_n1580_, new_n1580_);
  not g_15087 (not_new_n8032_, new_n8032_);
  not g_15088 (not_new_n9282_, new_n9282_);
  and g_15089 (new_n1325_, new_n2251_, new_n2250_);
  or g_15090 (new_n7161_, not_new_n720_, not_new_n7044_);
  not g_15091 (not_new_n6601_, new_n6601_);
  not g_15092 (not_new_n1605__2, new_n1605_);
  not g_15093 (not_new_n4165_, new_n4165_);
  not g_15094 (not_new_n6916_, new_n6916_);
  or g_15095 (new_n10032_, not_new_n1051__6782230728490, not_new_n647__16284135979104490);
  not g_15096 (not_new_n589__168070, new_n589_);
  not g_15097 (not_new_n3382_, new_n3382_);
  not g_15098 (not_new_n631__490, new_n631_);
  or g_15099 (new_n4755_, or_not_new_n4843__not_new_n4757_, not_new_n4760_);
  or g_15100 (new_n9749_, not_new_n9349_, not_new_n632__797922662976120010);
  not g_15101 (not_new_n4176_, new_n4176_);
  not g_15102 (not_new_n1018_, new_n1018_);
  not g_15103 (not_new_n10176_, new_n10176_);
  or g_15104 (new_n6758_, not_new_n6757_, not_new_n6545_);
  not g_15105 (not_new_n5596_, new_n5596_);
  or g_15106 (new_n3590_, not_new_n984_, not_pi161_0);
  not g_15107 (not_pi182_0, pi182);
  not g_15108 (not_new_n3054_, new_n3054_);
  and g_15109 (new_n4769_, new_n4862_, new_n4863_);
  or g_15110 (or_not_new_n2170__not_new_n2167_, not_new_n2167_, not_new_n2170_);
  and g_15111 (new_n1526_, new_n3077_, and_new_n3079__new_n998_);
  and g_15112 (new_n6599_, new_n6458_, new_n6737_);
  or g_15113 (new_n4959_, not_new_n648__3430, not_new_n1049__8);
  not g_15114 (not_new_n3702_, new_n3702_);
  or g_15115 (new_n4611_, not_new_n4426__0, not_pi167_3);
  or g_15116 (new_n9238_, not_new_n8849_, not_new_n1597__47475615099430);
  or g_15117 (new_n2131_, not_new_n588__403536070, not_pi117);
  not g_15118 (not_new_n1154_, new_n1154_);
  or g_15119 (new_n3460_, not_new_n1537__10, not_pi108_0);
  not g_15120 (not_new_n1039__2326305139872070, new_n1039_);
  not g_15121 (not_new_n4827__1, new_n4827_);
  not g_15122 (not_new_n3956_, new_n3956_);
  not g_15123 (not_new_n8145_, new_n8145_);
  or g_15124 (new_n4795_, not_new_n4797__0, not_new_n4829__0);
  not g_15125 (not_new_n581__6782230728490, new_n581_);
  or g_15126 (new_n5830_, not_new_n6122_, not_new_n6123_);
  or g_15127 (new_n2723_, not_new_n2720_, not_new_n3375__4);
  not g_15128 (not_po298_2, po298);
  not g_15129 (not_new_n3372__16284135979104490, new_n3372_);
  or g_15130 (or_or_not_new_n1787__not_new_n1788__not_new_n1790_, or_not_new_n1787__not_new_n1788_, not_new_n1790_);
  not g_15131 (not_new_n4116__2, new_n4116_);
  or g_15132 (new_n3835_, not_new_n631__70, not_new_n6443__3);
  or g_15133 (new_n2853_, not_new_n602__3430, not_new_n635__2);
  not g_15134 (not_new_n8837__0, new_n8837_);
  or g_15135 (new_n1694_, not_pi053, not_new_n1631__403536070);
  or g_15136 (new_n4458_, not_new_n4627_, not_new_n4628_);
  not g_15137 (not_new_n8655_, new_n8655_);
  not g_15138 (not_new_n7702_, new_n7702_);
  not g_15139 (not_new_n1537__968890104070, new_n1537_);
  not g_15140 (not_new_n3310__6, new_n3310_);
  not g_15141 (not_new_n9964__0, new_n9964_);
  xnor g_15142 (key_gate_116, key_116, not_new_n1631_);
  not g_15143 (not_po296_1577753820348458066150427430, po296);
  not g_15144 (not_new_n4670_, new_n4670_);
  not g_15145 (not_new_n7574_, new_n7574_);
  not g_15146 (not_pi226, pi226);
  not g_15147 (not_new_n8508_, new_n8508_);
  or g_15148 (new_n746_, not_new_n3200_, not_new_n3201_);
  not g_15149 (not_new_n7440_, new_n7440_);
  not g_15150 (not_new_n5276_, new_n5276_);
  not g_15151 (not_new_n629__9, new_n629_);
  not g_15152 (not_new_n3081_, new_n3081_);
  not g_15153 (not_new_n1065__8235430, new_n1065_);
  or g_15154 (new_n7870_, not_new_n7662__0, not_new_n7932_);
  not g_15155 (new_n4239_, new_n673_);
  not g_15156 (not_new_n5365_, new_n5365_);
  or g_15157 (new_n5251_, not_new_n5113_, not_new_n5082_);
  not g_15158 (not_new_n581__3119734822845423713013303218219760490, new_n581_);
  or g_15159 (new_n8736_, not_new_n8671_, or_not_new_n8595__not_new_n8593_);
  not g_15160 (not_new_n928__10, new_n928_);
  not g_15161 (not_new_n629__5, new_n629_);
  not g_15162 (not_new_n647__10, new_n647_);
  not g_15163 (not_new_n1536__3, new_n1536_);
  not g_15164 (not_new_n1612_, new_n1612_);
  not g_15165 (not_new_n7638_, new_n7638_);
  or g_15166 (or_not_new_n3155__not_new_n3154_, not_new_n3155_, not_new_n3154_);
  not g_15167 (not_new_n5813__0, new_n5813_);
  not g_15168 (not_new_n7895_, new_n7895_);
  not g_15169 (not_new_n602__0, new_n602_);
  and g_15170 (new_n8929_, new_n8800_, new_n9019_);
  or g_15171 (new_n5538_, not_new_n5500_, not_new_n5537_);
  not g_15172 (new_n4962_, new_n1057_);
  not g_15173 (not_new_n993_, new_n993_);
  or g_15174 (po180, not_new_n3587_, not_new_n3586_);
  not g_15175 (not_new_n724_, new_n724_);
  not g_15176 (not_new_n9969__0, new_n9969_);
  or g_15177 (new_n6535_, not_new_n6718_, not_new_n6720_);
  not g_15178 (not_new_n609__0, new_n609_);
  not g_15179 (not_new_n4330_, new_n4330_);
  or g_15180 (new_n3394_, not_pi032_0, not_new_n1536__3430);
  or g_15181 (new_n3391_, not_pi062_0, not_new_n1534__797922662976120010);
  not g_15182 (not_new_n8606_, new_n8606_);
  or g_15183 (new_n1536_, not_new_n3366_, not_new_n3369_);
  not g_15184 (not_new_n6521_, new_n6521_);
  not g_15185 (not_new_n1037__3, new_n1037_);
  not g_15186 (not_po296_125892552985318850263419623839875454447587430, po296);
  not g_15187 (not_new_n632__10, new_n632_);
  not g_15188 (not_new_n8545_, new_n8545_);
  and g_15189 (new_n9336_, new_n9614_, new_n9333_);
  not g_15190 (not_new_n1043__57648010, new_n1043_);
  or g_15191 (new_n8580_, not_new_n636__6782230728490, not_new_n8154__0);
  not g_15192 (not_new_n7451__1, new_n7451_);
  not g_15193 (not_new_n9454_, new_n9454_);
  not g_15194 (not_new_n6616_, new_n6616_);
  not g_15195 (not_new_n4260_, new_n4260_);
  not g_15196 (new_n4109_, pi247);
  not g_15197 (not_new_n9059__0, new_n9059_);
  not g_15198 (not_new_n1622_, new_n1622_);
  not g_15199 (not_new_n5078__1, new_n5078_);
  not g_15200 (not_new_n4343_, new_n4343_);
  not g_15201 (not_new_n639__47475615099430, new_n639_);
  not g_15202 (not_new_n7358_, new_n7358_);
  not g_15203 (new_n4925_, new_n1041_);
  not g_15204 (not_pi133_0, pi133);
  and g_15205 (new_n1297_, new_n2118_, new_n2117_);
  or g_15206 (new_n7242_, not_new_n7146_, not_new_n7082_);
  not g_15207 (not_new_n4987__0, new_n4987_);
  not g_15208 (not_new_n5568_, new_n5568_);
  not g_15209 (not_new_n6984__0, new_n6984_);
  not g_15210 (not_new_n6633__1, new_n6633_);
  not g_15211 (not_new_n5701_, new_n5701_);
  or g_15212 (new_n6714_, not_new_n1065__24010, not_new_n6531_);
  not g_15213 (not_new_n1023_, new_n1023_);
  not g_15214 (not_new_n10110_, new_n10110_);
  not g_15215 (not_new_n3232_, new_n3232_);
  or g_15216 (new_n2201_, not_new_n630_, not_new_n593__19773267430);
  or g_15217 (new_n10117_, new_n1604_, new_n640_);
  not g_15218 (not_pi064_5, pi064);
  not g_15219 (not_new_n3361_, new_n3361_);
  not g_15220 (not_new_n9906__0, new_n9906_);
  not g_15221 (not_new_n8233_, new_n8233_);
  not g_15222 (not_new_n9124_, new_n9124_);
  not g_15223 (not_new_n1714_, key_gate_33);
  not g_15224 (not_new_n1615__0, new_n1615_);
  not g_15225 (not_new_n3985_, new_n3985_);
  not g_15226 (not_new_n9344_, new_n9344_);
  or g_15227 (new_n5982_, not_new_n5716_, not_new_n5922_);
  not g_15228 (not_new_n6187_, new_n6187_);
  or g_15229 (new_n6665_, not_new_n6482__0, not_new_n6481_);
  not g_15230 (not_new_n5189_, new_n5189_);
  not g_15231 (not_new_n7936_, new_n7936_);
  or g_15232 (new_n7379_, not_new_n6976__2, not_new_n7020__0);
  not g_15233 (not_new_n994__19773267430, new_n994_);
  not g_15234 (not_new_n4902_, new_n4902_);
  and g_15235 (and_new_n4974__new_n5376_, new_n4974_, new_n5376_);
  not g_15236 (not_new_n9544_, new_n9544_);
  or g_15237 (new_n9758_, not_new_n9421_, not_new_n618__13410686196639649008070);
  not g_15238 (not_new_n598__0, new_n598_);
  not g_15239 (not_new_n5000_, new_n5000_);
  and g_15240 (new_n4302_, new_n4356_, new_n4355_);
  and g_15241 (new_n8967_, new_n9256_, new_n9257_);
  not g_15242 (not_new_n4692_, new_n4692_);
  not g_15243 (not_new_n10208_, new_n10208_);
  and g_15244 (new_n1382_, new_n2440_, new_n2441_);
  or g_15245 (new_n5277_, not_new_n5275_, not_new_n5164_);
  and g_15246 (new_n6571_, new_n6666_, new_n6667_);
  not g_15247 (not_new_n630__57648010, new_n630_);
  not g_15248 (new_n5469_, new_n1013_);
  not g_15249 (not_new_n7606_, new_n7606_);
  or g_15250 (new_n4606_, not_new_n4477__0, not_new_n4476_);
  or g_15251 (new_n6007_, not_new_n5805_, not_new_n1599__10);
  not g_15252 (not_new_n3311__0, new_n3311_);
  not g_15253 (not_new_n7035__0, new_n7035_);
  or g_15254 (po074, key_gate_99, not_new_n1201_);
  not g_15255 (new_n7134_, new_n717_);
  not g_15256 (not_new_n1045__0, new_n1045_);
  not g_15257 (new_n4319_, new_n649_);
  not g_15258 (not_new_n7013_, new_n7013_);
  and g_15259 (new_n6450_, new_n6732_, new_n6545_);
  not g_15260 (not_new_n9811_, new_n9811_);
  not g_15261 (not_new_n775__2, new_n775_);
  xnor g_15262 (key_gate_11, key_11, not_new_n1681_);
  not g_15263 (not_new_n4106_, new_n4106_);
  not g_15264 (not_new_n7940_, new_n7940_);
  or g_15265 (new_n727_, not_new_n3282_, not_new_n3281_);
  or g_15266 (or_or_or_not_new_n2497__not_new_n1568__not_new_n2498__not_new_n2500_, not_new_n2500_, or_or_not_new_n2497__not_new_n1568__not_new_n2498_);
  or g_15267 (new_n5996_, not_new_n5779_, not_new_n640__168070);
  or g_15268 (new_n3729_, not_new_n3727_, not_new_n3728_);
  or g_15269 (new_n7221_, not_new_n730_, not_new_n7035_);
  not g_15270 (not_new_n10273_, new_n10273_);
  not g_15271 (not_pi024, pi024);
  not g_15272 (not_new_n1069__57648010, new_n1069_);
  not g_15273 (not_new_n630__332329305696010, new_n630_);
  or g_15274 (new_n7031_, not_new_n7410_, not_new_n7411_);
  not g_15275 (not_new_n10071_, new_n10071_);
  not g_15276 (not_new_n2835_, new_n2835_);
  not g_15277 (not_new_n7106_, new_n7106_);
  or g_15278 (new_n8420_, not_new_n8271__1, not_new_n8213_);
  or g_15279 (new_n3478_, not_new_n1014__1, not_new_n1594__24010);
  not g_15280 (not_new_n7422_, new_n7422_);
  or g_15281 (new_n8871_, not_new_n9174_, not_new_n9061_);
  not g_15282 (not_new_n625__490, new_n625_);
  and g_15283 (new_n6457_, new_n6454_, new_n6710_);
  not g_15284 (not_new_n7320_, new_n7320_);
  or g_15285 (new_n6396_, not_new_n6295_, not_new_n626__19773267430);
  not g_15286 (not_new_n4126__1, new_n4126_);
  and g_15287 (new_n5738_, new_n6086_, new_n6080_);
  not g_15288 (not_new_n6631_, new_n6631_);
  or g_15289 (new_n2839_, not_new_n4123__2, not_new_n612__2);
  or g_15290 (new_n2261_, not_new_n1328_, not_new_n2256_);
  or g_15291 (new_n7041_, not_new_n7446_, not_new_n7447_);
  not g_15292 (not_new_n610__1176490, new_n610_);
  not g_15293 (new_n8890_, new_n622_);
  or g_15294 (new_n7478_, not_new_n7138__0, not_new_n7303_);
  or g_15295 (po262, not_new_n3710_, not_new_n3711_);
  or g_15296 (new_n9964_, not_new_n10299_, not_new_n10298_);
  not g_15297 (not_new_n4810_, new_n4810_);
  or g_15298 (new_n3614_, not_new_n984__70, not_pi173_0);
  not g_15299 (not_new_n593__6, new_n593_);
  or g_15300 (new_n2641_, not_new_n5479__0, not_new_n606__490);
  or g_15301 (new_n9295_, not_new_n9066__0, not_new_n9293_);
  and g_15302 (and_new_n2067__new_n2070_, new_n2067_, new_n2070_);
  or g_15303 (new_n5553_, not_pi139_1, not_new_n5452_);
  or g_15304 (new_n9826_, not_new_n9385__0, not_new_n638__4599865365447399609768010);
  not g_15305 (not_new_n6698_, new_n6698_);
  or g_15306 (new_n7532_, not_new_n7424__0, not_new_n730__0);
  or g_15307 (po137, not_new_n3501_, not_new_n3500_);
  not g_15308 (not_new_n1601__273687473400809163430, new_n1601_);
  not g_15309 (not_new_n6458_, new_n6458_);
  not g_15310 (not_new_n2936_, new_n2936_);
  or g_15311 (new_n1941_, not_new_n588__9, not_pi107);
  not g_15312 (new_n4019_, new_n3942_);
  or g_15313 (po158, not_new_n3543_, not_new_n3542_);
  or g_15314 (new_n6175_, not_new_n1035__9, not_new_n5752_);
  not g_15315 (not_new_n1436_, new_n1436_);
  not g_15316 (not_new_n10129_, new_n10129_);
  and g_15317 (new_n6628_, new_n6900_, new_n6899_);
  or g_15318 (new_n5384_, not_new_n4976_, not_new_n646__24010);
  or g_15319 (new_n1677_, not_pi017, not_po296_24010);
  not g_15320 (not_pi157, pi157);
  or g_15321 (new_n4067_, not_new_n3952_, not_pi049_3);
  not g_15322 (not_new_n1611__47475615099430, new_n1611_);
  or g_15323 (new_n9656_, not_new_n9654_, not_new_n9477_);
  not g_15324 (not_new_n641__138412872010, new_n641_);
  not g_15325 (not_new_n8130_, new_n8130_);
  not g_15326 (new_n2009_, new_n955_);
  or g_15327 (new_n1744_, not_pi088, not_new_n1728__490);
  not g_15328 (not_new_n10234_, new_n10234_);
  not g_15329 (not_new_n10043_, new_n10043_);
  not g_15330 (not_new_n8844_, new_n8844_);
  not g_15331 (not_new_n3942_, new_n3942_);
  not g_15332 (not_new_n6974__2326305139872070, new_n6974_);
  not g_15333 (not_pi018, pi018);
  not g_15334 (not_new_n9443_, new_n9443_);
  not g_15335 (not_new_n1603__6, new_n1603_);
  not g_15336 (not_new_n2613_, new_n2613_);
  not g_15337 (not_pi064_2824752490, pi064);
  not g_15338 (not_new_n1057__2824752490, new_n1057_);
  and g_15339 (new_n8815_, new_n9125_, new_n9128_);
  or g_15340 (new_n1789_, not_new_n586__1, not_pi161);
  not g_15341 (not_new_n1563_, new_n1563_);
  not g_15342 (new_n8870_, new_n643_);
  not g_15343 (not_new_n6206_, new_n6206_);
  not g_15344 (not_new_n1390_, new_n1390_);
  not g_15345 (not_new_n1014_, new_n1014_);
  or g_15346 (new_n3935_, not_new_n3959_, not_new_n3960_);
  not g_15347 (not_new_n2788_, new_n2788_);
  not g_15348 (not_new_n1596__8235430, new_n1596_);
  not g_15349 (not_new_n607__3, new_n607_);
  not g_15350 (po296, pi275);
  not g_15351 (not_new_n8781_, new_n8781_);
  not g_15352 (new_n4097_, pi254);
  buf g_15353 (po038, pi226);
  not g_15354 (not_new_n9085_, new_n9085_);
  not g_15355 (not_new_n4461__0, new_n4461_);
  not g_15356 (new_n5792_, new_n626_);
  not g_15357 (not_new_n6346_, new_n6346_);
  or g_15358 (new_n2946_, not_new_n3311__1176490, not_new_n1053__2);
  and g_15359 (new_n9469_, new_n9631_, new_n9507_);
  not g_15360 (not_new_n9028_, new_n9028_);
  not g_15361 (new_n6814_, new_n6642_);
  or g_15362 (new_n5107_, not_new_n634__3430, not_new_n5106_);
  not g_15363 (not_new_n8154__0, new_n8154_);
  not g_15364 (not_pi250_1, pi250);
  or g_15365 (new_n10188_, not_new_n10033_, not_new_n10184__0);
  or g_15366 (new_n3219_, not_new_n632__7, not_new_n589__168070);
  or g_15367 (new_n2411_, not_new_n597__10, not_new_n4808__0);
  or g_15368 (new_n6417_, or_or_or_not_new_n6226__not_new_n6323__not_new_n6324__not_new_n6242_, not_new_n1057__24010);
  not g_15369 (not_new_n9888__0, new_n9888_);
  or g_15370 (new_n3325_, not_new_n1534__4, not_pi042_0);
  or g_15371 (new_n5228_, not_new_n5226_, not_new_n5049_);
  or g_15372 (or_or_not_new_n9893__not_new_n9890__0_not_new_n10266_, not_new_n10266_, or_not_new_n9893__not_new_n9890__0);
  not g_15373 (not_new_n9964_, new_n9964_);
  not g_15374 (not_new_n644__8235430, new_n644_);
  or g_15375 (new_n9751_, not_new_n9487_, not_new_n619__19773267430);
  or g_15376 (new_n3162_, not_new_n928__47475615099430, not_new_n1059__3);
  not g_15377 (not_new_n7650_, new_n7650_);
  or g_15378 (new_n7815_, not_new_n7813_, not_new_n7702_);
  not g_15379 (not_new_n1158__1, new_n1158_);
  not g_15380 (not_new_n949_, new_n949_);
  not g_15381 (not_new_n596__490, key_gate_88);
  not g_15382 (not_new_n1538__113988951853731430, new_n1538_);
  and g_15383 (new_n6229_, new_n6240_, new_n6400_);
  not g_15384 (not_new_n5562_, new_n5562_);
  not g_15385 (not_new_n8999_, new_n8999_);
  not g_15386 (not_new_n9687_, new_n9687_);
  not g_15387 (not_new_n1216_, new_n1216_);
  not g_15388 (not_new_n5748_, new_n5748_);
  not g_15389 (not_new_n1291_, new_n1291_);
  not g_15390 (new_n7133_, new_n750_);
  or g_15391 (new_n1678_, key_gate_126, not_new_n596__24010);
  or g_15392 (new_n7891_, not_new_n7671_, not_new_n7769_);
  or g_15393 (new_n5185_, or_not_new_n5184__not_new_n5183_, not_new_n5182_);
  not g_15394 (not_new_n7536_, new_n7536_);
  and g_15395 (new_n1210_, new_n1719_, new_n1721_);
  not g_15396 (not_pi036_2, pi036);
  or g_15397 (new_n9961_, not_new_n10279_, not_new_n10280_);
  or g_15398 (new_n2071_, not_new_n2066_, not_new_n1288_);
  and g_15399 (po091, key_gate_101, pi070);
  not g_15400 (not_new_n7640_, new_n7640_);
  not g_15401 (new_n8630_, new_n1157_);
  or g_15402 (new_n9273_, not_new_n8880__0, not_new_n1603__968890104070);
  or g_15403 (new_n5302_, not_new_n4938__0, not_new_n634__168070);
  not g_15404 (not_new_n1055__24010, new_n1055_);
  or g_15405 (new_n3388_, not_new_n1534__113988951853731430, not_pi063_0);
  not g_15406 (not_new_n10219_, new_n10219_);
  not g_15407 (new_n5789_, new_n1059_);
  and g_15408 (new_n3992_, new_n4064_, new_n4063_);
  not g_15409 (not_new_n4467__0, new_n4467_);
  not g_15410 (not_new_n6613_, new_n6613_);
  not g_15411 (not_new_n3681_, new_n3681_);
  not g_15412 (not_new_n1002__1, new_n1002_);
  not g_15413 (not_new_n994_, new_n994_);
  not g_15414 (not_new_n6232__2, new_n6232_);
  not g_15415 (not_new_n586__8235430, new_n586_);
  not g_15416 (not_new_n4133__1, new_n4133_);
  and g_15417 (and_new_n3315__new_n923_, new_n923_, new_n3315_);
  or g_15418 (new_n10222_, not_new_n9879__1, not_new_n10052_);
  or g_15419 (new_n9115_, not_new_n8946_, not_new_n9113_);
  or g_15420 (po140, not_new_n3506_, not_new_n3507_);
  not g_15421 (not_new_n606__168070, new_n606_);
  not g_15422 (not_new_n1069__8, new_n1069_);
  or g_15423 (new_n2688_, not_new_n610__8235430, not_new_n4411__0);
  not g_15424 (not_new_n1615_, new_n1615_);
  or g_15425 (or_or_or_not_new_n6226__not_new_n6323__not_new_n6324__not_new_n6242_, not_new_n6242_, or_or_not_new_n6226__not_new_n6323__not_new_n6324_);
  not g_15426 (not_new_n1536__70, new_n1536_);
  or g_15427 (new_n3942_, not_new_n3913_, or_or_not_new_n3914__not_new_n3969__not_new_n4014_);
  not g_15428 (not_new_n1018__2, new_n1018_);
  or g_15429 (new_n8333_, not_new_n8285_, not_new_n8112__0);
  not g_15430 (not_new_n1061__4, new_n1061_);
  not g_15431 (not_new_n5416_, new_n5416_);
  not g_15432 (not_new_n6633__0, new_n6633_);
  not g_15433 (not_new_n7000_, new_n7000_);
  not g_15434 (not_new_n7645__0, new_n7645_);
  not g_15435 (not_new_n1063__332329305696010, new_n1063_);
  not g_15436 (not_new_n5195__0, new_n5195_);
  not g_15437 (not_new_n8561_, new_n8561_);
  not g_15438 (not_new_n2785_, new_n2785_);
  or g_15439 (new_n2817_, not_new_n626__3, not_new_n602__9);
  not g_15440 (not_new_n8924_, new_n8924_);
  not g_15441 (new_n8418_, new_n8161_);
  not g_15442 (not_new_n628__5, new_n628_);
  not g_15443 (not_new_n3437_, new_n3437_);
  or g_15444 (new_n8742_, not_new_n8740_, not_new_n8741_);
  not g_15445 (not_new_n9963__0, new_n9963_);
  not g_15446 (not_new_n9193_, new_n9193_);
  and g_15447 (new_n3931_, new_n3935_, new_n4010_);
  not g_15448 (not_new_n3579_, new_n3579_);
  or g_15449 (new_n2963_, or_not_new_n2962__not_new_n2961_, not_new_n2960_);
  or g_15450 (or_or_not_new_n2776__not_new_n2779__not_new_n2778_, not_new_n2778_, or_not_new_n2776__not_new_n2779_);
  and g_15451 (new_n1573_, new_n3817_, new_n3818_);
  not g_15452 (not_pi177_2, pi177);
  and g_15453 (new_n1438_, new_n2618_, new_n2619_);
  not g_15454 (not_new_n607__6, new_n607_);
  buf g_15455 (po040, pi224);
  and g_15456 (new_n9490_, new_n9759_, new_n9758_);
  or g_15457 (new_n6775_, not_new_n6524__1, not_new_n1055__57648010);
  not g_15458 (not_new_n7112_, new_n7112_);
  or g_15459 (new_n2676_, or_not_new_n2675__not_new_n2674_, not_new_n2673_);
  not g_15460 (not_new_n7669_, new_n7669_);
  and g_15461 (new_n1266_, new_n1968_, new_n1967_);
  or g_15462 (new_n5229_, new_n642_, new_n1035_);
  not g_15463 (not_new_n600__968890104070, new_n600_);
  or g_15464 (new_n6494_, not_new_n6491_, not_new_n6675_);
  or g_15465 (new_n8833_, not_new_n8994_, not_new_n8925_);
  not g_15466 (not_new_n598__403536070, new_n598_);
  not g_15467 (not_new_n1862_, new_n1862_);
  or g_15468 (new_n4581_, not_new_n4470_, not_new_n4579_);
  or g_15469 (new_n4117_, not_new_n4186_, not_new_n4185_);
  xor g_15470 (key_gate_39, key_39, not_new_n3928_);
  or g_15471 (new_n1773_, not_new_n1580__0, not_new_n6471_);
  not g_15472 (new_n7626_, new_n1600_);
  not g_15473 (not_new_n1293_, new_n1293_);
  not g_15474 (not_pi158, pi158);
  or g_15475 (new_n2301_, not_new_n586__16284135979104490, not_pi190);
  not g_15476 (not_po298_6, po298);
  or g_15477 (new_n1592_, not_new_n2349_, not_new_n1609_);
  not g_15478 (not_new_n638__10, new_n638_);
  not g_15479 (not_new_n4071__0, new_n4071_);
  not g_15480 (new_n9376_, new_n1597_);
  and g_15481 (new_n6578_, new_n6843_, new_n6655_);
  not g_15482 (not_new_n586__70, new_n586_);
  not g_15483 (new_n6483_, new_n1037_);
  not g_15484 (not_pi014_0, pi014);
  or g_15485 (new_n2985_, not_new_n595__2326305139872070, not_new_n6973_);
  not g_15486 (not_new_n4447__0, new_n4447_);
  not g_15487 (not_new_n4001_, new_n4001_);
  not g_15488 (not_new_n9024_, new_n9024_);
  not g_15489 (not_new_n6135_, new_n6135_);
  not g_15490 (not_new_n10317_, new_n10317_);
  not g_15491 (not_new_n1602__6, new_n1602_);
  not g_15492 (not_new_n946_, new_n946_);
  not g_15493 (not_new_n5750__0, new_n5750_);
  not g_15494 (not_new_n4161__1, new_n4161_);
  not g_15495 (not_new_n1613_, new_n1613_);
  not g_15496 (not_new_n9983_, new_n9983_);
  or g_15497 (new_n3378_, not_pi065, not_new_n1535_);
  not g_15498 (not_new_n7387_, new_n7387_);
  not g_15499 (not_new_n7588_, new_n7588_);
  not g_15500 (not_new_n4216_, new_n4216_);
  not g_15501 (not_new_n598__2326305139872070, new_n598_);
  not g_15502 (not_new_n10191_, new_n10191_);
  or g_15503 (po272, not_new_n2777_, or_or_or_not_new_n2776__not_new_n2779__not_new_n2778__not_new_n2780_);
  not g_15504 (not_new_n6974__3, new_n6974_);
  not g_15505 (not_new_n581__70, new_n581_);
  not g_15506 (not_new_n1047__8235430, new_n1047_);
  or g_15507 (new_n4415_, not_new_n1020__4, not_pi161_2);
  and g_15508 (and_new_n1745__new_n1744_, new_n1745_, new_n1744_);
  not g_15509 (not_new_n6486_, new_n6486_);
  not g_15510 (not_new_n593__8, new_n593_);
  or g_15511 (po287, or_or_or_not_new_n2910__not_new_n2913__not_new_n2912__not_new_n2914_, not_new_n2911_);
  and g_15512 (new_n8255_, new_n8512_, new_n8511_);
  not g_15513 (not_new_n8819_, new_n8819_);
  not g_15514 (not_new_n5449_, new_n5449_);
  not g_15515 (not_new_n4469_, new_n4469_);
  and g_15516 (new_n8932_, new_n9033_, new_n8798_);
  and g_15517 (new_n6316_, new_n6382_, new_n6369_);
  or g_15518 (new_n10139_, new_n621_, new_n1598_);
  not g_15519 (not_new_n631__8, new_n631_);
  not g_15520 (new_n9886_, new_n624_);
  or g_15521 (new_n4552_, not_pi172_1, not_new_n1018__2);
  or g_15522 (new_n9236_, not_new_n9234_, not_new_n9105_);
  not g_15523 (not_new_n1536__138412872010, new_n1536_);
  or g_15524 (or_not_new_n1546__not_new_n1362_, not_new_n1362_, not_new_n1546_);
  not g_15525 (not_pi269_2, pi269);
  not g_15526 (not_new_n1391_, new_n1391_);
  not g_15527 (not_new_n639__7, new_n639_);
  or g_15528 (new_n2391_, not_new_n597__6, not_new_n4728__0);
  not g_15529 (not_new_n6566_, new_n6566_);
  and g_15530 (new_n8819_, new_n9031_, new_n9034_);
  not g_15531 (not_new_n3199_, new_n3199_);
  not g_15532 (new_n1767_, new_n642_);
  not g_15533 (not_new_n3185__168070, new_n3185_);
  and g_15534 (new_n6600_, and_new_n6451__new_n6799_, new_n6756_);
  not g_15535 (not_new_n8811_, new_n8811_);
  or g_15536 (new_n5465_, not_new_n5567_, not_new_n5566_);
  not g_15537 (not_new_n1596__6782230728490, new_n1596_);
  or g_15538 (new_n4180_, not_new_n4078_, not_new_n4155__1);
  not g_15539 (not_new_n9683_, new_n9683_);
  or g_15540 (new_n6551_, not_new_n6892_, not_new_n6893_);
  not g_15541 (not_new_n621__1, new_n621_);
  or g_15542 (new_n2412_, not_new_n644__1, not_new_n603__70);
  xor g_15543 (key_gate_25, new_n1654_, key_25);
  not g_15544 (not_new_n629_, new_n629_);
  not g_15545 (not_new_n5668_, new_n5668_);
  or g_15546 (new_n3415_, not_pi099_0, not_new_n1537__1);
  not g_15547 (not_new_n3974_, new_n3974_);
  not g_15548 (not_new_n6443__7, new_n6443_);
  or g_15549 (new_n6640_, not_new_n6713_, or_not_new_n6817__not_new_n6788_);
  not g_15550 (not_new_n8473_, new_n8473_);
  not g_15551 (not_new_n3332_, new_n3332_);
  or g_15552 (new_n10293_, not_new_n10203_, not_new_n9947__0);
  not g_15553 (not_new_n583_, new_n583_);
  not g_15554 (not_new_n10147_, new_n10147_);
  or g_15555 (new_n8472_, not_new_n1045__332329305696010, not_new_n8118__2);
  not g_15556 (not_new_n8162__2, new_n8162_);
  or g_15557 (new_n5015_, not_new_n5382_, not_new_n5383_);
  not g_15558 (new_n4261_, new_n694_);
  or g_15559 (new_n6152_, not_new_n5768__0, not_new_n1600__70);
  and g_15560 (new_n6314_, new_n6384_, new_n6392_);
  or g_15561 (new_n3584_, not_new_n1538__16284135979104490, not_pi158_0);
  and g_15562 (new_n4726_, new_n4815_, new_n4821_);
  not g_15563 (not_new_n8596__2, new_n8596_);
  not g_15564 (not_new_n3384__0, new_n3384_);
  or g_15565 (new_n6197_, not_new_n6195_, not_new_n6196_);
  not g_15566 (not_new_n6804_, new_n6804_);
  not g_15567 (not_new_n9500_, new_n9500_);
  not g_15568 (not_new_n8213_, new_n8213_);
  not g_15569 (not_new_n8659_, new_n8659_);
  not g_15570 (not_new_n8322_, new_n8322_);
  not g_15571 (new_n6722_, new_n6535_);
  not g_15572 (not_new_n1039__9, new_n1039_);
  not g_15573 (not_new_n636__70, new_n636_);
  not g_15574 (not_new_n3565_, new_n3565_);
  not g_15575 (not_new_n8981_, new_n8981_);
  not g_15576 (not_new_n5454_, new_n5454_);
  not g_15577 (not_new_n4699_, new_n4699_);
  or g_15578 (new_n7843_, not_new_n7641_, not_new_n633__2824752490);
  not g_15579 (not_new_n9630_, new_n9630_);
  not g_15580 (new_n3976_, pi041);
  not g_15581 (new_n10120_, new_n9905_);
  not g_15582 (not_new_n1631__8235430, key_gate_76);
  or g_15583 (new_n7683_, not_new_n8068_, not_new_n8067_);
  not g_15584 (not_new_n7627__0, new_n7627_);
  or g_15585 (new_n4677_, not_pi176_3, not_new_n4444__0);
  or g_15586 (new_n3337_, not_new_n1534__10, not_pi036_0);
  or g_15587 (new_n7270_, not_new_n7138_, not_new_n7269_);
  not g_15588 (not_new_n1059__968890104070, new_n1059_);
  not g_15589 (not_new_n7897_, new_n7897_);
  or g_15590 (new_n9020_, not_new_n8929_, not_new_n9018_);
  or g_15591 (or_not_new_n2091__not_new_n2092_, not_new_n2092_, not_new_n2091_);
  or g_15592 (new_n6699_, not_new_n6698_, not_new_n6655__1);
  or g_15593 (new_n5132_, not_new_n4928__0, not_new_n5128_);
  and g_15594 (and_new_n2627__new_n2628_, new_n2627_, new_n2628_);
  or g_15595 (po055, key_gate_87, key_gate_28);
  not g_15596 (not_new_n9594__0, new_n9594_);
  not g_15597 (not_new_n3736_, new_n3736_);
  or g_15598 (new_n2728_, not_new_n3310_, not_new_n4132__2);
  not g_15599 (new_n4931_, new_n1031_);
  not g_15600 (not_new_n4443__0, new_n4443_);
  not g_15601 (new_n9924_, new_n1055_);
  not g_15602 (not_new_n8376__0, new_n8376_);
  not g_15603 (not_pi112_0, pi112);
  not g_15604 (not_new_n4994_, new_n4994_);
  or g_15605 (new_n2558_, not_new_n4465__0, not_new_n610__4);
  or g_15606 (new_n4404_, not_new_n4318_, not_new_n4402_);
  or g_15607 (new_n3224_, not_new_n3185__57648010, not_new_n1067__4);
  or g_15608 (new_n10076_, not_new_n10075_, not_new_n9983_);
  or g_15609 (new_n935_, not_new_n1768__1, not_new_n3384__1);
  or g_15610 (new_n1569_, not_new_n620_, not_new_n1344_);
  not g_15611 (not_new_n4228_, new_n4228_);
  or g_15612 (new_n8161_, not_new_n8341_, not_new_n8417_);
  not g_15613 (not_new_n4812_, new_n4812_);
  not g_15614 (not_new_n9771_, new_n9771_);
  not g_15615 (not_new_n8583_, new_n8583_);
  not g_15616 (not_new_n1063__1, new_n1063_);
  not g_15617 (not_new_n4465_, new_n4465_);
  not g_15618 (not_new_n9931_, new_n9931_);
  and g_15619 (new_n1506_, new_n1507_, new_n3034_);
  not g_15620 (not_new_n611_, new_n611_);
  or g_15621 (new_n3339_, not_new_n1534__70, not_pi035_0);
  not g_15622 (not_new_n640__1, new_n640_);
  not g_15623 (not_new_n5753__0, new_n5753_);
  not g_15624 (not_new_n5928__0, new_n5928_);
  not g_15625 (not_new_n4985__0, new_n4985_);
  not g_15626 (not_new_n6755_, new_n6755_);
  not g_15627 (not_new_n1327_, new_n1327_);
  not g_15628 (not_new_n4984__1, new_n4984_);
  or g_15629 (new_n8533_, not_new_n8386_, not_new_n8259_);
  or g_15630 (new_n3238_, not_new_n1053__5, not_new_n3185__47475615099430);
  or g_15631 (new_n4508_, not_new_n4543_, not_new_n4544_);
  not g_15632 (not_new_n6415_, new_n6415_);
  not g_15633 (not_new_n4197_, new_n4197_);
  not g_15634 (not_new_n1039__2824752490, new_n1039_);
  not g_15635 (new_n4817_, new_n4752_);
  not g_15636 (not_new_n8089_, new_n8089_);
  not g_15637 (not_new_n3878_, new_n3878_);
  not g_15638 (not_new_n3928_, new_n3928_);
  or g_15639 (or_or_not_new_n6240__not_new_n6330__not_new_n6331_, not_new_n6331_, or_not_new_n6240__not_new_n6330_);
  not g_15640 (not_new_n6443__9, new_n6443_);
  not g_15641 (not_new_n7010__0, new_n7010_);
  not g_15642 (not_new_n1061__70, new_n1061_);
  or g_15643 (new_n5639_, not_new_n5638_, not_new_n5637_);
  not g_15644 (not_new_n7614__0, new_n7614_);
  or g_15645 (new_n6785_, not_new_n6676_, not_new_n6453_);
  or g_15646 (new_n4534_, new_n1004_, pi168);
  or g_15647 (new_n3875_, not_new_n638__70, not_new_n6443__968890104070);
  not g_15648 (not_new_n8965_, new_n8965_);
  not g_15649 (not_new_n8392_, new_n8392_);
  or g_15650 (new_n2872_, not_new_n4122__1, not_new_n994__8235430);
  not g_15651 (not_new_n1037__138412872010, new_n1037_);
  or g_15652 (new_n5098_, not_new_n5024_, not_new_n4898__0);
  not g_15653 (not_new_n999_, new_n999_);
  not g_15654 (not_new_n5802_, new_n5802_);
  or g_15655 (new_n8198_, not_new_n8569_, not_new_n8568_);
  not g_15656 (not_pi034_1, pi034);
  not g_15657 (not_new_n628__1176490, new_n628_);
  or g_15658 (new_n664_, or_not_new_n3155__not_new_n3154_, not_new_n3153_);
  not g_15659 (not_pi162, pi162);
  not g_15660 (new_n6682_, new_n6613_);
  not g_15661 (not_new_n2035_, new_n2035_);
  not g_15662 (not_new_n775__7, new_n775_);
  or g_15663 (new_n3340_, not_pi064_70, not_new_n3929__0);
  or g_15664 (new_n6710_, not_new_n1057__168070, not_new_n6529_);
  not g_15665 (not_new_n7139__0, new_n7139_);
  or g_15666 (new_n6395_, not_new_n6311_, not_new_n6394_);
  or g_15667 (new_n2867_, not_new_n1616__3430, not_new_n2864_);
  not g_15668 (not_new_n2494_, new_n2494_);
  not g_15669 (new_n7766_, new_n7605_);
  not g_15670 (not_new_n3691_, new_n3691_);
  or g_15671 (new_n2955_, not_new_n613__6, not_new_n1601__1);
  not g_15672 (not_new_n8930_, new_n8930_);
  not g_15673 (not_new_n9383_, new_n9383_);
  not g_15674 (not_new_n8288_, new_n8288_);
  not g_15675 (not_new_n589__7490483309651862334944941026945644936490, new_n589_);
  not g_15676 (not_new_n7715_, new_n7715_);
  xnor g_15677 (key_gate_48, key_48, new_n1183_);
  not g_15678 (not_new_n5479__0, new_n5479_);
  not g_15679 (not_new_n1013__7, new_n1013_);
  not g_15680 (not_new_n602__168070, new_n602_);
  and g_15681 (new_n3921_, new_n4031_, new_n4039_);
  not g_15682 (not_new_n1588__3430, new_n1588_);
  not g_15683 (not_new_n1588__8235430, new_n1588_);
  not g_15684 (not_new_n1612__403536070, new_n1612_);
  or g_15685 (new_n9544_, not_new_n9543_, not_new_n9373__0);
  not g_15686 (not_new_n1397_, new_n1397_);
  not g_15687 (not_new_n1589__2, new_n1589_);
  or g_15688 (new_n3067_, not_new_n3372__113988951853731430, not_new_n643__4);
  not g_15689 (not_new_n922__0, new_n922_);
  or g_15690 (new_n4699_, not_new_n4698_, not_new_n4697_);
  not g_15691 (not_new_n9056__0, new_n9056_);
  or g_15692 (new_n5416_, not_new_n5414_, not_new_n5240__0);
  not g_15693 (not_new_n3819_, new_n3819_);
  or g_15694 (new_n7148_, not_new_n7081_, not_new_n7229_);
  not g_15695 (not_new_n8499_, new_n8499_);
  and g_15696 (new_n8702_, new_n8652_, new_n1156_);
  not g_15697 (not_new_n984__168070, new_n984_);
  or g_15698 (new_n2054_, not_pi145, not_new_n587__168070);
  not g_15699 (new_n4775_, new_n1601_);
  not g_15700 (not_new_n3087_, new_n3087_);
  not g_15701 (not_new_n9216_, new_n9216_);
  or g_15702 (new_n9797_, not_new_n9617_, not_new_n9795_);
  not g_15703 (not_new_n9965__0, new_n9965_);
  not g_15704 (not_new_n8423_, new_n8423_);
  not g_15705 (not_new_n631__138412872010, new_n631_);
  not g_15706 (new_n8868_, new_n644_);
  not g_15707 (not_new_n5280_, new_n5280_);
  or g_15708 (new_n3897_, not_new_n3899_, not_new_n10184_);
  not g_15709 (not_new_n5269_, new_n5269_);
  not g_15710 (not_po296_2326305139872070, po296);
  not g_15711 (not_new_n586__797922662976120010, new_n586_);
  not g_15712 (not_new_n9926__0, new_n9926_);
  and g_15713 (new_n9471_, new_n9339_, new_n9507_);
  not g_15714 (not_pi250_3, pi250);
  not g_15715 (not_new_n8141__0, new_n8141_);
  not g_15716 (not_new_n6615_, new_n6615_);
  or g_15717 (new_n4651_, not_new_n4490__0, not_pi180_2);
  not g_15718 (not_new_n1612__8, new_n1612_);
  not g_15719 (not_new_n3185__403536070, new_n3185_);
  not g_15720 (not_new_n7754__3, new_n7754_);
  not g_15721 (not_new_n9982_, new_n9982_);
  or g_15722 (new_n5278_, not_new_n4910_, not_new_n4999__1);
  not g_15723 (new_n8623_, new_n1069_);
  not g_15724 (not_new_n1065__6, new_n1065_);
  not g_15725 (not_new_n1432_, new_n1432_);
  not g_15726 (not_new_n2825_, new_n2825_);
  or g_15727 (new_n7434_, not_new_n7126_, not_new_n775__2824752490);
  not g_15728 (new_n8653_, new_n1156_);
  or g_15729 (new_n1167_, not_new_n3863_, not_new_n3864_);
  or g_15730 (new_n4885_, not_new_n4830_, not_new_n4794__0);
  not g_15731 (new_n8604_, new_n1045_);
  not g_15732 (not_new_n7663__1, new_n7663_);
  or g_15733 (new_n1161_, not_new_n3852_, not_new_n3851_);
  not g_15734 (not_new_n7643_, new_n7643_);
  not g_15735 (not_new_n2185__0, new_n2185_);
  not g_15736 (not_new_n968_, new_n968_);
  not g_15737 (not_pi020_0, pi020);
  and g_15738 (new_n8594_, new_n8766_, new_n8765_);
  not g_15739 (not_new_n6499__0, new_n6499_);
  or g_15740 (new_n5191_, not_new_n1602__8, not_new_n625__3430);
  not g_15741 (not_new_n635__968890104070, new_n635_);
  not g_15742 (not_new_n6689_, new_n6689_);
  not g_15743 (not_new_n1787_, new_n1787_);
  not g_15744 (not_new_n7845_, new_n7845_);
  not g_15745 (not_new_n626__13410686196639649008070, new_n626_);
  not g_15746 (not_new_n7678_, new_n7678_);
  not g_15747 (not_new_n10257_, new_n10257_);
  not g_15748 (not_new_n7020_, new_n7020_);
  not g_15749 (not_new_n8134_, new_n8134_);
  not g_15750 (not_new_n3918_, new_n3918_);
  not g_15751 (not_new_n9754_, new_n9754_);
  or g_15752 (or_or_not_new_n1283__not_new_n1281__not_new_n2040_, not_new_n2040_, or_not_new_n1283__not_new_n1281_);
  not g_15753 (new_n4252_, new_n666_);
  not g_15754 (not_new_n5767__2, new_n5767_);
  not g_15755 (not_new_n645__70, new_n645_);
  not g_15756 (new_n4264_, new_n660_);
  or g_15757 (new_n1668_, not_pi020, not_po296_70);
  not g_15758 (not_new_n3321_, new_n3321_);
  not g_15759 (not_new_n4829__0, new_n4829_);
  not g_15760 (not_new_n7074_, new_n7074_);
  not g_15761 (not_new_n10003_, new_n10003_);
  or g_15762 (po291, or_or_or_not_new_n2946__not_new_n2949__not_new_n2948__not_new_n2950_, not_new_n2947_);
  or g_15763 (new_n5370_, not_new_n639__24010, not_new_n4979_);
  and g_15764 (new_n4295_, and_new_n4344__new_n4343_, new_n4339_);
  not g_15765 (not_new_n589__1299348114471230201171721456984490, new_n589_);
  or g_15766 (new_n3762_, not_new_n3760_, not_new_n3761_);
  not g_15767 (not_new_n5791__2, new_n5791_);
  or g_15768 (new_n6946_, not_new_n6945_, not_new_n6816_);
  not g_15769 (not_new_n1009__0, new_n1009_);
  or g_15770 (or_or_not_new_n2740__not_new_n2743__not_new_n2742_, not_new_n2742_, or_not_new_n2740__not_new_n2743_);
  or g_15771 (or_not_new_n5266__not_new_n5206_, not_new_n5206_, not_new_n5266_);
  or g_15772 (new_n7992_, not_new_n7716_, not_new_n7744__0);
  not g_15773 (not_new_n5862_, new_n5862_);
  not g_15774 (not_new_n3678_, new_n3678_);
  not g_15775 (not_new_n1536__9, new_n1536_);
  not g_15776 (not_new_n596__0, key_gate_88);
  not g_15777 (not_new_n1396_, new_n1396_);
  not g_15778 (not_new_n4705_, new_n4705_);
  not g_15779 (not_new_n9106_, new_n9106_);
  or g_15780 (new_n8012_, not_new_n7627__2, not_new_n1601__968890104070);
  not g_15781 (not_new_n1612__2326305139872070, new_n1612_);
  not g_15782 (not_new_n1041__1, new_n1041_);
  not g_15783 (not_new_n4119_, new_n4119_);
  or g_15784 (or_or_not_new_n1939__not_new_n1940__not_new_n1942_, not_new_n1942_, or_not_new_n1939__not_new_n1940_);
  not g_15785 (not_new_n4128__1, new_n4128_);
  not g_15786 (not_new_n5702_, new_n5702_);
  not g_15787 (new_n8061_, new_n7730_);
  not g_15788 (not_new_n1035__1176490, new_n1035_);
  and g_15789 (new_n8242_, new_n8281_, new_n8586_);
  not g_15790 (not_new_n624__1, new_n624_);
  not g_15791 (not_new_n1534__10, key_gate_5);
  not g_15792 (not_new_n1069__138412872010, new_n1069_);
  or g_15793 (new_n7879_, not_new_n7722_, not_new_n7878_);
  or g_15794 (new_n3586_, not_new_n1538__113988951853731430, not_pi159_0);
  not g_15795 (not_new_n594__8, new_n594_);
  not g_15796 (not_new_n2300_, new_n2300_);
  or g_15797 (new_n5186_, new_n1069_, new_n646_);
  not g_15798 (not_new_n7080_, new_n7080_);
  not g_15799 (new_n6251_, new_n617_);
  not g_15800 (not_new_n7009_, new_n7009_);
  and g_15801 (and_new_n2404__new_n2403_, new_n2404_, new_n2403_);
  not g_15802 (not_new_n8481_, new_n8481_);
  not g_15803 (not_new_n775__3430, new_n775_);
  and g_15804 (and_new_n1460__new_n1466_, new_n1460_, new_n1466_);
  not g_15805 (not_new_n4427__0, new_n4427_);
  not g_15806 (not_new_n7339_, new_n7339_);
  not g_15807 (not_new_n1583__9, new_n1583_);
  not g_15808 (not_new_n9141_, new_n9141_);
  not g_15809 (not_new_n7771_, new_n7771_);
  not g_15810 (not_new_n1943_, new_n1943_);
  not g_15811 (not_new_n6531__0, new_n6531_);
  not g_15812 (not_new_n602__3430, new_n602_);
  and g_15813 (new_n7749_, new_n8019_, new_n8020_);
  not g_15814 (not_new_n2128__0, new_n2128_);
  not g_15815 (not_new_n8182_, new_n8182_);
  not g_15816 (new_n6187_, new_n5869_);
  or g_15817 (new_n9534_, not_new_n9365_, not_new_n9366_);
  not g_15818 (not_new_n1591__9, new_n1591_);
  not g_15819 (not_new_n5301_, new_n5301_);
  xor g_15820 (key_gate_97, key_97, not_new_n1645_);
  not g_15821 (not_new_n3553_, new_n3553_);
  not g_15822 (new_n4936_, new_n634_);
  or g_15823 (new_n5927_, not_new_n5899__1, not_new_n642__3430);
  not g_15824 (not_new_n8985_, new_n8985_);
  or g_15825 (new_n5363_, not_new_n625__24010, not_new_n4955_);
  or g_15826 (new_n6042_, not_new_n642__24010, not_new_n5898__0);
  or g_15827 (new_n4487_, not_new_n4488_, not_new_n4512_);
  not g_15828 (not_new_n596__47475615099430, key_gate_88);
  not g_15829 (not_new_n8355_, new_n8355_);
  not g_15830 (not_new_n7357__0, new_n7357_);
  not g_15831 (not_new_n9385__0, new_n9385_);
  or g_15832 (new_n2002_, not_new_n7683_, not_new_n1583__70);
  or g_15833 (new_n10157_, new_n1599_, new_n622_);
  not g_15834 (not_new_n10018__0, new_n10018_);
  not g_15835 (not_new_n3315__3430, new_n3315_);
  and g_15836 (new_n7076_, new_n7397_, and_new_n6983__new_n7398_);
  not g_15837 (not_new_n1600__332329305696010, new_n1600_);
  not g_15838 (not_new_n4789_, new_n4789_);
  or g_15839 (new_n3470_, not_pi110_0, not_new_n1537__490);
  and g_15840 (new_n3915_, new_n4047_, new_n4012_);
  not g_15841 (not_po296_12197604876358357001385738625629718207556152941312384010, po296);
  or g_15842 (new_n5970_, not_new_n5794_, not_new_n626__8235430);
  or g_15843 (new_n2984_, not_new_n1616__332329305696010, not_new_n2981_);
  not g_15844 (not_new_n7126_, new_n7126_);
  not g_15845 (not_new_n9129_, new_n9129_);
  not g_15846 (not_new_n1043__2824752490, new_n1043_);
  and g_15847 (new_n1531_, new_n1593_, new_n3183_);
  or g_15848 (new_n2452_, not_new_n603__403536070, not_new_n639__1);
  or g_15849 (new_n3495_, not_new_n1537__8235430, not_pi115_0);
  or g_15850 (new_n1840_, not_new_n593__2, not_new_n624_);
  or g_15851 (new_n9301_, not_new_n8975_, not_new_n8974_);
  not g_15852 (not_new_n8242_, new_n8242_);
  or g_15853 (new_n3621_, not_new_n958_, not_new_n1611__24010);
  not g_15854 (not_new_n2847_, new_n2847_);
  not g_15855 (not_new_n10165_, new_n10165_);
  not g_15856 (not_new_n5206_, new_n5206_);
  not g_15857 (not_new_n618__47475615099430, new_n618_);
  not g_15858 (not_pi167_2, pi167);
  not g_15859 (not_pi061_2, pi061);
  or g_15860 (new_n3816_, not_new_n3814_, not_new_n3815_);
  not g_15861 (not_new_n1055__6782230728490, new_n1055_);
  or g_15862 (new_n3646_, not_pi189_0, not_new_n984__2326305139872070);
  or g_15863 (new_n2862_, not_new_n602__24010, not_new_n633__3);
  not g_15864 (not_new_n643__3, new_n643_);
  not g_15865 (not_new_n1604__3, new_n1604_);
  not g_15866 (not_new_n3679_, new_n3679_);
  buf g_15867 (po002, pi195);
  not g_15868 (not_new_n625__797922662976120010, new_n625_);
  not g_15869 (not_new_n4656_, new_n4656_);
  not g_15870 (not_new_n1049__1, new_n1049_);
  not g_15871 (not_new_n1049__968890104070, new_n1049_);
  not g_15872 (not_new_n632__2326305139872070, new_n632_);
  not g_15873 (not_new_n4121__0, new_n4121_);
  or g_15874 (new_n8866_, not_new_n627__6782230728490, not_new_n1055__16284135979104490);
  and g_15875 (new_n8817_, new_n9115_, new_n9112_);
  not g_15876 (not_new_n631__5585458640832840070, new_n631_);
  not g_15877 (not_new_n9455_, new_n9455_);
  not g_15878 (not_new_n4979__0, new_n4979_);
  not g_15879 (not_new_n2893_, new_n2893_);
  not g_15880 (not_new_n2711_, new_n2711_);
  or g_15881 (new_n8789_, not_new_n1605__6, not_new_n8651_);
  not g_15882 (not_pi064_19773267430, pi064);
  not g_15883 (not_new_n9543_, new_n9543_);
  or g_15884 (new_n7810_, not_new_n631__47475615099430, not_new_n7599__0);
  not g_15885 (not_new_n9475_, new_n9475_);
  not g_15886 (not_new_n5794__0, new_n5794_);
  not g_15887 (not_new_n9425_, new_n9425_);
  not g_15888 (not_pi248_0, pi248);
  and g_15889 (new_n4916_, new_n5222_, new_n5220_);
  not g_15890 (not_new_n9691_, new_n9691_);
  not g_15891 (not_pi064_4, pi064);
  not g_15892 (not_new_n1043__4, new_n1043_);
  not g_15893 (not_new_n6232__5, new_n6232_);
  and g_15894 (new_n8661_, new_n1069_, new_n8624_);
  not g_15895 (not_new_n2939_, new_n2939_);
  not g_15896 (not_new_n622__8235430, new_n622_);
  not g_15897 (not_new_n1421_, new_n1421_);
  or g_15898 (po234, not_new_n3654_, not_new_n3655_);
  not g_15899 (not_new_n628__6, new_n628_);
  or g_15900 (new_n9215_, not_new_n9028__0, not_new_n9213_);
  not g_15901 (not_new_n8872_, new_n8872_);
  not g_15902 (not_new_n6232__4, new_n6232_);
  or g_15903 (new_n4515_, not_new_n4514_, not_new_n4487_);
  not g_15904 (not_new_n6825_, new_n6825_);
  not g_15905 (not_new_n8864_, new_n8864_);
  and g_15906 (new_n4728_, new_n4819_, new_n4752_);
  not g_15907 (not_new_n7638__0, new_n7638_);
  or g_15908 (new_n3818_, not_new_n1609__1, or_not_new_n1027__13410686196639649008070_not_new_n4227__0);
  or g_15909 (new_n5525_, not_new_n1009__5, not_pi131_1);
  or g_15910 (new_n2843_, not_new_n637__3, not_new_n604__70);
  not g_15911 (new_n6652_, new_n6545_);
  not g_15912 (not_new_n645__10, new_n645_);
  not g_15913 (not_new_n5456__0, new_n5456_);
  or g_15914 (new_n9438_, not_new_n9770_, not_new_n9771_);
  not g_15915 (not_new_n7797_, new_n7797_);
  not g_15916 (not_new_n638_, new_n638_);
  or g_15917 (new_n4877_, not_new_n1031__10, not_new_n4785_);
  not g_15918 (not_new_n1862__0, new_n1862_);
  and g_15919 (po113, key_gate_101, pi092);
  or g_15920 (new_n734_, not_new_n3296_, not_new_n3295_);
  or g_15921 (new_n6700_, not_new_n6490__0, not_new_n6673__0);
  or g_15922 (new_n4562_, new_n1015_, pi175);
  not g_15923 (not_new_n4210_, new_n4210_);
  not g_15924 (not_new_n10044_, new_n10044_);
  not g_15925 (not_new_n10242_, new_n10242_);
  and g_15926 (new_n6960_, new_n7172_, new_n7171_);
  not g_15927 (not_new_n4577_, new_n4577_);
  not g_15928 (not_new_n4956_, new_n4956_);
  or g_15929 (new_n5937_, not_new_n5713_, not_new_n5936_);
  not g_15930 (not_pi053_2, pi053);
  not g_15931 (not_new_n3178_, new_n3178_);
  not g_15932 (not_new_n5458__0, new_n5458_);
  not g_15933 (not_new_n10318_, new_n10318_);
  not g_15934 (not_new_n3917_, key_gate_70);
  or g_15935 (new_n2865_, not_new_n1065__1, not_new_n3311__10);
  not g_15936 (not_new_n1883_, new_n1883_);
  or g_15937 (new_n1658_, not_new_n1631__7, not_pi041);
  not g_15938 (not_new_n2351_, new_n2351_);
  and g_15939 (new_n8964_, new_n9237_, new_n9238_);
  or g_15940 (new_n9434_, not_new_n9743_, not_new_n9742_);
  not g_15941 (not_new_n6798_, new_n6798_);
  not g_15942 (not_new_n1039__10, new_n1039_);
  not g_15943 (not_pi262_0, pi262);
  not g_15944 (not_new_n1037__5, new_n1037_);
  not g_15945 (new_n8897_, new_n640_);
  or g_15946 (new_n3801_, not_new_n3800_, not_new_n3799_);
  and g_15947 (new_n1413_, new_n2506_, and_and_new_n2508__new_n2510__new_n2507_);
  or g_15948 (new_n2981_, or_not_new_n2980__not_new_n2979_, not_new_n2978_);
  not g_15949 (not_new_n1613__7, new_n1613_);
  not g_15950 (not_new_n3787_, new_n3787_);
  or g_15951 (new_n4053_, not_new_n4048_, not_new_n3980_);
  not g_15952 (not_pi178_0, pi178);
  not g_15953 (not_po298, po298);
  not g_15954 (not_new_n9082__0, new_n9082_);
  not g_15955 (not_new_n3925__0, key_gate_85);
  not g_15956 (not_new_n9612_, new_n9612_);
  not g_15957 (not_pi129_0, pi129);
  not g_15958 (not_pi121_0, pi121);
  not g_15959 (not_new_n9512__2, new_n9512_);
  not g_15960 (not_new_n1536__403536070, new_n1536_);
  not g_15961 (not_new_n5749__2, new_n5749_);
  not g_15962 (not_new_n8595__1, new_n8595_);
  not g_15963 (not_new_n1538__4, new_n1538_);
  not g_15964 (not_new_n7789_, new_n7789_);
  or g_15965 (new_n5315_, not_new_n5313_, not_new_n5128__0);
  not g_15966 (not_new_n3895_, new_n3895_);
  or g_15967 (new_n8345_, not_new_n8162_, not_new_n1065__138412872010);
  not g_15968 (not_new_n599__6782230728490, new_n599_);
  not g_15969 (not_new_n648__3, new_n648_);
  not g_15970 (not_new_n1624_, new_n1624_);
  not g_15971 (not_new_n619__8, new_n619_);
  or g_15972 (new_n3202_, not_new_n1597__4, not_new_n3185__7);
  not g_15973 (not_pi135_2, pi135);
  not g_15974 (not_new_n6473__1, new_n6473_);
  not g_15975 (not_new_n9269_, new_n9269_);
  and g_15976 (new_n1309_, new_n2175_, new_n2174_);
  or g_15977 (new_n2297_, not_new_n4766_, not_new_n591__2326305139872070);
  not g_15978 (not_new_n8954_, new_n8954_);
  not g_15979 (not_pi171_3, pi171);
  not g_15980 (new_n7635_, new_n645_);
  not g_15981 (new_n9897_, new_n647_);
  or g_15982 (new_n8401_, not_new_n8165__0, not_new_n8350__0);
  and g_15983 (and_and_not_pi056_1_not_pi055_1_not_pi054_1, not_pi054_1, and_not_pi056_1_not_pi055_1);
  not g_15984 (not_pi042_0, pi042);
  not g_15985 (not_new_n1537__168070, new_n1537_);
  not g_15986 (not_new_n1055__2824752490, new_n1055_);
  not g_15987 (not_new_n6476_, new_n6476_);
  not g_15988 (not_new_n8107_, new_n8107_);
  not g_15989 (not_new_n7569_, new_n7569_);
  or g_15990 (new_n4896_, not_new_n1053__8, not_new_n4810_);
  not g_15991 (not_new_n1534__5, key_gate_5);
  or g_15992 (new_n1938_, not_new_n1260_, not_new_n1933_);
  not g_15993 (not_new_n9087_, new_n9087_);
  not g_15994 (not_new_n8689_, new_n8689_);
  not g_15995 (not_new_n6286_, new_n6286_);
  or g_15996 (po150, not_new_n3526_, not_new_n3527_);
  not g_15997 (not_new_n3131_, new_n3131_);
  or g_15998 (new_n938_, not_new_n1578_, not_new_n3372__0);
  not g_15999 (not_new_n8502_, new_n8502_);
  not g_16000 (not_new_n7675_, new_n7675_);
  not g_16001 (not_new_n1053__3430, new_n1053_);
  not g_16002 (not_po296_85383234134508499009700170379408027452893070589186688070, po296);
  not g_16003 (not_new_n6620__0, new_n6620_);
  or g_16004 (po251, not_new_n3689_, not_new_n3688_);
  not g_16005 (not_pi071, pi071);
  or g_16006 (new_n10146_, not_new_n9993_, not_new_n10016_);
  not g_16007 (not_new_n3840_, new_n3840_);
  not g_16008 (not_new_n8552_, new_n8552_);
  not g_16009 (not_new_n726__0, new_n726_);
  and g_16010 (new_n1358_, new_n2380_, new_n2381_);
  not g_16011 (not_new_n4509_, new_n4509_);
  not g_16012 (not_new_n635__3, new_n635_);
  not g_16013 (not_new_n9379_, new_n9379_);
  not g_16014 (not_new_n928__332329305696010, new_n928_);
  not g_16015 (not_new_n1888_, new_n1888_);
  not g_16016 (not_new_n1061__6782230728490, new_n1061_);
  not g_16017 (not_new_n7691_, new_n7691_);
  or g_16018 (new_n4738_, not_new_n4809_, or_not_new_n4818__not_new_n4749_);
  not g_16019 (not_new_n1012__4, new_n1012_);
  or g_16020 (new_n2119_, not_new_n1581__8235430, not_new_n8186_);
  not g_16021 (not_new_n1061__47475615099430, new_n1061_);
  not g_16022 (not_new_n10192_, new_n10192_);
  not g_16023 (not_new_n7648__1, new_n7648_);
  not g_16024 (not_po296_52433383167563036344614587188619514555430, po296);
  not g_16025 (not_new_n8879_, new_n8879_);
  not g_16026 (not_new_n7288_, new_n7288_);
  not g_16027 (new_n7663_, new_n617_);
  or g_16028 (new_n6839_, not_new_n6689_, not_new_n6494__0);
  or g_16029 (new_n2367_, not_new_n603__2, not_new_n624__1);
  not g_16030 (new_n6479_, new_n1049_);
  not g_16031 (not_new_n7938_, new_n7938_);
  not g_16032 (not_new_n1599__6, new_n1599_);
  not g_16033 (not_new_n1606__4, new_n1606_);
  or g_16034 (new_n5222_, not_new_n5221_, not_new_n5374_);
  not g_16035 (not_new_n631__93874803376477543056490, new_n631_);
  or g_16036 (new_n7822_, not_new_n7650_, not_new_n627__2824752490);
  or g_16037 (new_n8049_, not_new_n637__19773267430, not_new_n7642__0);
  or g_16038 (new_n3883_, not_new_n627__70, not_new_n6443__2326305139872070);
  not g_16039 (not_new_n3475_, new_n3475_);
  or g_16040 (new_n8718_, not_new_n1163__0, not_new_n8648_);
  not g_16041 (not_new_n2615_, new_n2615_);
  not g_16042 (new_n3499_, new_n1071_);
  not g_16043 (not_new_n4102_, new_n4102_);
  not g_16044 (not_pi259_0, pi259);
  not g_16045 (not_new_n638__225393402906922580878632490, new_n638_);
  not g_16046 (not_new_n7362_, new_n7362_);
  not g_16047 (po298, new_n989_);
  not g_16048 (not_new_n4827__0, new_n4827_);
  or g_16049 (new_n2660_, not_new_n608__24010, not_new_n1007__0);
  and g_16050 (new_n3913_, not_pi057_1, and_and_not_pi060_1_not_pi059_1_not_pi058_1);
  not g_16051 (not_new_n4957__0, new_n4957_);
  or g_16052 (new_n8557_, not_new_n8267__0, not_new_n8235_);
  not g_16053 (not_new_n627__7, new_n627_);
  or g_16054 (new_n3794_, not_new_n636__10, not_new_n1057__6);
  not g_16055 (not_new_n6497__0, new_n6497_);
  not g_16056 (not_new_n636__7, new_n636_);
  not g_16057 (new_n4509_, new_n4488_);
  not g_16058 (not_new_n1728__10, new_n1728_);
  and g_16059 (new_n4920_, new_n5117_, new_n5120_);
  not g_16060 (not_new_n7827__0, new_n7827_);
  not g_16061 (not_new_n1317_, new_n1317_);
  not g_16062 (not_new_n3791_, new_n3791_);
  not g_16063 (new_n5807_, new_n1597_);
  not g_16064 (new_n3318_, new_n1001_);
  not g_16065 (not_pi255_3, pi255);
  not g_16066 (not_new_n1903_, new_n1903_);
  not g_16067 (not_new_n600__2, new_n600_);
  not g_16068 (not_new_n6641_, new_n6641_);
  not g_16069 (not_new_n7990_, new_n7990_);
  not g_16070 (not_new_n6974__3430, new_n6974_);
  not g_16071 (not_new_n7831_, new_n7831_);
  not g_16072 (not_new_n612__2, new_n612_);
  not g_16073 (not_new_n8910_, new_n8910_);
  not g_16074 (not_new_n9243_, new_n9243_);
  and g_16075 (and_new_n6977__new_n7377_, new_n6977_, new_n7377_);
  not g_16076 (not_new_n3286_, new_n3286_);
  not g_16077 (new_n8290_, new_n8121_);
  not g_16078 (not_new_n9862_, new_n9862_);
  not g_16079 (not_new_n8916_, new_n8916_);
  or g_16080 (new_n3674_, not_pi223, not_new_n989__9);
  not g_16081 (not_new_n1585__16284135979104490, new_n1585_);
  not g_16082 (not_new_n775__6782230728490, new_n775_);
  not g_16083 (not_new_n9955__0, new_n9955_);
  and g_16084 (new_n6612_, new_n6829_, new_n6828_);
  not g_16085 (not_new_n9422_, new_n9422_);
  not g_16086 (not_new_n593__47475615099430, new_n593_);
  not g_16087 (not_pi037_1, pi037);
  not g_16088 (not_new_n4959__0, new_n4959_);
  not g_16089 (not_new_n8151_, new_n8151_);
  not g_16090 (not_new_n5686__0, new_n5686_);
  or g_16091 (new_n5354_, not_new_n5066__0, not_new_n5260_);
  or g_16092 (new_n8710_, not_new_n8787_, not_new_n8788_);
  not g_16093 (not_new_n628__273687473400809163430, new_n628_);
  not g_16094 (not_new_n4990_, new_n4990_);
  not g_16095 (not_new_n4841__1, new_n4841_);
  or g_16096 (new_n741_, not_new_n3255_, not_new_n3256_);
  not g_16097 (not_new_n4728_, new_n4728_);
  or g_16098 (new_n6671_, not_new_n6655_, not_new_n6659_);
  not g_16099 (not_new_n5876_, new_n5876_);
  not g_16100 (not_new_n2988_, new_n2988_);
  not g_16101 (not_new_n8239_, new_n8239_);
  not g_16102 (not_pi135_1, pi135);
  not g_16103 (not_new_n602__57648010, new_n602_);
  not g_16104 (not_new_n1536__4, new_n1536_);
  not g_16105 (not_new_n3185__968890104070, new_n3185_);
  or g_16106 (new_n8403_, not_new_n8402_, not_new_n8443_);
  not g_16107 (not_new_n4932_, new_n4932_);
  not g_16108 (not_new_n6635__4, new_n6635_);
  not g_16109 (not_new_n5316_, new_n5316_);
  or g_16110 (new_n5580_, new_n1011_, pi147);
  not g_16111 (not_new_n633__7, new_n633_);
  not g_16112 (not_new_n742_, new_n742_);
  not g_16113 (not_new_n6448_, new_n6448_);
  or g_16114 (new_n1634_, key_gate_116, key_gate_81);
  not g_16115 (not_new_n9415_, new_n9415_);
  or g_16116 (new_n8373_, not_new_n8130_, not_new_n1599__1176490);
  or g_16117 (new_n9953_, not_new_n10321_, not_new_n10322_);
  not g_16118 (not_new_n5480_, new_n5480_);
  not g_16119 (not_new_n634__57648010, new_n634_);
  or g_16120 (new_n7229_, not_new_n6963_, not_new_n7016_);
  not g_16121 (not_pi011, pi011);
  not g_16122 (new_n5169_, new_n4984_);
  not g_16123 (not_new_n5826_, new_n5826_);
  not g_16124 (not_new_n10032_, new_n10032_);
  not g_16125 (new_n9352_, new_n628_);
  not g_16126 (not_new_n7775_, new_n7775_);
  or g_16127 (new_n4461_, not_new_n4659_, not_new_n4658_);
  not g_16128 (not_new_n3253_, new_n3253_);
  not g_16129 (not_new_n8276_, new_n8276_);
  or g_16130 (new_n2876_, not_new_n2873_, not_new_n1616__24010);
  not g_16131 (not_new_n3186_, new_n3186_);
  not g_16132 (not_new_n983_, new_n983_);
  not g_16133 (not_new_n599__1, new_n599_);
  not g_16134 (not_new_n588__5, new_n588_);
  or g_16135 (new_n2637_, not_new_n611__1176490, not_new_n2636_);
  not g_16136 (new_n7127_, new_n754_);
  or g_16137 (new_n2495_, not_new_n598__2326305139872070, not_new_n1596__0);
  not g_16138 (not_new_n603__4, new_n603_);
  not g_16139 (not_new_n10135_, new_n10135_);
  not g_16140 (not_new_n6981__0, new_n6981_);
  not g_16141 (not_new_n8012_, new_n8012_);
  not g_16142 (not_pi251, pi251);
  not g_16143 (not_new_n1768__0, new_n1768_);
  or g_16144 (new_n7205_, not_new_n6999_, not_new_n7418_);
  not g_16145 (not_new_n9406__0, new_n9406_);
  xnor g_16146 (key_gate_82, not_new_n1657_, key_82);
  not g_16147 (not_new_n3745_, new_n3745_);
  or g_16148 (new_n5083_, not_new_n636__24010, not_new_n1057__9);
  and g_16149 (and_new_n2998__new_n998_, new_n2998_, new_n998_);
  or g_16150 (new_n8908_, not_new_n9229_, not_new_n9228_);
  or g_16151 (new_n7588_, not_new_n7893_, not_new_n7890_);
  or g_16152 (new_n748_, not_new_n3205_, not_new_n3204_);
  or g_16153 (new_n4873_, not_new_n4780__1, not_new_n4835__1);
  not g_16154 (not_new_n1069__7, new_n1069_);
  or g_16155 (new_n7473_, not_new_n719__1, not_new_n7451__1);
  or g_16156 (new_n5307_, not_new_n4945__2, not_new_n5256_);
  not g_16157 (not_new_n9302_, new_n9302_);
  not g_16158 (not_new_n643__8, new_n643_);
  or g_16159 (new_n5907_, not_new_n5974_, not_new_n6069_);
  not g_16160 (new_n4251_, new_n667_);
  not g_16161 (not_new_n7754__0, new_n7754_);
  and g_16162 (and_new_n8104__new_n8464_, new_n8104_, new_n8464_);
  not g_16163 (not_new_n8436_, new_n8436_);
  not g_16164 (not_new_n6483_, new_n6483_);
  not g_16165 (not_new_n5132_, new_n5132_);
  or g_16166 (new_n1771_, not_new_n9430_, not_new_n1584_);
  not g_16167 (not_new_n3092_, new_n3092_);
  not g_16168 (not_new_n9541__0, new_n9541_);
  or g_16169 (or_not_new_n4410__not_new_n609_, not_new_n609_, not_new_n4410_);
  not g_16170 (not_new_n7694_, new_n7694_);
  and g_16171 (and_new_n5082__new_n5423_, new_n5423_, new_n5082_);
  not g_16172 (new_n1819_, new_n945_);
  not g_16173 (not_new_n3268_, new_n3268_);
  not g_16174 (not_new_n5974__0, new_n5974_);
  not g_16175 (not_new_n8292_, new_n8292_);
  not g_16176 (not_new_n1583__403536070, new_n1583_);
  not g_16177 (not_new_n4463__0, new_n4463_);
  not g_16178 (new_n7342_, new_n7023_);
  or g_16179 (new_n8837_, not_new_n1045__16284135979104490, not_new_n635__6782230728490);
  not g_16180 (not_new_n4474_, new_n4474_);
  or g_16181 (new_n2697_, not_new_n2696_, not_new_n611__138412872010);
  not g_16182 (not_new_n1534__3, key_gate_5);
  or g_16183 (new_n8460_, not_new_n647__968890104070, not_new_n8123__0);
  or g_16184 (new_n2866_, not_new_n4131__2, not_new_n3310__9);
  or g_16185 (new_n3548_, not_new_n1538__10, not_pi140_0);
  not g_16186 (not_pi256_1, pi256);
  or g_16187 (new_n7259_, not_new_n7451__0, not_new_n7013__0);
  not g_16188 (not_new_n3329_, new_n3329_);
  or g_16189 (new_n2112_, not_new_n588__57648010, not_pi116);
  and g_16190 (and_new_n6373__new_n6254_, new_n6373_, new_n6254_);
  or g_16191 (new_n2312_, not_new_n5009_, not_new_n1589__2326305139872070);
  not g_16192 (not_new_n594__9, new_n594_);
  or g_16193 (new_n9040_, not_new_n8830__1, not_new_n8833__0);
  not g_16194 (new_n7947_, new_n7754_);
  not g_16195 (not_new_n9105_, new_n9105_);
  not g_16196 (not_new_n7596_, new_n7596_);
  not g_16197 (not_new_n4126_, new_n4126_);
  or g_16198 (new_n1871_, not_new_n9347_, not_new_n1584__4);
  not g_16199 (not_new_n9461_, new_n9461_);
  not g_16200 (not_new_n2942_, new_n2942_);
  and g_16201 (new_n3930_, new_n4011_, new_n3939_);
  not g_16202 (not_new_n6474__0, new_n6474_);
  not g_16203 (not_new_n1584__47475615099430, new_n1584_);
  not g_16204 (not_new_n5113__0, new_n5113_);
  or g_16205 (new_n9626_, not_new_n9507_, not_new_n9515_);
  or g_16206 (or_not_new_n1243__not_new_n1241_, not_new_n1241_, not_new_n1243_);
  or g_16207 (new_n7974_, not_new_n1039__2824752490, not_new_n7606__2);
  or g_16208 (new_n2010_, not_new_n594__70, not_new_n9972_);
  not g_16209 (not_new_n625__4599865365447399609768010, new_n625_);
  and g_16210 (new_n5074_, new_n5397_, new_n5396_);
  not g_16211 (not_new_n1071__9, new_n1071_);
  not g_16212 (not_new_n3369__0, new_n3369_);
  not g_16213 (not_new_n597__2326305139872070, new_n597_);
  not g_16214 (not_new_n1728__113988951853731430, new_n1728_);
  or g_16215 (new_n2947_, not_new_n4137__2, not_new_n3310__168070);
  not g_16216 (not_pi134, pi134);
  not g_16217 (not_new_n2751_, new_n2751_);
  not g_16218 (not_new_n5739_, new_n5739_);
  not g_16219 (new_n6172_, new_n5866_);
  not g_16220 (not_new_n4997_, new_n4997_);
  not g_16221 (not_new_n10259_, new_n10259_);
  and g_16222 (new_n1326_, new_n2252_, new_n2253_);
  not g_16223 (not_new_n4016_, new_n4016_);
  or g_16224 (or_not_new_n1267__not_new_n1265_, not_new_n1265_, not_new_n1267_);
  not g_16225 (not_new_n3367_, new_n3367_);
  not g_16226 (new_n9418_, new_n622_);
  not g_16227 (not_new_n9904_, new_n9904_);
  not g_16228 (not_new_n8094_, new_n8094_);
  not g_16229 (not_new_n7109__1, new_n7109_);
  not g_16230 (not_new_n3182__0, new_n3182_);
  not g_16231 (not_new_n6895_, new_n6895_);
  not g_16232 (not_new_n4633_, new_n4633_);
  not g_16233 (not_new_n4122__1, new_n4122_);
  not g_16234 (not_new_n648__490, new_n648_);
  or g_16235 (new_n9563_, new_n624_, new_n1041_);
  not g_16236 (not_new_n1594__490, new_n1594_);
  not g_16237 (not_new_n2242__0, new_n2242_);
  not g_16238 (not_new_n595__4, new_n595_);
  not g_16239 (not_new_n7146__1, new_n7146_);
  not g_16240 (new_n3997_, pi045);
  not g_16241 (not_new_n5608_, new_n5608_);
  not g_16242 (not_new_n10225_, new_n10225_);
  not g_16243 (not_new_n4231_, new_n4231_);
  and g_16244 (new_n4140_, pi253, pi263);
  not g_16245 (not_pi239, pi239);
  or g_16246 (new_n703_, not_new_n2991_, not_new_n1487_);
  or g_16247 (new_n9082_, not_new_n9081_, not_new_n9080_);
  not g_16248 (not_new_n3489_, new_n3489_);
  not g_16249 (not_new_n2664_, new_n2664_);
  not g_16250 (not_new_n957_, new_n957_);
  or g_16251 (new_n2249_, not_new_n7675_, not_new_n1583__6782230728490);
  not g_16252 (not_pi142_0, pi142);
  not g_16253 (not_new_n4014__2, new_n4014_);
  not g_16254 (not_new_n9882_, new_n9882_);
  and g_16255 (new_n1277_, new_n2023_, new_n2022_);
  not g_16256 (not_new_n9188_, new_n9188_);
  not g_16257 (not_new_n730_, new_n730_);
  and g_16258 (new_n6621_, new_n6866_, new_n6867_);
  not g_16259 (not_new_n3311__4, new_n3311_);
  not g_16260 (not_new_n1631__47475615099430, key_gate_76);
  or g_16261 (new_n2429_, not_new_n599__24010, not_new_n9970__0);
  not g_16262 (not_new_n9610__0, new_n9610_);
  or g_16263 (new_n5561_, not_new_n1017__5, not_pi141_1);
  not g_16264 (not_new_n1604__490, new_n1604_);
  not g_16265 (not_new_n631__225393402906922580878632490, new_n631_);
  not g_16266 (not_new_n1584__5, new_n1584_);
  not g_16267 (not_new_n9430_, new_n9430_);
  and g_16268 (new_n9874_, new_n10079_, new_n10076_);
  or g_16269 (new_n3710_, not_pi241, not_new_n989__2326305139872070);
  not g_16270 (not_new_n643__968890104070, new_n643_);
  not g_16271 (not_new_n5306_, new_n5306_);
  not g_16272 (not_new_n1003_, new_n1003_);
  not g_16273 (not_new_n6541__1, new_n6541_);
  and g_16274 (and_and_not_pi044_1_not_pi043_1_not_pi046_1, and_not_pi044_1_not_pi043_1, not_pi046_1);
  not g_16275 (new_n5804_, new_n1599_);
  not g_16276 (not_new_n1580__4, new_n1580_);
  or g_16277 (new_n8906_, not_new_n9215_, not_new_n9214_);
  not g_16278 (not_new_n7433__0, new_n7433_);
  or g_16279 (or_not_new_n5441__not_new_n5617__1, not_new_n5441_, not_new_n5617__1);
  or g_16280 (new_n4077_, or_or_or_not_pi269_1_not_pi260_1_not_pi257_1_not_pi248_1, not_pi274_1);
  not g_16281 (not_new_n4456_, new_n4456_);
  not g_16282 (not_new_n1013__6, new_n1013_);
  not g_16283 (not_new_n7945_, new_n7945_);
  not g_16284 (not_new_n585__7, new_n585_);
  or g_16285 (new_n6911_, not_new_n6601_, not_new_n6632_);
  not g_16286 (not_new_n6469_, new_n6469_);
  not g_16287 (not_new_n7185_, new_n7185_);
  or g_16288 (new_n9675_, new_n1057_, new_n636_);
  not g_16289 (not_new_n6217_, new_n6217_);
  or g_16290 (or_not_new_n649__0_not_new_n4287_, not_new_n4287_, not_new_n649__0);
  not g_16291 (not_new_n628__7, new_n628_);
  or g_16292 (new_n5172_, not_new_n5169_, not_new_n1067__8);
  not g_16293 (not_new_n1069__6782230728490, new_n1069_);
  not g_16294 (new_n1630_, po297);
  not g_16295 (not_new_n3394_, new_n3394_);
  not g_16296 (not_pi085, pi085);
  not g_16297 (not_new_n7600_, new_n7600_);
  not g_16298 (not_new_n9343_, new_n9343_);
  or g_16299 (po257, not_new_n3701_, not_new_n3700_);
  not g_16300 (not_new_n6211_, new_n6211_);
  not g_16301 (not_new_n600__7, new_n600_);
  not g_16302 (not_new_n1004__3, new_n1004_);
  and g_16303 (new_n1492_, and_new_n3007__new_n998_, new_n3005_);
  or g_16304 (new_n2755_, not_new_n602__2, not_new_n645__2);
  not g_16305 (not_pi174_3, pi174);
  not g_16306 (not_new_n4272_, new_n4272_);
  or g_16307 (new_n3360_, not_pi064_19773267430, not_new_n3915__0);
  not g_16308 (not_new_n6500_, new_n6500_);
  not g_16309 (not_new_n4546_, new_n4546_);
  or g_16310 (new_n7954_, not_new_n1049__403536070, not_new_n7598__2);
  not g_16311 (not_new_n5350_, new_n5350_);
  not g_16312 (not_new_n1239_, new_n1239_);
  or g_16313 (new_n3513_, not_new_n1613__6782230728490, not_new_n2261_);
  not g_16314 (not_new_n7656__0, new_n7656_);
  or g_16315 (new_n4323_, or_not_new_n680__not_new_n4322_, not_new_n4321_);
  and g_16316 (new_n6575_, and_new_n6473__new_n6833_, new_n6832_);
  not g_16317 (new_n6787_, new_n6530_);
  not g_16318 (not_new_n4287_, new_n4287_);
  not g_16319 (not_new_n6999__0, new_n6999_);
  and g_16320 (new_n1362_, new_n2390_, new_n2391_);
  not g_16321 (not_new_n984__47475615099430, new_n984_);
  not g_16322 (not_new_n928__3430, new_n928_);
  not g_16323 (not_new_n596__332329305696010, key_gate_88);
  not g_16324 (not_new_n8842_, new_n8842_);
  not g_16325 (not_po298_968890104070, po298);
  not g_16326 (not_new_n9010_, new_n9010_);
  and g_16327 (new_n4756_, new_n4853_, new_n4852_);
  or g_16328 (new_n2896_, not_pi264, not_po296_725745515342319093317411710931737859674906464051430);
  not g_16329 (not_new_n7429_, new_n7429_);
  not g_16330 (not_new_n627__8, new_n627_);
  not g_16331 (not_new_n3582_, new_n3582_);
  or g_16332 (new_n8541_, not_new_n8432_, not_new_n8540_);
  and g_16333 (and_new_n1322__new_n2236_, new_n1322_, new_n2236_);
  or g_16334 (new_n2164_, not_new_n591__2824752490, not_new_n4784_);
  not g_16335 (not_new_n7427_, new_n7427_);
  not g_16336 (not_new_n7024__0, new_n7024_);
  not g_16337 (not_new_n4498_, new_n4498_);
  not g_16338 (not_new_n8123__0, new_n8123_);
  not g_16339 (not_new_n3491_, new_n3491_);
  or g_16340 (new_n1690_, not_new_n596__57648010, key_gate_53);
  not g_16341 (not_pi098, pi098);
  not g_16342 (new_n8294_, new_n8127_);
  or g_16343 (new_n4390_, not_new_n4313_, not_new_n4387_);
  or g_16344 (new_n7383_, not_new_n7360__0, not_new_n740__0);
  or g_16345 (new_n8901_, not_new_n9277_, not_new_n9278_);
  or g_16346 (new_n9122_, not_new_n9121_, not_new_n9274_);
  not g_16347 (not_new_n4412_, new_n4412_);
  or g_16348 (new_n9217_, not_new_n8824_, not_new_n1039__2326305139872070);
  not g_16349 (not_new_n1049__1176490, new_n1049_);
  or g_16350 (new_n5145_, not_new_n5088_, not_new_n4901_);
  not g_16351 (not_pi113, pi113);
  not g_16352 (not_new_n4135_, new_n4135_);
  not g_16353 (not_pi125, pi125);
  not g_16354 (not_new_n7184_, new_n7184_);
  and g_16355 (new_n7579_, new_n7571_, new_n7801_);
  not g_16356 (not_new_n5570_, new_n5570_);
  not g_16357 (not_new_n1616__24010, new_n1616_);
  not g_16358 (not_new_n9986_, new_n9986_);
  or g_16359 (new_n4398_, not_new_n4283_, not_new_n683_);
  not g_16360 (not_new_n2865_, new_n2865_);
  not g_16361 (not_new_n7476_, new_n7476_);
  not g_16362 (not_new_n5197__0, new_n5197_);
  or g_16363 (new_n2533_, not_new_n609__2, not_new_n4463_);
  not g_16364 (not_new_n7602__0, new_n7602_);
  or g_16365 (new_n10238_, not_new_n10237_, not_new_n10236_);
  or g_16366 (new_n2927_, or_not_new_n2926__not_new_n2925_, not_new_n2924_);
  or g_16367 (new_n3905_, not_new_n10028_, not_new_n10027_);
  or g_16368 (new_n7614_, not_new_n7601_, not_new_n624__2824752490);
  not g_16369 (not_new_n7707_, new_n7707_);
  not g_16370 (not_new_n1581__16284135979104490, new_n1581_);
  not g_16371 (not_pi064_3430, pi064);
  not g_16372 (new_n2247_, new_n621_);
  not g_16373 (not_new_n1537__70, new_n1537_);
  or g_16374 (new_n8277_, not_new_n8265__0, not_new_n8264_);
  not g_16375 (not_new_n8823_, new_n8823_);
  not g_16376 (not_new_n589__1070069044235980333563563003849377848070, new_n589_);
  not g_16377 (not_new_n5828_, new_n5828_);
  not g_16378 (not_new_n1045__968890104070, new_n1045_);
  not g_16379 (not_new_n3372__2824752490, new_n3372_);
  or g_16380 (or_not_new_n4461__not_new_n609__0, not_new_n4461_, not_new_n609__0);
  or g_16381 (new_n6701_, not_new_n6580_, not_new_n6823_);
  not g_16382 (not_pi126, pi126);
  or g_16383 (or_or_not_new_n6226__not_new_n6323__not_new_n6324_, or_not_new_n6226__not_new_n6323_, not_new_n6324_);
  or g_16384 (po239, not_new_n3665_, not_new_n3664_);
  not g_16385 (not_new_n7609_, new_n7609_);
  not g_16386 (not_new_n6518__0, new_n6518_);
  or g_16387 (new_n4634_, not_new_n4485__0, not_new_n4484_);
  or g_16388 (new_n8916_, not_new_n9288_, not_new_n9287_);
  not g_16389 (not_new_n5936_, new_n5936_);
  not g_16390 (not_new_n621__3430, new_n621_);
  not g_16391 (not_new_n1603__9, new_n1603_);
  or g_16392 (new_n2386_, not_new_n597__5, not_new_n4727__0);
  and g_16393 (new_n1280_, new_n2031_, and_and_new_n2029__new_n2032__new_n2030_);
  not g_16394 (not_new_n4433_, new_n4433_);
  not g_16395 (not_new_n1009__6, new_n1009_);
  not g_16396 (not_new_n1061__403536070, new_n1061_);
  or g_16397 (or_not_new_n3118__not_new_n3119_, not_new_n3119_, not_new_n3118_);
  not g_16398 (not_new_n3184__403536070, new_n3184_);
  not g_16399 (not_new_n1023__0, new_n1023_);
  not g_16400 (not_new_n597__24010, new_n597_);
  not g_16401 (not_new_n646__16284135979104490, new_n646_);
  not g_16402 (not_new_n3183_, new_n3183_);
  or g_16403 (new_n8342_, not_new_n636__968890104070, not_new_n8154_);
  not g_16404 (not_new_n5343_, new_n5343_);
  not g_16405 (not_new_n8928_, new_n8928_);
  or g_16406 (new_n2511_, not_po296_5585458640832840070, not_pi268);
  or g_16407 (new_n5203_, new_n617_, new_n1597_);
  or g_16408 (new_n10080_, new_n624_, new_n1041_);
  not g_16409 (not_new_n5008_, new_n5008_);
  and g_16410 (new_n5041_, new_n5079_, new_n5203_);
  or g_16411 (new_n4536_, not_pi168_1, not_new_n1004__2);
  not g_16412 (not_new_n6503__0, new_n6503_);
  not g_16413 (not_new_n5107_, new_n5107_);
  not g_16414 (not_new_n6533_, new_n6533_);
  or g_16415 (new_n2607_, not_new_n2606_, not_new_n611__3430);
  not g_16416 (not_new_n8613_, new_n8613_);
  not g_16417 (not_new_n2566_, new_n2566_);
  not g_16418 (new_n8107_, new_n1045_);
  not g_16419 (not_new_n8865_, new_n8865_);
  and g_16420 (new_n1394_, new_n2470_, new_n2471_);
  not g_16421 (not_new_n630__5, new_n630_);
  not g_16422 (not_new_n6405_, new_n6405_);
  not g_16423 (not_new_n6952_, new_n6952_);
  or g_16424 (new_n10315_, not_new_n1603__16284135979104490, not_new_n9911_);
  or g_16425 (new_n1893_, not_new_n8905_, not_new_n1591__5);
  or g_16426 (new_n4118_, not_new_n4187_, not_new_n4188_);
  not g_16427 (not_new_n8120_, new_n8120_);
  or g_16428 (new_n3070_, not_new_n644__4, not_new_n3372__797922662976120010);
  not g_16429 (not_new_n5313_, new_n5313_);
  not g_16430 (new_n4271_, new_n657_);
  not g_16431 (new_n9881_, new_n1037_);
  or g_16432 (new_n1708_, key_gate_117, not_new_n596__6782230728490);
  not g_16433 (not_new_n4104_, new_n4104_);
  or g_16434 (new_n3760_, not_new_n1597__6, not_new_n617__10);
  not g_16435 (not_new_n9267_, new_n9267_);
  not g_16436 (not_new_n4013_, new_n4013_);
  or g_16437 (new_n5596_, not_new_n5447__0, not_pi137_2);
  or g_16438 (new_n8239_, not_new_n8574_, not_new_n8575_);
  not g_16439 (new_n10218_, new_n9931_);
  not g_16440 (not_new_n1013__2, new_n1013_);
  not g_16441 (not_pi064_24010, pi064);
  or g_16442 (new_n6903_, not_new_n6505__0, not_new_n1603__168070);
  and g_16443 (and_new_n3064__new_n998_, new_n998_, new_n3064_);
  and g_16444 (new_n5043_, new_n4911_, new_n5079_);
  not g_16445 (not_new_n627__2824752490, new_n627_);
  or g_16446 (new_n3599_, not_new_n947_, not_new_n1611__3);
  not g_16447 (not_new_n4283_, new_n4283_);
  or g_16448 (new_n4743_, or_not_new_n4833__not_new_n4782_, not_new_n4787_);
  not g_16449 (not_new_n8799_, new_n8799_);
  or g_16450 (new_n6433_, or_or_or_not_new_n6239__not_new_n6350__not_new_n6232__3_not_new_n6317__0, not_new_n1037__3430);
  or g_16451 (new_n2136_, not_new_n1585__57648010, not_new_n5821_);
  not g_16452 (not_new_n3988_, new_n3988_);
  not g_16453 (not_new_n6196_, new_n6196_);
  or g_16454 (new_n3118_, not_new_n581__77309937197074445241370944070, not_new_n617__6);
  or g_16455 (new_n8376_, not_new_n8217_, not_new_n8256__0);
  or g_16456 (new_n1700_, not_pi055, not_new_n1631__19773267430);
  not g_16457 (not_new_n9494__0, new_n9494_);
  not g_16458 (new_n6305_, new_n1606_);
  not g_16459 (not_new_n7857_, new_n7857_);
  not g_16460 (not_new_n5013_, new_n5013_);
  not g_16461 (not_new_n1580__3, new_n1580_);
  or g_16462 (new_n4352_, not_new_n667_, not_new_n4248_);
  not g_16463 (not_new_n994__4, new_n994_);
  not g_16464 (not_new_n1055__10, new_n1055_);
  not g_16465 (not_new_n2244_, new_n2244_);
  not g_16466 (not_new_n4118__2, new_n4118_);
  not g_16467 (not_new_n728_, new_n728_);
  or g_16468 (new_n7973_, not_new_n628__6782230728490, not_new_n7610__0);
  not g_16469 (not_new_n3060_, new_n3060_);
  not g_16470 (not_new_n1604__968890104070, new_n1604_);
  or g_16471 (new_n7679_, not_new_n8036_, not_new_n8037_);
  not g_16472 (not_new_n2623_, new_n2623_);
  not g_16473 (not_new_n8905_, new_n8905_);
  or g_16474 (new_n2892_, not_new_n613__4, not_new_n1603__1);
  or g_16475 (new_n5758_, not_new_n5939_, not_new_n5937_);
  not g_16476 (new_n8109_, new_n1047_);
  not g_16477 (new_n4963_, new_n636_);
  or g_16478 (new_n1043_, not_new_n3428_, not_new_n3427_);
  not g_16479 (not_new_n8169_, new_n8169_);
  not g_16480 (not_new_n3733_, new_n3733_);
  or g_16481 (new_n8412_, not_new_n646__138412872010, not_new_n8167_);
  not g_16482 (not_new_n7381_, new_n7381_);
  or g_16483 (new_n5668_, not_new_n1013__7, not_new_n5468__0);
  or g_16484 (new_n8318_, not_new_n8287_, not_new_n8125_);
  or g_16485 (new_n6709_, not_new_n6707_, not_new_n6708_);
  and g_16486 (new_n1318_, new_n2214_, new_n2215_);
  or g_16487 (or_not_new_n2953__not_new_n2952_, not_new_n2953_, not_new_n2952_);
  not g_16488 (new_n4231_, new_n710_);
  not g_16489 (new_n9906_, new_n1604_);
  not g_16490 (not_new_n5769__0, new_n5769_);
  not g_16491 (not_new_n5242_, new_n5242_);
  or g_16492 (new_n8711_, not_new_n8716_, not_new_n8793_);
  or g_16493 (new_n4602_, not_pi168_2, not_new_n4428_);
  not g_16494 (not_new_n9421_, new_n9421_);
  not g_16495 (not_new_n3983_, new_n3983_);
  not g_16496 (not_new_n5392_, new_n5392_);
  or g_16497 (new_n9518_, new_n624_, new_n1041_);
  not g_16498 (not_new_n8851_, new_n8851_);
  not g_16499 (not_new_n5407_, new_n5407_);
  not g_16500 (not_new_n9932_, new_n9932_);
  not g_16501 (not_new_n3992__0, key_gate_56);
  not g_16502 (not_new_n1599__968890104070, new_n1599_);
  or g_16503 (new_n2840_, not_new_n1616__10, not_new_n2837_);
  not g_16504 (not_new_n3189_, new_n3189_);
  and g_16505 (new_n8694_, new_n8774_, new_n8775_);
  not g_16506 (not_new_n5505_, new_n5505_);
  or g_16507 (or_or_not_new_n2557__not_new_n2561__not_new_n1427_, or_not_new_n2557__not_new_n2561_, not_new_n1427_);
  and g_16508 (and_and_new_n3792__new_n3795__new_n3801_, and_new_n3792__new_n3795_, new_n3801_);
  or g_16509 (new_n3192_, not_new_n3185__2, not_new_n1045__4);
  or g_16510 (new_n7893_, not_new_n7728_, not_new_n7891_);
  not g_16511 (not_new_n1594__8235430, new_n1594_);
  not g_16512 (not_new_n2803_, new_n2803_);
  not g_16513 (not_new_n6041_, new_n6041_);
  and g_16514 (new_n8680_, new_n1177_, new_n8617_);
  not g_16515 (not_new_n632__2, new_n632_);
  or g_16516 (or_not_new_n6590__not_new_n6589_, not_new_n6589_, not_new_n6590_);
  not g_16517 (not_new_n994__16284135979104490, new_n994_);
  and g_16518 (new_n1194_, new_n1673_, new_n1671_);
  and g_16519 (new_n4478_, new_n4609_, new_n4608_);
  or g_16520 (new_n3622_, not_new_n984__168070, not_pi177_0);
  not g_16521 (not_new_n5443__0, new_n5443_);
  and g_16522 (and_new_n6365__new_n6439_, new_n6365_, new_n6439_);
  and g_16523 (new_n589_, new_n3180_, new_n922_);
  not g_16524 (not_new_n4303_, new_n4303_);
  not g_16525 (not_new_n9331_, new_n9331_);
  or g_16526 (or_not_pi269_2_not_pi248_2, not_pi269_2, not_pi248_2);
  or g_16527 (new_n661_, or_not_new_n3145__not_new_n3146_, not_new_n3144_);
  or g_16528 (new_n5598_, not_pi137_3, not_new_n5447__1);
  or g_16529 (new_n9744_, not_new_n628__1915812313805664144010, not_new_n9351_);
  not g_16530 (not_new_n3198_, new_n3198_);
  or g_16531 (new_n10074_, new_n624_, new_n1041_);
  not g_16532 (not_new_n1031__0, new_n1031_);
  not g_16533 (not_new_n9919_, new_n9919_);
  or g_16534 (new_n5669_, not_new_n5469__0, not_pi145_3);
  or g_16535 (new_n4891_, not_new_n4802__1, not_new_n4827__1);
  not g_16536 (not_new_n6806_, new_n6806_);
  not g_16537 (not_new_n6638_, new_n6638_);
  not g_16538 (not_pi001, pi001);
  not g_16539 (not_new_n7610__1, new_n7610_);
  or g_16540 (or_not_new_n4812__not_new_n4736_, not_new_n4812_, not_new_n4736_);
  or g_16541 (new_n8421_, not_new_n8355_, not_new_n8353_);
  or g_16542 (new_n2732_, not_new_n622__2, not_new_n604__0);
  not g_16543 (new_n6088_, new_n5900_);
  not g_16544 (not_new_n1905_, new_n1905_);
  or g_16545 (new_n2051_, not_new_n1588__24010, not_new_n1061_);
  not g_16546 (not_new_n4286_, new_n4286_);
  not g_16547 (not_new_n2971_, new_n2971_);
  not g_16548 (not_new_n3185__9, new_n3185_);
  not g_16549 (not_new_n608__10, new_n608_);
  or g_16550 (new_n6022_, not_new_n5905__0, not_new_n5984_);
  not g_16551 (not_new_n6510_, new_n6510_);
  or g_16552 (new_n9491_, not_new_n9716_, not_new_n9470_);
  not g_16553 (new_n1581_, new_n933_);
  not g_16554 (not_new_n7514_, new_n7514_);
  or g_16555 (new_n4005_, not_new_n4003_, not_new_n3976_);
  not g_16556 (not_new_n6835_, new_n6835_);
  not g_16557 (not_new_n634__8, new_n634_);
  or g_16558 (new_n8018_, not_new_n7748_, not_new_n7876__0);
  not g_16559 (not_new_n9950__1, new_n9950_);
  not g_16560 (not_new_n3823_, new_n3823_);
  or g_16561 (new_n2350_, not_new_n584__0, not_new_n1346_);
  not g_16562 (not_new_n8855_, new_n8855_);
  not g_16563 (not_new_n8256__1, new_n8256_);
  not g_16564 (not_new_n8112__1, new_n8112_);
  or g_16565 (new_n9075_, new_n1604_, new_n640_);
  or g_16566 (new_n3555_, not_new_n1612__3430, not_new_n2052__0);
  not g_16567 (not_new_n644__3, new_n644_);
  not g_16568 (not_pi184_0, pi184);
  not g_16569 (not_new_n5720__0, new_n5720_);
  or g_16570 (new_n5211_, not_new_n4994_, not_new_n5210_);
  not g_16571 (not_new_n630__19773267430, new_n630_);
  or g_16572 (new_n9143_, not_new_n8952_, not_new_n9142_);
  not g_16573 (not_new_n1597__9, new_n1597_);
  not g_16574 (not_new_n1600__70, new_n1600_);
  not g_16575 (not_new_n610__57648010, new_n610_);
  not g_16576 (not_new_n9740_, new_n9740_);
  not g_16577 (not_new_n2052_, new_n2052_);
  not g_16578 (not_new_n1055__2, new_n1055_);
  not g_16579 (not_new_n4476_, new_n4476_);
  buf g_16580 (po015, pi208);
  or g_16581 (new_n3116_, not_new_n3315__10, not_new_n617__5);
  not g_16582 (not_new_n2567_, new_n2567_);
  not g_16583 (not_new_n8720__0, new_n8720_);
  and g_16584 (and_new_n6388__new_n6313_, new_n6388_, new_n6313_);
  not g_16585 (new_n7436_, new_n7038_);
  or g_16586 (new_n2273_, not_new_n1591__47475615099430, not_new_n8817_);
  not g_16587 (not_new_n3072_, new_n3072_);
  or g_16588 (new_n2128_, not_new_n2123_, not_new_n1300_);
  not g_16589 (not_new_n7754_, new_n7754_);
  and g_16590 (new_n9871_, new_n10169_, new_n10167_);
  or g_16591 (new_n7318_, not_new_n6989_, not_new_n7187_);
  or g_16592 (new_n6770_, not_new_n6534__0, not_new_n6719__0);
  or g_16593 (new_n7211_, not_new_n7209_, not_new_n7078_);
  or g_16594 (new_n8100_, not_new_n8328_, not_new_n8325_);
  not g_16595 (not_new_n607__1, new_n607_);
  not g_16596 (not_pi146_0, pi146);
  or g_16597 (new_n2980_, not_new_n994__113988951853731430, not_new_n4115__1);
  not g_16598 (not_new_n7671__0, new_n7671_);
  not g_16599 (not_new_n5156_, new_n5156_);
  and g_16600 (and_new_n4295__new_n4334_, new_n4334_, new_n4295_);
  not g_16601 (not_new_n1055__8, new_n1055_);
  not g_16602 (not_new_n1051__490, new_n1051_);
  and g_16603 (new_n5503_, new_n5636_, new_n5635_);
  not g_16604 (not_new_n719_, new_n719_);
  not g_16605 (not_new_n6954_, new_n6954_);
  not g_16606 (not_new_n1053__5, new_n1053_);
  not g_16607 (not_new_n621__19773267430, new_n621_);
  or g_16608 (new_n5155_, not_new_n5153_, not_new_n5038_);
  not g_16609 (not_new_n9315_, new_n9315_);
  or g_16610 (new_n10298_, not_new_n10204_, not_new_n10016__1);
  not g_16611 (not_new_n4124_, new_n4124_);
  not g_16612 (not_new_n6368_, new_n6368_);
  or g_16613 (or_or_not_new_n2072__not_new_n2073__not_new_n2075_, or_not_new_n2072__not_new_n2073_, not_new_n2075_);
  not g_16614 (not_new_n591__2824752490, new_n591_);
  or g_16615 (new_n6200_, not_new_n5813__0, not_new_n6031_);
  not g_16616 (not_new_n3317_, new_n3317_);
  or g_16617 (new_n10203_, not_new_n10163_, not_new_n10034__0);
  not g_16618 (not_new_n4807__1, new_n4807_);
  not g_16619 (not_new_n6925_, new_n6925_);
  or g_16620 (new_n8752_, not_new_n8595__2, not_new_n8676_);
  or g_16621 (new_n3848_, not_new_n1576__9, not_new_n618__70);
  not g_16622 (not_new_n8371_, new_n8371_);
  not g_16623 (not_new_n4219_, new_n4219_);
  or g_16624 (new_n7447_, not_new_n751_, not_new_n6974__968890104070);
  or g_16625 (new_n8273_, not_new_n8444_, not_new_n8340_);
  or g_16626 (new_n5915_, not_new_n1053__490, not_new_n5792_);
  not g_16627 (not_new_n4942_, new_n4942_);
  or g_16628 (new_n1811_, not_new_n642__0, not_new_n601__0);
  not g_16629 (not_new_n8558_, new_n8558_);
  or g_16630 (new_n9228_, not_new_n8961_, not_new_n8960_);
  not g_16631 (not_new_n8434_, new_n8434_);
  or g_16632 (po157, not_new_n3541_, not_new_n3540_);
  not g_16633 (not_new_n989__403536070, new_n989_);
  xor g_16634 (key_gate_118, not_new_n1672_, key_118);
  not g_16635 (not_new_n9981_, new_n9981_);
  not g_16636 (not_new_n635__113988951853731430, new_n635_);
  not g_16637 (not_new_n642__332329305696010, new_n642_);
  and g_16638 (new_n5877_, new_n6091_, new_n6092_);
  or g_16639 (new_n8282_, not_new_n1063__8235430, not_new_n8163_);
  not g_16640 (not_new_n9901_, new_n9901_);
  or g_16641 (new_n3257_, not_new_n1039__5, not_new_n589__1915812313805664144010);
  not g_16642 (not_new_n5452__0, new_n5452_);
  and g_16643 (new_n9975_, new_n1037_, new_n632_);
  not g_16644 (not_new_n7544_, new_n7544_);
  not g_16645 (not_new_n10126_, new_n10126_);
  or g_16646 (new_n8727_, not_new_n1047__403536070, not_new_n8634_);
  or g_16647 (new_n2192_, not_new_n1583__19773267430, not_new_n7690_);
  not g_16648 (not_pi064_1, pi064);
  not g_16649 (not_new_n9140_, new_n9140_);
  and g_16650 (new_n1196_, new_n1679_, new_n1677_);
  or g_16651 (new_n6928_, not_new_n6517__0, not_new_n633__403536070);
  not g_16652 (not_new_n9930__0, new_n9930_);
  or g_16653 (new_n9266_, not_new_n8856__0, not_new_n1602__6782230728490);
  or g_16654 (new_n3063_, not_new_n1173_, not_new_n1027__2326305139872070);
  not g_16655 (new_n10113_, new_n9915_);
  or g_16656 (new_n7902_, not_new_n7732_, not_new_n7900_);
  not g_16657 (not_new_n1538__5, new_n1538_);
  not g_16658 (not_pi064_70, pi064);
  not g_16659 (not_new_n3375__5, new_n3375_);
  not g_16660 (not_new_n3372__4, new_n3372_);
  or g_16661 (new_n4064_, not_new_n4032__1, not_new_n3991__0);
  or g_16662 (new_n9315_, not_new_n8900__0, not_new_n9164_);
  or g_16663 (new_n2219_, not_new_n594__138412872010, not_new_n9965_);
  not g_16664 (not_new_n7031_, new_n7031_);
  or g_16665 (new_n5481_, not_new_n5627_, not_new_n5628_);
  or g_16666 (new_n7336_, not_new_n7018__1, not_new_n6988_);
  not g_16667 (not_new_n5052_, new_n5052_);
  or g_16668 (new_n3265_, not_new_n1599__5, not_new_n589__4599865365447399609768010);
  not g_16669 (not_new_n7143_, new_n7143_);
  or g_16670 (new_n8067_, not_new_n8066_, not_new_n7936_);
  or g_16671 (new_n1774_, not_new_n1591_, not_new_n8902_);
  not g_16672 (not_pi104_0, pi104);
  and g_16673 (and_new_n1543__new_n2376_, new_n1543_, new_n2376_);
  not g_16674 (not_new_n7603_, new_n7603_);
  not g_16675 (not_new_n4662_, new_n4662_);
  or g_16676 (new_n7963_, not_new_n7962_, not_new_n7961_);
  not g_16677 (not_new_n7759__1, new_n7759_);
  not g_16678 (not_new_n6859_, new_n6859_);
  not g_16679 (not_new_n5972_, new_n5972_);
  not g_16680 (not_new_n2862_, new_n2862_);
  or g_16681 (po195, not_new_n1374_, or_or_not_new_n1552__not_new_n2419__not_new_n1373_);
  and g_16682 (new_n6355_, new_n1067_, new_n6224_);
  or g_16683 (new_n6144_, not_new_n621__8235430, not_new_n5806__0);
  not g_16684 (new_n1962_, new_n627_);
  not g_16685 (not_new_n8633_, new_n8633_);
  or g_16686 (new_n8036_, not_new_n7947_, not_new_n8035_);
  not g_16687 (new_n4272_, new_n656_);
  not g_16688 (not_new_n6307_, new_n6307_);
  and g_16689 (new_n7096_, new_n6962_, new_n7298_);
  not g_16690 (not_new_n2303_, new_n2303_);
  or g_16691 (new_n8511_, not_new_n1598__403536070, not_new_n8168__0);
  and g_16692 (new_n4311_, new_n4383_, new_n4382_);
  not g_16693 (not_new_n6047_, new_n6047_);
  not g_16694 (not_new_n589__3, new_n589_);
  or g_16695 (new_n7025_, not_new_n7350_, not_new_n7349_);
  or g_16696 (new_n1059_, not_new_n3468_, not_new_n3467_);
  not g_16697 (not_new_n4597_, new_n4597_);
  or g_16698 (new_n3516_, not_new_n1537__332329305696010, not_pi124_0);
  not g_16699 (not_new_n1538__2824752490, new_n1538_);
  not g_16700 (not_new_n8207_, new_n8207_);
  not g_16701 (not_pi138_1, pi138);
  or g_16702 (new_n728_, not_new_n3284_, not_new_n3283_);
  not g_16703 (not_new_n2535_, new_n2535_);
  not g_16704 (not_new_n10158_, new_n10158_);
  not g_16705 (not_new_n1602__403536070, new_n1602_);
  not g_16706 (not_pi114, pi114);
  not g_16707 (not_new_n1868_, new_n1868_);
  and g_16708 (new_n1259_, new_n1931_, and_new_n1258__new_n1932_);
  not g_16709 (not_new_n1612__7, new_n1612_);
  or g_16710 (new_n7568_, not_new_n7027__0, not_new_n7567_);
  not g_16711 (new_n7323_, new_n7111_);
  not g_16712 (new_n3981_, pi063);
  not g_16713 (not_new_n8258_, new_n8258_);
  not g_16714 (not_new_n5799_, new_n5799_);
  not g_16715 (not_new_n1028__490, new_n1028_);
  and g_16716 (new_n1397_, new_n2477_, new_n2478_);
  not g_16717 (new_n7277_, new_n7015_);
  or g_16718 (new_n985_, or_not_new_n3375__2_not_new_n3387__1, not_new_n1577_);
  and g_16719 (and_and_new_n1043__new_n6232__new_n6229_, and_new_n1043__new_n6232_, new_n6229_);
  not g_16720 (not_new_n1600__47475615099430, new_n1600_);
  or g_16721 (new_n1024_, not_new_n3374_, not_new_n3373_);
  not g_16722 (not_new_n609__7, new_n609_);
  not g_16723 (new_n7010_, new_n720_);
  not g_16724 (not_new_n640__24010, new_n640_);
  or g_16725 (new_n10209_, not_new_n10100__0, not_new_n9926__0);
  or g_16726 (po175, not_new_n3577_, not_new_n3576_);
  not g_16727 (not_new_n4434_, new_n4434_);
  and g_16728 (new_n5852_, new_n6055_, new_n6006_);
  not g_16729 (not_new_n1687_, key_gate_103);
  or g_16730 (new_n2975_, not_new_n2972_, not_new_n1616__47475615099430);
  not g_16731 (not_new_n7454__0, new_n7454_);
  not g_16732 (not_new_n1728__9, new_n1728_);
  or g_16733 (new_n4353_, not_new_n666_, not_new_n4253_);
  not g_16734 (not_new_n8427_, new_n8427_);
  or g_16735 (or_not_new_n8833__not_new_n8830__0, not_new_n8830__0, not_new_n8833_);
  or g_16736 (new_n7945_, not_new_n7605__1, not_new_n7781_);
  not g_16737 (not_pi047_3, pi047);
  and g_16738 (new_n1234_, new_n1815_, new_n1816_);
  not g_16739 (not_new_n603__19773267430, new_n603_);
  not g_16740 (not_new_n6673_, new_n6673_);
  or g_16741 (new_n7185_, not_new_n7184_, not_new_n7021_);
  not g_16742 (not_new_n7342__0, new_n7342_);
  not g_16743 (new_n6252_, new_n624_);
  not g_16744 (not_new_n647__19773267430, new_n647_);
  or g_16745 (new_n5813_, not_new_n5801_, not_new_n6022_);
  not g_16746 (not_new_n4828_, new_n4828_);
  or g_16747 (new_n4345_, not_new_n4242_, not_new_n702_);
  not g_16748 (not_new_n5620_, new_n5620_);
  not g_16749 (not_new_n4417__0, new_n4417_);
  or g_16750 (new_n7066_, not_new_n7545_, not_new_n7544_);
  or g_16751 (new_n10137_, not_new_n630__797922662976120010, not_new_n1601__1915812313805664144010);
  not g_16752 (not_new_n6625_, new_n6625_);
  or g_16753 (new_n4675_, not_pi176_2, not_new_n4444_);
  not g_16754 (not_new_n984__1, new_n984_);
  not g_16755 (not_new_n5914_, new_n5914_);
  not g_16756 (not_new_n9854__0, new_n9854_);
  not g_16757 (not_new_n1049__7, new_n1049_);
  and g_16758 (new_n8205_, new_n8416_, new_n8204_);
  and g_16759 (new_n5495_, new_n5589_, new_n5590_);
  not g_16760 (not_new_n627__6, new_n627_);
  and g_16761 (new_n4798_, new_n4886_, new_n4887_);
  or g_16762 (new_n7214_, not_new_n7213_, not_new_n7211_);
  or g_16763 (new_n6407_, not_new_n642__1176490, not_new_n6281_);
  or g_16764 (new_n9748_, not_new_n9746_, not_new_n9565_);
  or g_16765 (new_n2998_, not_new_n3372__6, not_new_n634__4);
  or g_16766 (or_or_not_new_n2227__not_new_n2224__not_new_n2225_, or_not_new_n2227__not_new_n2224_, not_new_n2225_);
  or g_16767 (new_n5593_, not_new_n5592_, not_new_n5591_);
  or g_16768 (new_n9259_, not_new_n1601__797922662976120010, not_new_n8887__0);
  or g_16769 (new_n3107_, not_new_n581__32199057558131797268376070, not_new_n623__1);
  not g_16770 (not_new_n5531_, new_n5531_);
  or g_16771 (new_n5111_, new_n1049_, new_n648_);
  not g_16772 (not_pi244, pi244);
  not g_16773 (new_n9917_, new_n1063_);
  and g_16774 (new_n5719_, new_n5999_, new_n5998_);
  not g_16775 (not_new_n8520_, new_n8520_);
  not g_16776 (not_new_n3837_, new_n3837_);
  not g_16777 (not_pi015, pi015);
  or g_16778 (new_n2383_, not_new_n4116__0, not_new_n600__5);
  not g_16779 (not_new_n4126__0, new_n4126_);
  not g_16780 (not_new_n8595__3, new_n8595_);
  not g_16781 (not_new_n9536_, new_n9536_);
  not g_16782 (not_new_n5140_, new_n5140_);
  or g_16783 (new_n3721_, not_new_n1605__3, not_new_n620__3);
  not g_16784 (not_new_n3032_, new_n3032_);
  not g_16785 (not_new_n2614_, new_n2614_);
  or g_16786 (new_n1692_, not_pi012_0, not_po296_403536070);
  or g_16787 (new_n2643_, not_new_n4457_, not_new_n609__3430);
  or g_16788 (or_or_not_new_n4246__not_new_n4350__not_new_n669_, or_not_new_n4246__not_new_n4350_, not_new_n669_);
  not g_16789 (not_new_n1995__0, new_n1995_);
  or g_16790 (po210, not_new_n1404_, or_or_not_new_n1567__not_new_n2494__not_new_n1403_);
  or g_16791 (new_n3155_, not_new_n638__5, not_new_n3315__968890104070);
  or g_16792 (new_n7904_, not_new_n7903_, not_new_n7768__0);
  not g_16793 (not_new_n3921__0, key_gate_75);
  not g_16794 (not_pi183_0, pi183);
  not g_16795 (not_new_n1037__968890104070, new_n1037_);
  not g_16796 (not_new_n589__8235430, new_n589_);
  not g_16797 (not_new_n5033_, new_n5033_);
  or g_16798 (or_or_not_new_n6337__not_new_n6373__6_not_new_n6338_, not_new_n6338_, or_not_new_n6337__not_new_n6373__6);
  not g_16799 (new_n4760_, new_n1607_);
  and g_16800 (new_n590_, pi275, new_n614_);
  or g_16801 (new_n7483_, not_new_n7139__1, not_new_n7304_);
  not g_16802 (not_new_n1051__138412872010, new_n1051_);
  or g_16803 (po292, not_new_n2956_, or_or_or_not_new_n2955__not_new_n2958__not_new_n2957__not_new_n2959_);
  not g_16804 (not_new_n8303_, new_n8303_);
  or g_16805 (new_n6562_, not_new_n6850_, not_new_n6851_);
  or g_16806 (new_n1680_, not_po296_168070, not_pi016);
  or g_16807 (new_n3749_, not_new_n965_, not_new_n2152_);
  not g_16808 (new_n6520_, new_n1061_);
  not g_16809 (not_new_n1057__47475615099430, new_n1057_);
  and g_16810 (and_new_n8304__new_n8299_, new_n8304_, new_n8299_);
  or g_16811 (new_n9688_, not_new_n9382__0, not_new_n9627__0);
  or g_16812 (new_n6824_, not_new_n6636_, not_new_n6727_);
  or g_16813 (new_n9305_, not_new_n643__113988951853731430, not_new_n8869__0);
  not g_16814 (not_po296_77309937197074445241370944070, po296);
  not g_16815 (not_new_n1613__3430, new_n1613_);
  not g_16816 (not_new_n1051__70, new_n1051_);
  or g_16817 (new_n1974_, not_new_n591__10, not_new_n4811_);
  not g_16818 (not_new_n7424__0, new_n7424_);
  or g_16819 (new_n3240_, not_new_n1035__4, not_new_n3185__332329305696010);
  or g_16820 (new_n2396_, not_new_n4753__0, not_new_n597__7);
  not g_16821 (not_new_n6613__1, new_n6613_);
  not g_16822 (not_new_n5746__0, new_n5746_);
  not g_16823 (new_n6761_, new_n6546_);
  not g_16824 (not_new_n634__9, new_n634_);
  not g_16825 (not_new_n5781_, new_n5781_);
  not g_16826 (not_new_n10204_, new_n10204_);
  or g_16827 (new_n7328_, not_new_n7155_, not_new_n7205_);
  or g_16828 (new_n8306_, not_new_n8248_, not_new_n8083_);
  not g_16829 (not_new_n4322__0, new_n4322_);
  not g_16830 (new_n8889_, new_n1599_);
  not g_16831 (not_new_n3516_, new_n3516_);
  not g_16832 (not_new_n5733__0, new_n5733_);
  not g_16833 (not_new_n9083_, new_n9083_);
  not g_16834 (not_new_n1598__1, new_n1598_);
  not g_16835 (not_new_n5550_, new_n5550_);
  or g_16836 (new_n3285_, not_new_n589__1299348114471230201171721456984490, not_new_n1065__5);
  or g_16837 (new_n5891_, not_new_n5852_, not_new_n6065_);
  or g_16838 (new_n1627_, not_new_n940_, not_new_n614_);
  not g_16839 (not_new_n6517_, new_n6517_);
  not g_16840 (not_pi133_3, pi133);
  not g_16841 (not_new_n3463_, new_n3463_);
  not g_16842 (not_new_n7753_, new_n7753_);
  not g_16843 (not_new_n1057__6, new_n1057_);
  not g_16844 (not_new_n9873_, new_n9873_);
  not g_16845 (not_new_n7599_, new_n7599_);
  not g_16846 (not_new_n5808__1, new_n5808_);
  not g_16847 (not_new_n1231_, new_n1231_);
  not g_16848 (not_new_n9373__1, new_n9373_);
  not g_16849 (not_new_n6443__16284135979104490, new_n6443_);
  or g_16850 (new_n6122_, not_new_n5967_, not_new_n5763__1);
  or g_16851 (new_n7687_, not_new_n7971_, not_new_n7970_);
  or g_16852 (new_n5521_, not_new_n5520_, not_new_n1010__4);
  not g_16853 (not_new_n3897_, new_n3897_);
  not g_16854 (not_new_n4963_, new_n4963_);
  not g_16855 (not_new_n6994__0, new_n6994_);
  not g_16856 (not_new_n6580_, new_n6580_);
  and g_16857 (new_n1270_, new_n1987_, new_n1986_);
  not g_16858 (not_new_n605__3, new_n605_);
  not g_16859 (not_new_n637__1, new_n637_);
  not g_16860 (not_new_n655_, new_n655_);
  not g_16861 (not_new_n3120_, new_n3120_);
  or g_16862 (new_n4325_, not_new_n678_, not_new_n4231_);
  or g_16863 (po248, not_new_n3683_, not_new_n3682_);
  not g_16864 (not_new_n3416_, new_n3416_);
  and g_16865 (new_n1481_, new_n2832_, new_n2833_);
  not g_16866 (not_new_n5474__0, new_n5474_);
  or g_16867 (new_n8508_, not_new_n8129__1, not_new_n617__16284135979104490);
  not g_16868 (not_new_n3654_, new_n3654_);
  not g_16869 (not_new_n4129__1, new_n4129_);
  or g_16870 (new_n2078_, not_new_n1583__168070, not_new_n7588_);
  or g_16871 (new_n3603_, not_new_n1611__5, not_new_n949_);
  or g_16872 (new_n2672_, not_new_n2509__168070, not_pi209);
  not g_16873 (not_new_n1597__1, new_n1597_);
  not g_16874 (not_new_n7960_, new_n7960_);
  not g_16875 (not_new_n602__5, new_n602_);
  not g_16876 (not_new_n1013__5, new_n1013_);
  not g_16877 (not_new_n5335_, new_n5335_);
  or g_16878 (new_n4083_, not_new_n4139_, not_new_n4157_);
  not g_16879 (not_new_n7629__0, new_n7629_);
  or g_16880 (new_n5963_, not_new_n5742__1, not_new_n631__57648010);
  not g_16881 (not_pi058_3, pi058);
  not g_16882 (not_new_n646__10, new_n646_);
  not g_16883 (new_n8009_, new_n7720_);
  or g_16884 (new_n8888_, not_new_n8940_, not_new_n9182_);
  not g_16885 (not_pi255_0, pi255);
  not g_16886 (not_new_n1583__6, new_n1583_);
  not g_16887 (not_new_n3311__3, new_n3311_);
  and g_16888 (new_n1402_, new_n2491_, new_n2490_);
  not g_16889 (not_new_n8711_, new_n8711_);
  not g_16890 (not_new_n8206_, new_n8206_);
  or g_16891 (new_n2276_, not_new_n9872_, not_new_n594__47475615099430);
  not g_16892 (not_new_n739__0, new_n739_);
  and g_16893 (new_n1473_, new_n987_, and_new_n1575__new_n938_);
  or g_16894 (new_n2557_, not_new_n2556_, not_new_n611__8);
  not g_16895 (new_n4256_, new_n664_);
  or g_16896 (new_n7824_, not_new_n7571_, not_new_n7778_);
  not g_16897 (not_new_n9411_, new_n9411_);
  not g_16898 (not_new_n1039__6, new_n1039_);
  and g_16899 (new_n6968_, new_n7296_, new_n7299_);
  not g_16900 (not_po298_403536070, po298);
  or g_16901 (new_n1963_, not_new_n647__0, not_new_n601__8);
  or g_16902 (or_not_new_n2890__not_new_n2889_, not_new_n2890_, not_new_n2889_);
  not g_16903 (not_new_n3570_, new_n3570_);
  not g_16904 (not_new_n9848_, new_n9848_);
  not g_16905 (not_new_n1581__1176490, new_n1581_);
  not g_16906 (not_new_n1602__138412872010, new_n1602_);
  not g_16907 (new_n8633_, new_n1152_);
  or g_16908 (new_n9356_, not_new_n1041__138412872010, not_new_n624__332329305696010);
  or g_16909 (new_n8276_, not_new_n8253_, not_new_n8219_);
  or g_16910 (new_n3389_, not_pi064_113988951853731430, not_new_n3982__0);
  not g_16911 (not_new_n7211_, new_n7211_);
  or g_16912 (new_n4820_, not_new_n4815_, not_new_n1045__7);
  not g_16913 (not_new_n9489_, new_n9489_);
  or g_16914 (new_n8512_, not_new_n8128__0, not_new_n621__6782230728490);
  not g_16915 (not_new_n3428_, new_n3428_);
  not g_16916 (not_new_n5493_, new_n5493_);
  not g_16917 (not_new_n3879_, new_n3879_);
  or g_16918 (new_n4037_, not_new_n4036_, not_pi054_3);
  not g_16919 (not_new_n9399_, new_n9399_);
  not g_16920 (not_new_n1597__2824752490, new_n1597_);
  not g_16921 (not_new_n7913_, new_n7913_);
  or g_16922 (new_n3843_, not_new_n628__70, not_new_n6443__7);
  or g_16923 (new_n3311_, not_new_n1618_, not_new_n3309_);
  or g_16924 (new_n2055_, not_new_n588__168070, not_pi113);
  not g_16925 (not_new_n8271__2, new_n8271_);
  not g_16926 (not_new_n6608_, new_n6608_);
  or g_16927 (new_n4009_, not_new_n4000_, not_new_n3978_);
  and g_16928 (new_n9855_, new_n10041_, new_n10042_);
  and g_16929 (new_n8208_, new_n8076_, new_n8327_);
  not g_16930 (not_new_n9280_, new_n9280_);
  not g_16931 (new_n7204_, new_n7155_);
  not g_16932 (new_n5751_, new_n1031_);
  not g_16933 (not_new_n2263_, new_n2263_);
  and g_16934 (new_n8678_, new_n8677_, new_n8742_);
  not g_16935 (not_new_n5905__2, new_n5905_);
  not g_16936 (not_new_n1009__4, new_n1009_);
  or g_16937 (new_n8746_, not_new_n8745_, not_new_n8674_);
  or g_16938 (new_n10079_, not_new_n10077_, not_new_n9984_);
  not g_16939 (not_new_n3185__47475615099430, new_n3185_);
  or g_16940 (new_n7487_, not_new_n722__1, not_new_n7448__1);
  not g_16941 (not_new_n3826_, new_n3826_);
  and g_16942 (new_n5729_, new_n6128_, new_n6127_);
  or g_16943 (new_n5801_, not_new_n5787_, not_new_n643__57648010);
  not g_16944 (not_pi018_0, pi018);
  and g_16945 (and_new_n8874__new_n9276_, new_n9276_, new_n8874_);
  not g_16946 (not_new_n8808_, new_n8808_);
  not g_16947 (not_new_n3803_, new_n3803_);
  not g_16948 (new_n5471_, new_n1012_);
  not g_16949 (not_new_n2903_, new_n2903_);
  or g_16950 (new_n4616_, not_pi166_2, not_new_n4424_);
  or g_16951 (new_n4208_, not_new_n4166__0, not_new_n4095_);
  not g_16952 (not_new_n644__113988951853731430, new_n644_);
  not g_16953 (not_new_n599__7, new_n599_);
  not g_16954 (not_new_n3439_, new_n3439_);
  not g_16955 (not_new_n10015_, new_n10015_);
  not g_16956 (not_new_n3427_, new_n3427_);
  or g_16957 (new_n3530_, not_pi131_0, not_new_n1538__1);
  or g_16958 (new_n1985_, not_new_n1584__10, not_new_n9449_);
  or g_16959 (new_n5342_, not_new_n5064_, not_new_n5065_);
  or g_16960 (new_n9707_, not_new_n9424_, not_new_n9336_);
  not g_16961 (not_new_n587__332329305696010, new_n587_);
  not g_16962 (not_new_n1594__7, new_n1594_);
  not g_16963 (not_new_n642__70, new_n642_);
  not g_16964 (not_new_n1589__57648010, new_n1589_);
  not g_16965 (not_new_n1589__968890104070, new_n1589_);
  not g_16966 (not_new_n1163_, new_n1163_);
  not g_16967 (not_new_n6530_, new_n6530_);
  or g_16968 (new_n3579_, not_new_n2280__0, not_new_n1612__47475615099430);
  not g_16969 (not_new_n1295_, new_n1295_);
  or g_16970 (new_n3061_, not_new_n3372__2326305139872070, not_new_n637__4);
  not g_16971 (not_new_n8244__2, new_n8244_);
  not g_16972 (not_new_n663_, new_n663_);
  not g_16973 (not_new_n3657_, new_n3657_);
  not g_16974 (not_new_n624__70, new_n624_);
  not g_16975 (new_n4032_, new_n3948_);
  and g_16976 (po114, key_gate_101, pi093);
  not g_16977 (not_new_n3298_, new_n3298_);
  not g_16978 (not_new_n1588__7, new_n1588_);
  and g_16979 (new_n9986_, new_n10032_, new_n10091_);
  not g_16980 (not_new_n635__332329305696010, new_n635_);
  not g_16981 (new_n9349_, new_n1037_);
  not g_16982 (not_new_n2509__8, new_n2509_);
  not g_16983 (not_new_n8653_, new_n8653_);
  not g_16984 (not_new_n4769_, new_n4769_);
  not g_16985 (not_new_n648__5, new_n648_);
  not g_16986 (not_new_n6883_, new_n6883_);
  or g_16987 (new_n7523_, not_new_n7147_, not_new_n7148__0);
  not g_16988 (new_n2047_, new_n957_);
  or g_16989 (new_n980_, not_new_n2305_, or_or_not_new_n1339__not_new_n1337__not_new_n2306_);
  or g_16990 (new_n7597_, not_new_n634__19773267430, not_new_n7602_);
  or g_16991 (new_n6406_, not_new_n6405_, not_new_n641__24010);
  not g_16992 (not_new_n4807_, new_n4807_);
  not g_16993 (not_new_n1599__3, new_n1599_);
  or g_16994 (new_n2300_, not_new_n585__16284135979104490, not_new_n4072_);
  or g_16995 (new_n4364_, not_new_n4258_, not_new_n663_);
  not g_16996 (not_new_n7403_, new_n7403_);
  not g_16997 (not_pi127_0, pi127);
  not g_16998 (not_pi076, pi076);
  or g_16999 (new_n3184_, not_new_n3183_, not_new_n3182_);
  or g_17000 (or_or_not_new_n6327__not_new_n6373__2_not_new_n1051__490, or_not_new_n6327__not_new_n6373__2, not_new_n1051__490);
  not g_17001 (not_new_n8929_, new_n8929_);
  not g_17002 (not_new_n8738_, new_n8738_);
  or g_17003 (new_n3336_, not_new_n3979__0, not_pi064_9);
  not g_17004 (not_new_n744_, new_n744_);
  not g_17005 (not_new_n3269_, new_n3269_);
  not g_17006 (not_new_n3680_, new_n3680_);
  or g_17007 (new_n7476_, not_new_n7044__0, not_new_n7010__2);
  or g_17008 (new_n2221_, not_new_n4776_, not_new_n591__968890104070);
  not g_17009 (not_new_n6373__6, new_n6373_);
  not g_17010 (not_new_n601__3430, new_n601_);
  or g_17011 (new_n4358_, not_new_n665_, not_new_n4254_);
  or g_17012 (new_n5564_, not_pi142_1, not_new_n5459_);
  and g_17013 (and_new_n8884__new_n9290_, new_n8884_, new_n9290_);
  not g_17014 (not_new_n7488_, new_n7488_);
  and g_17015 (new_n1296_, and_and_new_n2105__new_n2108__new_n2106_, new_n2107_);
  not g_17016 (not_new_n1049__57648010, new_n1049_);
  or g_17017 (new_n3805_, not_new_n3414_, not_new_n1786_);
  not g_17018 (not_new_n4725_, new_n4725_);
  or g_17019 (new_n7465_, not_new_n7156_, or_not_new_n7046__not_new_n7265_);
  not g_17020 (not_new_n9757_, new_n9757_);
  not g_17021 (not_new_n6175_, new_n6175_);
  not g_17022 (not_new_n8101_, new_n8101_);
  and g_17023 (new_n9857_, new_n10089_, new_n10088_);
  not g_17024 (not_new_n1601__13410686196639649008070, new_n1601_);
  or g_17025 (new_n4682_, not_pi175_2, not_new_n4442_);
  and g_17026 (new_n5070_, new_n5371_, new_n5370_);
  not g_17027 (not_new_n4745_, new_n4745_);
  or g_17028 (new_n992_, not_new_n1467_, not_new_n1468_);
  or g_17029 (new_n1781_, not_new_n1776_, not_new_n1216_);
  or g_17030 (new_n6158_, not_new_n5773__0, not_new_n630__8235430);
  not g_17031 (not_new_n1041__7, new_n1041_);
  not g_17032 (not_new_n4510__0, new_n4510_);
  not g_17033 (not_new_n4837__0, new_n4837_);
  not g_17034 (not_new_n1553_, new_n1553_);
  not g_17035 (not_new_n2541_, new_n2541_);
  not g_17036 (not_new_n4192_, new_n4192_);
  or g_17037 (new_n5659_, not_new_n1012__6, not_new_n5470_);
  or g_17038 (new_n9680_, not_new_n626__4599865365447399609768010, not_new_n1053__47475615099430);
  not g_17039 (not_new_n5547_, new_n5547_);
  or g_17040 (new_n3181_, not_new_n935_, or_or_not_new_n934__not_new_n933__0_not_new_n941__0);
  or g_17041 (new_n2224_, not_pi186, not_new_n586__6782230728490);
  not g_17042 (not_new_n1938_, new_n1938_);
  or g_17043 (new_n925_, not_new_n999__0, not_new_n3324_);
  or g_17044 (new_n2563_, not_new_n4466_, not_new_n609__5);
  not g_17045 (not_new_n8255_, new_n8255_);
  not g_17046 (new_n6244_, new_n618_);
  not g_17047 (not_new_n7180_, new_n7180_);
  or g_17048 (new_n4362_, not_new_n695_, not_new_n4259_);
  and g_17049 (and_new_n1330__new_n2274_, new_n2274_, new_n1330_);
  or g_17050 (new_n8305_, not_new_n8118__0, not_new_n1045__6782230728490);
  and g_17051 (and_and_and_new_n1460__new_n1466__new_n1458__new_n1459_, new_n1459_, and_and_new_n1460__new_n1466__new_n1458_);
  not g_17052 (not_new_n4446__0, new_n4446_);
  or g_17053 (new_n2370_, not_new_n598__2, not_new_n1039__0);
  not g_17054 (not_new_n926_, new_n926_);
  not g_17055 (not_new_n9959_, new_n9959_);
  or g_17056 (new_n7267_, not_new_n7139__0, not_new_n7258_);
  not g_17057 (not_new_n6117_, new_n6117_);
  not g_17058 (new_n5753_, new_n1039_);
  not g_17059 (not_new_n6977__0, new_n6977_);
  not g_17060 (not_new_n1059_, new_n1059_);
  or g_17061 (new_n3342_, not_pi064_490, not_new_n3957__0);
  or g_17062 (new_n3688_, not_new_n989__1176490, not_pi230);
  or g_17063 (new_n7555_, not_new_n7554_, not_new_n7553_);
  not g_17064 (not_new_n9966_, new_n9966_);
  or g_17065 (new_n7637_, not_new_n645__2824752490, not_new_n7638_);
  not g_17066 (not_new_n636__47475615099430, new_n636_);
  and g_17067 (new_n8081_, new_n8363_, new_n8176_);
  not g_17068 (not_new_n3458_, new_n3458_);
  not g_17069 (not_new_n7653__0, new_n7653_);
  not g_17070 (not_new_n3936_, new_n3936_);
  or g_17071 (new_n7377_, not_new_n7021__1, not_new_n6978__1);
  not g_17072 (not_new_n10185_, new_n10185_);
  not g_17073 (not_new_n7146__0, new_n7146_);
  not g_17074 (not_new_n8899__0, new_n8899_);
  not g_17075 (not_new_n4759__0, new_n4759_);
  or g_17076 (new_n3939_, not_new_n3940_, not_new_n3999_);
  or g_17077 (new_n9220_, not_new_n9037_, not_new_n9218_);
  not g_17078 (not_new_n8080_, new_n8080_);
  or g_17079 (new_n2902_, not_new_n3310__70, not_pi265_3);
  or g_17080 (new_n7979_, not_new_n7820_, not_new_n7620__1);
  not g_17081 (not_new_n4144_, new_n4144_);
  or g_17082 (new_n9736_, not_new_n9530__0, not_new_n9734_);
  or g_17083 (new_n5151_, new_n644_, new_n1059_);
  not g_17084 (not_new_n10029__2, new_n10029_);
  not g_17085 (not_new_n7602_, new_n7602_);
  not g_17086 (not_new_n626__968890104070, new_n626_);
  not g_17087 (not_new_n1597__16284135979104490, new_n1597_);
  or g_17088 (new_n8010_, not_new_n8009_, not_new_n7928_);
  or g_17089 (new_n6163_, not_new_n625__57648010, not_new_n5774__1);
  not g_17090 (not_new_n1045__9, new_n1045_);
  not g_17091 (not_new_n2186_, new_n2186_);
  not g_17092 (not_new_n647__9, new_n647_);
  or g_17093 (new_n2174_, not_new_n1585__2824752490, not_new_n5833_);
  not g_17094 (new_n6268_, new_n637_);
  or g_17095 (new_n2972_, or_not_new_n2971__not_new_n2970_, not_new_n2969_);
  or g_17096 (new_n9717_, not_new_n9709_, not_new_n9631__0);
  or g_17097 (new_n2413_, not_new_n600__70, not_new_n4135__0);
  not g_17098 (not_new_n1605_, new_n1605_);
  not g_17099 (not_new_n5851_, new_n5851_);
  not g_17100 (not_new_n6482__1, new_n6482_);
  or g_17101 (new_n2804_, not_new_n612__1, not_new_n4127__2);
  or g_17102 (new_n2739_, not_new_n985__0, not_new_n2738_);
  not g_17103 (not_new_n6875_, new_n6875_);
  not g_17104 (not_new_n4507_, new_n4507_);
  or g_17105 (new_n4031_, not_new_n3951_, not_new_n4030__0);
  or g_17106 (new_n9031_, not_new_n9030_, not_new_n8931_);
  not g_17107 (new_n9949_, new_n640_);
  or g_17108 (new_n2144_, not_new_n593__57648010, not_new_n640_);
  not g_17109 (new_n7645_, new_n644_);
  or g_17110 (po294, not_new_n2974_, or_or_or_not_new_n2973__not_new_n2976__not_new_n2975__not_new_n2977_);
  not g_17111 (not_new_n8330_, new_n8330_);
  or g_17112 (new_n10338_, not_new_n9951__2, not_new_n10207_);
  not g_17113 (not_new_n3136_, new_n3136_);
  or g_17114 (new_n3290_, not_new_n643__8, not_new_n3184__19773267430);
  or g_17115 (new_n1902_, not_pi137, not_new_n587__7);
  or g_17116 (new_n6221_, not_new_n5814__0, not_new_n6040_);
  and g_17117 (new_n7708_, new_n7843_, new_n7915_);
  not g_17118 (not_new_n6488_, new_n6488_);
  or g_17119 (or_or_not_new_n2617__not_new_n2621__not_new_n1439_, or_not_new_n2617__not_new_n2621_, not_new_n1439_);
  not g_17120 (not_new_n6235__0, new_n6235_);
  or g_17121 (new_n6553_, not_new_n6915_, not_new_n6916_);
  or g_17122 (new_n2785_, not_new_n613__0, not_new_n1602__1);
  or g_17123 (new_n3842_, not_new_n1576__6, not_new_n623__4);
  or g_17124 (new_n4570_, pi177, new_n1013_);
  not g_17125 (not_new_n9885_, new_n9885_);
  or g_17126 (new_n9087_, new_n1603_, new_n639_);
  not g_17127 (not_new_n9421__0, new_n9421_);
  not g_17128 (new_n8629_, new_n1168_);
  not g_17129 (not_new_n5812_, new_n5812_);
  or g_17130 (new_n2833_, not_pi257_0, not_po296_881247870897231951843937366879128181133112010);
  not g_17131 (not_new_n4735__0, new_n4735_);
  not g_17132 (not_pi043_3, pi043);
  or g_17133 (new_n9178_, not_new_n8899__1, not_new_n8810_);
  or g_17134 (new_n5656_, not_new_n5654_, not_new_n5655_);
  not g_17135 (not_new_n609__1, new_n609_);
  not g_17136 (not_new_n4726__0, new_n4726_);
  or g_17137 (new_n1746_, not_new_n1728__24010, not_pi090);
  not g_17138 (new_n4322_, new_n712_);
  or g_17139 (new_n3715_, not_new_n623__2, not_po298_797922662976120010);
  or g_17140 (new_n9745_, not_new_n1039__797922662976120010, not_new_n9352_);
  not g_17141 (not_new_n10276_, new_n10276_);
  not g_17142 (not_new_n6983_, new_n6983_);
  or g_17143 (new_n8226_, not_new_n8521_, not_new_n8520_);
  not g_17144 (not_new_n1488_, new_n1488_);
  not g_17145 (not_new_n6200_, new_n6200_);
  or g_17146 (new_n5311_, not_new_n624__24010, not_new_n4925_);
  or g_17147 (new_n5402_, not_new_n5400_, not_new_n5163_);
  not g_17148 (not_new_n8376_, new_n8376_);
  not g_17149 (not_new_n6513_, new_n6513_);
  or g_17150 (new_n5462_, not_new_n5564_, not_new_n5563_);
  not g_17151 (new_n6192_, new_n5870_);
  not g_17152 (not_new_n967_, new_n967_);
  not g_17153 (new_n1619_, new_n993_);
  not g_17154 (not_new_n9326__1, new_n9326_);
  not g_17155 (not_new_n642__1176490, new_n642_);
  not g_17156 (not_new_n1534__2, key_gate_5);
  not g_17157 (not_new_n8980_, new_n8980_);
  not g_17158 (not_new_n6740_, new_n6740_);
  not g_17159 (not_new_n1576__47475615099430, new_n1576_);
  or g_17160 (new_n10186_, not_new_n9952__0, not_new_n10185_);
  not g_17161 (not_new_n6017_, new_n6017_);
  not g_17162 (not_new_n3991__0, new_n3991_);
  not g_17163 (not_new_n7513_, new_n7513_);
  not g_17164 (not_new_n5976_, new_n5976_);
  not g_17165 (not_new_n6993__1, new_n6993_);
  not g_17166 (not_new_n4563_, new_n4563_);
  not g_17167 (not_new_n8222_, new_n8222_);
  not g_17168 (not_new_n3916__0, new_n3916_);
  not g_17169 (not_new_n5551_, new_n5551_);
  or g_17170 (or_not_new_n8941__not_new_n8811_, not_new_n8811_, not_new_n8941_);
  and g_17171 (new_n8254_, new_n8510_, new_n8509_);
  not g_17172 (not_new_n9512__0, new_n9512_);
  not g_17173 (not_new_n3862_, new_n3862_);
  and g_17174 (and_new_n6369__new_n6320_, new_n6369_, new_n6320_);
  or g_17175 (new_n7735_, not_new_n7909_, not_new_n7699_);
  or g_17176 (new_n3231_, not_new_n643__7, not_new_n589__19773267430);
  not g_17177 (not_new_n587__968890104070, new_n587_);
  or g_17178 (new_n3368_, not_pi064_6782230728490, not_new_n3985__0);
  not g_17179 (not_new_n10121_, new_n10121_);
  not g_17180 (not_new_n6264_, new_n6264_);
  and g_17181 (new_n5865_, new_n6018_, new_n5719_);
  and g_17182 (new_n1282_, new_n2043_, new_n2044_);
  not g_17183 (not_new_n5317_, new_n5317_);
  or g_17184 (new_n6721_, not_new_n6455_, not_new_n6640_);
  not g_17185 (not_new_n602__332329305696010, new_n602_);
  or g_17186 (po166, not_new_n3559_, not_new_n3558_);
  or g_17187 (new_n4645_, not_new_n4643_, not_new_n4644_);
  or g_17188 (new_n2512_, not_new_n608_, not_new_n1028__5);
  not g_17189 (not_new_n8503_, new_n8503_);
  not g_17190 (not_new_n3310__70, new_n3310_);
  or g_17191 (new_n3227_, not_new_n589__403536070, not_new_n637__7);
  not g_17192 (not_new_n4351_, new_n4351_);
  or g_17193 (new_n8159_, not_new_n8123_, not_new_n647__138412872010);
  not g_17194 (not_new_n1071__57648010, new_n1071_);
  not g_17195 (not_new_n1045__5585458640832840070, new_n1045_);
  or g_17196 (new_n7669_, not_new_n7916_, not_new_n7849_);
  not g_17197 (not_new_n1428_, new_n1428_);
  or g_17198 (new_n1858_, not_new_n594__3, not_new_n9958_);
  not g_17199 (not_new_n5898__0, new_n5898_);
  not g_17200 (not_new_n597__138412872010, new_n597_);
  or g_17201 (new_n8186_, not_new_n8556_, not_new_n8557_);
  not g_17202 (not_new_n6945_, new_n6945_);
  not g_17203 (not_pi004_0, pi004);
  or g_17204 (new_n7145_, not_new_n7166_, not_new_n6987_);
  or g_17205 (new_n8019_, not_new_n1603__8235430, not_new_n7629__0);
  not g_17206 (not_new_n6534_, new_n6534_);
  not g_17207 (not_new_n604__19773267430, new_n604_);
  not g_17208 (not_new_n625__57648010, new_n625_);
  or g_17209 (new_n5810_, not_new_n6053_, not_new_n6004_);
  not g_17210 (not_new_n9373_, new_n9373_);
  or g_17211 (new_n1954_, not_new_n593__8, not_new_n626_);
  not g_17212 (not_new_n1534__1176490, key_gate_5);
  or g_17213 (new_n2482_, not_new_n603__47475615099430, not_new_n617__1);
  or g_17214 (new_n1955_, not_new_n591__9, not_new_n4750_);
  not g_17215 (not_new_n2778_, new_n2778_);
  or g_17216 (new_n7903_, not_new_n7651__1, not_new_n626__16284135979104490);
  or g_17217 (new_n5282_, not_new_n5039_, not_new_n4999__2);
  not g_17218 (not_new_n1585__2, new_n1585_);
  not g_17219 (not_new_n641_, new_n641_);
  not g_17220 (not_new_n602__7, new_n602_);
  or g_17221 (new_n2027_, not_new_n4913_, not_new_n1589__490);
  not g_17222 (not_new_n5794__2, new_n5794_);
  not g_17223 (not_new_n3184__7, new_n3184_);
  or g_17224 (new_n2103_, not_new_n4914_, not_new_n1589__1176490);
  or g_17225 (new_n1922_, not_pi106, not_new_n588__8);
  or g_17226 (new_n6016_, not_new_n5764_, not_new_n618__1176490);
  buf g_17227 (po050, pi214);
  not g_17228 (not_new_n5286__0, new_n5286_);
  or g_17229 (new_n2303_, not_pi126, not_new_n588__16284135979104490);
  not g_17230 (not_pi157_0, pi157);
  not g_17231 (not_new_n1015__0, new_n1015_);
  or g_17232 (new_n7467_, not_new_n7014__1, not_new_n7045__1);
  not g_17233 (not_new_n3185__2326305139872070, new_n3185_);
  not g_17234 (not_new_n9495_, new_n9495_);
  or g_17235 (new_n3541_, not_new_n1612__6, not_new_n1919__0);
  not g_17236 (not_new_n10036_, new_n10036_);
  not g_17237 (not_new_n6683__0, new_n6683_);
  or g_17238 (new_n7528_, not_new_n6992__2, not_new_n7028__0);
  or g_17239 (new_n3486_, not_new_n1613__168070, not_new_n2090_);
  not g_17240 (not_new_n7286_, new_n7286_);
  not g_17241 (not_new_n643__8235430, new_n643_);
  not g_17242 (not_new_n4733__0, new_n4733_);
  or g_17243 (new_n9300_, not_new_n9299_, not_new_n9298_);
  or g_17244 (new_n4389_, not_new_n4277_, not_new_n654_);
  or g_17245 (new_n2768_, not_pi250_3, not_new_n3310__2);
  not g_17246 (not_new_n1585__3430, new_n1585_);
  not g_17247 (new_n9370_, new_n647_);
  not g_17248 (new_n6992_, new_n729_);
  or g_17249 (new_n3300_, not_new_n642__7, not_new_n3184__332329305696010);
  not g_17250 (not_new_n3784_, new_n3784_);
  and g_17251 (and_new_n1334__new_n2293_, new_n1334_, new_n2293_);
  and g_17252 (new_n9498_, new_n9799_, new_n9798_);
  not g_17253 (not_new_n8001_, new_n8001_);
  or g_17254 (new_n7207_, not_new_n7412_, not_new_n6998_);
  or g_17255 (new_n4947_, not_new_n5123_, not_new_n5122_);
  not g_17256 (not_new_n2768_, new_n2768_);
  not g_17257 (not_new_n3749_, new_n3749_);
  not g_17258 (not_new_n5353_, new_n5353_);
  not g_17259 (not_new_n928__16284135979104490, new_n928_);
  not g_17260 (new_n9395_, new_n1059_);
  not g_17261 (not_new_n630__1, new_n630_);
  not g_17262 (not_new_n1604__19773267430, new_n1604_);
  not g_17263 (not_new_n7196_, new_n7196_);
  not g_17264 (not_new_n7630__0, new_n7630_);
  not g_17265 (not_new_n4552_, new_n4552_);
  not g_17266 (not_new_n9844_, new_n9844_);
  or g_17267 (new_n3438_, not_new_n1004__1, not_new_n1594__6);
  not g_17268 (new_n4169_, new_n4100_);
  or g_17269 (new_n5704_, not_new_n5702_, not_new_n5554_);
  not g_17270 (not_new_n8856_, new_n8856_);
  not g_17271 (not_new_n4780_, new_n4780_);
  not g_17272 (not_new_n4117__1, new_n4117_);
  not g_17273 (new_n6297_, new_n1041_);
  not g_17274 (not_new_n9954__0, new_n9954_);
  not g_17275 (not_new_n1013__1, new_n1013_);
  and g_17276 (new_n5499_, new_n5609_, new_n5610_);
  and g_17277 (new_n1542_, new_n3597_, new_n3596_);
  not g_17278 (not_new_n599__403536070, new_n599_);
  not g_17279 (not_new_n5679_, new_n5679_);
  not g_17280 (not_new_n3656_, new_n3656_);
  or g_17281 (new_n8311_, not_new_n8310_, not_new_n8110_);
  not g_17282 (not_new_n7043__0, new_n7043_);
  and g_17283 (new_n8952_, new_n9310_, and_new_n8983__new_n9311_);
  not g_17284 (not_pi143_2, pi143);
  not g_17285 (not_new_n10313_, new_n10313_);
  not g_17286 (not_new_n1043__138412872010, new_n1043_);
  not g_17287 (not_new_n10034__0, new_n10034_);
  not g_17288 (not_new_n1576__8, new_n1576_);
  or g_17289 (new_n5892_, not_new_n6061_, not_new_n6054_);
  not g_17290 (not_new_n1600__0, new_n1600_);
  not g_17291 (not_new_n7029__0, new_n7029_);
  or g_17292 (new_n3549_, not_new_n1995__0, not_new_n1612__10);
  and g_17293 (and_new_n1540__new_n2361_, new_n2361_, new_n1540_);
  not g_17294 (not_new_n1576__10, new_n1576_);
  not g_17295 (not_new_n7604__0, new_n7604_);
  and g_17296 (and_new_n8982__new_n9323_, new_n8982_, new_n9323_);
  not g_17297 (new_n5192_, new_n4988_);
  not g_17298 (not_new_n589__39098210485829880490, new_n589_);
  not g_17299 (not_new_n6882_, new_n6882_);
  not g_17300 (not_new_n640__7, new_n640_);
  or g_17301 (new_n6434_, not_new_n6263_, not_new_n1603__3430);
  or g_17302 (new_n7246_, not_new_n7245_, not_new_n7143_);
  xor g_17303 (key_gate_16, not_new_n3916_, key_16);
  or g_17304 (new_n4855_, not_new_n4844_, not_new_n4757__0);
  not g_17305 (new_n1876_, new_n948_);
  and g_17306 (and_and_new_n6385__new_n6386__new_n6241_, and_new_n6385__new_n6386_, new_n6241_);
  not g_17307 (not_new_n3372__93874803376477543056490, new_n3372_);
  or g_17308 (new_n9966_, not_new_n10313_, not_new_n10312_);
  and g_17309 (new_n1442_, and_new_n2637__new_n2638_, new_n2639_);
  not g_17310 (not_new_n1013__4, new_n1013_);
  or g_17311 (new_n5377_, not_new_n5093_, not_new_n5072_);
  not g_17312 (new_n3980_, pi064);
  not g_17313 (new_n4940_, new_n1049_);
  or g_17314 (new_n2587_, not_new_n2586_, not_new_n611__70);
  not g_17315 (not_pi174_2, pi174);
  or g_17316 (new_n10185_, new_n1057_, new_n636_);
  or g_17317 (new_n9023_, not_new_n1037__19773267430, not_new_n632__47475615099430);
  or g_17318 (new_n9104_, not_new_n1597__6782230728490, not_new_n617__113988951853731430);
  not g_17319 (not_new_n1584__3430, new_n1584_);
  not g_17320 (not_new_n6827_, new_n6827_);
  buf g_17321 (po047, pi217);
  not g_17322 (not_pi247_0, pi247);
  not g_17323 (not_new_n8005_, new_n8005_);
  or g_17324 (new_n3041_, not_new_n1027__2824752490, not_new_n1166_);
  not g_17325 (not_new_n1168_, new_n1168_);
  not g_17326 (not_new_n8710_, new_n8710_);
  not g_17327 (not_new_n4221_, new_n4221_);
  or g_17328 (new_n9844_, not_new_n9668__0, not_new_n9842_);
  not g_17329 (not_new_n6157_, new_n6157_);
  or g_17330 (new_n7235_, not_new_n7436_, not_new_n7007_);
  not g_17331 (not_new_n7663_, new_n7663_);
  not g_17332 (not_new_n7169_, new_n7169_);
  or g_17333 (new_n2177_, not_new_n6566_, not_new_n1580__19773267430);
  not g_17334 (not_new_n587__7, new_n587_);
  not g_17335 (new_n4549_, new_n4506_);
  not g_17336 (not_new_n8185_, new_n8185_);
  not g_17337 (not_new_n1616__8, new_n1616_);
  not g_17338 (not_new_n8887__0, new_n8887_);
  not g_17339 (not_new_n5469__0, new_n5469_);
  or g_17340 (new_n7027_, not_new_n7346_, not_new_n7347_);
  not g_17341 (not_new_n928__6, new_n928_);
  not g_17342 (not_new_n617__19773267430, new_n617_);
  not g_17343 (not_new_n5903_, new_n5903_);
  not g_17344 (not_new_n1380_, new_n1380_);
  or g_17345 (po187, or_not_new_n1544__not_new_n1358_, not_new_n1357_);
  not g_17346 (not_new_n9970_, new_n9970_);
  not g_17347 (not_new_n618__13410686196639649008070, new_n618_);
  not g_17348 (not_new_n5044_, new_n5044_);
  not g_17349 (not_new_n8291_, new_n8291_);
  not g_17350 (new_n6266_, new_n646_);
  not g_17351 (not_new_n1585__2326305139872070, new_n1585_);
  not g_17352 (not_new_n6258_, new_n6258_);
  not g_17353 (not_new_n8377_, new_n8377_);
  not g_17354 (not_new_n9379__0, new_n9379_);
  not g_17355 (not_new_n3196_, new_n3196_);
  not g_17356 (not_new_n4083_, new_n4083_);
  not g_17357 (not_new_n1613__490, new_n1613_);
  not g_17358 (not_pi025_0, pi025);
  not g_17359 (not_new_n1726_, key_gate_23);
  or g_17360 (new_n8002_, not_new_n1599__168070, not_new_n7623__0);
  not g_17361 (not_new_n4929_, new_n4929_);
  or g_17362 (new_n2827_, not_new_n4118__1, not_new_n994__490);
  or g_17363 (new_n675_, not_new_n3098_, or_not_new_n3100__not_new_n3099_);
  not g_17364 (not_new_n5683_, new_n5683_);
  not g_17365 (not_new_n585__4, new_n585_);
  not g_17366 (not_new_n2227_, new_n2227_);
  and g_17367 (new_n6455_, new_n6448_, new_n6719_);
  or g_17368 (new_n2781_, not_new_n639__2, not_new_n604__5);
  not g_17369 (new_n9946_, new_n1596_);
  not g_17370 (new_n4772_, new_n1600_);
  or g_17371 (new_n2475_, not_new_n598__968890104070, not_new_n1600__0);
  or g_17372 (new_n4211_, not_pi259_1, not_new_n4149_);
  not g_17373 (not_new_n1536__10, new_n1536_);
  not g_17374 (new_n4426_, new_n1005_);
  or g_17375 (new_n3908_, not_new_n643__3430, not_new_n9929_);
  and g_17376 (new_n1412_, pi275, new_n998_);
  not g_17377 (not_new_n1631__6782230728490, key_gate_76);
  or g_17378 (new_n4554_, new_n1017_, pi173);
  not g_17379 (not_new_n4189_, new_n4189_);
  and g_17380 (new_n1364_, new_n2396_, new_n2395_);
  and g_17381 (new_n8698_, new_n8777_, new_n8778_);
  or g_17382 (new_n5954_, not_new_n5921__0, not_new_n5740__1);
  not g_17383 (not_new_n1602__16284135979104490, new_n1602_);
  not g_17384 (not_new_n4723_, new_n4723_);
  not g_17385 (not_new_n9712_, new_n9712_);
  or g_17386 (new_n5893_, not_new_n5771_, not_new_n1602__70);
  not g_17387 (not_new_n609__5, new_n609_);
  or g_17388 (po131, not_new_n3471_, not_new_n3470_);
  not g_17389 (not_new_n1583__47475615099430, new_n1583_);
  not g_17390 (not_new_n1067__332329305696010, new_n1067_);
  not g_17391 (not_new_n1537__2326305139872070, new_n1537_);
  not g_17392 (new_n1596_, new_n979_);
  or g_17393 (new_n7394_, not_new_n7393_, not_new_n7392_);
  not g_17394 (not_new_n6975_, new_n6975_);
  not g_17395 (not_new_n9240_, new_n9240_);
  not g_17396 (not_new_n2854_, new_n2854_);
  or g_17397 (or_not_new_n2625__not_new_n2624_, not_new_n2624_, not_new_n2625_);
  not g_17398 (not_new_n7133_, new_n7133_);
  not g_17399 (not_new_n3472_, new_n3472_);
  not g_17400 (not_new_n1580__10, new_n1580_);
  not g_17401 (not_new_n1881_, new_n1881_);
  not g_17402 (new_n4013_, new_n3955_);
  not g_17403 (not_new_n632__24010, new_n632_);
  not g_17404 (not_new_n7550_, new_n7550_);
  or g_17405 (new_n7498_, not_new_n7496_, not_new_n7244_);
  or g_17406 (new_n4454_, not_new_n4600_, not_new_n4599_);
  not g_17407 (not_new_n4831__1, new_n4831_);
  not g_17408 (not_new_n5664_, new_n5664_);
  or g_17409 (new_n3199_, not_new_n589__5, not_new_n628__7);
  not g_17410 (not_pi200, pi200);
  or g_17411 (new_n5327_, not_new_n5326_, not_new_n5325_);
  not g_17412 (not_new_n5015_, new_n5015_);
  not g_17413 (not_new_n1053__0, new_n1053_);
  not g_17414 (not_new_n1536_, new_n1536_);
  or g_17415 (new_n1641_, not_pi029, not_po296_2);
  or g_17416 (new_n3604_, not_pi168_0, not_new_n984__6);
  not g_17417 (not_new_n9870_, new_n9870_);
  and g_17418 (new_n7577_, and_new_n7791__new_n7786_, new_n7773_);
  or g_17419 (new_n1827_, not_pi101, not_new_n588__3);
  or g_17420 (new_n9123_, new_n645_, new_n1071_);
  and g_17421 (new_n1457_, new_n2700_, and_new_n2702__new_n2701_);
  or g_17422 (new_n4739_, or_not_new_n4825__not_new_n4804_, not_new_n4807_);
  not g_17423 (not_new_n10009_, new_n10009_);
  or g_17424 (new_n5283_, not_new_n5190_, not_new_n4995_);
  not g_17425 (not_po296_3, po296);
  not g_17426 (not_new_n6561_, new_n6561_);
  not g_17427 (not_new_n2340_, new_n2340_);
  not g_17428 (not_new_n9386_, new_n9386_);
  or g_17429 (new_n9755_, not_new_n9754_, not_new_n9753_);
  not g_17430 (not_new_n637__2, new_n637_);
  not g_17431 (not_new_n3685_, new_n3685_);
  not g_17432 (not_new_n8277_, new_n8277_);
  not g_17433 (not_new_n5318_, new_n5318_);
  not g_17434 (not_new_n5211_, new_n5211_);
  not g_17435 (not_new_n10138_, new_n10138_);
  or g_17436 (new_n3757_, not_new_n1600__6, not_new_n629__10);
  or g_17437 (new_n6771_, not_new_n6527__0, not_new_n626__968890104070);
  not g_17438 (not_new_n5919__0, new_n5919_);
  not g_17439 (not_new_n589__26517308458596534717790233816010, new_n589_);
  not g_17440 (not_new_n586__16284135979104490, new_n586_);
  not g_17441 (not_new_n2784_, new_n2784_);
  or g_17442 (or_not_new_n9103__not_new_n8987__0, not_new_n8987__0, not_new_n9103_);
  or g_17443 (new_n9394_, not_new_n627__332329305696010, not_new_n1055__797922662976120010);
  or g_17444 (new_n2035_, not_pi144, not_new_n587__24010);
  and g_17445 (new_n1460_, and_and_new_n3792__new_n3795__new_n3801_, new_n3798_);
  not g_17446 (not_new_n2696_, new_n2696_);
  not g_17447 (not_new_n1602__490, new_n1602_);
  not g_17448 (not_new_n1002__6, new_n1002_);
  not g_17449 (not_new_n1576__168070, new_n1576_);
  not g_17450 (not_new_n1596__2824752490, new_n1596_);
  not g_17451 (not_new_n5597__0, new_n5597_);
  not g_17452 (not_new_n7867_, new_n7867_);
  or g_17453 (new_n1053_, not_new_n3453_, not_new_n3452_);
  not g_17454 (not_new_n1642_, key_gate_100);
  or g_17455 (new_n3610_, not_pi171_0, not_new_n984__9);
  not g_17456 (not_new_n4424__0, new_n4424_);
  not g_17457 (not_new_n4749_, new_n4749_);
  not g_17458 (not_new_n7995_, new_n7995_);
  not g_17459 (not_new_n10283_, new_n10283_);
  or g_17460 (new_n3538_, not_pi135_0, not_new_n1538__5);
  or g_17461 (new_n2935_, not_new_n4071__1, not_new_n994__6782230728490);
  not g_17462 (not_new_n6885_, new_n6885_);
  not g_17463 (not_new_n1053__490, new_n1053_);
  not g_17464 (not_new_n10186_, new_n10186_);
  not g_17465 (not_new_n6872_, new_n6872_);
  not g_17466 (not_new_n8140__0, new_n8140_);
  or g_17467 (new_n2135_, not_new_n7679_, not_new_n1583__57648010);
  or g_17468 (new_n3626_, not_new_n984__8235430, not_pi179_0);
  or g_17469 (new_n5732_, not_new_n6089_, or_or_not_new_n6160__not_new_n6161__not_new_n6090_);
  not g_17470 (not_new_n593__9, new_n593_);
  not g_17471 (not_new_n989__9, new_n989_);
  and g_17472 (and_and_new_n2048__new_n2051__new_n2049_, new_n2049_, and_new_n2048__new_n2051_);
  or g_17473 (new_n9258_, not_new_n8886__0, not_new_n630__332329305696010);
  not g_17474 (not_pi040, pi040);
  not g_17475 (not_new_n633__39098210485829880490, new_n633_);
  not g_17476 (not_new_n1616__332329305696010, new_n1616_);
  not g_17477 (not_new_n3438_, new_n3438_);
  not g_17478 (not_new_n10007_, new_n10007_);
  not g_17479 (not_new_n8828_, new_n8828_);
  not g_17480 (new_n8883_, new_n633_);
  or g_17481 (new_n7667_, not_new_n7859_, not_new_n7920_);
  not g_17482 (not_new_n638__138412872010, new_n638_);
  or g_17483 (new_n5921_, not_new_n5739_, not_new_n1047__70);
  not g_17484 (not_new_n8244__3, new_n8244_);
  and g_17485 (new_n1468_, new_n1461_, and_and_and_new_n1460__new_n1466__new_n1458__new_n1459_);
  or g_17486 (new_n10234_, not_new_n9991_, not_new_n9951__1);
  and g_17487 (and_new_n3768__new_n3771_, new_n3771_, new_n3768_);
  not g_17488 (not_new_n587__8, new_n587_);
  or g_17489 (new_n6759_, not_new_n6508__0, not_new_n6737__0);
  not g_17490 (not_new_n8799__1, new_n8799_);
  or g_17491 (new_n10006_, not_new_n10223_, not_new_n10213_);
  not g_17492 (new_n8307_, new_n8122_);
  or g_17493 (new_n2968_, not_pi272_0, not_po296_4183778472590916451475308348590993345191760458870147715430);
  or g_17494 (new_n3297_, not_new_n1053__6, not_new_n589__152867006319425761937651857692768264010);
  not g_17495 (not_new_n5231_, new_n5231_);
  not g_17496 (not_new_n7004__1, new_n7004_);
  not g_17497 (not_new_n701_, new_n701_);
  not g_17498 (not_new_n1004__6, new_n1004_);
  or g_17499 (new_n2589_, not_po296_32199057558131797268376070, not_pi251);
  or g_17500 (new_n10274_, not_new_n9946_, not_new_n618__32199057558131797268376070);
  not g_17501 (not_new_n3718_, new_n3718_);
  not g_17502 (not_new_n4748_, new_n4748_);
  not g_17503 (not_new_n603__10, new_n603_);
  or g_17504 (new_n4610_, not_new_n1005__4, not_new_n4425__0);
  or g_17505 (new_n7237_, not_new_n6964_, not_new_n7163_);
  not g_17506 (new_n8117_, new_n1039_);
  or g_17507 (new_n9690_, not_new_n9406__0, not_new_n9614__0);
  not g_17508 (not_new_n3975_, new_n3975_);
  or g_17509 (new_n4186_, not_new_n4075_, not_new_n4153_);
  or g_17510 (new_n700_, not_new_n3072_, not_new_n1524_);
  or g_17511 (new_n9051_, new_n644_, new_n1059_);
  not g_17512 (not_new_n1600__4, new_n1600_);
  not g_17513 (not_new_n4175_, new_n4175_);
  not g_17514 (not_new_n3372__3, new_n3372_);
  not g_17515 (not_new_n8338_, new_n8338_);
  not g_17516 (not_new_n1594__10, new_n1594_);
  not g_17517 (not_new_n7657__0, new_n7657_);
  not g_17518 (not_new_n1012__2, new_n1012_);
  not g_17519 (not_new_n6498_, new_n6498_);
  not g_17520 (not_new_n7683_, new_n7683_);
  and g_17521 (new_n1359_, new_n2382_, and_new_n2384__new_n2383_);
  not g_17522 (not_new_n7475_, new_n7475_);
  not g_17523 (not_new_n629__8235430, new_n629_);
  or g_17524 (new_n3598_, not_pi165_0, not_new_n984__3);
  not g_17525 (not_new_n630__403536070, new_n630_);
  not g_17526 (new_n8612_, new_n1063_);
  not g_17527 (not_new_n8830__1, new_n8830_);
  not g_17528 (not_new_n9390_, new_n9390_);
  not g_17529 (not_new_n1600__1, new_n1600_);
  not g_17530 (not_new_n3931__0, key_gate_6);
  not g_17531 (not_new_n1601__57648010, new_n1601_);
  not g_17532 (not_new_n3250_, new_n3250_);
  or g_17533 (new_n7955_, not_new_n648__6782230728490, not_new_n7603__1);
  not g_17534 (new_n9889_, new_n1043_);
  not g_17535 (not_new_n8410_, new_n8410_);
  not g_17536 (not_new_n1580__403536070, new_n1580_);
  and g_17537 (new_n1432_, new_n2589_, new_n2588_);
  not g_17538 (not_new_n5746__1, new_n5746_);
  and g_17539 (and_new_n2379__new_n2378_, new_n2378_, new_n2379_);
  not g_17540 (not_new_n6995__1, new_n6995_);
  or g_17541 (new_n3344_, not_pi064_3430, not_new_n3921__0);
  not g_17542 (not_pi132_2, pi132);
  not g_17543 (not_new_n2275_, new_n2275_);
  or g_17544 (new_n2340_, not_pi160, not_new_n587__797922662976120010);
  not g_17545 (new_n10009_, new_n1607_);
  not g_17546 (not_new_n1158_, new_n1158_);
  not g_17547 (new_n7101_, new_n773_);
  or g_17548 (new_n9190_, not_new_n8851_, not_new_n8984__1);
  or g_17549 (new_n8365_, not_new_n8138_, not_new_n625__2326305139872070);
  not g_17550 (not_new_n5491__0, new_n5491_);
  not g_17551 (not_new_n5796__0, new_n5796_);
  not g_17552 (not_new_n581__2824752490, new_n581_);
  or g_17553 (or_not_new_n1295__not_new_n1293_, not_new_n1295_, not_new_n1293_);
  or g_17554 (or_or_not_new_n6334__not_new_n6232__0_not_new_n6235__0, not_new_n6235__0, or_not_new_n6334__not_new_n6232__0);
  not g_17555 (not_new_n7480_, new_n7480_);
  not g_17556 (not_new_n8835_, new_n8835_);
  not g_17557 (not_new_n9347_, new_n9347_);
  not g_17558 (not_new_n8107__0, new_n8107_);
  not g_17559 (not_new_n1426_, new_n1426_);
  not g_17560 (not_new_n3779_, new_n3779_);
  not g_17561 (not_new_n3372__24010, new_n3372_);
  or g_17562 (new_n2146_, not_new_n1071_, not_new_n1588__403536070);
  not g_17563 (not_new_n3884_, new_n3884_);
  and g_17564 (new_n5863_, new_n6002_, new_n5727_);
  not g_17565 (not_new_n9846_, new_n9846_);
  not g_17566 (not_new_n1538__138412872010, new_n1538_);
  not g_17567 (not_new_n7203_, new_n7203_);
  not g_17568 (not_new_n638__4599865365447399609768010, new_n638_);
  not g_17569 (not_new_n2504_, new_n2504_);
  xor g_17570 (key_gate_126, not_new_n3919_, key_126);
  not g_17571 (not_new_n3185__332329305696010, new_n3185_);
  not g_17572 (not_new_n10145_, new_n10145_);
  or g_17573 (new_n3420_, not_new_n1537__2, not_pi100_0);
  not g_17574 (new_n4830_, new_n4795_);
  or g_17575 (new_n4198_, not_new_n4105_, not_new_n4171__0);
  not g_17576 (not_new_n628__2326305139872070, new_n628_);
  and g_17577 (new_n1260_, and_and_new_n1934__new_n1937__new_n1935_, new_n1936_);
  not g_17578 (not_new_n587__403536070, new_n587_);
  not g_17579 (new_n4419_, pi164);
  not g_17580 (not_new_n7108_, new_n7108_);
  and g_17581 (new_n1519_, new_n3056_, and_new_n3058__new_n998_);
  not g_17582 (not_new_n648__332329305696010, new_n648_);
  not g_17583 (not_new_n3725_, new_n3725_);
  not g_17584 (new_n4561_, new_n4500_);
  or g_17585 (new_n3289_, not_new_n589__63668057609090279857414351392240010, not_new_n1061__5);
  not g_17586 (not_new_n6496__1, new_n6496_);
  and g_17587 (and_new_n9905__new_n10320_, new_n9905_, new_n10320_);
  and g_17588 (new_n6456_, new_n6737_, new_n6450_);
  not g_17589 (not_new_n617__1176490, new_n617_);
  or g_17590 (new_n1891_, not_new_n8100_, not_new_n1581__5);
  not g_17591 (not_new_n10336_, new_n10336_);
  and g_17592 (new_n1501_, new_n3024_, new_n998_);
  or g_17593 (new_n9572_, new_n626_, new_n1053_);
  or g_17594 (new_n9321_, not_new_n9050_, not_new_n9319_);
  and g_17595 (new_n9340_, new_n9678_, new_n9681_);
  not g_17596 (not_pi003, pi003);
  not g_17597 (not_new_n6814_, new_n6814_);
  not g_17598 (not_new_n6774_, new_n6774_);
  not g_17599 (not_new_n631__2326305139872070, new_n631_);
  or g_17600 (new_n5200_, new_n621_, new_n1598_);
  not g_17601 (not_new_n9923_, new_n9923_);
  not g_17602 (not_new_n1607__5, new_n1607_);
  not g_17603 (not_new_n633__403536070, new_n633_);
  or g_17604 (new_n5292_, not_new_n4943_, not_new_n647__24010);
  not g_17605 (new_n8164_, new_n643_);
  or g_17606 (new_n2439_, not_new_n599__1176490, not_new_n9869__0);
  not g_17607 (not_new_n9556_, new_n9556_);
  not g_17608 (not_new_n631__19773267430, new_n631_);
  not g_17609 (not_new_n8114_, new_n8114_);
  not g_17610 (not_new_n4485__0, new_n4485_);
  or g_17611 (new_n10246_, not_new_n634__273687473400809163430, not_new_n9880__0);
  not g_17612 (not_new_n630__6, new_n630_);
  not g_17613 (not_new_n5885_, new_n5885_);
  not g_17614 (not_new_n8290_, new_n8290_);
  or g_17615 (new_n4056_, not_new_n3981__1, not_new_n4019__1);
  or g_17616 (new_n9027_, not_new_n1039__47475615099430, not_new_n628__113988951853731430);
  not g_17617 (not_new_n622__1, new_n622_);
  or g_17618 (new_n10263_, not_new_n10007_, not_new_n10202_);
  not g_17619 (not_new_n2056_, new_n2056_);
  not g_17620 (not_pi253_1, pi253);
  not g_17621 (not_new_n1071__0, new_n1071_);
  and g_17622 (new_n1213_, new_n1769_, new_n1770_);
  not g_17623 (not_new_n8424_, new_n8424_);
  not g_17624 (not_new_n648__39098210485829880490, new_n648_);
  or g_17625 (new_n8029_, not_new_n7752__1, not_new_n642__138412872010);
  not g_17626 (not_new_n1055__0, new_n1055_);
  and g_17627 (and_new_n2707__new_n2708_, new_n2707_, new_n2708_);
  not g_17628 (not_new_n1063__0, new_n1063_);
  or g_17629 (or_or_not_new_n1882__not_new_n1883__not_new_n1885_, or_not_new_n1882__not_new_n1883_, not_new_n1885_);
  not g_17630 (not_new_n5947_, new_n5947_);
  not g_17631 (not_new_n586__2824752490, new_n586_);
  not g_17632 (not_pi177, pi177);
  not g_17633 (not_new_n3853_, new_n3853_);
  or g_17634 (new_n9034_, not_new_n8932_, not_new_n9032_);
  not g_17635 (not_new_n638__2326305139872070, new_n638_);
  not g_17636 (not_new_n581__21838143759917965991093122527538323430, new_n581_);
  or g_17637 (new_n5179_, not_new_n1604__8, not_new_n5178_);
  or g_17638 (new_n2546_, or_not_new_n2545__not_new_n2544_, not_new_n2543_);
  not g_17639 (not_new_n2419_, new_n2419_);
  not g_17640 (not_pi270, pi270);
  or g_17641 (or_not_new_n2827__not_new_n2826_, not_new_n2826_, not_new_n2827_);
  or g_17642 (new_n5969_, not_new_n627__1176490, not_new_n5793_);
  or g_17643 (new_n1008_, not_new_n3338_, not_new_n3337_);
  not g_17644 (not_new_n1071__7, new_n1071_);
  or g_17645 (new_n8463_, not_new_n8105__1, not_new_n1049__19773267430);
  not g_17646 (not_new_n6976__1, new_n6976_);
  not g_17647 (not_new_n6994__1, new_n6994_);
  not g_17648 (new_n8834_, new_n1045_);
  or g_17649 (new_n7773_, not_new_n1043__168070, not_new_n7612_);
  or g_17650 (po156, not_new_n3538_, not_new_n3539_);
  and g_17651 (new_n582_, new_n1023_, new_n1578_);
  or g_17652 (new_n7504_, not_new_n7305_, not_new_n7015__0);
  not g_17653 (new_n6298_, new_n1037_);
  not g_17654 (not_new_n1631__5, key_gate_76);
  not g_17655 (not_new_n7040__1, new_n7040_);
  not g_17656 (not_pi006_0, pi006);
  or g_17657 (new_n7817_, not_new_n7773__1, not_new_n7816_);
  or g_17658 (new_n8069_, not_new_n1055__968890104070, not_new_n7648__2);
  or g_17659 (new_n8195_, not_new_n8514_, not_new_n8513_);
  or g_17660 (new_n9909_, not_new_n646__16284135979104490, not_new_n1069__6782230728490);
  or g_17661 (new_n3461_, not_new_n1613__10, not_new_n1995_);
  not g_17662 (not_new_n7454__1, new_n7454_);
  not g_17663 (not_new_n1589__9, new_n1589_);
  not g_17664 (not_new_n9707_, new_n9707_);
  or g_17665 (new_n4854_, not_new_n4758_, not_new_n1606__4);
  and g_17666 (and_new_n2086__new_n2089_, new_n2089_, new_n2086_);
  or g_17667 (new_n8343_, not_new_n8152_, not_new_n1059__403536070);
  not g_17668 (not_new_n646__1, new_n646_);
  not g_17669 (not_new_n7415__0, new_n7415_);
  not g_17670 (not_new_n589__13410686196639649008070, new_n589_);
  not g_17671 (not_new_n4460_, new_n4460_);
  or g_17672 (new_n3746_, not_new_n975_, not_new_n2247_);
  or g_17673 (new_n5590_, not_pi138_2, not_new_n5450_);
  or g_17674 (new_n6563_, not_new_n6860_, not_new_n6859_);
  or g_17675 (or_not_new_n3397__not_new_n3398_, not_new_n3397_, not_new_n3398_);
  buf g_17676 (po003, pi196);
  or g_17677 (new_n2453_, not_new_n4127__0, not_new_n600__403536070);
  and g_17678 (new_n1289_, new_n2079_, new_n2080_);
  not g_17679 (not_pi126_0, pi126);
  not g_17680 (new_n9400_, new_n1071_);
  and g_17681 (new_n1286_, new_n2062_, new_n2063_);
  or g_17682 (new_n8784_, not_new_n8713__0, not_new_n8702_);
  or g_17683 (new_n5177_, new_n1603_, new_n639_);
  or g_17684 (new_n3119_, not_new_n621__5, not_new_n3315__70);
  or g_17685 (new_n5573_, not_new_n5513_, not_new_n5572_);
  or g_17686 (new_n4394_, not_new_n653_, not_new_n4278_);
  not g_17687 (not_new_n8796_, new_n8796_);
  or g_17688 (new_n6550_, not_new_n6888_, not_new_n6887_);
  and g_17689 (new_n1513_, new_n998_, new_n3042_);
  xor g_17690 (key_gate_30, key_30, not_new_n3920_);
  not g_17691 (not_new_n1067__6, new_n1067_);
  not g_17692 (not_new_n3548_, new_n3548_);
  or g_17693 (po136, not_new_n3496_, not_new_n3495_);
  not g_17694 (not_new_n4800_, new_n4800_);
  not g_17695 (not_new_n609__6, new_n609_);
  and g_17696 (and_and_new_n6227__new_n6232__new_n6229_, new_n6229_, and_new_n6227__new_n6232_);
  not g_17697 (not_new_n10002_, new_n10002_);
  or g_17698 (new_n7181_, not_new_n6978_, not_new_n7363_);
  not g_17699 (not_new_n4129_, new_n4129_);
  not g_17700 (not_new_n4607_, new_n4607_);
  not g_17701 (not_new_n6519_, new_n6519_);
  not g_17702 (not_new_n1536__8, new_n1536_);
  or g_17703 (new_n7755_, not_new_n7708_, not_new_n7914_);
  not g_17704 (new_n4840_, new_n4768_);
  not g_17705 (not_new_n7656_, new_n7656_);
  not g_17706 (not_new_n1990_, new_n1990_);
  not g_17707 (not_new_n5308_, new_n5308_);
  not g_17708 (not_new_n4933_, new_n4933_);
  not g_17709 (new_n4438_, new_n1017_);
  not g_17710 (not_new_n1922_, new_n1922_);
  not g_17711 (not_new_n6067_, new_n6067_);
  or g_17712 (new_n10313_, not_new_n10311_, not_new_n10235_);
  and g_17713 (new_n1312_, and_and_new_n2181__new_n2184__new_n2182_, new_n2183_);
  not g_17714 (not_new_n3414_, new_n3414_);
  not g_17715 (not_new_n3574_, new_n3574_);
  not g_17716 (not_pi121, pi121);
  and g_17717 (new_n7721_, new_n7881_, new_n7576_);
  or g_17718 (new_n9724_, not_new_n9722_, not_new_n9541__0);
  or g_17719 (new_n962_, not_new_n2134_, or_or_not_new_n1303__not_new_n1301__not_new_n2135_);
  not g_17720 (not_new_n638__6, new_n638_);
  not g_17721 (not_new_n6691_, new_n6691_);
  not g_17722 (not_new_n8597_, new_n8597_);
  not g_17723 (not_new_n7801__0, new_n7801_);
  or g_17724 (new_n7803_, not_new_n7597__0, not_new_n7795_);
  not g_17725 (not_new_n3876_, new_n3876_);
  or g_17726 (new_n3138_, not_new_n1604__3, not_new_n928__8235430);
  or g_17727 (or_not_new_n9893__not_new_n9890__0, not_new_n9890__0, not_new_n9893_);
  not g_17728 (not_new_n7825_, new_n7825_);
  not g_17729 (not_new_n1059__47475615099430, new_n1059_);
  not g_17730 (not_new_n8023_, new_n8023_);
  not g_17731 (not_new_n8063_, new_n8063_);
  not g_17732 (not_new_n7312_, new_n7312_);
  or g_17733 (new_n622_, or_or_not_new_n2227__not_new_n2224__not_new_n2225_, not_new_n2226_);
  not g_17734 (new_n5815_, new_n641_);
  or g_17735 (new_n2873_, not_new_n2870_, or_not_new_n2872__not_new_n2871_);
  not g_17736 (not_new_n2439_, new_n2439_);
  not g_17737 (not_new_n9371_, new_n9371_);
  not g_17738 (not_new_n6223__0, new_n6223_);
  or g_17739 (new_n4691_, not_pi174_3, not_new_n4440__0);
  or g_17740 (or_or_not_new_n1247__not_new_n1245__not_new_n1869_, or_not_new_n1247__not_new_n1245_, not_new_n1869_);
  or g_17741 (or_not_new_n6348__not_new_n6232__2, not_new_n6232__2, not_new_n6348_);
  not g_17742 (not_pi183, pi183);
  or g_17743 (new_n9955_, not_new_n10239_, not_new_n10240_);
  or g_17744 (or_or_not_new_n1239__not_new_n1237__not_new_n1831_, not_new_n1831_, or_not_new_n1239__not_new_n1237_);
  not g_17745 (not_new_n7928_, new_n7928_);
  not g_17746 (not_new_n4155__0, new_n4155_);
  not g_17747 (not_pi062_0, pi062);
  not g_17748 (not_new_n7315_, new_n7315_);
  or g_17749 (new_n10190_, not_new_n10188_, not_new_n10003_);
  not g_17750 (not_new_n1043__7, new_n1043_);
  not g_17751 (not_new_n638__19773267430, new_n638_);
  not g_17752 (new_n4982_, new_n637_);
  not g_17753 (not_new_n1914_, new_n1914_);
  or g_17754 (new_n4591_, not_new_n4589_, not_new_n4590_);
  not g_17755 (not_pi035_2, pi035);
  not g_17756 (not_new_n6478__0, new_n6478_);
  or g_17757 (new_n5586_, new_n1011_, pi147);
  or g_17758 (new_n2812_, not_new_n3311__5, not_new_n1031__4);
  not g_17759 (not_new_n8168_, new_n8168_);
  or g_17760 (new_n9603_, new_n1604_, new_n640_);
  not g_17761 (not_new_n4215_, new_n4215_);
  and g_17762 (and_new_n10034__new_n10289_, new_n10289_, new_n10034_);
  not g_17763 (not_new_n7372_, new_n7372_);
  not g_17764 (not_new_n6089_, new_n6089_);
  not g_17765 (not_new_n3387__0, new_n3387_);
  not g_17766 (not_new_n9305_, new_n9305_);
  or g_17767 (new_n3539_, not_new_n1612__5, not_new_n1900__0);
  not g_17768 (not_new_n9801_, new_n9801_);
  not g_17769 (not_new_n2318__0, new_n2318_);
  or g_17770 (new_n9888_, not_new_n1041__6782230728490, not_new_n624__16284135979104490);
  not g_17771 (not_pi190, pi190);
  not g_17772 (not_new_n3310__1, new_n3310_);
  or g_17773 (new_n3260_, not_new_n3184__6, not_new_n618__7);
  not g_17774 (not_new_n3422_, new_n3422_);
  not g_17775 (not_new_n640__2, new_n640_);
  and g_17776 (new_n1186_, new_n1649_, new_n1647_);
  not g_17777 (not_new_n8386_, new_n8386_);
  not g_17778 (not_new_n2850_, new_n2850_);
  not g_17779 (not_new_n1016__4, new_n1016_);
  not g_17780 (not_new_n8477_, new_n8477_);
  not g_17781 (not_new_n9652_, new_n9652_);
  not g_17782 (not_new_n8593_, new_n8593_);
  or g_17783 (new_n9324_, not_new_n641__403536070, not_new_n8831_);
  or g_17784 (new_n7551_, not_new_n7308_, not_new_n7017__0);
  or g_17785 (new_n4609_, not_new_n4426_, not_pi167_2);
  not g_17786 (not_pi147, pi147);
  not g_17787 (not_new_n3512_, new_n3512_);
  or g_17788 (new_n672_, or_not_new_n3091__not_new_n3090_, not_new_n3089_);
  not g_17789 (not_new_n776_, new_n776_);
  not g_17790 (not_new_n589__47475615099430, new_n589_);
  not g_17791 (not_new_n7326_, new_n7326_);
  not g_17792 (not_new_n7634__0, new_n7634_);
  not g_17793 (not_new_n6865_, new_n6865_);
  or g_17794 (new_n3264_, not_new_n621__8, not_new_n3184__8);
  not g_17795 (new_n10046_, new_n9890_);
  not g_17796 (not_new_n1602__0, new_n1602_);
  not g_17797 (not_new_n1053__3, new_n1053_);
  not g_17798 (not_new_n8896_, new_n8896_);
  not g_17799 (not_new_n8746_, new_n8746_);
  not g_17800 (not_pi166_0, pi166);
  not g_17801 (not_new_n7641_, new_n7641_);
  not g_17802 (not_new_n1027__138412872010, new_n1027_);
  not g_17803 (not_new_n928__24010, new_n928_);
  and g_17804 (and_and_new_n1820__new_n1823__new_n1821_, and_new_n1820__new_n1823_, new_n1821_);
  not g_17805 (new_n1607_, new_n981_);
  or g_17806 (new_n2365_, not_new_n1037__0, not_new_n598__1);
  not g_17807 (not_new_n587__3430, new_n587_);
  not g_17808 (not_new_n3372__70, new_n3372_);
  or g_17809 (new_n4344_, not_new_n4245_, not_new_n670_);
  not g_17810 (not_new_n9952__0, new_n9952_);
  not g_17811 (not_new_n582_, new_n582_);
  not g_17812 (not_new_n10134_, new_n10134_);
  or g_17813 (new_n9269_, not_new_n9089_, not_new_n9267_);
  not g_17814 (not_po296_6, po296);
  not g_17815 (not_new_n3705_, new_n3705_);
  and g_17816 (new_n9464_, new_n9700_, new_n9577_);
  or g_17817 (new_n6402_, not_new_n6288_, not_new_n628__403536070);
  or g_17818 (new_n2813_, not_new_n2810_, not_pi255_2);
  not g_17819 (not_new_n1340_, new_n1340_);
  and g_17820 (and_new_n1731__new_n1732_, new_n1731_, new_n1732_);
  or g_17821 (new_n8561_, not_new_n8354_, not_new_n8560_);
  not g_17822 (not_new_n633__24010, new_n633_);
  not g_17823 (not_new_n5004_, new_n5004_);
  and g_17824 (new_n4723_, new_n4847_, new_n4729_);
  not g_17825 (not_new_n1598_, new_n1598_);
  not g_17826 (not_new_n8105_, new_n8105_);
  not g_17827 (not_new_n4962_, new_n4962_);
  not g_17828 (not_new_n4124__0, new_n4124_);
  or g_17829 (new_n7977_, not_new_n1037__8235430, not_new_n7604__0);
  not g_17830 (new_n2322_, new_n623_);
  not g_17831 (not_new_n1472_, new_n1472_);
  or g_17832 (new_n7308_, not_new_n7300_, not_new_n7159__0);
  not g_17833 (not_pi263, pi263);
  not g_17834 (not_new_n9492_, new_n9492_);
  or g_17835 (new_n7894_, not_new_n638__2326305139872070, not_new_n7643__1);
  not g_17836 (not_new_n626__24010, new_n626_);
  not g_17837 (not_new_n9448_, new_n9448_);
  not g_17838 (new_n6289_, new_n1071_);
  not g_17839 (not_new_n608__70, new_n608_);
  or g_17840 (new_n5701_, not_new_n5456__0, not_pi140_3);
  not g_17841 (not_new_n5844_, new_n5844_);
  not g_17842 (not_new_n3666_, new_n3666_);
  not g_17843 (not_new_n4530_, new_n4530_);
  not g_17844 (not_new_n1581__490, new_n1581_);
  or g_17845 (new_n8272_, not_new_n8446_, not_new_n8161_);
  not g_17846 (not_new_n3184__19773267430, new_n3184_);
  not g_17847 (new_n9089_, new_n8969_);
  not g_17848 (new_n8151_, new_n1061_);
  not g_17849 (not_new_n9915__1, new_n9915_);
  or g_17850 (new_n2820_, not_new_n3311__6, not_new_n1051__1);
  or g_17851 (new_n7552_, not_new_n7550_, not_new_n7293__0);
  not g_17852 (not_new_n2805_, new_n2805_);
  or g_17853 (new_n10051_, not_new_n1043__332329305696010, not_new_n10031_);
  or g_17854 (new_n8371_, not_new_n8132_, not_new_n1600__57648010);
  not g_17855 (not_new_n1597__19773267430, new_n1597_);
  not g_17856 (not_new_n2128_, new_n2128_);
  not g_17857 (not_new_n610__10, new_n610_);
  not g_17858 (not_new_n1009_, new_n1009_);
  not g_17859 (not_new_n7884_, new_n7884_);
  not g_17860 (not_new_n1240_, new_n1240_);
  or g_17861 (new_n8732_, not_new_n8630_, not_new_n1039__6782230728490);
  or g_17862 (new_n1723_, key_gate_32, not_new_n596__113988951853731430);
  not g_17863 (not_new_n1001_, new_n1001_);
  not g_17864 (not_new_n5850_, new_n5850_);
  not g_17865 (not_new_n1043__5, new_n1043_);
  not g_17866 (not_new_n3869_, new_n3869_);
  not g_17867 (not_new_n4920_, new_n4920_);
  not g_17868 (not_new_n7125_, new_n7125_);
  and g_17869 (and_new_n6481__new_n6853_, new_n6481_, new_n6853_);
  not g_17870 (not_new_n3686_, new_n3686_);
  not g_17871 (not_new_n1602__113988951853731430, new_n1602_);
  not g_17872 (not_new_n596_, key_gate_88);
  not g_17873 (not_new_n6182_, new_n6182_);
  not g_17874 (not_new_n8156__0, new_n8156_);
  not g_17875 (not_new_n1591__5, new_n1591_);
  not g_17876 (not_new_n4009_, new_n4009_);
  not g_17877 (not_new_n630__2824752490, new_n630_);
  or g_17878 (new_n2156_, not_new_n9343_, not_new_n1584__403536070);
  or g_17879 (new_n5356_, not_new_n630__24010, not_new_n4986_);
  or g_17880 (new_n7437_, not_new_n7127_, not_new_n775__19773267430);
  or g_17881 (new_n5017_, not_new_n5394_, not_new_n5395_);
  not g_17882 (not_new_n8699_, new_n8699_);
  not g_17883 (not_new_n8798__0, new_n8798_);
  not g_17884 (not_new_n1603__47475615099430, new_n1603_);
  not g_17885 (not_new_n8373_, new_n8373_);
  or g_17886 (new_n10302_, not_new_n9934__0, not_new_n630__39098210485829880490);
  not g_17887 (not_new_n4844_, new_n4844_);
  or g_17888 (new_n9275_, not_new_n640__47475615099430, not_new_n8875__0);
  not g_17889 (not_new_n1249_, new_n1249_);
  or g_17890 (new_n1793_, not_new_n7678_, not_new_n1583__0);
  or g_17891 (po213, not_new_n2503_, or_not_new_n1571__not_new_n2504_);
  not g_17892 (not_new_n619__57648010, new_n619_);
  not g_17893 (not_new_n8813_, new_n8813_);
  not g_17894 (not_new_n5806_, new_n5806_);
  not g_17895 (not_new_n10120_, new_n10120_);
  not g_17896 (not_new_n1049__403536070, new_n1049_);
  or g_17897 (or_not_new_n6250__not_new_n6371_, not_new_n6250_, not_new_n6371_);
  not g_17898 (not_new_n581__332329305696010, new_n581_);
  or g_17899 (new_n3736_, not_new_n3424_, not_new_n1829_);
  or g_17900 (new_n2422_, not_new_n603__3430, not_new_n638__1);
  not g_17901 (not_new_n5326_, new_n5326_);
  not g_17902 (not_new_n4181_, new_n4181_);
  or g_17903 (new_n3682_, not_pi227, not_new_n989__3430);
  not g_17904 (not_new_n5762__0, new_n5762_);
  or g_17905 (new_n7838_, not_new_n7655__0, not_new_n1065__403536070);
  or g_17906 (new_n7925_, not_new_n7583_, not_new_n7754__0);
  not g_17907 (not_new_n8978_, new_n8978_);
  not g_17908 (not_new_n581__2569235775210588780886114772242356213216070, new_n581_);
  not g_17909 (not_new_n8957_, new_n8957_);
  not g_17910 (not_new_n9227_, new_n9227_);
  not g_17911 (not_new_n4945__1, new_n4945_);
  not g_17912 (not_new_n737_, new_n737_);
  and g_17913 (new_n1384_, new_n2445_, new_n2446_);
  not g_17914 (not_new_n633__797922662976120010, new_n633_);
  not g_17915 (new_n8843_, new_n1051_);
  or g_17916 (new_n3491_, not_new_n1613__1176490, not_new_n2109_);
  and g_17917 (new_n5026_, and_new_n5097__new_n5098_, new_n5100_);
  not g_17918 (not_new_n6720_, new_n6720_);
  not g_17919 (not_new_n8725_, new_n8725_);
  or g_17920 (new_n2928_, not_new_n3311__24010, not_new_n1071__1);
  not g_17921 (not_new_n1591__8235430, new_n1591_);
  or g_17922 (new_n8187_, not_new_n8562_, not_new_n8561_);
  or g_17923 (new_n10047_, not_new_n9854_, not_new_n9974_);
  not g_17924 (not_new_n6063_, new_n6063_);
  not g_17925 (not_new_n4827_, new_n4827_);
  not g_17926 (not_new_n8580_, new_n8580_);
  not g_17927 (not_new_n6656__0, new_n6656_);
  or g_17928 (new_n9770_, not_new_n9493_, not_new_n9492_);
  not g_17929 (new_n6272_, new_n1057_);
  or g_17930 (new_n6404_, not_new_n6235_, or_or_not_new_n6318__not_new_n6373__0_not_new_n6319_);
  not g_17931 (not_new_n581__8, new_n581_);
  not g_17932 (not_new_n6679_, new_n6679_);
  not g_17933 (not_new_n1043__8, new_n1043_);
  not g_17934 (not_new_n4113__1, new_n4113_);
  or g_17935 (new_n4566_, new_n1014_, pi176);
  not g_17936 (not_new_n6559_, new_n6559_);
  not g_17937 (not_new_n8996__0, new_n8996_);
  or g_17938 (new_n9536_, not_new_n9533_, not_new_n1047__968890104070);
  or g_17939 (new_n4150_, not_new_n4161__0, not_pi272_1);
  not g_17940 (not_new_n6443__2824752490, new_n6443_);
  not g_17941 (not_new_n1536__3430, new_n1536_);
  not g_17942 (not_new_n5277_, new_n5277_);
  or g_17943 (new_n5331_, not_new_n4992_, not_new_n1596__10);
  or g_17944 (new_n628_, or_or_not_new_n1806__not_new_n1807__not_new_n1809_, not_new_n1808_);
  or g_17945 (new_n1844_, not_pi166, not_new_n586__4);
  or g_17946 (new_n5651_, not_new_n5649_, not_new_n5650_);
  not g_17947 (not_new_n4792__1, new_n4792_);
  or g_17948 (new_n3027_, not_new_n1598__2, not_new_n581__490);
  not g_17949 (not_new_n8067_, new_n8067_);
  not g_17950 (not_new_n644__7, new_n644_);
  not g_17951 (not_new_n9130_, new_n9130_);
  not g_17952 (not_new_n1584__968890104070, new_n1584_);
  not g_17953 (not_new_n599__1176490, new_n599_);
  not g_17954 (not_new_n9620_, new_n9620_);
  not g_17955 (not_new_n1063_, new_n1063_);
  not g_17956 (not_new_n2994_, new_n2994_);
  or g_17957 (new_n2790_, not_new_n604__6, not_new_n636__3);
  or g_17958 (new_n3793_, not_new_n3464_, not_new_n1981_);
  not g_17959 (not_new_n1012__5, new_n1012_);
  or g_17960 (new_n2034_, not_new_n586__24010, not_pi176);
  not g_17961 (not_new_n9542_, new_n9542_);
  not g_17962 (not_new_n4119__0, new_n4119_);
  and g_17963 (and_new_n6983__new_n7398_, new_n6983_, new_n7398_);
  not g_17964 (not_new_n8200_, new_n8200_);
  not g_17965 (not_new_n7622_, new_n7622_);
  not g_17966 (not_new_n1017_, new_n1017_);
  not g_17967 (not_new_n4808_, new_n4808_);
  not g_17968 (not_new_n7701_, new_n7701_);
  not g_17969 (not_new_n1537__490, new_n1537_);
  and g_17970 (new_n9458_, new_n9553_, new_n9555_);
  not g_17971 (new_n6807_, new_n6626_);
  not g_17972 (new_n2285_, new_n618_);
  not g_17973 (not_po296_103677930763188441902487387275962551382129494864490, po296);
  not g_17974 (not_new_n3360_, new_n3360_);
  and g_17975 (and_new_n1991__new_n1994_, new_n1991_, new_n1994_);
  not g_17976 (not_new_n1065__2, new_n1065_);
  not g_17977 (not_new_n619__2824752490, new_n619_);
  not g_17978 (not_new_n636__10, new_n636_);
  not g_17979 (not_new_n4744_, new_n4744_);
  xnor g_17980 (key_gate_4, not_pi032, key_4);
  not g_17981 (not_new_n613__4, new_n613_);
  not g_17982 (not_new_n9251_, new_n9251_);
  or g_17983 (new_n3873_, not_new_n637__70, not_new_n6443__138412872010);
  not g_17984 (not_pi163, pi163);
  or g_17985 (new_n2664_, not_new_n1008_, not_new_n607__3430);
  or g_17986 (new_n7808_, not_new_n7791_, not_new_n7739__0);
  not g_17987 (not_new_n5552_, new_n5552_);
  not g_17988 (not_new_n593__1176490, new_n593_);
  not g_17989 (not_new_n8266__0, new_n8266_);
  not g_17990 (not_new_n617__1, new_n617_);
  not g_17991 (not_new_n1063__168070, new_n1063_);
  not g_17992 (not_new_n2147_, new_n2147_);
  not g_17993 (not_new_n2133_, new_n2133_);
  not g_17994 (not_new_n6727_, new_n6727_);
  or g_17995 (new_n9829_, not_new_n9503_, not_new_n9502_);
  or g_17996 (new_n8716_, not_new_n8794_, not_new_n8699_);
  not g_17997 (not_new_n621__4, new_n621_);
  not g_17998 (not_new_n3168_, new_n3168_);
  or g_17999 (new_n8738_, not_new_n8618_, not_new_n1175__0);
  or g_18000 (new_n3514_, not_new_n1537__47475615099430, not_pi123_0);
  not g_18001 (not_new_n3423_, new_n3423_);
  or g_18002 (new_n7505_, not_new_n7503_, not_new_n7277__0);
  not g_18003 (not_new_n10166_, new_n10166_);
  not g_18004 (not_new_n7033__1, new_n7033_);
  not g_18005 (not_new_n646__7, new_n646_);
  or g_18006 (new_n1898_, not_new_n591__6, not_new_n4727_);
  or g_18007 (new_n1802_, not_new_n593__0, not_new_n632_);
  not g_18008 (not_new_n1580__5, new_n1580_);
  and g_18009 (and_and_new_n2029__new_n2032__new_n2030_, and_new_n2029__new_n2032_, new_n2030_);
  not g_18010 (not_new_n4527_, new_n4527_);
  not g_18011 (not_new_n4291_, new_n4291_);
  not g_18012 (new_n4927_, new_n631_);
  not g_18013 (not_new_n7661__0, new_n7661_);
  not g_18014 (not_new_n5061_, new_n5061_);
  not g_18015 (not_new_n3279_, new_n3279_);
  not g_18016 (not_new_n8525_, new_n8525_);
  not g_18017 (not_new_n9607_, new_n9607_);
  not g_18018 (not_new_n3275_, new_n3275_);
  not g_18019 (not_new_n4784_, new_n4784_);
  not g_18020 (not_new_n1037__0, new_n1037_);
  not g_18021 (not_new_n3417_, new_n3417_);
  not g_18022 (not_pi108_0, pi108);
  or g_18023 (new_n2626_, or_not_new_n2625__not_new_n2624_, not_new_n2623_);
  not g_18024 (not_new_n6087_, new_n6087_);
  and g_18025 (and_not_pi040_1_not_pi039_1, not_pi039_1, not_pi040_1);
  not g_18026 (not_new_n9353_, new_n9353_);
  or g_18027 (new_n4043_, not_pi047_4, not_new_n3941_);
  or g_18028 (new_n8032_, not_new_n7724_, not_new_n7753__2);
  not g_18029 (not_new_n629__2, new_n629_);
  or g_18030 (new_n3568_, not_pi150_0, not_new_n1538__2824752490);
  not g_18031 (not_new_n5557_, new_n5557_);
  not g_18032 (not_new_n4627_, new_n4627_);
  not g_18033 (not_new_n5043_, new_n5043_);
  not g_18034 (not_new_n3384__1, new_n3384_);
  or g_18035 (new_n2467_, not_new_n629__1, not_new_n603__138412872010);
  not g_18036 (not_new_n622__490, new_n622_);
  not g_18037 (not_new_n5782__0, new_n5782_);
  not g_18038 (not_new_n581__797922662976120010, new_n581_);
  not g_18039 (not_new_n9601_, new_n9601_);
  not g_18040 (not_new_n1598__8, new_n1598_);
  not g_18041 (not_new_n3217_, new_n3217_);
  not g_18042 (not_new_n1591__6782230728490, new_n1591_);
  and g_18043 (new_n7144_, new_n7507_, new_n7506_);
  not g_18044 (not_new_n4146_, new_n4146_);
  or g_18045 (new_n3322_, not_pi058_0, not_new_n1534__3);
  or g_18046 (new_n8779_, not_new_n8776_, not_new_n8698_);
  or g_18047 (new_n1808_, not_pi100, not_new_n588__2);
  not g_18048 (new_n7424_, new_n7035_);
  and g_18049 (new_n1251_, new_n1893_, and_new_n1250__new_n1894_);
  and g_18050 (new_n4296_, new_n4241_, new_n703_);
  not g_18051 (not_new_n4529_, new_n4529_);
  not g_18052 (not_new_n7911_, new_n7911_);
  not g_18053 (not_new_n611__57648010, new_n611_);
  not g_18054 (new_n7847_, new_n7637_);
  or g_18055 (new_n2848_, not_new_n4130__2, not_new_n3310__7);
  not g_18056 (not_new_n6919_, new_n6919_);
  not g_18057 (not_new_n7835_, new_n7835_);
  or g_18058 (new_n9576_, new_n626_, new_n1053_);
  not g_18059 (not_new_n637__8235430, new_n637_);
  not g_18060 (not_new_n928__70, new_n928_);
  not g_18061 (new_n6514_, new_n1071_);
  not g_18062 (not_new_n7128_, new_n7128_);
  or g_18063 (or_or_or_not_new_n2727__not_new_n2730__not_new_n2729__not_new_n2731_, or_or_not_new_n2727__not_new_n2730__not_new_n2729_, not_new_n2731_);
  or g_18064 (new_n7048_, not_new_n7368_, not_new_n7367_);
  or g_18065 (new_n6910_, not_new_n6801_, not_new_n6909_);
  or g_18066 (new_n1806_, not_new_n586__2, not_pi164);
  or g_18067 (new_n9242_, not_new_n8964_, not_new_n8965_);
  or g_18068 (new_n729_, not_new_n3285_, not_new_n3286_);
  not g_18069 (not_new_n8175_, new_n8175_);
  or g_18070 (new_n5237_, not_new_n5235_, not_new_n5051_);
  not g_18071 (not_new_n1626_, new_n1626_);
  not g_18072 (not_new_n9509_, new_n9509_);
  or g_18073 (new_n1741_, not_pi085, not_new_n1728__9);
  not g_18074 (new_n1625_, new_n925_);
  not g_18075 (not_new_n625__2, new_n625_);
  not g_18076 (not_new_n5532_, new_n5532_);
  or g_18077 (new_n9296_, not_new_n638__1915812313805664144010, not_new_n8857_);
  not g_18078 (not_new_n1805_, new_n1805_);
  not g_18079 (not_new_n634__4, new_n634_);
  and g_18080 (and_and_new_n1739__new_n1740__new_n1742_, and_new_n1739__new_n1740_, new_n1742_);
  not g_18081 (not_new_n3808_, new_n3808_);
  or g_18082 (new_n8072_, not_new_n1053__8235430, not_new_n7649__0);
  or g_18083 (new_n1977_, not_new_n586__70, not_pi173);
  not g_18084 (not_new_n6841_, new_n6841_);
  not g_18085 (not_new_n5498__0, new_n5498_);
  or g_18086 (new_n2491_, not_new_n597__332329305696010, not_new_n4766__0);
  or g_18087 (new_n5993_, not_new_n5778_, not_new_n1071__10);
  not g_18088 (not_new_n9338_, new_n9338_);
  or g_18089 (new_n10050_, not_new_n631__4599865365447399609768010, not_new_n10049_);
  not g_18090 (not_new_n7364_, new_n7364_);
  or g_18091 (new_n5600_, not_new_n5596_, or_not_new_n5448__not_new_n5597__1);
  or g_18092 (new_n3206_, not_new_n1599__4, not_new_n3185__9);
  not g_18093 (not_new_n7671_, new_n7671_);
  or g_18094 (new_n4653_, not_new_n1011__3, not_new_n4449_);
  not g_18095 (not_new_n1584__6, new_n1584_);
  or g_18096 (new_n5262_, not_new_n4978__0, not_new_n5186__0);
  and g_18097 (new_n8213_, new_n8355_, new_n8086_);
  not g_18098 (not_new_n3308_, new_n3308_);
  not g_18099 (not_new_n1607__1176490, new_n1607_);
  not g_18100 (new_n10165_, new_n9950_);
  not g_18101 (not_new_n6726_, new_n6726_);
  or g_18102 (new_n2690_, not_new_n1010__0, not_new_n608__8235430);
  not g_18103 (not_new_n1027__2326305139872070, new_n1027_);
  or g_18104 (new_n4460_, not_new_n4641_, not_new_n4642_);
  not g_18105 (new_n5449_, pi137);
  not g_18106 (not_new_n1007_, new_n1007_);
  not g_18107 (not_pi102, pi102);
  not g_18108 (not_new_n7919_, new_n7919_);
  not g_18109 (new_n7102_, new_n774_);
  not g_18110 (not_new_n6514__0, new_n6514_);
  not g_18111 (not_new_n9962__0, new_n9962_);
  not g_18112 (not_new_n10125_, new_n10125_);
  not g_18113 (not_new_n6677__0, new_n6677_);
  not g_18114 (not_new_n9991_, new_n9991_);
  or g_18115 (new_n2773_, not_new_n602__4, not_new_n636__2);
  or g_18116 (new_n8755_, not_new_n8680_, not_new_n8595__5);
  or g_18117 (new_n3576_, not_new_n1538__6782230728490, not_pi154_0);
  not g_18118 (not_new_n3457_, new_n3457_);
  not g_18119 (not_new_n2564_, new_n2564_);
  not g_18120 (not_new_n4982_, new_n4982_);
  not g_18121 (not_new_n1607__8235430, new_n1607_);
  or g_18122 (new_n9235_, not_new_n8962_, not_new_n8963__1);
  not g_18123 (not_new_n4818_, new_n4818_);
  and g_18124 (new_n1354_, and_new_n1542__new_n2371_, new_n2370_);
  not g_18125 (not_new_n3406_, new_n3406_);
  not g_18126 (not_new_n9733_, new_n9733_);
  not g_18127 (not_new_n5786__2, new_n5786_);
  or g_18128 (or_not_new_n9327__0_not_new_n9524__0, not_new_n9524__0, not_new_n9327__0);
  not g_18129 (not_new_n737__0, new_n737_);
  not g_18130 (not_new_n4454_, new_n4454_);
  and g_18131 (new_n8088_, new_n8085_, new_n8341_);
  or g_18132 (new_n9655_, not_new_n640__332329305696010, not_new_n1604__47475615099430);
  not g_18133 (not_new_n9507_, new_n9507_);
  not g_18134 (not_new_n1055__47475615099430, new_n1055_);
  not g_18135 (not_new_n1616__47475615099430, new_n1616_);
  not g_18136 (not_pi064_1176490, pi064);
  not g_18137 (not_new_n2556_, new_n2556_);
  not g_18138 (not_new_n1031__3430, new_n1031_);
  not g_18139 (not_new_n603__9, new_n603_);
  not g_18140 (not_new_n648__57648010, new_n648_);
  not g_18141 (not_pi231, pi231);
  not g_18142 (not_new_n4806_, new_n4806_);
  not g_18143 (not_new_n7433_, new_n7433_);
  not g_18144 (not_new_n1045__24010, new_n1045_);
  or g_18145 (new_n8324_, not_new_n8322_, not_new_n8323_);
  not g_18146 (not_new_n741__1, new_n741_);
  not g_18147 (new_n7610_, new_n1039_);
  or g_18148 (new_n3624_, not_new_n984__1176490, not_pi178_0);
  not g_18149 (not_new_n4540_, new_n4540_);
  not g_18150 (new_n7457_, new_n7042_);
  or g_18151 (or_not_new_n1563__not_new_n2474_, not_new_n2474_, not_new_n1563_);
  not g_18152 (not_new_n647__403536070, new_n647_);
  not g_18153 (not_new_n1789_, new_n1789_);
  or g_18154 (new_n2245_, not_pi123, not_new_n588__47475615099430);
  or g_18155 (new_n5897_, not_new_n5780_, not_new_n6057_);
  not g_18156 (not_new_n1444_, new_n1444_);
  or g_18157 (new_n2554_, not_new_n607__2, not_new_n1015_);
  not g_18158 (not_new_n1619_, new_n1619_);
  or g_18159 (new_n7413_, not_new_n7119_, not_new_n775__3430);
  or g_18160 (new_n9237_, not_new_n8848_, not_new_n617__797922662976120010);
  not g_18161 (new_n1924_, new_n647_);
  not g_18162 (not_new_n2807_, new_n2807_);
  or g_18163 (new_n1761_, not_new_n3387__3, not_new_n3384__4);
  not g_18164 (not_new_n5577_, new_n5577_);
  not g_18165 (not_new_n1599__2, new_n1599_);
  not g_18166 (not_pi177_0, pi177);
  not g_18167 (not_new_n9211_, new_n9211_);
  not g_18168 (not_new_n7577_, new_n7577_);
  or g_18169 (new_n3331_, not_new_n1534__7, not_pi039_0);
  not g_18170 (not_new_n2831_, new_n2831_);
  or g_18171 (new_n5005_, not_new_n5308_, not_new_n5307_);
  or g_18172 (new_n2616_, or_not_new_n2615__not_new_n2614_, not_new_n2613_);
  not g_18173 (not_new_n9100_, new_n9100_);
  not g_18174 (not_new_n638__8, new_n638_);
  not g_18175 (not_new_n1468_, new_n1468_);
  not g_18176 (new_n5526_, new_n5435_);
  not g_18177 (not_pi064_138412872010, pi064);
  or g_18178 (new_n5617_, not_new_n5442_, not_new_n5533_);
  not g_18179 (not_new_n632__39098210485829880490, new_n632_);
  or g_18180 (new_n5139_, not_new_n5321_, or_or_not_new_n4933__not_new_n4930__0_not_new_n5322_);
  or g_18181 (new_n7411_, not_new_n761_, not_new_n6974__70);
  not g_18182 (not_new_n588__8235430, new_n588_);
  not g_18183 (not_new_n4813_, new_n4813_);
  and g_18184 (new_n9460_, new_n9326_, new_n9561_);
  not g_18185 (not_new_n612__3, new_n612_);
  not g_18186 (not_new_n8858_, new_n8858_);
  not g_18187 (not_new_n10031_, new_n10031_);
  not g_18188 (not_new_n984__2326305139872070, new_n984_);
  or g_18189 (new_n4893_, not_new_n4804__0, not_new_n4826_);
  not g_18190 (not_new_n775__57648010, new_n775_);
  not g_18191 (new_n4250_, new_n668_);
  not g_18192 (not_new_n646__2824752490, new_n646_);
  or g_18193 (new_n724_, not_new_n3273_, not_new_n3274_);
  or g_18194 (new_n3072_, not_new_n1176_, not_new_n1027__797922662976120010);
  not g_18195 (not_new_n6507_, new_n6507_);
  not g_18196 (not_new_n7045__2, new_n7045_);
  or g_18197 (new_n3901_, not_new_n9922_, not_new_n636__3430);
  not g_18198 (not_new_n9350_, new_n9350_);
  or g_18199 (new_n6104_, not_new_n5754__2, not_new_n1045__3430);
  not g_18200 (not_new_n10024_, new_n10024_);
  or g_18201 (new_n1822_, not_new_n4723_, not_new_n591__2);
  not g_18202 (not_new_n10184_, new_n10184_);
  or g_18203 (new_n1969_, not_new_n8812_, not_new_n1591__9);
  not g_18204 (new_n3991_, pi053);
  not g_18205 (not_new_n593__24010, new_n593_);
  not g_18206 (not_new_n5339_, new_n5339_);
  not g_18207 (not_new_n974_, new_n974_);
  or g_18208 (new_n4623_, not_new_n4422_, not_pi165_2);
  not g_18209 (not_pi052_1, pi052);
  not g_18210 (not_new_n4501_, new_n4501_);
  not g_18211 (not_new_n4172__0, new_n4172_);
  not g_18212 (not_pi131_2, pi131);
  not g_18213 (not_pi191, pi191);
  or g_18214 (new_n8495_, not_new_n8250__0, not_new_n619__57648010);
  not g_18215 (new_n8155_, new_n627_);
  not g_18216 (new_n7596_, new_n634_);
  or g_18217 (new_n2198_, not_new_n1589__19773267430, not_new_n5014_);
  not g_18218 (not_new_n2509__168070, new_n2509_);
  not g_18219 (not_new_n8671_, new_n8671_);
  not g_18220 (not_new_n7457_, new_n7457_);
  or g_18221 (new_n3068_, not_new_n1059__2, not_new_n581__332329305696010);
  not g_18222 (not_new_n1589__332329305696010, new_n1589_);
  not g_18223 (new_n4955_, new_n1602_);
  not g_18224 (not_new_n2663_, new_n2663_);
  not g_18225 (not_new_n6123_, new_n6123_);
  not g_18226 (new_n6510_, new_n640_);
  not g_18227 (not_new_n704_, new_n704_);
  not g_18228 (not_new_n5988_, new_n5988_);
  not g_18229 (not_new_n1328_, new_n1328_);
  or g_18230 (new_n6863_, not_new_n6620__0, not_new_n1607__70);
  or g_18231 (new_n5435_, not_new_n5525_, not_new_n5524_);
  not g_18232 (not_new_n5240_, new_n5240_);
  not g_18233 (not_new_n643__9, new_n643_);
  not g_18234 (not_new_n617__13410686196639649008070, new_n617_);
  or g_18235 (new_n7203_, not_new_n7109__0, not_new_n736_);
  not g_18236 (not_new_n1047__9, new_n1047_);
  not g_18237 (not_new_n2626_, new_n2626_);
  not g_18238 (not_new_n647__57648010, new_n647_);
  not g_18239 (not_new_n602__2326305139872070, new_n602_);
  not g_18240 (not_new_n641__1, new_n641_);
  not g_18241 (not_new_n1344_, new_n1344_);
  not g_18242 (not_new_n591__797922662976120010, new_n591_);
  not g_18243 (not_new_n7027__0, new_n7027_);
  or g_18244 (new_n9044_, new_n626_, new_n1053_);
  not g_18245 (not_new_n1017__4, new_n1017_);
  or g_18246 (new_n4618_, not_new_n4424__0, not_pi166_3);
  or g_18247 (new_n8748_, not_new_n1151__0, not_new_n8602_);
  not g_18248 (new_n4278_, new_n685_);
  or g_18249 (or_or_not_new_n2749__not_new_n2752__not_new_n2751_, not_new_n2751_, or_not_new_n2749__not_new_n2752_);
  or g_18250 (new_n6427_, not_new_n1604__3430, or_or_not_new_n6339__not_new_n6232__1_not_new_n6242__3);
  not g_18251 (not_new_n5473__0, new_n5473_);
  not g_18252 (not_new_n8076_, new_n8076_);
  not g_18253 (not_new_n1601__16284135979104490, new_n1601_);
  not g_18254 (not_new_n1588_, new_n1588_);
  or g_18255 (new_n635_, or_or_not_new_n1863__not_new_n1864__not_new_n1866_, not_new_n1865_);
  not g_18256 (not_po296_63668057609090279857414351392240010, po296);
  and g_18257 (and_new_n6244__new_n6372_, new_n6372_, new_n6244_);
  not g_18258 (not_new_n633__4, new_n633_);
  not g_18259 (not_new_n9300_, new_n9300_);
  not g_18260 (new_n4445_, pi177);
  not g_18261 (not_new_n648__3430, new_n648_);
  or g_18262 (new_n5424_, not_new_n4931_, not_new_n641__490);
  not g_18263 (not_new_n1581__3430, new_n1581_);
  not g_18264 (not_new_n5548_, new_n5548_);
  or g_18265 (new_n4888_, not_new_n1061__9, not_new_n4800_);
  not g_18266 (not_new_n9368_, new_n9368_);
  not g_18267 (not_new_n642__3, new_n642_);
  not g_18268 (not_new_n7662_, new_n7662_);
  not g_18269 (not_new_n1636_, key_gate_71);
  not g_18270 (new_n9930_, new_n643_);
  not g_18271 (not_new_n5689_, new_n5689_);
  not g_18272 (not_new_n9609_, new_n9609_);
  or g_18273 (new_n2401_, not_new_n597__8, not_new_n4750__0);
  or g_18274 (or_or_not_new_n2607__not_new_n2611__not_new_n1437_, or_not_new_n2607__not_new_n2611_, not_new_n1437_);
  not g_18275 (not_new_n604__0, new_n604_);
  or g_18276 (new_n9116_, new_n1599_, new_n622_);
  or g_18277 (new_n939_, not_new_n3372__1, not_new_n1028__2);
  not g_18278 (not_new_n2970_, new_n2970_);
  or g_18279 (new_n3591_, not_new_n942_, not_new_n1611_);
  not g_18280 (not_new_n638__7, new_n638_);
  not g_18281 (not_new_n9699_, new_n9699_);
  or g_18282 (new_n7658_, not_new_n643__968890104070, not_new_n7644_);
  not g_18283 (not_new_n8450_, new_n8450_);
  not g_18284 (not_new_n7421_, new_n7421_);
  not g_18285 (not_new_n5502_, new_n5502_);
  not g_18286 (not_new_n7729_, new_n7729_);
  or g_18287 (new_n8347_, not_new_n8150_, not_new_n638__113988951853731430);
  not g_18288 (not_new_n1602__3430, new_n1602_);
  or g_18289 (new_n6431_, or_or_not_new_n6348__not_new_n6232__2_not_new_n6234__1, not_new_n1049__3430);
  not g_18290 (not_new_n1039__138412872010, new_n1039_);
  not g_18291 (not_new_n9940__0, new_n9940_);
  not g_18292 (not_new_n4510_, new_n4510_);
  not g_18293 (not_pi049_1, pi049);
  not g_18294 (not_new_n1604__1, new_n1604_);
  not g_18295 (not_new_n9144_, new_n9144_);
  not g_18296 (not_new_n5591_, new_n5591_);
  buf g_18297 (po001, pi194);
  and g_18298 (new_n4901_, new_n5144_, new_n5143_);
  not g_18299 (not_new_n4554_, new_n4554_);
  and g_18300 (new_n1507_, new_n998_, new_n3033_);
  or g_18301 (new_n7884_, not_new_n7770__0, not_new_n7883_);
  or g_18302 (new_n7595_, not_new_n7905_, not_new_n7753_);
  not g_18303 (not_new_n1599__8, new_n1599_);
  or g_18304 (po147, not_new_n3520_, not_new_n3521_);
  not g_18305 (not_new_n3772_, new_n3772_);
  not g_18306 (not_new_n5261_, new_n5261_);
  not g_18307 (not_new_n6184_, new_n6184_);
  not g_18308 (not_new_n1569__0, new_n1569_);
  or g_18309 (new_n4683_, not_new_n1015__4, not_new_n4441__0);
  or g_18310 (new_n3906_, not_new_n3907_, not_new_n3908_);
  and g_18311 (new_n1393_, new_n2467_, new_n2468_);
  or g_18312 (new_n2130_, not_pi149, not_new_n587__403536070);
  not g_18313 (not_new_n10137_, new_n10137_);
  not g_18314 (not_new_n3167_, new_n3167_);
  or g_18315 (new_n2714_, not_pi275_3, not_new_n2712_);
  not g_18316 (not_new_n775__138412872010, new_n775_);
  not g_18317 (not_new_n3655_, new_n3655_);
  or g_18318 (new_n738_, not_new_n3250_, not_new_n3249_);
  or g_18319 (new_n9899_, not_new_n9919_, not_new_n10060_);
  not g_18320 (not_new_n7005_, new_n7005_);
  and g_18321 (new_n1371_, new_n2412_, and_new_n2414__new_n2413_);
  or g_18322 (or_not_new_n1549__not_new_n1368_, not_new_n1368_, not_new_n1549_);
  or g_18323 (new_n2691_, not_new_n5427__0, not_new_n606__8235430);
  and g_18324 (new_n8201_, new_n8285_, new_n8295_);
  and g_18325 (new_n7581_, new_n7575_, new_n7855_);
  not g_18326 (not_new_n639__1176490, new_n639_);
  or g_18327 (new_n2933_, not_new_n632__3, not_new_n604__19773267430);
  not g_18328 (not_new_n2747_, new_n2747_);
  not g_18329 (not_new_n1027__2, new_n1027_);
  not g_18330 (not_new_n5401_, new_n5401_);
  not g_18331 (not_new_n4002_, new_n4002_);
  not g_18332 (not_new_n7100_, new_n7100_);
  not g_18333 (new_n1728_, new_n927_);
  not g_18334 (not_new_n989__3430, new_n989_);
  not g_18335 (not_new_n7613_, new_n7613_);
  or g_18336 (new_n5104_, new_n1045_, new_n635_);
  or g_18337 (new_n6675_, not_new_n6452_, not_new_n6617_);
  not g_18338 (not_new_n1538__70, new_n1538_);
  not g_18339 (not_new_n1603__24010, new_n1603_);
  not g_18340 (not_new_n6034_, new_n6034_);
  not g_18341 (not_new_n740_, new_n740_);
  not g_18342 (not_new_n8360_, new_n8360_);
  or g_18343 (new_n3254_, not_new_n631__8, not_new_n3184__3);
  or g_18344 (new_n1031_, not_new_n3395_, not_new_n3394_);
  or g_18345 (new_n3376_, not_new_n1001__0, not_new_n926__0);
  not g_18346 (not_new_n9917_, new_n9917_);
  not g_18347 (not_new_n4970_, new_n4970_);
  not g_18348 (not_new_n720__0, new_n720_);
  not g_18349 (not_new_n1067__4, new_n1067_);
  or g_18350 (new_n4637_, not_pi163_2, not_new_n4418_);
  or g_18351 (new_n2226_, not_pi122, not_new_n588__6782230728490);
  not g_18352 (new_n6278_, new_n630_);
  or g_18353 (new_n1067_, not_new_n3487_, not_new_n3488_);
  or g_18354 (new_n7966_, not_new_n7619__0, not_new_n7817_);
  not g_18355 (not_new_n8845_, new_n8845_);
  not g_18356 (not_new_n5502__0, new_n5502_);
  or g_18357 (new_n8790_, or_not_new_n1159__0_not_new_n8794__0, not_new_n8708_);
  or g_18358 (new_n3237_, not_new_n627__7, not_new_n589__6782230728490);
  not g_18359 (not_new_n1588__113988951853731430, new_n1588_);
  not g_18360 (not_new_n647_, new_n647_);
  or g_18361 (new_n5295_, not_new_n5254_, not_new_n4944__0);
  not g_18362 (not_new_n7971_, new_n7971_);
  not g_18363 (not_new_n8307_, new_n8307_);
  or g_18364 (new_n2262_, not_new_n586__332329305696010, not_pi188);
  not g_18365 (not_pi048_0, pi048);
  or g_18366 (new_n3178_, not_new_n581__6168735096280623662907561568153897267931784070, not_new_n641__4);
  not g_18367 (not_new_n9666_, new_n9666_);
  or g_18368 (new_n10049_, not_new_n9888_, not_new_n9889_);
  and g_18369 (new_n4492_, new_n4653_, new_n4654_);
  not g_18370 (not_new_n3349_, new_n3349_);
  or g_18371 (new_n3605_, not_new_n950_, not_new_n1611__6);
  not g_18372 (not_new_n2730_, new_n2730_);
  not g_18373 (not_new_n4548_, new_n4548_);
  not g_18374 (not_new_n624__9, new_n624_);
  not g_18375 (not_pi178_3, pi178);
  not g_18376 (new_n3454_, new_n1053_);
  not g_18377 (not_new_n1514_, new_n1514_);
  not g_18378 (new_n5081_, new_n4928_);
  not g_18379 (not_new_n6012_, new_n6012_);
  not g_18380 (new_n5113_, new_n4944_);
  and g_18381 (and_and_new_n1754__new_n1755__new_n1757_, and_new_n1754__new_n1755_, new_n1757_);
  not g_18382 (new_n6288_, new_n1039_);
  or g_18383 (new_n6067_, not_new_n5948__0, not_new_n5878_);
  not g_18384 (not_new_n1039__332329305696010, new_n1039_);
  or g_18385 (new_n7258_, not_new_n7457_, not_new_n7011_);
  or g_18386 (new_n1721_, not_pi062, not_new_n1631__16284135979104490);
  or g_18387 (new_n2894_, not_new_n2891_, not_new_n1616__1176490);
  not g_18388 (not_new_n8081_, new_n8081_);
  not g_18389 (not_new_n8894_, new_n8894_);
  not g_18390 (not_new_n597__70, new_n597_);
  not g_18391 (not_new_n5890__2, new_n5890_);
  not g_18392 (not_new_n6985__0, new_n6985_);
  not g_18393 (new_n3986_, pi057);
  not g_18394 (not_new_n7780_, new_n7780_);
  or g_18395 (new_n8786_, or_or_not_new_n1158__0_not_new_n8713__1_not_new_n8785_, not_new_n8707__0);
  not g_18396 (new_n9175_, new_n8871_);
  not g_18397 (not_new_n6991_, new_n6991_);
  not g_18398 (not_new_n8173_, new_n8173_);
  not g_18399 (not_new_n626__2, new_n626_);
  not g_18400 (not_new_n2817_, new_n2817_);
  not g_18401 (not_new_n618__7, new_n618_);
  not g_18402 (not_new_n7038__0, new_n7038_);
  not g_18403 (new_n5773_, new_n1601_);
  or g_18404 (new_n3909_, not_new_n9930__0, not_new_n1061__8);
  not g_18405 (not_new_n2976_, new_n2976_);
  not g_18406 (not_new_n603__6, new_n603_);
  not g_18407 (not_po296_445676403263631959001900459745680070, po296);
  or g_18408 (new_n9059_, not_new_n9055_, not_new_n9057_);
  not g_18409 (not_new_n647__1, new_n647_);
  not g_18410 (not_new_n8577_, new_n8577_);
  not g_18411 (not_pi254_0, pi254);
  not g_18412 (new_n7625_, new_n629_);
  not g_18413 (new_n4942_, new_n647_);
  not g_18414 (not_new_n9088_, new_n9088_);
  or g_18415 (or_or_not_new_n6335__not_new_n6373__4_not_new_n1071__490, not_new_n1071__490, or_not_new_n6335__not_new_n6373__4);
  not g_18416 (not_new_n3976_, new_n3976_);
  or g_18417 (new_n2772_, not_new_n626__2, not_new_n604__4);
  or g_18418 (new_n4022_, not_pi062_2, not_new_n4018_);
  or g_18419 (new_n6893_, not_new_n6595_, not_new_n6627_);
  not g_18420 (not_new_n627_, new_n627_);
  not g_18421 (not_new_n10015__0, new_n10015_);
  not g_18422 (not_new_n5619_, new_n5619_);
  not g_18423 (not_new_n4030__0, new_n4030_);
  or g_18424 (new_n8756_, not_new_n8618__0, not_new_n1175__1);
  or g_18425 (or_or_or_not_new_n2919__not_new_n2922__not_new_n2921__not_new_n2923_, or_or_not_new_n2919__not_new_n2922__not_new_n2921_, not_new_n2923_);
  or g_18426 (new_n8359_, not_new_n1071__8235430, not_new_n8142_);
  not g_18427 (not_new_n617__332329305696010, new_n617_);
  or g_18428 (new_n2786_, not_new_n4125__2, not_new_n612__0);
  or g_18429 (new_n7462_, not_new_n7087_, not_new_n7135_);
  or g_18430 (new_n2988_, not_new_n2987_, not_new_n1021_);
  or g_18431 (new_n6651_, not_new_n6532_, not_new_n1063__3430);
  not g_18432 (not_new_n1021__0, new_n1021_);
  not g_18433 (not_new_n4314_, new_n4314_);
  not g_18434 (not_new_n7631__2, new_n7631_);
  and g_18435 (new_n4305_, new_n4365_, new_n4364_);
  not g_18436 (new_n7631_, new_n1602_);
  or g_18437 (new_n2634_, not_new_n607__10, not_new_n1005_);
  or g_18438 (new_n1663_, not_new_n596__9, key_gate_26);
  or g_18439 (new_n3243_, not_new_n641__5, not_new_n589__2326305139872070);
  or g_18440 (new_n2406_, not_new_n4811__0, not_new_n597__9);
  not g_18441 (not_new_n1864_, new_n1864_);
  or g_18442 (new_n8470_, not_new_n8125__0, not_new_n8320_);
  not g_18443 (not_new_n5282_, new_n5282_);
  not g_18444 (not_pi252_0, pi252);
  or g_18445 (new_n5524_, not_new_n5504_, not_new_n5523_);
  or g_18446 (new_n2835_, not_new_n602__70, not_new_n622__3);
  not g_18447 (not_new_n4814__0, new_n4814_);
  not g_18448 (not_pi136_0, pi136);
  not g_18449 (not_new_n9593_, new_n9593_);
  or g_18450 (new_n6092_, not_new_n5759__0, not_new_n647__1176490);
  not g_18451 (not_new_n4242_, new_n4242_);
  or g_18452 (new_n3190_, not_new_n1047__4, not_new_n3185__1);
  not g_18453 (not_new_n625__19773267430, new_n625_);
  buf g_18454 (po028, pi236);
  not g_18455 (not_new_n7406__2, new_n7406_);
  not g_18456 (not_new_n9266_, new_n9266_);
  or g_18457 (new_n5285_, not_new_n1598__9, not_new_n5197__0);
  or g_18458 (or_or_or_not_new_n6897__not_new_n6798__not_new_n6826__not_new_n6827_, or_or_not_new_n6897__not_new_n6798__not_new_n6826_, not_new_n6827_);
  not g_18459 (not_new_n1043__2, new_n1043_);
  or g_18460 (new_n7868_, not_new_n7665_, not_new_n1596__57648010);
  not g_18461 (not_new_n2742_, new_n2742_);
  not g_18462 (not_pi229, pi229);
  not g_18463 (not_new_n721__0, new_n721_);
  or g_18464 (new_n7866_, not_new_n7765_, not_new_n617__968890104070);
  not g_18465 (not_new_n6366_, new_n6366_);
  or g_18466 (new_n7472_, not_new_n7262_, not_new_n7470_);
  not g_18467 (not_new_n1057__2, new_n1057_);
  not g_18468 (not_new_n1456_, new_n1456_);
  and g_18469 (new_n7715_, new_n7869_, new_n7586_);
  not g_18470 (not_new_n5485_, new_n5485_);
  or g_18471 (new_n3888_, not_new_n1576__113988951853731430, not_new_n642__70);
  not g_18472 (not_new_n7665__0, new_n7665_);
  not g_18473 (not_new_n1598__138412872010, new_n1598_);
  or g_18474 (new_n1906_, not_new_n635__0, not_new_n601__5);
  not g_18475 (not_new_n2722_, new_n2722_);
  not g_18476 (not_new_n8328_, new_n8328_);
  not g_18477 (new_n9377_, new_n617_);
  not g_18478 (not_new_n9507__0, new_n9507_);
  or g_18479 (new_n4535_, not_new_n4477_, not_new_n4534_);
  not g_18480 (not_new_n8853_, new_n8853_);
  or g_18481 (new_n4612_, not_new_n4610_, not_new_n4611_);
  not g_18482 (not_new_n7918_, new_n7918_);
  or g_18483 (new_n5515_, not_new_n5557_, not_new_n5556_);
  not g_18484 (not_new_n581__7490483309651862334944941026945644936490, new_n581_);
  and g_18485 (new_n4304_, new_n4361_, new_n4362_);
  not g_18486 (not_new_n617__797922662976120010, new_n617_);
  or g_18487 (new_n2573_, not_new_n4467_, not_new_n609__6);
  or g_18488 (new_n1729_, not_new_n3318_, not_new_n925_);
  or g_18489 (new_n5072_, not_new_n5229_, not_new_n4930_);
  and g_18490 (new_n8705_, new_n8790_, new_n8704_);
  or g_18491 (new_n10171_, not_new_n10170_, not_new_n9950__0);
  not g_18492 (not_new_n7021__0, new_n7021_);
  or g_18493 (or_or_or_not_new_n2758__not_new_n2761__not_new_n2760__not_new_n2762_, or_or_not_new_n2758__not_new_n2761__not_new_n2760_, not_new_n2762_);
  not g_18494 (not_new_n9977_, new_n9977_);
  not g_18495 (not_new_n6788_, new_n6788_);
  or g_18496 (new_n8404_, not_new_n8242_, not_new_n8403_);
  not g_18497 (not_new_n9994_, new_n9994_);
  not g_18498 (not_new_n5818_, new_n5818_);
  not g_18499 (not_new_n8248__2, new_n8248_);
  not g_18500 (not_new_n3584_, new_n3584_);
  not g_18501 (not_new_n5543_, new_n5543_);
  not g_18502 (not_new_n1273_, new_n1273_);
  or g_18503 (new_n10048_, not_new_n9854__0, not_new_n9976_);
  not g_18504 (not_new_n6768_, new_n6768_);
  not g_18505 (not_new_n3887_, new_n3887_);
  not g_18506 (not_new_n5482_, new_n5482_);
  not g_18507 (not_new_n5881_, new_n5881_);
  or g_18508 (new_n7744_, not_new_n7863_, not_new_n7712_);
  or g_18509 (new_n8005_, not_new_n8004_, not_new_n7930_);
  and g_18510 (new_n3918_, new_n4043_, new_n4015_);
  not g_18511 (not_new_n598__5, new_n598_);
  not g_18512 (not_new_n2154_, new_n2154_);
  not g_18513 (not_new_n5712_, new_n5712_);
  not g_18514 (not_new_n5166_, new_n5166_);
  not g_18515 (not_new_n1773_, new_n1773_);
  not g_18516 (not_new_n2509__9, new_n2509_);
  or g_18517 (new_n5309_, not_new_n4929__0, not_new_n631__168070);
  or g_18518 (new_n9038_, not_new_n1039__332329305696010, not_new_n628__797922662976120010);
  or g_18519 (new_n4605_, not_new_n4603_, not_new_n4604_);
  not g_18520 (new_n3387_, new_n1027_);
  not g_18521 (not_new_n1631__0, key_gate_76);
  not g_18522 (not_new_n10240_, new_n10240_);
  not g_18523 (not_new_n5908_, new_n5908_);
  not g_18524 (not_new_n3710_, new_n3710_);
  not g_18525 (new_n5522_, new_n5504_);
  and g_18526 (new_n5894_, new_n6162_, new_n6163_);
  or g_18527 (or_not_new_n680__not_new_n4322_, not_new_n680_, not_new_n4322_);
  not g_18528 (not_new_n1613__332329305696010, new_n1613_);
  not g_18529 (not_new_n7725_, new_n7725_);
  or g_18530 (new_n5246_, not_new_n5053_, not_new_n5244_);
  or g_18531 (new_n2791_, not_new_n643__3, not_new_n602__6);
  not g_18532 (not_new_n8084_, new_n8084_);
  not g_18533 (new_n7876_, new_n7670_);
  not g_18534 (not_new_n1067__1, new_n1067_);
  or g_18535 (new_n1653_, not_po296_6, not_pi025);
  or g_18536 (or_or_not_new_n1158__0_not_new_n8713__1_not_new_n8785_, not_new_n8785_, or_not_new_n1158__0_not_new_n8713__1);
  not g_18537 (not_new_n7648__0, new_n7648_);
  not g_18538 (not_new_n4153_, new_n4153_);
  not g_18539 (not_new_n9954_, new_n9954_);
  not g_18540 (not_new_n8153_, new_n8153_);
  not g_18541 (not_new_n608__24010, new_n608_);
  not g_18542 (not_new_n5600_, new_n5600_);
  and g_18543 (and_new_n1278__new_n2027_, new_n1278_, new_n2027_);
  not g_18544 (not_new_n1039__5585458640832840070, new_n1039_);
  not g_18545 (not_new_n5406_, new_n5406_);
  and g_18546 (new_n6330_, new_n6271_, new_n6373_);
  or g_18547 (new_n9064_, new_n1063_, new_n638_);
  not g_18548 (not_new_n1601__0, new_n1601_);
  not g_18549 (not_new_n4503_, new_n4503_);
  and g_18550 (and_and_new_n1877__new_n1880__new_n1878_, and_new_n1877__new_n1880_, new_n1878_);
  not g_18551 (not_new_n601__168070, new_n601_);
  or g_18552 (new_n7319_, not_new_n7206_, not_new_n6966_);
  or g_18553 (new_n2012_, not_new_n4806_, not_new_n591__490);
  or g_18554 (new_n2886_, not_new_n595__1176490, not_new_n7067_);
  not g_18555 (not_new_n3184__70, new_n3184_);
  or g_18556 (new_n3700_, not_pi236, not_new_n989__138412872010);
  not g_18557 (new_n7779_, new_n7753_);
  or g_18558 (new_n3249_, not_new_n589__797922662976120010, not_new_n1047__5);
  or g_18559 (new_n2382_, not_new_n603__5, not_new_n634__1);
  or g_18560 (new_n9840_, not_new_n636__16284135979104490, not_new_n9390_);
  not g_18561 (not_new_n1584__8, new_n1584_);
  or g_18562 (new_n9248_, not_new_n9246_, not_new_n9247_);
  not g_18563 (not_new_n4040_, new_n4040_);
  and g_18564 (new_n8084_, new_n8309_, new_n8287_);
  not g_18565 (not_new_n7666_, new_n7666_);
  or g_18566 (new_n711_, not_new_n3081_, not_new_n1527_);
  or g_18567 (new_n9106_, not_new_n8963__0, not_new_n1596__6782230728490);
  not g_18568 (not_new_n10110__0, new_n10110_);
  or g_18569 (new_n2720_, not_new_n930_, or_not_new_n929__not_new_n931_);
  not g_18570 (not_pi064_7, pi064);
  not g_18571 (not_new_n4815_, new_n4815_);
  not g_18572 (not_new_n618__4599865365447399609768010, new_n618_);
  not g_18573 (not_new_n7114_, new_n7114_);
  and g_18574 (and_new_n1318__new_n2217_, new_n2217_, new_n1318_);
  not g_18575 (not_new_n5208_, new_n5208_);
  not g_18576 (not_new_n994__10, new_n994_);
  not g_18577 (not_new_n1017__3, new_n1017_);
  not g_18578 (not_new_n636__138412872010, new_n636_);
  or g_18579 (new_n3131_, not_new_n3315__168070, not_new_n625__5);
  not g_18580 (not_new_n1281_, new_n1281_);
  not g_18581 (not_new_n775__4, new_n775_);
  or g_18582 (new_n7961_, not_new_n1045__138412872010, not_new_n7611__2);
  not g_18583 (not_new_n1588__2326305139872070, new_n1588_);
  not g_18584 (not_new_n3929_, key_gate_36);
  or g_18585 (new_n9145_, not_new_n1059__968890104070, not_new_n644__2326305139872070);
  not g_18586 (new_n9364_, new_n634_);
  not g_18587 (not_new_n9023_, new_n9023_);
  not g_18588 (not_new_n1728__8235430, new_n1728_);
  not g_18589 (not_new_n4794__0, new_n4794_);
  not g_18590 (not_new_n7001_, new_n7001_);
  not g_18591 (not_new_n1824_, new_n1824_);
  or g_18592 (new_n4685_, not_new_n4683_, not_new_n4684_);
  not g_18593 (not_new_n7022__0, new_n7022_);
  not g_18594 (not_new_n5455__0, new_n5455_);
  not g_18595 (not_new_n5815_, new_n5815_);
  not g_18596 (not_new_n9383__0, new_n9383_);
  not g_18597 (not_new_n8912_, new_n8912_);
  not g_18598 (not_new_n5519__0, new_n5519_);
  not g_18599 (new_n5786_, new_n1063_);
  or g_18600 (new_n2702_, not_new_n2509__57648010, not_pi212);
  not g_18601 (not_new_n10295_, new_n10295_);
  not g_18602 (not_new_n1580__0, new_n1580_);
  not g_18603 (not_new_n5402_, new_n5402_);
  and g_18604 (and_new_n1314__new_n2198_, new_n2198_, new_n1314_);
  not g_18605 (not_new_n7774__0, new_n7774_);
  not g_18606 (not_new_n9192_, new_n9192_);
  or g_18607 (new_n6595_, not_new_n6889_, not_new_n6890_);
  not g_18608 (not_new_n7415_, new_n7415_);
  or g_18609 (new_n3662_, not_new_n989__3, not_pi217);
  not g_18610 (not_new_n2925_, new_n2925_);
  not g_18611 (not_new_n1051__3430, new_n1051_);
  not g_18612 (not_new_n6932_, new_n6932_);
  or g_18613 (new_n4212_, not_new_n4090_, not_new_n4164_);
  or g_18614 (new_n2748_, not_new_n2745_, or_not_new_n2747__not_new_n2746_);
  not g_18615 (not_new_n618__32199057558131797268376070, new_n618_);
  or g_18616 (new_n3416_, not_new_n1613__1, not_new_n1824_);
  not g_18617 (not_new_n10328_, new_n10328_);
  not g_18618 (new_n7354_, new_n7024_);
  not g_18619 (not_new_n6592_, new_n6592_);
  not g_18620 (not_new_n1015__3, new_n1015_);
  not g_18621 (not_pi064_168070, pi064);
  and g_18622 (new_n6319_, new_n6230_, new_n1035_);
  or g_18623 (po224, not_new_n1436_, or_or_not_new_n2607__not_new_n2611__not_new_n1437_);
  or g_18624 (new_n6821_, not_new_n6496__0, not_new_n6654__0);
  not g_18625 (not_pi139_3, pi139);
  not g_18626 (not_new_n5614_, new_n5614_);
  not g_18627 (not_new_n637__7, new_n637_);
  not g_18628 (not_po298_19773267430, po298);
  not g_18629 (not_new_n8030_, new_n8030_);
  not g_18630 (new_n4951_, new_n1598_);
  not g_18631 (not_new_n4120_, new_n4120_);
  and g_18632 (new_n8934_, new_n9046_, new_n8982_);
  not g_18633 (not_new_n3098_, new_n3098_);
  or g_18634 (new_n9970_, not_new_n3912_, not_new_n3911_);
  not g_18635 (not_new_n3880_, new_n3880_);
  not g_18636 (new_n4969_, new_n1061_);
  or g_18637 (new_n1896_, not_new_n9957_, not_new_n594__5);
  not g_18638 (new_n1595_, new_n994_);
  not g_18639 (not_new_n4502_, new_n4502_);
  not g_18640 (not_new_n3658_, new_n3658_);
  or g_18641 (new_n6799_, not_new_n6737__1, not_new_n6544__0);
  not g_18642 (not_new_n638__1, new_n638_);
  not g_18643 (not_new_n3138_, new_n3138_);
  or g_18644 (new_n3188_, not_new_n3185__0, not_new_n1049__4);
  not g_18645 (new_n5912_, new_n5766_);
  not g_18646 (not_new_n3978__0, new_n3978_);
  and g_18647 (and_new_n2409__new_n2408_, new_n2409_, new_n2408_);
  or g_18648 (new_n4411_, not_new_n4489_, not_new_n4586_);
  not g_18649 (not_new_n8114__0, new_n8114_);
  or g_18650 (new_n1847_, not_new_n4117_, not_new_n585__4);
  not g_18651 (not_new_n624__10, new_n624_);
  not g_18652 (not_new_n1576__70, new_n1576_);
  and g_18653 (new_n8667_, new_n8760_, new_n8759_);
  not g_18654 (not_new_n9855__1, new_n9855_);
  not g_18655 (not_new_n9221_, new_n9221_);
  or g_18656 (new_n9589_, new_n643_, new_n1061_);
  or g_18657 (or_or_not_new_n1275__not_new_n1273__not_new_n2002_, or_not_new_n1275__not_new_n1273_, not_new_n2002_);
  not g_18658 (not_new_n6524__1, new_n6524_);
  or g_18659 (new_n4642_, not_new_n4640_, not_new_n4513_);
  or g_18660 (new_n7032_, not_new_n7407_, not_new_n7408_);
  or g_18661 (new_n8758_, not_new_n8739_, not_new_n8660_);
  not g_18662 (new_n9487_, new_n1607_);
  or g_18663 (new_n4939_, not_new_n5108_, not_new_n5107_);
  not g_18664 (not_new_n7052_, new_n7052_);
  or g_18665 (new_n3742_, not_new_n622__10, not_new_n1599__6);
  not g_18666 (not_new_n7455_, new_n7455_);
  or g_18667 (new_n3058_, not_new_n633__4, not_new_n3372__332329305696010);
  not g_18668 (not_new_n9366_, new_n9366_);
  not g_18669 (not_new_n9095__0, new_n9095_);
  not g_18670 (not_new_n10128__0, new_n10128_);
  not g_18671 (not_new_n6019_, new_n6019_);
  not g_18672 (not_new_n627__24010, new_n627_);
  not g_18673 (not_new_n6820_, new_n6820_);
  or g_18674 (new_n4397_, not_new_n4280_, not_new_n684_);
  not g_18675 (not_new_n9327__0, new_n9327_);
  not g_18676 (not_new_n1065__1176490, new_n1065_);
  or g_18677 (new_n936_, not_new_n1582_, not_new_n3375__0);
  or g_18678 (new_n1843_, not_new_n1240_, not_new_n1838_);
  not g_18679 (new_n9928_, new_n644_);
  not g_18680 (not_new_n10237_, new_n10237_);
  or g_18681 (new_n3558_, not_pi145_0, not_new_n1538__168070);
  or g_18682 (new_n7392_, not_new_n7342__1, not_new_n741__1);
  not g_18683 (not_new_n619__10, new_n619_);
  not g_18684 (not_new_n3160_, new_n3160_);
  and g_18685 (new_n9866_, new_n10105_, new_n9864_);
  or g_18686 (new_n4342_, not_new_n4296_, not_new_n4344__0);
  not g_18687 (not_pi051, pi051);
  or g_18688 (new_n2094_, not_new_n4129_, not_new_n585__8235430);
  not g_18689 (not_new_n7138_, new_n7138_);
  or g_18690 (new_n9484_, not_new_n9697_, not_new_n9537_);
  or g_18691 (or_not_new_n9631__not_new_n9515__0, not_new_n9515__0, not_new_n9631_);
  not g_18692 (not_new_n722__1, new_n722_);
  not g_18693 (not_new_n7412__0, new_n7412_);
  not g_18694 (new_n9389_, new_n626_);
  not g_18695 (not_pi047_4, pi047);
  or g_18696 (new_n9661_, not_new_n9427__0, not_new_n9660_);
  and g_18697 (new_n8693_, new_n8771_, new_n8773_);
  not g_18698 (not_new_n5960_, new_n5960_);
  not g_18699 (not_new_n750_, new_n750_);
  not g_18700 (new_n5774_, new_n1602_);
  not g_18701 (not_new_n5684_, new_n5684_);
  not g_18702 (not_new_n775__6, new_n775_);
  not g_18703 (not_new_n10020__0, new_n10020_);
  or g_18704 (new_n1758_, not_new_n1728__332329305696010, not_pi072);
  not g_18705 (not_new_n929_, new_n929_);
  or g_18706 (new_n7547_, not_new_n7031__1, not_new_n6998__1);
  not g_18707 (not_new_n639__5585458640832840070, new_n639_);
  or g_18708 (new_n4080_, not_new_n4138_, not_new_n4155_);
  not g_18709 (not_new_n5001_, new_n5001_);
  not g_18710 (not_new_n8956__0, new_n8956_);
  not g_18711 (not_new_n630__138412872010, new_n630_);
  not g_18712 (not_new_n621__2824752490, new_n621_);
  or g_18713 (new_n4069_, not_new_n3955_, not_pi045_2);
  not g_18714 (new_n8614_, new_n1057_);
  not g_18715 (not_new_n8485_, new_n8485_);
  not g_18716 (not_new_n646__1176490, new_n646_);
  not g_18717 (not_new_n2759_, new_n2759_);
  not g_18718 (new_n8131_, new_n1599_);
  or g_18719 (new_n941_, not_new_n1027__2, not_new_n3375__1);
  not g_18720 (not_new_n3157_, new_n3157_);
  not g_18721 (not_new_n1597__3430, new_n1597_);
  not g_18722 (not_new_n5017_, new_n5017_);
  and g_18723 (new_n3965_, not_pi045_1, and_and_not_pi044_1_not_pi043_1_not_pi046_1);
  or g_18724 (new_n9809_, not_new_n9807_, not_new_n9808_);
  buf g_18725 (po020, pi244);
  and g_18726 (new_n5064_, new_n5337_, new_n5338_);
  not g_18727 (not_new_n5788_, new_n5788_);
  or g_18728 (new_n6837_, not_new_n6472__0, not_new_n1047__24010);
  or g_18729 (new_n6943_, not_new_n1059__1176490, not_new_n6521__0);
  not g_18730 (not_new_n984__0, new_n984_);
  not g_18731 (not_new_n5795__0, new_n5795_);
  not g_18732 (not_pi043_2, pi043);
  or g_18733 (new_n10191_, new_n1057_, new_n636_);
  not g_18734 (new_n7934_, new_n7672_);
  not g_18735 (not_new_n6793_, new_n6793_);
  not g_18736 (not_new_n10170_, new_n10170_);
  or g_18737 (new_n2562_, not_pi198, not_new_n2509__4);
  or g_18738 (new_n6898_, not_new_n6461_, not_new_n6658__0);
  not g_18739 (not_new_n9219_, new_n9219_);
  not g_18740 (not_new_n9360_, new_n9360_);
  not g_18741 (not_new_n602_, new_n602_);
  not g_18742 (not_new_n8317_, new_n8317_);
  xnor g_18743 (key_gate_100, key_100, new_n1642_);
  not g_18744 (not_po296_168070, po296);
  not g_18745 (not_new_n1576_, new_n1576_);
  not g_18746 (not_new_n5743__0, new_n5743_);
  not g_18747 (not_new_n9468_, new_n9468_);
  not g_18748 (not_new_n669_, new_n669_);
  not g_18749 (not_new_n4430__0, new_n4430_);
  not g_18750 (not_new_n596__2326305139872070, key_gate_88);
  not g_18751 (not_new_n2449_, new_n2449_);
  not g_18752 (not_new_n586__57648010, new_n586_);
  or g_18753 (new_n3004_, not_new_n3372__8, not_new_n631__4);
  not g_18754 (not_new_n5192__0, new_n5192_);
  not g_18755 (new_n8985_, new_n8866_);
  or g_18756 (new_n983_, not_pi001, not_new_n1536__10);
  not g_18757 (not_new_n7030__0, new_n7030_);
  or g_18758 (new_n2088_, not_new_n4796_, not_new_n591__1176490);
  not g_18759 (not_new_n3409_, new_n3409_);
  not g_18760 (not_new_n3442_, new_n3442_);
  not g_18761 (not_new_n1717_, key_gate_10);
  or g_18762 (new_n1892_, not_new_n6469_, not_new_n1580__6);
  not g_18763 (not_new_n601__332329305696010, new_n601_);
  not g_18764 (not_new_n1602__5, new_n1602_);
  and g_18765 (new_n1272_, and_and_new_n1991__new_n1994__new_n1992_, new_n1993_);
  or g_18766 (new_n5226_, not_new_n4974__0, not_new_n5218_);
  or g_18767 (new_n2384_, not_new_n9957__0, not_new_n599__5);
  or g_18768 (new_n5112_, not_new_n5056_, not_new_n5111_);
  or g_18769 (new_n8121_, not_new_n624__138412872010, not_new_n8108_);
  or g_18770 (new_n976_, not_new_n2267_, or_or_not_new_n1331__not_new_n1329__not_new_n2268_);
  not g_18771 (not_new_n8251_, new_n8251_);
  not g_18772 (not_new_n1607__19773267430, new_n1607_);
  or g_18773 (new_n3055_, not_new_n3372__47475615099430, not_new_n646__4);
  or g_18774 (new_n6690_, not_new_n6673_, not_new_n6617__0);
  not g_18775 (not_new_n1043__16284135979104490, new_n1043_);
  or g_18776 (new_n4937_, not_new_n1045__8, not_new_n635__3430);
  not g_18777 (not_new_n1347_, new_n1347_);
  not g_18778 (not_new_n625__403536070, new_n625_);
  not g_18779 (not_new_n9314_, new_n9314_);
  or g_18780 (new_n2906_, not_new_n604__57648010, not_new_n634__3);
  not g_18781 (not_new_n597__2824752490, new_n597_);
  not g_18782 (not_new_n7424__1, new_n7424_);
  not g_18783 (not_new_n6787_, new_n6787_);
  not g_18784 (not_pi089, pi089);
  not g_18785 (not_new_n4125_, new_n4125_);
  not g_18786 (not_new_n6533__0, new_n6533_);
  not g_18787 (not_new_n1061__7, new_n1061_);
  or g_18788 (new_n6704_, not_new_n6526_, not_new_n627__57648010);
  not g_18789 (not_new_n7148__0, new_n7148_);
  or g_18790 (new_n2438_, not_new_n600__1176490, not_new_n4130__0);
  or g_18791 (new_n9735_, not_new_n9373__2, not_new_n9684_);
  not g_18792 (not_new_n4760_, new_n4760_);
  buf g_18793 (po007, pi200);
  or g_18794 (new_n2521_, not_new_n606__0, not_new_n5484__0);
  or g_18795 (new_n9561_, not_new_n1043__6782230728490, not_new_n631__93874803376477543056490);
  or g_18796 (new_n2780_, not_po296_7490483309651862334944941026945644936490, not_pi251_0);
  or g_18797 (new_n5505_, not_pi130_1, not_new_n5519_);
  not g_18798 (not_new_n3260_, new_n3260_);
  or g_18799 (or_not_new_n2527__not_new_n2531_, not_new_n2531_, not_new_n2527_);
  not g_18800 (not_new_n6097_, new_n6097_);
  not g_18801 (not_new_n2531_, new_n2531_);
  or g_18802 (new_n2281_, not_pi189, not_new_n586__2326305139872070);
  or g_18803 (new_n3000_, not_new_n1152_, not_new_n1027__6);
  or g_18804 (new_n8332_, not_new_n8211_, not_new_n8454_);
  not g_18805 (not_new_n8838_, new_n8838_);
  not g_18806 (not_new_n1370_, new_n1370_);
  not g_18807 (not_new_n7807_, new_n7807_);
  or g_18808 (new_n3521_, not_new_n1613__16284135979104490, not_new_n2338_);
  not g_18809 (not_new_n5430__0, new_n5430_);
  not g_18810 (not_new_n5899__0, new_n5899_);
  not g_18811 (not_new_n8407_, new_n8407_);
  not g_18812 (not_new_n7616__0, new_n7616_);
  or g_18813 (new_n3984_, not_new_n3946_, not_new_n4025_);
  not g_18814 (not_pi275_2, pi275);
  not g_18815 (not_new_n8180_, new_n8180_);
  not g_18816 (new_n5746_, new_n1049_);
  not g_18817 (not_new_n9688_, new_n9688_);
  or g_18818 (new_n7507_, not_new_n7026__0, not_new_n6985__0);
  or g_18819 (new_n2859_, not_new_n7051_, not_new_n595__3430);
  not g_18820 (not_pi046_0, pi046);
  or g_18821 (new_n2931_, not_new_n7062_, not_new_n595__19773267430);
  or g_18822 (new_n8499_, not_new_n1596__968890104070, not_new_n8172__1);
  not g_18823 (not_new_n5328_, new_n5328_);
  not g_18824 (new_n8646_, new_n1164_);
  not g_18825 (not_new_n8569_, new_n8569_);
  not g_18826 (new_n5428_, pi129);
  not g_18827 (not_new_n9920_, new_n9920_);
  or g_18828 (new_n7417_, not_new_n764_, not_new_n6974__3430);
  not g_18829 (not_new_n632__403536070, new_n632_);
  not g_18830 (not_new_n9373__0, new_n9373_);
  and g_18831 (and_and_new_n6251__new_n6371__new_n1597_, new_n1597_, and_new_n6251__new_n6371_);
  not g_18832 (not_new_n632__8235430, new_n632_);
  not g_18833 (not_new_n9190_, new_n9190_);
  not g_18834 (not_new_n4442_, new_n4442_);
  not g_18835 (not_new_n7829_, new_n7829_);
  not g_18836 (not_new_n7837_, new_n7837_);
  or g_18837 (or_not_new_n3122__not_new_n3121_, not_new_n3121_, not_new_n3122_);
  not g_18838 (not_new_n4415_, new_n4415_);
  not g_18839 (not_new_n2949_, new_n2949_);
  not g_18840 (not_new_n4525_, new_n4525_);
  or g_18841 (new_n5175_, new_n1604_, new_n640_);
  not g_18842 (not_new_n3263_, new_n3263_);
  not g_18843 (not_new_n6475__2, new_n6475_);
  not g_18844 (not_new_n636__8235430, new_n636_);
  or g_18845 (new_n1823_, not_new_n1037_, not_new_n1588__2);
  not g_18846 (not_new_n1588__19773267430, new_n1588_);
  or g_18847 (new_n629_, or_or_not_new_n2208__not_new_n2205__not_new_n2206_, not_new_n2207_);
  not g_18848 (not_new_n589__2, new_n589_);
  not g_18849 (not_new_n7598__2, new_n7598_);
  and g_18850 (new_n1529_, new_n3372_, new_n3375_);
  not g_18851 (not_new_n3185__1176490, new_n3185_);
  not g_18852 (not_new_n602__968890104070, new_n602_);
  or g_18853 (new_n6206_, not_new_n1059__3430, not_new_n5788__0);
  not g_18854 (not_new_n630__16284135979104490, new_n630_);
  not g_18855 (new_n4240_, new_n672_);
  or g_18856 (new_n3704_, not_new_n989__6782230728490, not_pi238);
  not g_18857 (not_new_n7661_, new_n7661_);
  buf g_18858 (po032, pi232);
  or g_18859 (new_n3128_, not_new_n3315__24010, not_new_n630__5);
  or g_18860 (new_n3276_, not_new_n640__8, not_new_n3184__24010);
  not g_18861 (not_new_n4300_, new_n4300_);
  or g_18862 (new_n10225_, not_new_n9900__0, not_new_n10063_);
  not g_18863 (not_new_n1047__6782230728490, new_n1047_);
  or g_18864 (new_n9551_, not_new_n1037__6782230728490, not_new_n632__16284135979104490);
  not g_18865 (not_new_n1037__168070, new_n1037_);
  or g_18866 (new_n8505_, not_new_n8129__0, not_new_n617__2326305139872070);
  not g_18867 (not_new_n2704_, new_n2704_);
  not g_18868 (not_new_n6617__2, new_n6617_);
  or g_18869 (or_not_new_n2129__not_new_n2130_, not_new_n2129_, not_new_n2130_);
  not g_18870 (new_n1867_, new_n635_);
  or g_18871 (new_n6184_, not_new_n5900__4, not_new_n5868_);
  or g_18872 (new_n5574_, not_new_n1013__5, not_pi145_1);
  or g_18873 (or_or_not_new_n6339__not_new_n6232__1_not_new_n6242__3, or_not_new_n6339__not_new_n6232__1, not_new_n6242__3);
  or g_18874 (new_n5394_, not_new_n4999__3, not_new_n5263_);
  not g_18875 (not_new_n7046_, new_n7046_);
  not g_18876 (not_pi116_0, pi116);
  not g_18877 (not_new_n1596__168070, new_n1596_);
  not g_18878 (not_new_n6826_, new_n6826_);
  not g_18879 (not_new_n5490_, new_n5490_);
  or g_18880 (new_n6626_, not_new_n6796_, not_new_n6806_);
  not g_18881 (not_new_n1534__4, key_gate_5);
  not g_18882 (not_new_n1631__113988951853731430, key_gate_76);
  or g_18883 (new_n8487_, not_new_n8486_, not_new_n8485_);
  xnor g_18884 (key_gate_85, new_n3925_, key_85);
  not g_18885 (not_new_n3312_, new_n3312_);
  not g_18886 (not_po298_3, po298);
  or g_18887 (new_n7989_, not_new_n7664__1, not_new_n618__47475615099430);
  not g_18888 (not_new_n954_, new_n954_);
  or g_18889 (new_n3862_, not_new_n1576__1176490, not_new_n639__490);
  or g_18890 (or_or_not_new_n1295__not_new_n1293__not_new_n2097_, or_not_new_n1295__not_new_n1293_, not_new_n2097_);
  not g_18891 (not_new_n8984__2, new_n8984_);
  or g_18892 (new_n5820_, not_new_n6179_, not_new_n6178_);
  not g_18893 (not_new_n8500_, new_n8500_);
  or g_18894 (new_n2089_, not_new_n1588__1176490, not_new_n1065_);
  or g_18895 (new_n5215_, not_new_n5213_, not_new_n5046_);
  or g_18896 (new_n6465_, or_or_or_not_new_n6897__not_new_n6798__not_new_n6826__not_new_n6827_, not_new_n6898_);
  not g_18897 (not_new_n7402_, new_n7402_);
  not g_18898 (not_new_n5680__0, new_n5680_);
  and g_18899 (new_n9868_, new_n10187_, new_n10190_);
  and g_18900 (new_n6226_, new_n6225_, new_n6314_);
  not g_18901 (not_new_n7212_, new_n7212_);
  and g_18902 (new_n1449_, and_new_n2667__new_n2668_, new_n2669_);
  not g_18903 (not_new_n928__2326305139872070, new_n928_);
  or g_18904 (po282, or_or_or_not_new_n2865__not_new_n2868__not_new_n2867__not_new_n2869_, not_new_n2866_);
  or g_18905 (or_not_new_n1558__not_new_n2449_, not_new_n2449_, not_new_n1558_);
  or g_18906 (new_n3948_, not_new_n4030_, not_new_n3972_);
  not g_18907 (not_new_n648__4, new_n648_);
  not g_18908 (not_new_n1612__10, new_n1612_);
  or g_18909 (new_n1175_, not_new_n3879_, not_new_n3880_);
  not g_18910 (not_new_n8150__2, new_n8150_);
  or g_18911 (new_n3532_, not_pi132_0, not_new_n1538__2);
  or g_18912 (new_n9061_, new_n643_, new_n1061_);
  or g_18913 (new_n10133_, not_new_n1602__16284135979104490, not_new_n625__93874803376477543056490);
  xor g_18914 (key_gate_93, key_93, not_new_n3934_);
  not g_18915 (not_new_n1031__10, new_n1031_);
  not g_18916 (not_new_n8353_, new_n8353_);
  not g_18917 (not_new_n9896_, new_n9896_);
  not g_18918 (not_new_n8119__0, new_n8119_);
  not g_18919 (not_pi144_0, pi144);
  not g_18920 (not_new_n9482_, new_n9482_);
  not g_18921 (not_new_n706_, new_n706_);
  not g_18922 (not_new_n2870_, new_n2870_);
  or g_18923 (new_n4996_, not_new_n5172_, not_new_n5171_);
  or g_18924 (new_n2538_, not_new_n4463__0, not_new_n610__2);
  not g_18925 (not_new_n4767__0, new_n4767_);
  not g_18926 (new_n4517_, new_n4485_);
  not g_18927 (not_pi148_0, pi148);
  not g_18928 (not_new_n9657_, new_n9657_);
  not g_18929 (not_new_n7039__0, new_n7039_);
  or g_18930 (new_n1862_, not_new_n1244_, not_new_n1857_);
  not g_18931 (not_po296_968890104070, po296);
  or g_18932 (new_n3526_, not_pi129_1, not_new_n1538_);
  not g_18933 (not_new_n594__6, new_n594_);
  or g_18934 (new_n2194_, not_new_n9442_, not_new_n1584__19773267430);
  or g_18935 (new_n10310_, not_new_n9933__0, not_new_n1602__797922662976120010);
  not g_18936 (not_new_n5230_, new_n5230_);
  not g_18937 (not_new_n8876_, new_n8876_);
  not g_18938 (not_new_n775__5, new_n775_);
  not g_18939 (not_new_n8829_, new_n8829_);
  not g_18940 (new_n6294_, new_n1061_);
  or g_18941 (new_n3453_, not_new_n1594__9, not_new_n1019__1);
  or g_18942 (new_n6681_, not_new_n6649_, not_new_n648__403536070);
  or g_18943 (new_n4040_, not_new_n3995_, not_new_n4016_);
  or g_18944 (new_n6636_, not_new_n6583_, not_new_n6789_);
  not g_18945 (not_new_n3470_, new_n3470_);
  or g_18946 (new_n5314_, not_new_n4946__0, not_new_n5257_);
  or g_18947 (new_n7964_, not_new_n7612__0, not_new_n1043__1176490);
  and g_18948 (and_new_n9510__new_n9851_, new_n9510_, new_n9851_);
  or g_18949 (new_n2970_, not_new_n602__332329305696010, not_new_n618__2);
  not g_18950 (not_new_n2112_, new_n2112_);
  not g_18951 (not_new_n6996__0, new_n6996_);
  or g_18952 (new_n5597_, not_new_n5449_, not_new_n5544_);
  not g_18953 (not_new_n6650__0, new_n6650_);
  or g_18954 (new_n2490_, not_new_n1597__0, not_new_n598__332329305696010);
  or g_18955 (new_n7028_, not_new_n7429_, not_new_n7428_);
  not g_18956 (not_pi273, pi273);
  not g_18957 (not_new_n3979_, new_n3979_);
  or g_18958 (new_n7508_, not_new_n7345__1, not_new_n744__1);
  not g_18959 (not_new_n9984_, new_n9984_);
  not g_18960 (not_new_n8598_, new_n8598_);
  or g_18961 (new_n5943_, not_new_n1049__10, not_new_n5741_);
  or g_18962 (new_n2229_, not_new_n630__0, not_new_n601__138412872010);
  or g_18963 (new_n5513_, not_new_n5570_, not_new_n5569_);
  not g_18964 (not_new_n4132__1, new_n4132_);
  and g_18965 (new_n6971_, new_n7271_, new_n7274_);
  or g_18966 (new_n9720_, not_new_n647__2326305139872070, not_new_n9371_);
  not g_18967 (not_new_n5513_, new_n5513_);
  not g_18968 (not_pi180, pi180);
  not g_18969 (not_new_n6658_, new_n6658_);
  not g_18970 (not_new_n626__4599865365447399609768010, new_n626_);
  or g_18971 (new_n2548_, not_new_n610__3, not_new_n4464__0);
  or g_18972 (new_n9574_, not_new_n1053__6782230728490, not_new_n626__657123623635342801395430);
  not g_18973 (not_new_n628__113988951853731430, new_n628_);
  or g_18974 (new_n3861_, not_new_n639__70, not_new_n6443__1176490);
  not g_18975 (not_new_n1597__0, new_n1597_);
  not g_18976 (not_new_n3665_, new_n3665_);
  not g_18977 (new_n7752_, new_n1035_);
  or g_18978 (new_n10092_, not_new_n10090_, not_new_n9986_);
  or g_18979 (new_n5683_, not_new_n5679_, or_not_new_n5463__not_new_n5680__1);
  or g_18980 (new_n5427_, not_new_n5588_, not_new_n5506_);
  or g_18981 (new_n3808_, not_new_n3429_, not_new_n1848_);
  or g_18982 (po174, not_new_n3574_, not_new_n3575_);
  and g_18983 (po110, pi089, key_gate_101);
  not g_18984 (not_pi180_0, pi180);
  not g_18985 (new_n4979_, new_n1603_);
  not g_18986 (not_new_n6507__1, new_n6507_);
  or g_18987 (new_n5602_, not_new_n1004__6, not_new_n5445_);
  not g_18988 (not_new_n617__70, new_n617_);
  or g_18989 (new_n2825_, not_new_n604__9, not_new_n628__3);
  not g_18990 (not_new_n9563_, new_n9563_);
  not g_18991 (not_new_n1352_, new_n1352_);
  and g_18992 (new_n6223_, new_n6381_, new_n6380_);
  not g_18993 (not_new_n984__3, new_n984_);
  or g_18994 (new_n2595_, not_new_n605__8, not_new_n5492_);
  or g_18995 (new_n4377_, not_new_n658_, not_new_n4269_);
  not g_18996 (not_new_n5470_, new_n5470_);
  not g_18997 (not_pi047_2, pi047);
  or g_18998 (new_n2816_, not_new_n648__2, not_new_n604__8);
  not g_18999 (not_new_n603__70, new_n603_);
  not g_19000 (not_new_n5731_, new_n5731_);
  or g_19001 (new_n5260_, not_new_n4954__0, not_new_n5199__0);
  not g_19002 (not_new_n10269_, new_n10269_);
  or g_19003 (new_n9590_, not_new_n1061__47475615099430, not_new_n643__797922662976120010);
  or g_19004 (new_n5587_, not_new_n5585_, not_new_n5494_);
  or g_19005 (new_n5605_, not_new_n5446__0, not_pi136_3);
  not g_19006 (not_new_n7955_, new_n7955_);
  not g_19007 (not_new_n5058__0, new_n5058_);
  or g_19008 (new_n4600_, not_new_n4598_, not_new_n4537_);
  not g_19009 (not_new_n5387_, new_n5387_);
  or g_19010 (new_n5149_, not_new_n5147_, not_new_n5148_);
  not g_19011 (not_new_n6684_, new_n6684_);
  not g_19012 (not_new_n6447_, new_n6447_);
  not g_19013 (not_new_n4988_, new_n4988_);
  not g_19014 (not_new_n8830__0, new_n8830_);
  not g_19015 (not_new_n6363_, new_n6363_);
  not g_19016 (not_new_n5209__0, new_n5209_);
  or g_19017 (new_n1964_, not_new_n7694_, not_new_n1583__9);
  not g_19018 (not_new_n6511_, new_n6511_);
  or g_19019 (new_n10173_, not_new_n10165_, not_new_n9905__0);
  not g_19020 (not_new_n9157_, new_n9157_);
  or g_19021 (or_or_not_new_n2758__not_new_n2761__not_new_n2760_, not_new_n2760_, or_not_new_n2758__not_new_n2761_);
  and g_19022 (new_n8682_, new_n8612_, new_n1173_);
  or g_19023 (new_n2267_, not_new_n622__0, not_new_n601__6782230728490);
  not g_19024 (not_new_n9538_, new_n9538_);
  not g_19025 (not_new_n6736_, new_n6736_);
  not g_19026 (not_new_n10061_, new_n10061_);
  not g_19027 (not_new_n9239_, new_n9239_);
  not g_19028 (not_pi048_1, pi048);
  or g_19029 (new_n2316_, not_new_n4764_, not_new_n591__16284135979104490);
  not g_19030 (not_new_n1009__1, new_n1009_);
  or g_19031 (or_not_new_n3363__not_new_n583__0, not_new_n3363_, not_new_n583__0);
  or g_19032 (new_n2718_, not_new_n994_, not_new_n4132__1);
  not g_19033 (not_new_n4481_, new_n4481_);
  not g_19034 (not_new_n7693_, new_n7693_);
  not g_19035 (not_new_n644__490, new_n644_);
  not g_19036 (not_new_n4804__0, new_n4804_);
  or g_19037 (new_n4406_, not_new_n681_, not_new_n4319_);
  not g_19038 (not_new_n8199_, new_n8199_);
  or g_19039 (new_n2995_, not_new_n3372__5, not_new_n648__4);
  or g_19040 (new_n9673_, not_new_n644__797922662976120010, not_new_n1059__332329305696010);
  or g_19041 (new_n3789_, not_new_n3787_, not_new_n3788_);
  not g_19042 (not_new_n7758_, new_n7758_);
  not g_19043 (not_new_n1037__7, new_n1037_);
  not g_19044 (not_new_n632_, new_n632_);
  not g_19045 (not_new_n1538__1, new_n1538_);
  not g_19046 (new_n2161_, new_n964_);
  not g_19047 (new_n6485_, new_n642_);
  not g_19048 (not_new_n9988_, new_n9988_);
  or g_19049 (new_n5761_, not_new_n5940_, not_new_n5758_);
  not g_19050 (new_n4273_, new_n688_);
  not g_19051 (not_new_n3003_, new_n3003_);
  not g_19052 (not_new_n5471__0, new_n5471_);
  not g_19053 (not_new_n594__2, new_n594_);
  not g_19054 (new_n9911_, new_n639_);
  or g_19055 (new_n4763_, not_new_n4765__0, not_new_n4841__0);
  not g_19056 (not_new_n7305_, new_n7305_);
  not g_19057 (not_new_n1019__4, new_n1019_);
  not g_19058 (not_new_n5111_, new_n5111_);
  not g_19059 (not_new_n589__19773267430, new_n589_);
  and g_19060 (new_n1338_, new_n2309_, new_n2310_);
  not g_19061 (not_new_n3711_, new_n3711_);
  or g_19062 (new_n7453_, not_new_n6974__47475615099430, not_new_n749_);
  not g_19063 (not_new_n589__0, new_n589_);
  and g_19064 (new_n7695_, new_n7772_, new_n7782_);
  or g_19065 (new_n2042_, not_new_n9447_, not_new_n1584__3430);
  not g_19066 (not_new_n3820_, new_n3820_);
  or g_19067 (new_n6871_, not_new_n6870_, not_new_n6749_);
  or g_19068 (new_n3803_, not_new_n633__10, not_new_n1067__6);
  not g_19069 (not_new_n3325_, new_n3325_);
  or g_19070 (new_n2433_, not_new_n4131__0, not_new_n600__168070);
  not g_19071 (not_new_n7115_, new_n7115_);
  or g_19072 (new_n9285_, not_new_n1069__19773267430, not_new_n8877_);
  not g_19073 (new_n7164_, new_n7012_);
  not g_19074 (not_new_n7412_, new_n7412_);
  not g_19075 (not_new_n10258_, new_n10258_);
  not g_19076 (not_new_n1151_, new_n1151_);
  not g_19077 (not_new_n7066_, new_n7066_);
  not g_19078 (not_new_n645__6, new_n645_);
  or g_19079 (new_n5890_, not_new_n6008_, not_new_n6009_);
  not g_19080 (not_new_n9377__0, new_n9377_);
  or g_19081 (new_n7549_, not_new_n6995__2, not_new_n7030__0);
  not g_19082 (not_new_n6370__1, new_n6370_);
  not g_19083 (not_new_n3132_, new_n3132_);
  not g_19084 (not_new_n5716_, new_n5716_);
  not g_19085 (not_new_n1053__2326305139872070, new_n1053_);
  not g_19086 (not_new_n7882_, new_n7882_);
  not g_19087 (not_pi053, pi053);
  not g_19088 (not_new_n8986_, new_n8986_);
  not g_19089 (not_new_n6975__1, new_n6975_);
  or g_19090 (new_n4387_, not_new_n4312_, not_new_n4384_);
  not g_19091 (not_new_n4460__0, new_n4460_);
  not g_19092 (new_n5207_, new_n5061_);
  xor g_19093 (key_gate_122, key_122, new_n1182_);
  not g_19094 (not_new_n7410_, new_n7410_);
  not g_19095 (not_new_n619__8235430, new_n619_);
  or g_19096 (new_n5201_, not_new_n5286_, not_new_n5043_);
  or g_19097 (new_n7538_, not_new_n7536_, not_new_n7218_);
  not g_19098 (not_new_n3069_, new_n3069_);
  not g_19099 (not_new_n585__6, new_n585_);
  or g_19100 (new_n2945_, or_not_new_n2944__not_new_n2943_, not_new_n2942_);
  not g_19101 (not_new_n9319_, new_n9319_);
  or g_19102 (new_n6103_, not_new_n5879_, not_new_n5942__0);
  not g_19103 (not_new_n4169__0, new_n4169_);
  or g_19104 (new_n5223_, new_n645_, new_n1071_);
  not g_19105 (not_new_n2015_, new_n2015_);
  or g_19106 (new_n9431_, not_new_n9724_, not_new_n9723_);
  not g_19107 (not_new_n4440__0, new_n4440_);
  not g_19108 (not_pi065, pi065);
  not g_19109 (not_new_n4449__0, new_n4449_);
  not g_19110 (not_new_n3372__8235430, new_n3372_);
  or g_19111 (new_n5672_, not_new_n5571_, not_new_n5670_);
  not g_19112 (not_new_n5352_, new_n5352_);
  or g_19113 (new_n3108_, not_new_n1039__3, not_new_n928__7);
  or g_19114 (new_n8408_, not_new_n626__39098210485829880490, not_new_n8158__1);
  or g_19115 (new_n7674_, not_new_n7991_, not_new_n7992_);
  not g_19116 (not_new_n8907_, new_n8907_);
  not g_19117 (not_new_n6493__0, new_n6493_);
  not g_19118 (not_pi266, pi266);
  not g_19119 (not_pi057_0, pi057);
  and g_19120 (new_n6593_, new_n6653_, new_n6625_);
  or g_19121 (new_n2658_, not_new_n4458__0, not_new_n610__24010);
  not g_19122 (new_n9386_, new_n638_);
  or g_19123 (new_n10178_, new_n645_, new_n1071_);
  or g_19124 (new_n3733_, not_new_n3454_, not_new_n1943_);
  not g_19125 (not_new_n2776_, new_n2776_);
  not g_19126 (not_new_n7529_, new_n7529_);
  not g_19127 (not_new_n6792_, new_n6792_);
  or g_19128 (new_n1638_, not_pi030, not_po296_1);
  not g_19129 (not_new_n8314__0, new_n8314_);
  or g_19130 (new_n9047_, not_new_n8934_, not_new_n9045_);
  not g_19131 (not_new_n7860_, new_n7860_);
  not g_19132 (not_pi034, pi034);
  not g_19133 (not_new_n1612__332329305696010, new_n1612_);
  not g_19134 (new_n5095_, new_n4933_);
  or g_19135 (new_n8769_, not_new_n1071__403536070, not_new_n8622_);
  not g_19136 (not_po296_11044276742439206463052992010, po296);
  not g_19137 (not_new_n5729_, new_n5729_);
  or g_19138 (new_n8783_, or_or_not_new_n8781__not_new_n8701__not_new_n8780_, not_new_n8712_);
  or g_19139 (new_n5000_, not_new_n5239_, not_new_n4966_);
  or g_19140 (new_n3807_, not_new_n3805_, not_new_n3806_);
  or g_19141 (new_n2145_, not_new_n4788_, not_new_n591__403536070);
  not g_19142 (not_new_n1584__70, new_n1584_);
  not g_19143 (not_new_n4533_, new_n4533_);
  not g_19144 (new_n8157_, new_n1055_);
  or g_19145 (or_not_new_n1315__not_new_n1313_, not_new_n1315_, not_new_n1313_);
  not g_19146 (not_new_n585__2, new_n585_);
  not g_19147 (not_new_n2090__0, new_n2090_);
  not g_19148 (not_new_n5284_, new_n5284_);
  or g_19149 (or_not_new_n1239__not_new_n1237_, not_new_n1239_, not_new_n1237_);
  not g_19150 (not_po298_2824752490, po298);
  not g_19151 (not_new_n9879__1, new_n9879_);
  not g_19152 (new_n4416_, new_n1010_);
  not g_19153 (not_new_n8308__0, new_n8308_);
  or g_19154 (new_n1765_, not_pi098, not_new_n588_);
  not g_19155 (not_new_n980_, new_n980_);
  not g_19156 (not_new_n596__7, key_gate_88);
  or g_19157 (new_n4933_, not_new_n5025_, not_new_n5094_);
  not g_19158 (not_new_n589__3119734822845423713013303218219760490, new_n589_);
  or g_19159 (new_n7676_, not_new_n8011_, not_new_n8010_);
  not g_19160 (not_new_n1031__138412872010, new_n1031_);
  not g_19161 (new_n6929_, new_n6605_);
  not g_19162 (not_new_n6134_, new_n6134_);
  not g_19163 (not_new_n9099_, new_n9099_);
  not g_19164 (not_new_n4054_, new_n4054_);
  not g_19165 (not_new_n7038__1, new_n7038_);
  and g_19166 (new_n9328_, new_n9531_, new_n9532_);
  not g_19167 (not_new_n7719_, new_n7719_);
  and g_19168 (and_and_new_n8723__new_n1174__new_n8719_, new_n8719_, and_new_n8723__new_n1174_);
  not g_19169 (not_new_n6978_, new_n6978_);
  or g_19170 (new_n2395_, not_new_n598__7, not_new_n1049__0);
  not g_19171 (not_new_n589__273687473400809163430, new_n589_);
  or g_19172 (new_n4672_, not_new_n4496__0, not_new_n4495_);
  not g_19173 (not_new_n1041__70, new_n1041_);
  not g_19174 (not_new_n598__6, new_n598_);
  not g_19175 (not_new_n9861_, new_n9861_);
  not g_19176 (not_new_n1585__70, new_n1585_);
  not g_19177 (not_new_n6491_, new_n6491_);
  or g_19178 (new_n8022_, not_new_n7749_, not_new_n7926_);
  not g_19179 (not_new_n1599__6782230728490, new_n1599_);
  not g_19180 (not_new_n737__1, new_n737_);
  or g_19181 (new_n4681_, not_new_n1015__3, not_new_n4441_);
  or g_19182 (or_or_not_new_n2874__not_new_n2877__not_new_n2876_, or_not_new_n2874__not_new_n2877_, not_new_n2876_);
  not g_19183 (not_new_n3659_, new_n3659_);
  not g_19184 (not_new_n984__19773267430, new_n984_);
  or g_19185 (new_n2775_, or_not_new_n2774__not_new_n2773_, not_new_n2772_);
  not g_19186 (not_new_n3310__2, new_n3310_);
  not g_19187 (not_new_n9428__0, new_n9428_);
  not g_19188 (not_new_n3797_, new_n3797_);
  or g_19189 (new_n4732_, not_new_n4733_, or_not_new_n4816__not_new_n4751_);
  not g_19190 (not_new_n5742__2, new_n5742_);
  not g_19191 (not_new_n6462_, new_n6462_);
  or g_19192 (new_n6809_, not_new_n6584_, not_new_n6635__4);
  not g_19193 (not_new_n9053_, new_n9053_);
  not g_19194 (not_new_n636__9, new_n636_);
  not g_19195 (not_new_n1448_, new_n1448_);
  or g_19196 (new_n5709_, not_new_n5705_, or_not_new_n5453__not_new_n5706__1);
  and g_19197 (new_n10025_, new_n10341_, new_n10340_);
  or g_19198 (new_n8433_, not_new_n8266__0, not_new_n8089_);
  not g_19199 (not_new_n5695_, new_n5695_);
  or g_19200 (po132, not_new_n3475_, not_new_n3476_);
  or g_19201 (new_n8532_, not_new_n8260_, not_new_n8389_);
  not g_19202 (not_new_n6443__47475615099430, new_n6443_);
  or g_19203 (new_n2763_, not_new_n604__3, not_new_n642__2);
  not g_19204 (not_new_n8931_, new_n8931_);
  not g_19205 (not_new_n1071__2, new_n1071_);
  or g_19206 (new_n6670_, not_new_n631__2824752490, not_new_n6475_);
  not g_19207 (not_new_n641__0, new_n641_);
  not g_19208 (not_new_n7768__0, new_n7768_);
  not g_19209 (not_new_n1607__2824752490, new_n1607_);
  not g_19210 (not_new_n1022_, new_n1022_);
  not g_19211 (not_new_n3084_, new_n3084_);
  not g_19212 (not_new_n7394_, new_n7394_);
  not g_19213 (new_n8163_, new_n638_);
  xnor g_19214 (key_gate_114, key_114, new_n3998_);
  not g_19215 (not_new_n3145_, new_n3145_);
  not g_19216 (not_new_n586__403536070, new_n586_);
  not g_19217 (not_new_n638__797922662976120010, new_n638_);
  not g_19218 (not_new_n3833_, new_n3833_);
  or g_19219 (new_n9714_, not_new_n9623__0, not_new_n9620_);
  not g_19220 (not_new_n6535_, new_n6535_);
  not g_19221 (new_n7011_, new_n721_);
  or g_19222 (or_not_new_n2575__not_new_n2574_, not_new_n2575_, not_new_n2574_);
  not g_19223 (not_new_n645__168070, new_n645_);
  not g_19224 (new_n8153_, new_n1059_);
  not g_19225 (not_new_n604__24010, new_n604_);
  not g_19226 (new_n2190_, new_n630_);
  not g_19227 (not_new_n6554_, new_n6554_);
  not g_19228 (new_n6213_, new_n5874_);
  not g_19229 (not_new_n1012__1, new_n1012_);
  not g_19230 (new_n8656_, new_n1160_);
  or g_19231 (new_n9638_, new_n1599_, new_n622_);
  or g_19232 (new_n3253_, not_new_n1043__5, not_new_n589__39098210485829880490);
  or g_19233 (new_n7855_, not_new_n1603__1176490, not_new_n7629_);
  not g_19234 (not_new_n5680_, new_n5680_);
  or g_19235 (new_n4218_, not_new_n4088_, not_new_n4161__1);
  or g_19236 (new_n5584_, not_new_n1011__6, not_pi147_2);
  or g_19237 (new_n3175_, not_new_n642__5, not_new_n581__881247870897231951843937366879128181133112010);
  not g_19238 (not_new_n5078__2, new_n5078_);
  not g_19239 (not_new_n1047__6, new_n1047_);
  not g_19240 (not_new_n8846_, new_n8846_);
  not g_19241 (not_new_n7754__2, new_n7754_);
  and g_19242 (and_new_n10032__new_n580_, new_n10032_, new_n580_);
  or g_19243 (new_n9554_, not_new_n9375_, not_new_n9519_);
  not g_19244 (not_new_n6763_, new_n6763_);
  not g_19245 (not_new_n631__403536070, new_n631_);
  or g_19246 (new_n9282_, not_new_n9161_, not_new_n8898__1);
  not g_19247 (not_new_n9943_, new_n9943_);
  not g_19248 (not_new_n5426__0, new_n5426_);
  or g_19249 (new_n8428_, not_new_n8173_, not_new_n8373_);
  not g_19250 (new_n2066_, new_n958_);
  or g_19251 (new_n6645_, not_new_n6588_, not_new_n6622_);
  not g_19252 (not_new_n7113__1, new_n7113_);
  or g_19253 (new_n9289_, not_new_n633__332329305696010, not_new_n8885__0);
  not g_19254 (not_new_n608__4, new_n608_);
  not g_19255 (not_new_n7044_, new_n7044_);
  and g_19256 (new_n8668_, and_new_n8667__new_n8666_, new_n8758_);
  not g_19257 (not_new_n5400_, new_n5400_);
  and g_19258 (and_and_new_n8724__new_n8726__new_n8728_, new_n8728_, and_new_n8724__new_n8726_);
  not g_19259 (not_new_n1009__5, new_n1009_);
  or g_19260 (new_n8966_, not_new_n9095_, not_new_n9094_);
  not g_19261 (not_new_n2147__0, new_n2147_);
  or g_19262 (new_n3417_, not_new_n1536__1176490, not_pi029_0);
  not g_19263 (not_new_n8329_, new_n8329_);
  not g_19264 (not_new_n618__8, new_n618_);
  not g_19265 (not_new_n613__5, new_n613_);
  not g_19266 (not_new_n6450_, new_n6450_);
  and g_19267 (and_new_n1446__new_n2659_, new_n1446_, new_n2659_);
  not g_19268 (not_new_n627__968890104070, new_n627_);
  not g_19269 (not_new_n10123_, new_n10123_);
  not g_19270 (not_new_n641__7, new_n641_);
  or g_19271 (new_n6746_, not_new_n6538_, not_new_n6539__0);
  and g_19272 (and_and_new_n4298__new_n4341__new_n4345_, and_new_n4298__new_n4341_, new_n4345_);
  or g_19273 (new_n5399_, not_new_n1063__10, not_new_n4958__0);
  not g_19274 (not_new_n9726_, new_n9726_);
  or g_19275 (or_or_not_new_n8528__not_new_n8429__not_new_n8457_, not_new_n8457_, or_not_new_n8528__not_new_n8429_);
  or g_19276 (new_n9131_, new_n645_, new_n1071_);
  not g_19277 (not_new_n4966_, new_n4966_);
  not g_19278 (not_new_n1202_, new_n1202_);
  not g_19279 (not_new_n8054_, new_n8054_);
  not g_19280 (not_new_n3075_, new_n3075_);
  not g_19281 (not_new_n1604__7, new_n1604_);
  not g_19282 (not_new_n645__9, new_n645_);
  or g_19283 (new_n9905_, not_new_n645__16284135979104490, not_new_n1071__6782230728490);
  not g_19284 (not_new_n3200_, new_n3200_);
  and g_19285 (po105, key_gate_101, pi084);
  or g_19286 (new_n9737_, not_new_n9357__0, not_new_n631__657123623635342801395430);
  or g_19287 (new_n933_, not_new_n1028__1, not_new_n1623_);
  not g_19288 (not_new_n9058_, new_n9058_);
  not g_19289 (not_new_n4568_, new_n4568_);
  or g_19290 (new_n3048_, not_new_n1168_, not_new_n1027__138412872010);
  not g_19291 (not_new_n8573_, new_n8573_);
  and g_19292 (new_n8080_, new_n8346_, new_n8347_);
  not g_19293 (not_new_n3519_, new_n3519_);
  not g_19294 (not_new_n1534__403536070, key_gate_5);
  not g_19295 (not_new_n1045__5, new_n1045_);
  not g_19296 (not_new_n1161__0, new_n1161_);
  or g_19297 (new_n1013_, not_new_n3348_, not_new_n3347_);
  not g_19298 (not_new_n611__403536070, new_n611_);
  or g_19299 (new_n4578_, new_n1011_, pi179);
  not g_19300 (not_new_n5495_, new_n5495_);
  not g_19301 (not_new_n7347_, new_n7347_);
  or g_19302 (new_n657_, not_new_n3129_, or_not_new_n3130__not_new_n3131_);
  or g_19303 (new_n8014_, not_new_n8012_, not_new_n8013_);
  and g_19304 (new_n8936_, new_n9049_, new_n9172_);
  or g_19305 (new_n5274_, not_new_n5162_, not_new_n5159__0);
  not g_19306 (not_new_n3576_, new_n3576_);
  not g_19307 (not_new_n6745__0, new_n6745_);
  not g_19308 (not_new_n9979_, new_n9979_);
  and g_19309 (and_and_new_n6369__new_n6320__new_n6230_, new_n6230_, and_new_n6369__new_n6320_);
  and g_19310 (new_n1246_, new_n1872_, new_n1873_);
  or g_19311 (new_n3212_, not_new_n3185__490, not_new_n1602__4);
  or g_19312 (or_or_not_new_n1773__not_new_n1213__not_new_n1214_, not_new_n1214_, or_not_new_n1773__not_new_n1213_);
  not g_19313 (not_new_n1599__403536070, new_n1599_);
  not g_19314 (not_new_n9424_, new_n9424_);
  not g_19315 (not_new_n8159_, new_n8159_);
  not g_19316 (not_new_n4791_, new_n4791_);
  or g_19317 (new_n4500_, not_new_n4560_, not_new_n4559_);
  not g_19318 (not_new_n9644_, new_n9644_);
  not g_19319 (not_new_n3372__797922662976120010, new_n3372_);
  or g_19320 (new_n8356_, not_new_n8148_, not_new_n633__138412872010);
  not g_19321 (not_new_n1065__47475615099430, new_n1065_);
  not g_19322 (not_new_n630__24010, new_n630_);
  not g_19323 (not_new_n8104__0, new_n8104_);
  or g_19324 (new_n3785_, not_new_n1031__9, not_new_n641__8);
  not g_19325 (not_new_n1548_, new_n1548_);
  or g_19326 (new_n6367_, or_not_new_n6373__not_new_n6413_, not_new_n6232_);
  not g_19327 (not_new_n6908_, new_n6908_);
  or g_19328 (new_n6698_, not_new_n631__138412872010, not_new_n6475__1);
  or g_19329 (new_n2686_, or_not_new_n2685__not_new_n2684_, not_new_n2683_);
  not g_19330 (not_new_n1071__3430, new_n1071_);
  or g_19331 (new_n7668_, not_new_n7857_, not_new_n7918_);
  not g_19332 (not_new_n3560_, new_n3560_);
  not g_19333 (not_new_n7007_, new_n7007_);
  not g_19334 (not_new_n6057_, new_n6057_);
  not g_19335 (not_new_n8653__0, new_n8653_);
  not g_19336 (not_new_n626__57648010, new_n626_);
  or g_19337 (new_n3023_, not_new_n1160_, not_new_n1027__24010);
  not g_19338 (not_pi257_3, pi257);
  or g_19339 (new_n2926_, not_new_n4128__1, not_new_n994__968890104070);
  not g_19340 (not_new_n4275_, new_n4275_);
  not g_19341 (not_new_n3802_, new_n3802_);
  and g_19342 (new_n1550_, new_n3613_, new_n3612_);
  not g_19343 (not_new_n612__7, new_n612_);
  not g_19344 (not_new_n2772_, new_n2772_);
  and g_19345 (new_n1486_, new_n2940_, new_n2941_);
  not g_19346 (not_new_n1065__168070, new_n1065_);
  not g_19347 (not_new_n4319__0, new_n4319_);
  not g_19348 (not_new_n1538__168070, new_n1538_);
  or g_19349 (or_not_pi245_0_not_new_n1625_, not_pi245_0, not_new_n1625_);
  not g_19350 (not_new_n4282_, new_n4282_);
  or g_19351 (new_n8192_, not_new_n8478_, not_new_n8477_);
  not g_19352 (not_new_n2284_, new_n2284_);
  or g_19353 (new_n2974_, not_new_n612__7, not_new_n4120__2);
  not g_19354 (not_new_n10004_, new_n10004_);
  not g_19355 (new_n1590_, new_n1575_);
  not g_19356 (not_new_n600__10, new_n600_);
  not g_19357 (not_new_n6575_, new_n6575_);
  not g_19358 (not_new_n8685_, new_n8685_);
  not g_19359 (not_new_n3388_, new_n3388_);
  not g_19360 (not_new_n603__7, new_n603_);
  not g_19361 (not_new_n4936_, new_n4936_);
  not g_19362 (new_n8651_, new_n1155_);
  not g_19363 (new_n5434_, new_n1009_);
  or g_19364 (new_n7355_, not_new_n7105_, not_new_n775__6);
  and g_19365 (new_n5840_, new_n5945_, new_n5946_);
  not g_19366 (not_new_n5798__0, new_n5798_);
  not g_19367 (not_new_n3663_, new_n3663_);
  or g_19368 (new_n7174_, not_new_n7025_, not_new_n7173_);
  or g_19369 (new_n9176_, not_new_n8937_, not_new_n8978__2);
  not g_19370 (not_new_n8271__1, new_n8271_);
  or g_19371 (new_n678_, not_new_n3141_, or_not_new_n3143__not_new_n3142_);
  not g_19372 (not_new_n4673_, new_n4673_);
  not g_19373 (not_new_n1588__39098210485829880490, new_n1588_);
  not g_19374 (not_new_n8859_, new_n8859_);
  not g_19375 (new_n8434_, new_n8262_);
  not g_19376 (not_pi210, pi210);
  not g_19377 (not_new_n1604__113988951853731430, new_n1604_);
  not g_19378 (not_new_n3125_, new_n3125_);
  not g_19379 (new_n4258_, new_n695_);
  not g_19380 (not_new_n594__138412872010, new_n594_);
  or g_19381 (new_n9485_, not_new_n9552_, not_new_n9564_);
  or g_19382 (new_n1011_, not_new_n3344_, not_new_n3343_);
  or g_19383 (new_n7915_, not_new_n7842_, not_new_n7840_);
  or g_19384 (new_n5520_, not_new_n5432_, not_new_n5431_);
  or g_19385 (or_or_or_not_new_n2820__not_new_n2823__not_new_n2822__not_new_n2824_, not_new_n2824_, or_or_not_new_n2820__not_new_n2823__not_new_n2822_);
  and g_19386 (new_n6307_, new_n6279_, new_n1599_);
  not g_19387 (not_new_n2718_, new_n2718_);
  not g_19388 (new_n4421_, pi165);
  not g_19389 (not_new_n618__9, new_n618_);
  not g_19390 (not_new_n1591__1, new_n1591_);
  or g_19391 (new_n2657_, not_new_n611__57648010, not_new_n2656_);
  not g_19392 (not_new_n1775_, new_n1775_);
  not g_19393 (not_new_n7366__1, new_n7366_);
  and g_19394 (new_n6344_, new_n6232_, new_n6384_);
  not g_19395 (not_new_n1406_, new_n1406_);
  not g_19396 (not_new_n10027_, new_n10027_);
  not g_19397 (not_new_n5511_, new_n5511_);
  not g_19398 (not_new_n6212_, new_n6212_);
  not g_19399 (not_new_n8097_, new_n8097_);
  not g_19400 (not_new_n5459_, new_n5459_);
  not g_19401 (not_new_n6526_, new_n6526_);
  or g_19402 (new_n6958_, not_new_n6547__0, not_new_n6778_);
  not g_19403 (not_new_n5079_, new_n5079_);
  not g_19404 (not_new_n9829_, new_n9829_);
  not g_19405 (not_new_n4112_, new_n4112_);
  or g_19406 (new_n7030_, not_new_n7414_, not_new_n7413_);
  not g_19407 (not_new_n1431_, new_n1431_);
  not g_19408 (not_new_n8869_, new_n8869_);
  not g_19409 (not_new_n8816_, new_n8816_);
  not g_19410 (not_new_n594__3, new_n594_);
  and g_19411 (and_and_new_n1801__new_n1804__new_n1802_, and_new_n1801__new_n1804_, new_n1802_);
  not g_19412 (not_new_n1604__332329305696010, new_n1604_);
  or g_19413 (new_n658_, not_new_n3132_, or_not_new_n3134__not_new_n3133_);
  not g_19414 (not_new_n637__6, new_n637_);
  or g_19415 (or_not_new_n1564__not_new_n2479_, not_new_n1564_, not_new_n2479_);
  not g_19416 (new_n5782_, new_n646_);
  not g_19417 (not_new_n648__797922662976120010, new_n648_);
  and g_19418 (and_new_n2424__new_n2423_, new_n2424_, new_n2423_);
  not g_19419 (not_new_n601__3, new_n601_);
  or g_19420 (new_n993_, not_new_n1588_, not_new_n590__0);
  not g_19421 (not_new_n10075_, new_n10075_);
  not g_19422 (not_new_n611__19773267430, new_n611_);
  or g_19423 (new_n9685_, not_new_n9356__1, not_new_n9563_);
  not g_19424 (not_pi275_3, pi275);
  buf g_19425 (po036, pi228);
  not g_19426 (not_new_n1043__1176490, new_n1043_);
  not g_19427 (not_new_n8934_, new_n8934_);
  not g_19428 (not_new_n7454_, new_n7454_);
  or g_19429 (new_n3323_, not_new_n3925__0, not_pi064_3);
  not g_19430 (not_new_n7728_, new_n7728_);
  and g_19431 (new_n3966_, and_not_pi034_2_not_pi033_4, not_pi035_2);
  not g_19432 (not_new_n7129_, new_n7129_);
  not g_19433 (not_new_n9835_, new_n9835_);
  not g_19434 (not_pi238, pi238);
  and g_19435 (new_n6448_, new_n6714_, new_n6651_);
  or g_19436 (new_n9416_, not_new_n9710_, not_new_n9468_);
  or g_19437 (or_not_new_n5430__0_not_pi130_2, not_pi130_2, not_new_n5430__0);
  not g_19438 (not_pi116, pi116);
  xnor g_19439 (key_gate_15, new_n3932_, key_15);
  or g_19440 (new_n3186_, not_new_n3185_, not_new_n1051__4);
  buf g_19441 (po048, pi216);
  or g_19442 (new_n4370_, not_new_n661_, not_new_n4262_);
  or g_19443 (new_n9627_, new_n1600_, new_n629_);
  or g_19444 (new_n4746_, not_new_n4770_, or_not_new_n4839__not_new_n4767_);
  not g_19445 (not_new_n581_, new_n581_);
  not g_19446 (not_new_n7024_, new_n7024_);
  or g_19447 (or_not_new_n2617__not_new_n2621_, not_new_n2621_, not_new_n2617_);
  not g_19448 (new_n10152_, new_n10013_);
  not g_19449 (not_new_n4125__0, new_n4125_);
  not g_19450 (not_new_n643__113988951853731430, new_n643_);
  or g_19451 (po268, or_or_or_not_new_n2740__not_new_n2743__not_new_n2742__not_new_n2744_, not_new_n2741_);
  not g_19452 (not_new_n9487__0, new_n9487_);
  and g_19453 (new_n6466_, new_n6752_, new_n6783_);
  not g_19454 (not_new_n984__6, new_n984_);
  not g_19455 (not_new_n624__57648010, new_n624_);
  or g_19456 (or_not_new_n2765__not_new_n2764_, not_new_n2764_, not_new_n2765_);
  not g_19457 (not_new_n6639_, new_n6639_);
  not g_19458 (not_new_n5759_, new_n5759_);
  not g_19459 (not_new_n2264_, new_n2264_);
  or g_19460 (new_n1915_, not_new_n9875_, not_new_n594__6);
  not g_19461 (not_new_n630__6782230728490, new_n630_);
  not g_19462 (not_new_n6529_, new_n6529_);
  or g_19463 (new_n9587_, not_new_n9583_, not_new_n9585_);
  or g_19464 (new_n9711_, not_new_n9423_, not_new_n9618_);
  not g_19465 (new_n4977_, new_n646_);
  and g_19466 (new_n4902_, new_n5151_, new_n5152_);
  not g_19467 (not_new_n7008__1, new_n7008_);
  or g_19468 (new_n6865_, not_new_n6863_, not_new_n6864_);
  or g_19469 (new_n3583_, not_new_n2318__0, not_new_n1612__2326305139872070);
  not g_19470 (not_new_n7067_, new_n7067_);
  not g_19471 (not_new_n7887_, new_n7887_);
  not g_19472 (not_new_n3949_, new_n3949_);
  not g_19473 (not_new_n8618_, new_n8618_);
  or g_19474 (new_n8768_, not_new_n8662_, not_new_n8722_);
  or g_19475 (new_n3578_, not_new_n1538__47475615099430, not_pi155_0);
  not g_19476 (not_new_n8854__0, new_n8854_);
  not g_19477 (not_new_n1438_, new_n1438_);
  not g_19478 (not_new_n8572_, new_n8572_);
  or g_19479 (new_n8062_, not_new_n7938_, not_new_n8061_);
  not g_19480 (new_n3414_, new_n1037_);
  or g_19481 (po144, not_new_n3515_, not_new_n3514_);
  not g_19482 (not_new_n2684_, new_n2684_);
  not g_19483 (not_new_n621__24010, new_n621_);
  not g_19484 (not_new_n5734_, new_n5734_);
  not g_19485 (not_pi247, pi247);
  not g_19486 (not_new_n589__70, new_n589_);
  not g_19487 (not_new_n581__1915812313805664144010, new_n581_);
  not g_19488 (not_new_n1067__490, new_n1067_);
  not g_19489 (not_pi054_0, pi054);
  not g_19490 (not_new_n5508_, new_n5508_);
  not g_19491 (not_new_n636__1, new_n636_);
  not g_19492 (not_new_n6586_, new_n6586_);
  or g_19493 (new_n2427_, not_new_n637__1, not_new_n603__24010);
  and g_19494 (new_n7703_, new_n7773_, new_n7963_);
  not g_19495 (not_new_n6983__1, new_n6983_);
  not g_19496 (not_new_n9900__1, new_n9900_);
  not g_19497 (not_new_n4989_, new_n4989_);
  not g_19498 (not_new_n9506__2, new_n9506_);
  or g_19499 (new_n7407_, not_new_n7117_, not_new_n775__70);
  or g_19500 (new_n9186_, not_new_n9092_, not_new_n9095__0);
  not g_19501 (not_new_n2945_, new_n2945_);
  not g_19502 (not_new_n8848__0, new_n8848_);
  and g_19503 (new_n610_, new_n592_, new_n583_);
  not g_19504 (not_new_n4448_, new_n4448_);
  not g_19505 (not_new_n639__273687473400809163430, new_n639_);
  or g_19506 (new_n5359_, not_new_n4987__0, not_new_n1601__10);
  not g_19507 (not_new_n8177__0, new_n8177_);
  or g_19508 (new_n3198_, not_new_n3185__5, not_new_n1039__4);
  not g_19509 (not_new_n594__2326305139872070, new_n594_);
  or g_19510 (new_n4120_, not_new_n4191_, not_new_n4192_);
  not g_19511 (not_new_n7600__0, new_n7600_);
  not g_19512 (not_new_n4756_, new_n4756_);
  and g_19513 (new_n8211_, new_n8285_, new_n8487_);
  not g_19514 (not_new_n3372__273687473400809163430, new_n3372_);
  or g_19515 (new_n5376_, not_new_n1604__10, not_new_n4997__0);
  not g_19516 (not_new_n2484_, new_n2484_);
  or g_19517 (new_n3492_, not_pi014_0, not_new_n1536__5585458640832840070);
  not g_19518 (not_new_n6309_, new_n6309_);
  or g_19519 (new_n10288_, not_new_n9941_, not_new_n621__273687473400809163430);
  not g_19520 (not_pi164, pi164);
  not g_19521 (not_new_n5192_, new_n5192_);
  and g_19522 (new_n6359_, new_n6421_, new_n6420_);
  not g_19523 (not_new_n6341_, new_n6341_);
  not g_19524 (not_new_n5995_, new_n5995_);
  or g_19525 (new_n4892_, not_new_n4805_, not_new_n1057__8);
  or g_19526 (new_n9067_, new_n1067_, new_n633_);
  not g_19527 (not_new_n1604__403536070, new_n1604_);
  not g_19528 (not_po298_138412872010, po298);
  not g_19529 (not_new_n634__332329305696010, new_n634_);
  not g_19530 (not_new_n621__490, new_n621_);
  not g_19531 (not_new_n1537__57648010, new_n1537_);
  not g_19532 (new_n7442_, new_n7037_);
  not g_19533 (not_new_n648__1176490, new_n648_);
  not g_19534 (new_n5947_, new_n5878_);
  not g_19535 (not_new_n2636_, new_n2636_);
  not g_19536 (not_new_n604__403536070, new_n604_);
  not g_19537 (not_new_n4506_, new_n4506_);
  not g_19538 (not_new_n622__138412872010, new_n622_);
  not g_19539 (new_n8861_, new_n626_);
  not g_19540 (not_new_n1051__0, new_n1051_);
  or g_19541 (new_n5100_, not_new_n5099_, not_new_n631__3430);
  not g_19542 (not_new_n604__3, new_n604_);
  not g_19543 (not_new_n4877_, new_n4877_);
  not g_19544 (not_new_n581__1, new_n581_);
  not g_19545 (not_new_n732__1, new_n732_);
  not g_19546 (not_new_n5799__0, new_n5799_);
  or g_19547 (new_n1150_, not_new_n3830_, not_new_n3829_);
  not g_19548 (not_pi062, pi062);
  not g_19549 (not_new_n6158_, new_n6158_);
  not g_19550 (not_new_n3448_, new_n3448_);
  or g_19551 (new_n10267_, not_new_n619__968890104070, not_new_n10009_);
  not g_19552 (not_new_n5539_, new_n5539_);
  and g_19553 (new_n7710_, new_n7861_, new_n7922_);
  not g_19554 (not_new_n8536_, new_n8536_);
  or g_19555 (new_n5099_, not_new_n4929_, not_new_n4928_);
  not g_19556 (not_new_n4809__0, new_n4809_);
  not g_19557 (not_new_n1065__138412872010, new_n1065_);
  not g_19558 (new_n3393_, new_n1030_);
  not g_19559 (not_new_n2334_, new_n2334_);
  or g_19560 (or_not_new_n3094__not_new_n3093_, not_new_n3094_, not_new_n3093_);
  or g_19561 (new_n7865_, not_new_n7864_, not_new_n7622_);
  or g_19562 (new_n1736_, not_new_n1728__4, not_pi080);
  or g_19563 (new_n3283_, not_new_n589__185621159210175743024531636712070, not_new_n1067__5);
  not g_19564 (not_new_n5537_, new_n5537_);
  or g_19565 (new_n6165_, not_new_n5894_, not_new_n6064__0);
  not g_19566 (not_new_n2338_, new_n2338_);
  not g_19567 (not_new_n5478__0, new_n5478_);
  not g_19568 (not_new_n5510_, new_n5510_);
  or g_19569 (new_n7927_, not_new_n7754__1, not_new_n7584_);
  not g_19570 (not_pi094, pi094);
  or g_19571 (new_n2445_, not_new_n598__8235430, not_new_n1069__0);
  or g_19572 (new_n9581_, not_new_n9330_, not_new_n9513_);
  not g_19573 (not_new_n625__138412872010, new_n625_);
  not g_19574 (not_new_n5615_, new_n5615_);
  not g_19575 (new_n9398_, new_n643_);
  not g_19576 (not_new_n9970__0, new_n9970_);
  not g_19577 (not_new_n4296_, new_n4296_);
  not g_19578 (not_new_n2246_, new_n2246_);
  not g_19579 (new_n7002_, new_n730_);
  not g_19580 (not_new_n9171_, new_n9171_);
  not g_19581 (not_new_n8681_, new_n8681_);
  not g_19582 (not_pi138, pi138);
  or g_19583 (new_n9187_, or_not_new_n9103__not_new_n8987__0, not_new_n8979__0);
  not g_19584 (not_new_n3184__5, new_n3184_);
  not g_19585 (not_new_n648__0, new_n648_);
  not g_19586 (not_new_n1365_, new_n1365_);
  not g_19587 (not_new_n6492__0, new_n6492_);
  not g_19588 (not_new_n632__1176490, new_n632_);
  or g_19589 (po139, not_new_n3504_, not_new_n3505_);
  or g_19590 (new_n1575_, not_new_n1580_, not_new_n3372__2);
  not g_19591 (not_new_n625__113988951853731430, new_n625_);
  not g_19592 (not_new_n8713__1, new_n8713_);
  not g_19593 (not_new_n5513__0, new_n5513_);
  not g_19594 (not_new_n1536__5585458640832840070, new_n1536_);
  or g_19595 (new_n8023_, not_new_n1604__8235430, not_new_n7634__0);
  not g_19596 (not_new_n5278_, new_n5278_);
  not g_19597 (new_n5749_, new_n628_);
  not g_19598 (not_new_n4191_, new_n4191_);
  not g_19599 (not_new_n8845__0, new_n8845_);
  not g_19600 (not_new_n3528_, new_n3528_);
  xnor g_19601 (key_gate_49, key_49, new_n1648_);
  not g_19602 (not_new_n7951_, new_n7951_);
  not g_19603 (not_new_n639__19773267430, new_n639_);
  not g_19604 (not_pi169, pi169);
  not g_19605 (not_new_n693_, new_n693_);
  not g_19606 (not_new_n8958__0, new_n8958_);
  not g_19607 (not_new_n4028_, new_n4028_);
  not g_19608 (not_new_n3185__6782230728490, new_n3185_);
  or g_19609 (new_n4871_, not_new_n4777__0, not_new_n4836_);
  or g_19610 (new_n3601_, not_new_n948_, not_new_n1611__4);
  or g_19611 (new_n10087_, not_new_n9985_, not_new_n10085_);
  or g_19612 (new_n8007_, not_new_n7625__0, not_new_n1600__8235430);
  not g_19613 (not_new_n9693_, new_n9693_);
  or g_19614 (new_n3854_, not_new_n1576__490, not_new_n622__490);
  not g_19615 (not_po298_57648010, po298);
  not g_19616 (not_new_n1041__4, new_n1041_);
  or g_19617 (new_n3189_, not_new_n648__7, not_new_n589__0);
  or g_19618 (new_n9584_, new_n627_, new_n1055_);
  not g_19619 (not_new_n3041_, new_n3041_);
  not g_19620 (not_new_n7801_, new_n7801_);
  not g_19621 (not_new_n1053__10, new_n1053_);
  not g_19622 (not_new_n8267_, new_n8267_);
  or g_19623 (new_n4889_, not_new_n4799__0, not_new_n4828_);
  or g_19624 (new_n9731_, not_new_n9364_, not_new_n1047__47475615099430);
  not g_19625 (not_new_n5773_, new_n5773_);
  not g_19626 (not_new_n5372_, new_n5372_);
  not g_19627 (not_new_n4468_, new_n4468_);
  or g_19628 (new_n4852_, not_new_n4755_, not_new_n1605__4);
  or g_19629 (new_n4485_, not_new_n4515_, not_new_n4516_);
  and g_19630 (new_n1388_, new_n2455_, new_n2456_);
  and g_19631 (new_n6447_, new_n6704_, new_n6705_);
  not g_19632 (not_new_n6094_, new_n6094_);
  not g_19633 (not_new_n4410__0, new_n4410_);
  or g_19634 (new_n6015_, not_new_n5808_, not_new_n1596__490);
  not g_19635 (not_new_n3311__8235430, new_n3311_);
  not g_19636 (not_new_n4930__1, new_n4930_);
  not g_19637 (not_new_n4431_, new_n4431_);
  or g_19638 (new_n8383_, not_new_n8224_, not_new_n8275_);
  not g_19639 (not_new_n1027__7, new_n1027_);
  not g_19640 (new_n7248_, new_n7141_);
  or g_19641 (new_n1672_, not_new_n596__490, key_gate_84);
  not g_19642 (not_new_n9365__0, new_n9365_);
  not g_19643 (not_new_n1604__10, new_n1604_);
  and g_19644 (new_n7696_, new_n7785_, new_n7784_);
  not g_19645 (not_new_n7250_, new_n7250_);
  not g_19646 (not_new_n3915__0, key_gate_66);
  not g_19647 (not_new_n6232_, new_n6232_);
  and g_19648 (new_n9870_, new_n10172_, new_n10175_);
  not g_19649 (not_new_n1419_, new_n1419_);
  not g_19650 (not_new_n7929_, new_n7929_);
  or g_19651 (or_or_or_not_new_n1773__not_new_n1213__not_new_n1214__not_new_n1775_, not_new_n1775_, or_or_not_new_n1773__not_new_n1213__not_new_n1214_);
  not g_19652 (not_new_n632__2824752490, new_n632_);
  not g_19653 (not_new_n928__6782230728490, new_n928_);
  not g_19654 (not_new_n1071__8, new_n1071_);
  and g_19655 (new_n6353_, new_n6266_, and_new_n6373__new_n6389_);
  not g_19656 (not_new_n4131_, new_n4131_);
  or g_19657 (new_n9323_, not_new_n1053__968890104070, not_new_n8861_);
  or g_19658 (new_n4221_, not_pi263_2, not_new_n4083_);
  not g_19659 (not_new_n10081_, new_n10081_);
  not g_19660 (not_new_n7626__0, new_n7626_);
  not g_19661 (not_new_n7592_, new_n7592_);
  not g_19662 (not_new_n1055__9, new_n1055_);
  or g_19663 (new_n2359_, not_new_n9953__0, not_new_n599__0);
  not g_19664 (not_new_n6505_, new_n6505_);
  not g_19665 (new_n4412_, pi161);
  not g_19666 (not_new_n3763_, new_n3763_);
  or g_19667 (new_n4706_, not_new_n4705_, not_new_n4704_);
  or g_19668 (new_n1720_, key_gate_39, not_new_n596__16284135979104490);
  or g_19669 (new_n2291_, not_new_n6466_, not_new_n1580__2326305139872070);
  or g_19670 (new_n2470_, not_new_n598__138412872010, not_new_n1601__0);
  or g_19671 (new_n6386_, not_new_n639__57648010, not_new_n6299_);
  not g_19672 (not_new_n626__3430, new_n626_);
  not g_19673 (not_new_n1045__273687473400809163430, new_n1045_);
  or g_19674 (new_n1851_, not_new_n1585__3, not_new_n5829_);
  or g_19675 (new_n3402_, not_new_n3312_, not_new_n927__1);
  or g_19676 (new_n6688_, not_new_n6687_, not_new_n6575_);
  or g_19677 (new_n9802_, not_new_n9801_, not_new_n9800_);
  or g_19678 (new_n9030_, not_new_n9029_, not_new_n8846_);
  or g_19679 (new_n7998_, not_new_n1598__8235430, not_new_n7661__0);
  not g_19680 (new_n8836_, new_n634_);
  not g_19681 (not_new_n3255_, new_n3255_);
  not g_19682 (not_new_n702_, new_n702_);
  not g_19683 (new_n7599_, new_n1043_);
  not g_19684 (not_new_n609__10, new_n609_);
  or g_19685 (new_n1618_, not_new_n590__3, not_new_n1587_);
  not g_19686 (not_new_n1581__6782230728490, new_n1581_);
  not g_19687 (not_new_n2824_, new_n2824_);
  and g_19688 (new_n3928_, new_n3942_, new_n4022_);
  and g_19689 (and_new_n6395__new_n6396_, new_n6396_, new_n6395_);
  or g_19690 (new_n5775_, not_new_n5776_, not_new_n639__1176490);
  not g_19691 (not_new_n5767__1, new_n5767_);
  not g_19692 (not_new_n1613__19773267430, new_n1613_);
  not g_19693 (not_new_n4843__0, new_n4843_);
  not g_19694 (not_new_n7154_, new_n7154_);
  not g_19695 (not_new_n9729_, new_n9729_);
  or g_19696 (new_n10042_, new_n1037_, new_n632_);
  or g_19697 (new_n2996_, not_new_n1047__2, not_new_n581__2);
  or g_19698 (or_not_new_n7046__not_new_n7265_, not_new_n7046_, not_new_n7265_);
  not g_19699 (not_new_n3372__47475615099430, new_n3372_);
  or g_19700 (new_n997_, not_new_n1028__4, not_new_n3375__3);
  not g_19701 (not_new_n8836_, new_n8836_);
  not g_19702 (not_new_n5677_, new_n5677_);
  not g_19703 (not_new_n631__10, new_n631_);
  or g_19704 (new_n3804_, not_new_n3802_, not_new_n3803_);
  or g_19705 (or_not_new_n5041__not_new_n4911_, not_new_n5041_, not_new_n4911_);
  not g_19706 (not_new_n7617_, new_n7617_);
  or g_19707 (new_n5581_, not_new_n5580_, not_new_n5474_);
  or g_19708 (po281, not_new_n2856_, or_or_not_new_n1482__not_new_n2858__not_new_n2857_);
  not g_19709 (not_new_n8656_, new_n8656_);
  or g_19710 (new_n8579_, not_new_n8160__0, not_new_n1057__2824752490);
  not g_19711 (not_new_n6870_, new_n6870_);
  not g_19712 (not_new_n596__10, key_gate_88);
  not g_19713 (not_new_n6687_, new_n6687_);
  not g_19714 (not_new_n7842_, new_n7842_);
  and g_19715 (new_n8931_, and_new_n8828__new_n9210_, new_n9209_);
  or g_19716 (new_n2233_, not_new_n8182_, not_new_n1581__968890104070);
  or g_19717 (new_n3208_, not_new_n3185__10, not_new_n1600__4);
  not g_19718 (not_new_n6539_, new_n6539_);
  not g_19719 (not_new_n5756__0, new_n5756_);
  not g_19720 (not_new_n1028__3, new_n1028_);
  or g_19721 (new_n1959_, not_new_n587__10, not_pi140);
  not g_19722 (not_new_n1043__9, new_n1043_);
  not g_19723 (not_new_n1002_, new_n1002_);
  not g_19724 (not_new_n5500_, new_n5500_);
  or g_19725 (new_n5582_, not_new_n1011__5, not_pi147_1);
  not g_19726 (not_new_n627__332329305696010, new_n627_);
  or g_19727 (or_or_not_new_n1299__not_new_n1297__not_new_n2116_, not_new_n2116_, or_not_new_n1299__not_new_n1297_);
  not g_19728 (not_new_n4487__0, new_n4487_);
  not g_19729 (not_new_n1584__0, new_n1584_);
  not g_19730 (not_new_n10144__0, new_n10144_);
  xor g_19731 (key_gate_91, key_91, not_new_n1687_);
  or g_19732 (new_n9317_, not_new_n627__47475615099430, not_new_n8864_);
  or g_19733 (new_n5710_, not_new_n5708_, not_new_n1019__6);
  not g_19734 (not_new_n618__70, new_n618_);
  not g_19735 (not_new_n5564_, new_n5564_);
  not g_19736 (not_new_n7777_, new_n7777_);
  not g_19737 (not_new_n1383_, new_n1383_);
  not g_19738 (not_new_n4330__0, new_n4330_);
  or g_19739 (new_n8891_, or_not_new_n9191__not_new_n9190_, not_new_n9100_);
  or g_19740 (new_n10144_, new_n1600_, new_n629_);
  or g_19741 (new_n3087_, not_new_n581__39098210485829880490, not_new_n647__5);
  or g_19742 (new_n4638_, not_new_n4417__0, not_new_n1009__4);
  or g_19743 (new_n9203_, not_new_n8836_, not_new_n1047__138412872010);
  or g_19744 (new_n7261_, not_new_n7259_, not_new_n7257_);
  not g_19745 (not_new_n1607__6, new_n1607_);
  and g_19746 (new_n1407_, new_n929_, and_new_n933__new_n935_);
  not g_19747 (not_new_n4751__0, new_n4751_);
  not g_19748 (not_new_n1589__138412872010, new_n1589_);
  not g_19749 (not_new_n10294_, new_n10294_);
  or g_19750 (new_n2577_, not_new_n611__10, not_new_n2576_);
  not g_19751 (not_new_n3941_, new_n3941_);
  not g_19752 (not_new_n638__6782230728490, new_n638_);
  not g_19753 (not_new_n635__7, new_n635_);
  not g_19754 (not_new_n646__968890104070, new_n646_);
  not g_19755 (not_pi132_0, pi132);
  not g_19756 (new_n6509_, new_n1603_);
  or g_19757 (new_n7682_, not_new_n8062_, not_new_n8063_);
  not g_19758 (new_n3459_, new_n1055_);
  not g_19759 (not_new_n3430_, new_n3430_);
  not g_19760 (not_new_n581__19773267430, new_n581_);
  not g_19761 (not_new_n1939_, new_n1939_);
  or g_19762 (or_not_new_n2675__not_new_n2674_, not_new_n2674_, not_new_n2675_);
  not g_19763 (not_new_n4719_, new_n4719_);
  or g_19764 (new_n2526_, or_not_new_n2525__not_new_n2524_, not_new_n2523_);
  not g_19765 (not_new_n8396_, new_n8396_);
  not g_19766 (not_new_n4911_, new_n4911_);
  or g_19767 (new_n6413_, not_new_n6412_, not_new_n6411_);
  or g_19768 (new_n3170_, not_new_n626__5, not_new_n3315__16284135979104490);
  not g_19769 (new_n7463_, new_n7046_);
  not g_19770 (new_n9357_, new_n1043_);
  not g_19771 (not_new_n625__7, new_n625_);
  not g_19772 (not_new_n5270_, new_n5270_);
  or g_19773 (new_n2017_, not_pi111, not_new_n588__3430);
  not g_19774 (not_new_n3372__57648010, new_n3372_);
  or g_19775 (po269, or_or_or_not_new_n2749__not_new_n2752__not_new_n2751__not_new_n2753_, not_new_n2750_);
  not g_19776 (not_new_n631__1, new_n631_);
  or g_19777 (new_n2369_, not_new_n9959__0, not_new_n599__2);
  not g_19778 (new_n9391_, new_n636_);
  or g_19779 (new_n2163_, not_new_n593__403536070, not_new_n639_);
  not g_19780 (not_new_n2304_, new_n2304_);
  and g_19781 (new_n7705_, new_n7772_, new_n7976_);
  buf g_19782 (po024, pi240);
  not g_19783 (not_new_n4014__4, new_n4014_);
  and g_19784 (new_n7574_, new_n7833_, new_n7834_);
  not g_19785 (not_new_n6007_, new_n6007_);
  not g_19786 (new_n1601_, new_n969_);
  not g_19787 (not_new_n10278_, new_n10278_);
  or g_19788 (new_n6410_, not_new_n6322_, not_new_n6321_);
  or g_19789 (new_n6867_, not_new_n6540__0, or_not_new_n618__19773267430_not_new_n6865_);
  not g_19790 (not_new_n3315__70, new_n3315_);
  not g_19791 (not_new_n8952_, new_n8952_);
  or g_19792 (new_n1688_, not_pi051, not_new_n1631__8235430);
  not g_19793 (not_pi006, pi006);
  or g_19794 (new_n6740_, not_new_n6501_, not_new_n1600__24010);
  or g_19795 (new_n3713_, not_po298_113988951853731430, not_new_n619__4);
  not g_19796 (not_new_n9391_, new_n9391_);
  not g_19797 (not_new_n625__3430, new_n625_);
  or g_19798 (new_n2178_, not_new_n1591__2824752490, not_new_n8816_);
  not g_19799 (new_n5087_, new_n4954_);
  not g_19800 (not_new_n2607_, new_n2607_);
  or g_19801 (new_n4710_, not_pi171_2, not_new_n4434_);
  or g_19802 (new_n5339_, not_new_n617__168070, not_new_n4948__0);
  and g_19803 (new_n6343_, new_n6373_, new_n6269_);
  or g_19804 (new_n6991_, or_not_new_n7313__not_new_n7314_, not_new_n7169_);
  not g_19805 (not_new_n9169_, new_n9169_);
  not g_19806 (not_new_n4502__0, new_n4502_);
  or g_19807 (new_n6440_, not_new_n6370_, or_not_new_n6373__9_not_new_n6237_);
  and g_19808 (and_and_and_not_pi051_1_not_pi050_1_not_pi049_1_not_pi048_1, and_and_not_pi051_1_not_pi050_1_not_pi049_1, not_pi048_1);
  and g_19809 (new_n1458_, and_and_new_n3768__new_n3771__new_n3777_, new_n3774_);
  not g_19810 (not_new_n3206_, new_n3206_);
  not g_19811 (not_new_n5430_, new_n5430_);
  not g_19812 (not_new_n2036_, new_n2036_);
  not g_19813 (not_pi117, pi117);
  or g_19814 (or_or_not_pi269_1_not_pi260_1_not_pi257_1, not_pi257_1, or_not_pi269_1_not_pi260_1);
  or g_19815 (new_n4523_, not_new_n4522_, not_new_n4483_);
  or g_19816 (new_n5293_, not_new_n4942_, not_new_n1051__9);
  or g_19817 (new_n2172_, not_new_n640__0, not_new_n601__403536070);
  or g_19818 (new_n3508_, not_pi120_0, not_new_n1537__138412872010);
  not g_19819 (not_new_n8701_, new_n8701_);
  and g_19820 (new_n591_, new_n3372_, and_new_n3375__new_n3387_);
  or g_19821 (new_n5294_, not_new_n5293_, not_new_n5292_);
  or g_19822 (new_n3812_, not_new_n1039__6, not_new_n628__10);
  not g_19823 (not_pi058, pi058);
  or g_19824 (new_n2484_, not_new_n599__47475615099430, not_new_n9872__0);
  or g_19825 (new_n5204_, not_new_n617__3430, not_new_n1597__8);
  or g_19826 (new_n2124_, not_new_n9968_, not_new_n594__8235430);
  not g_19827 (not_new_n4707_, new_n4707_);
  not g_19828 (not_new_n6539__1, new_n6539_);
  not g_19829 (not_new_n619__968890104070, new_n619_);
  not g_19830 (new_n5124_, new_n4947_);
  not g_19831 (not_new_n5041_, new_n5041_);
  or g_19832 (new_n6733_, not_new_n630__57648010, not_new_n6506_);
  or g_19833 (or_or_not_new_n6160__not_new_n6161__not_new_n6090_, or_not_new_n6160__not_new_n6161_, not_new_n6090_);
  not g_19834 (not_new_n4805_, new_n4805_);
  or g_19835 (new_n4639_, not_pi163_3, not_new_n4418__0);
  or g_19836 (new_n5347_, not_new_n1599__9, not_new_n4990_);
  not g_19837 (not_new_n5760_, new_n5760_);
  not g_19838 (not_new_n6993__0, new_n6993_);
  or g_19839 (new_n737_, not_new_n3247_, not_new_n3248_);
  not g_19840 (not_new_n1006__6, new_n1006_);
  not g_19841 (not_new_n621__3, new_n621_);
  not g_19842 (not_new_n4575_, new_n4575_);
  or g_19843 (new_n9440_, not_new_n9782_, not_new_n9783_);
  or g_19844 (new_n5641_, not_new_n5639_, not_new_n5522_);
  or g_19845 (or_or_not_new_n1251__not_new_n1249__not_new_n1888_, or_not_new_n1251__not_new_n1249_, not_new_n1888_);
  or g_19846 (new_n1759_, not_new_n1728__2326305139872070, not_pi073);
  not g_19847 (not_new_n1581__19773267430, new_n1581_);
  not g_19848 (not_new_n1063__968890104070, new_n1063_);
  not g_19849 (not_new_n9959__0, new_n9959_);
  or g_19850 (new_n1695_, not_pi011_0, not_po296_2824752490);
  or g_19851 (new_n7842_, not_new_n1067__168070, not_new_n7640_);
  or g_19852 (new_n6046_, not_new_n5974__0, not_new_n5976_);
  not g_19853 (not_new_n3310__10, new_n3310_);
  not g_19854 (not_new_n626__225393402906922580878632490, new_n626_);
  and g_19855 (new_n1240_, and_and_new_n1839__new_n1842__new_n1840_, new_n1841_);
  not g_19856 (new_n8631_, new_n1154_);
  or g_19857 (new_n6706_, not_new_n6660_, not_new_n6446_);
  not g_19858 (not_new_n1826_, new_n1826_);
  not g_19859 (new_n4082_, pi270);
  not g_19860 (not_new_n6038_, new_n6038_);
  not g_19861 (not_new_n3193_, new_n3193_);
  not g_19862 (not_new_n8713__0, new_n8713_);
  not g_19863 (not_new_n9484_, new_n9484_);
  or g_19864 (new_n4197_, not_pi258_1, not_new_n4104_);
  not g_19865 (not_new_n6039_, new_n6039_);
  not g_19866 (not_new_n5882__1, new_n5882_);
  not g_19867 (not_new_n4905_, new_n4905_);
  not g_19868 (not_new_n5112_, new_n5112_);
  or g_19869 (new_n5995_, not_new_n5777_, not_new_n1604__70);
  or g_19870 (new_n8041_, not_new_n7844_, not_new_n8040_);
  or g_19871 (new_n3711_, not_new_n618__8, not_po298_16284135979104490);
  not g_19872 (not_new_n1597__6782230728490, new_n1597_);
  not g_19873 (not_new_n1067_, new_n1067_);
  not g_19874 (not_new_n1065__70, new_n1065_);
  or g_19875 (new_n6017_, not_new_n5766__0, not_new_n5918__0);
  not g_19876 (not_new_n739_, new_n739_);
  not g_19877 (not_new_n4238_, new_n4238_);
  not g_19878 (not_new_n648_, new_n648_);
  or g_19879 (new_n5135_, new_n624_, new_n1041_);
  or g_19880 (po164, not_new_n3554_, not_new_n3555_);
  not g_19881 (new_n6261_, new_n638_);
  not g_19882 (not_new_n8158__0, new_n8158_);
  not g_19883 (not_new_n1063__1176490, new_n1063_);
  not g_19884 (not_new_n647__24010, new_n647_);
  and g_19885 (and_new_n1250__new_n1894_, new_n1250_, new_n1894_);
  not g_19886 (not_new_n625__3, new_n625_);
  and g_19887 (and_new_n5268__new_n5267_, new_n5267_, new_n5268_);
  not g_19888 (new_n5444_, new_n1005_);
  not g_19889 (new_n8640_, new_n1173_);
  not g_19890 (not_new_n7894_, new_n7894_);
  or g_19891 (new_n3567_, not_new_n1612__403536070, not_new_n2166__0);
  not g_19892 (not_pi064_5585458640832840070, pi064);
  or g_19893 (new_n7202_, not_new_n6982__1, not_new_n7354__1);
  not g_19894 (not_new_n8139__1, new_n8139_);
  not g_19895 (not_new_n1569_, new_n1569_);
  not g_19896 (not_new_n8662_, new_n8662_);
  or g_19897 (new_n8196_, not_new_n8532_, not_new_n8533_);
  not g_19898 (not_new_n3947_, new_n3947_);
  or g_19899 (new_n3441_, not_new_n1919_, not_new_n1613__6);
  not g_19900 (not_new_n7444_, new_n7444_);
  not g_19901 (not_new_n591__8, new_n591_);
  or g_19902 (new_n5004_, not_new_n5301_, not_new_n5300_);
  not g_19903 (not_new_n3960_, new_n3960_);
  or g_19904 (po208, or_or_not_new_n1565__not_new_n2484__not_new_n1399_, not_new_n1400_);
  or g_19905 (new_n4199_, not_pi271_1, not_new_n4102_);
  not g_19906 (not_new_n731__1, new_n731_);
  not g_19907 (new_n9130_, new_n8972_);
  or g_19908 (new_n3400_, not_new_n927__0, not_new_n1730__0);
  not g_19909 (not_new_n1596__10, new_n1596_);
  and g_19910 (new_n6570_, new_n6654_, new_n6664_);
  or g_19911 (new_n9084_, not_new_n639__47475615099430, not_new_n1603__19773267430);
  or g_19912 (new_n2522_, not_pi194, not_new_n2509__0);
  not g_19913 (not_new_n3924_, new_n3924_);
  not g_19914 (new_n7609_, new_n642_);
  and g_19915 (new_n1191_, new_n1664_, new_n1662_);
  not g_19916 (not_new_n1504_, new_n1504_);
  not g_19917 (not_new_n603__8, new_n603_);
  not g_19918 (not_new_n7385_, new_n7385_);
  not g_19919 (not_new_n1267_, new_n1267_);
  not g_19920 (not_new_n741_, new_n741_);
  not g_19921 (not_new_n596__1176490, key_gate_88);
  not g_19922 (not_new_n633__16284135979104490, new_n633_);
  and g_19923 (new_n1253_, new_n1908_, new_n1909_);
  not g_19924 (not_new_n9402__0, new_n9402_);
  not g_19925 (not_new_n3890_, new_n3890_);
  not g_19926 (not_new_n591__0, new_n591_);
  not g_19927 (not_new_n642__9, new_n642_);
  not g_19928 (not_new_n7975_, new_n7975_);
  not g_19929 (not_new_n5846_, new_n5846_);
  not g_19930 (new_n8829_, new_n1043_);
  not g_19931 (not_new_n639__70, new_n639_);
  not g_19932 (not_new_n1069__0, new_n1069_);
  or g_19933 (new_n2632_, not_new_n2509__70, not_pi205);
  not g_19934 (not_pi135_3, pi135);
  or g_19935 (new_n6146_, not_new_n6010_, not_new_n5889_);
  or g_19936 (new_n6508_, not_new_n6509_, not_new_n639__403536070);
  or g_19937 (new_n3705_, not_new_n622__9, not_po298_47475615099430);
  not g_19938 (not_new_n3805_, new_n3805_);
  not g_19939 (not_new_n628__9, new_n628_);
  not g_19940 (not_new_n1564_, new_n1564_);
  and g_19941 (and_new_n6417__new_n6418_, new_n6418_, new_n6417_);
  not g_19942 (not_new_n1596__1915812313805664144010, new_n1596_);
  not g_19943 (not_new_n1613__6782230728490, new_n1613_);
  or g_19944 (new_n7038_, not_new_n7435_, not_new_n7434_);
  not g_19945 (not_new_n5555_, new_n5555_);
  not g_19946 (not_new_n1567_, new_n1567_);
  not g_19947 (not_new_n5519_, new_n5519_);
  or g_19948 (new_n8297_, not_new_n8117_, not_new_n8296_);
  not g_19949 (new_n6072_, new_n5906_);
  not g_19950 (not_new_n1538__24010, new_n1538_);
  or g_19951 (new_n10223_, not_new_n9856_, not_new_n9900_);
  or g_19952 (new_n2090_, not_new_n2085_, not_new_n1292_);
  or g_19953 (new_n9800_, not_new_n9407__0, not_new_n639__797922662976120010);
  not g_19954 (new_n5764_, new_n1596_);
  or g_19955 (new_n4042_, not_pi048_4, not_new_n4015_);
  or g_19956 (or_not_new_n7316__not_new_n7186_, not_new_n7316_, not_new_n7186_);
  not g_19957 (not_new_n638__0, new_n638_);
  or g_19958 (new_n8271_, not_new_n8344_, or_not_new_n8448__not_new_n8419_);
  not g_19959 (not_new_n5724_, new_n5724_);
  or g_19960 (new_n7480_, not_new_n721__0, not_new_n7457__0);
  not g_19961 (not_new_n1611__490, new_n1611_);
  not g_19962 (not_new_n9876_, new_n9876_);
  not g_19963 (not_new_n5477__0, new_n5477_);
  or g_19964 (new_n8060_, not_new_n7646__0, not_new_n644__968890104070);
  not g_19965 (not_new_n4835__1, new_n4835_);
  not g_19966 (not_new_n598__2, new_n598_);
  not g_19967 (not_new_n989__8, new_n989_);
  or g_19968 (new_n1704_, not_pi008_0, not_po296_968890104070);
  not g_19969 (not_new_n754_, new_n754_);
  and g_19970 (new_n7110_, new_n7370_, new_n7369_);
  not g_19971 (not_pi165_1, pi165);
  or g_19972 (new_n8525_, not_new_n8134__2, not_new_n1601__2326305139872070);
  not g_19973 (not_new_n3672_, new_n3672_);
  not g_19974 (not_new_n4462__0, new_n4462_);
  not g_19975 (not_new_n1616__70, new_n1616_);
  or g_19976 (new_n7313_, not_new_n7070_, not_new_n7315_);
  not g_19977 (new_n8449_, new_n8271_);
  not g_19978 (not_pi176_0, pi176);
  not g_19979 (not_new_n1028__9, new_n1028_);
  not g_19980 (not_new_n9874_, new_n9874_);
  not g_19981 (not_new_n8322__0, new_n8322_);
  not g_19982 (not_new_n7735__2, new_n7735_);
  not g_19983 (new_n7135_, new_n746_);
  and g_19984 (new_n8686_, new_n1167_, new_n8628_);
  or g_19985 (new_n1832_, not_new_n1585__2, not_new_n5734_);
  not g_19986 (not_new_n613__3, new_n613_);
  not g_19987 (not_pi039_4, pi039);
  or g_19988 (new_n10260_, not_new_n628__657123623635342801395430, not_new_n9883_);
  or g_19989 (or_not_new_n9084__not_new_n9083_, not_new_n9084_, not_new_n9083_);
  not g_19990 (not_new_n5475__0, new_n5475_);
  not g_19991 (not_new_n2123_, new_n2123_);
  not g_19992 (not_new_n634__24010, new_n634_);
  not g_19993 (not_pi101_0, pi101);
  not g_19994 (not_new_n8629_, new_n8629_);
  or g_19995 (or_or_or_not_new_n2955__not_new_n2958__not_new_n2957__not_new_n2959_, or_or_not_new_n2955__not_new_n2958__not_new_n2957_, not_new_n2959_);
  or g_19996 (new_n5126_, not_new_n5091_, not_new_n4947_);
  or g_19997 (new_n2151_, not_new_n4126_, not_new_n585__2824752490);
  not g_19998 (not_new_n7139__1, new_n7139_);
  not g_19999 (not_new_n3315__4, new_n3315_);
  or g_20000 (new_n9046_, not_new_n626__1915812313805664144010, not_new_n1053__19773267430);
  or g_20001 (new_n6603_, not_new_n6917_, not_new_n6918_);
  not g_20002 (new_n5794_, new_n1053_);
  not g_20003 (not_new_n1031__168070, new_n1031_);
  or g_20004 (new_n4558_, new_n1016_, pi174);
  not g_20005 (not_new_n7564_, new_n7564_);
  not g_20006 (not_new_n5743_, new_n5743_);
  not g_20007 (not_new_n6476__0, new_n6476_);
  or g_20008 (new_n7593_, not_new_n7815_, not_new_n7812_);
  not g_20009 (not_new_n7699_, new_n7699_);
  not g_20010 (not_new_n1010__1, new_n1010_);
  or g_20011 (new_n8011_, not_new_n7747_, not_new_n7720_);
  or g_20012 (new_n7040_, not_new_n7443_, not_new_n7444_);
  and g_20013 (new_n1512_, new_n1513_, new_n3043_);
  not g_20014 (not_new_n728__1, new_n728_);
  not g_20015 (not_new_n1999_, new_n1999_);
  not g_20016 (not_new_n4097_, new_n4097_);
  not g_20017 (not_new_n9292_, new_n9292_);
  not g_20018 (not_new_n1808_, new_n1808_);
  not g_20019 (new_n8824_, new_n628_);
  not g_20020 (not_new_n1616__6, new_n1616_);
  not g_20021 (not_new_n607__10, new_n607_);
  not g_20022 (not_new_n4906_, new_n4906_);
  not g_20023 (not_new_n2876_, new_n2876_);
  not g_20024 (not_po296_0, po296);
  not g_20025 (not_po296_13410686196639649008070, po296);
  not g_20026 (not_new_n604__332329305696010, new_n604_);
  or g_20027 (new_n2407_, not_new_n603__10, not_new_n636__1);
  or g_20028 (new_n3505_, not_new_n1613__2824752490, not_new_n2185_);
  not g_20029 (not_new_n675_, new_n675_);
  not g_20030 (not_new_n922_, new_n922_);
  or g_20031 (new_n662_, not_new_n3147_, or_not_new_n3149__not_new_n3148_);
  not g_20032 (not_new_n7026_, new_n7026_);
  or g_20033 (new_n8562_, not_new_n8236_, not_new_n8268_);
  not g_20034 (not_new_n9084_, new_n9084_);
  not g_20035 (not_new_n6644__0, new_n6644_);
  or g_20036 (new_n1679_, not_pi048, not_new_n1631__24010);
  not g_20037 (not_new_n2748_, new_n2748_);
  not g_20038 (not_new_n621__8235430, new_n621_);
  or g_20039 (new_n1661_, not_pi042, not_new_n1631__8);
  and g_20040 (new_n3973_, not_pi054_2, not_pi053_2);
  and g_20041 (new_n5051_, new_n4903_, new_n5236_);
  and g_20042 (and_new_n6375__new_n6382_, new_n6382_, new_n6375_);
  not g_20043 (not_new_n4162_, new_n4162_);
  and g_20044 (new_n1206_, new_n1709_, new_n1707_);
  or g_20045 (new_n927_, not_new_n3376_, or_not_new_n999__1_not_new_n3377_);
  or g_20046 (or_not_new_n2567__not_new_n2571_, not_new_n2571_, not_new_n2567_);
  not g_20047 (not_new_n7497_, new_n7497_);
  or g_20048 (new_n5141_, not_new_n632__24010, not_new_n1037__9);
  or g_20049 (new_n9159_, not_new_n8984__0, not_new_n9116_);
  or g_20050 (new_n4604_, not_new_n4428__0, not_pi168_3);
  and g_20051 (and_new_n1542__new_n2371_, new_n1542_, new_n2371_);
  not g_20052 (not_new_n9661_, new_n9661_);
  not g_20053 (not_new_n1192_, new_n1192_);
  not g_20054 (not_pi249_2, pi249);
  and g_20055 (new_n8976_, new_n9303_, new_n9304_);
  not g_20056 (not_new_n1047__47475615099430, new_n1047_);
  or g_20057 (new_n2908_, not_new_n994__19773267430, not_new_n4114__1);
  not g_20058 (not_new_n4090_, new_n4090_);
  not g_20059 (not_pi057_1, pi057);
  not g_20060 (not_new_n4435__0, new_n4435_);
  not g_20061 (not_new_n6509__0, new_n6509_);
  or g_20062 (or_or_not_new_n2820__not_new_n2823__not_new_n2822_, not_new_n2822_, or_not_new_n2820__not_new_n2823_);
  or g_20063 (new_n9147_, new_n1057_, new_n636_);
  or g_20064 (or_not_new_n2973__not_new_n2976_, not_new_n2976_, not_new_n2973_);
  not g_20065 (not_new_n7170__0, new_n7170_);
  not g_20066 (not_pi052, pi052);
  not g_20067 (not_new_n6033_, new_n6033_);
  not g_20068 (not_new_n631__39098210485829880490, new_n631_);
  not g_20069 (new_n4446_, new_n1013_);
  not g_20070 (not_new_n8009_, new_n8009_);
  not g_20071 (not_new_n4276_, new_n4276_);
  or g_20072 (new_n6202_, not_new_n5800__0, not_new_n1061__24010);
  not g_20073 (not_new_n9065_, new_n9065_);
  not g_20074 (not_new_n609__24010, new_n609_);
  not g_20075 (not_new_n8595__4, new_n8595_);
  not g_20076 (not_new_n9513_, new_n9513_);
  and g_20077 (new_n8807_, new_n9056_, new_n8802_);
  or g_20078 (new_n1872_, not_new_n8192_, not_new_n1581__4);
  not g_20079 (new_n5280_, new_n4995_);
  not g_20080 (not_new_n9714_, new_n9714_);
  not g_20081 (not_new_n596__24010, key_gate_88);
  not g_20082 (not_new_n6659_, new_n6659_);
  not g_20083 (not_new_n627__168070, new_n627_);
  not g_20084 (new_n6803_, new_n6631_);
  and g_20085 (new_n8685_, new_n1171_, new_n8626_);
  not g_20086 (not_new_n581__490, new_n581_);
  not g_20087 (not_new_n3436_, new_n3436_);
  or g_20088 (new_n5407_, not_new_n5406_, not_new_n5405_);
  or g_20089 (new_n5080_, not_new_n5063_, not_new_n618__490);
  not g_20090 (not_new_n8632_, new_n8632_);
  or g_20091 (new_n3573_, not_new_n2223__0, not_new_n1612__138412872010);
  not g_20092 (not_new_n1603__5, new_n1603_);
  not g_20093 (not_new_n5304_, new_n5304_);
  not g_20094 (not_new_n4136__0, new_n4136_);
  or g_20095 (new_n6435_, not_new_n1602__3430, not_new_n6259_);
  not g_20096 (not_new_n6331_, new_n6331_);
  or g_20097 (new_n7509_, not_new_n6985__1, not_new_n7026__1);
  not g_20098 (not_new_n4271_, new_n4271_);
  not g_20099 (not_new_n7409__0, new_n7409_);
  not g_20100 (not_new_n1728__403536070, new_n1728_);
  and g_20101 (new_n1454_, and_new_n2687__new_n2688_, new_n2689_);
  not g_20102 (not_new_n6950_, new_n6950_);
  not g_20103 (not_new_n2166__0, new_n2166_);
  not g_20104 (new_n8436_, new_n8258_);
  and g_20105 (new_n4489_, new_n4647_, new_n4646_);
  not g_20106 (not_new_n5457_, new_n5457_);
  not g_20107 (not_new_n10324_, new_n10324_);
  not g_20108 (not_new_n10173_, new_n10173_);
  not g_20109 (not_new_n2732_, new_n2732_);
  and g_20110 (new_n8202_, new_n8297_, new_n8298_);
  or g_20111 (new_n4641_, not_new_n4487__0, not_new_n4486_);
  not g_20112 (not_new_n5626_, new_n5626_);
  or g_20113 (new_n5290_, not_new_n4951_, not_new_n5084__1);
  not g_20114 (not_new_n9821_, new_n9821_);
  not g_20115 (new_n6659_, new_n6490_);
  not g_20116 (not_new_n628__5585458640832840070, new_n628_);
  not g_20117 (not_new_n7449_, new_n7449_);
  or g_20118 (new_n9973_, not_new_n3893_, not_new_n3892_);
  not g_20119 (not_new_n1600__2, new_n1600_);
  or g_20120 (new_n7468_, not_new_n718__2, not_new_n7406__2);
  or g_20121 (new_n8191_, not_new_n8471_, not_new_n8470_);
  not g_20122 (new_n4429_, pi169);
  not g_20123 (not_new_n8104__1, new_n8104_);
  or g_20124 (new_n9041_, not_new_n632__332329305696010, not_new_n1037__138412872010);
  not g_20125 (not_new_n6375_, new_n6375_);
  not g_20126 (not_pi007_0, pi007);
  not g_20127 (not_new_n1774_, new_n1774_);
  not g_20128 (not_new_n2075_, new_n2075_);
  not g_20129 (not_new_n638__1176490, new_n638_);
  or g_20130 (new_n3281_, not_new_n589__26517308458596534717790233816010, not_new_n1069__5);
  not g_20131 (new_n7942_, new_n7739_);
  not g_20132 (not_new_n10073__0, new_n10073_);
  or g_20133 (or_not_new_n4839__not_new_n4767_, not_new_n4839_, not_new_n4767_);
  not g_20134 (not_po296_35561530251773635572553173835655155124070416738520070, po296);
  or g_20135 (new_n2394_, not_new_n599__7, not_new_n9956__0);
  or g_20136 (new_n3955_, not_new_n3975_, not_new_n4004_);
  or g_20137 (new_n3433_, not_new_n1594__5, not_new_n1005__1);
  or g_20138 (new_n8909_, not_new_n9236_, not_new_n9235_);
  not g_20139 (not_new_n597__4, new_n597_);
  not g_20140 (not_new_n4638_, new_n4638_);
  or g_20141 (new_n3223_, not_new_n646__7, not_new_n589__8235430);
  not g_20142 (not_new_n1781_, new_n1781_);
  not g_20143 (not_new_n628__16284135979104490, new_n628_);
  not g_20144 (not_new_n1957_, new_n1957_);
  not g_20145 (not_new_n1200_, new_n1200_);
  not g_20146 (not_new_n7002_, new_n7002_);
  not g_20147 (not_new_n7433__1, new_n7433_);
  not g_20148 (not_new_n9050_, new_n9050_);
  not g_20149 (not_new_n7103_, new_n7103_);
  not g_20150 (not_new_n8959_, new_n8959_);
  not g_20151 (new_n1604_, new_n963_);
  not g_20152 (not_new_n4456__0, new_n4456_);
  or g_20153 (new_n8304_, not_new_n8120_, not_new_n1041__8235430);
  or g_20154 (new_n9501_, not_new_n9698_, not_new_n9601_);
  not g_20155 (not_new_n597__57648010, new_n597_);
  or g_20156 (new_n3296_, not_new_n3184__6782230728490, not_new_n627__8);
  not g_20157 (not_new_n1537__16284135979104490, new_n1537_);
  not g_20158 (not_new_n7089_, new_n7089_);
  not g_20159 (not_new_n5754__2, new_n5754_);
  not g_20160 (not_new_n2830_, new_n2830_);
  not g_20161 (not_new_n3918__0, new_n3918_);
  or g_20162 (new_n3866_, not_new_n1576__57648010, not_new_n632__490);
  not g_20163 (not_new_n639__6782230728490, new_n639_);
  or g_20164 (new_n2195_, not_new_n1581__19773267430, not_new_n8196_);
  not g_20165 (not_new_n1153__0, new_n1153_);
  not g_20166 (not_new_n7155__1, new_n7155_);
  and g_20167 (new_n9982_, new_n10072_, new_n10070_);
  or g_20168 (new_n2147_, not_new_n2142_, not_new_n1304_);
  or g_20169 (new_n4379_, not_new_n690_, not_new_n4268_);
  or g_20170 (new_n7730_, not_new_n8060_, not_new_n8059_);
  not g_20171 (not_new_n1039__2, new_n1039_);
  or g_20172 (new_n945_, or_or_not_new_n1235__not_new_n1233__not_new_n1812_, not_new_n1811_);
  or g_20173 (new_n6405_, not_new_n714_, not_new_n1031__24010);
  or g_20174 (new_n3570_, not_new_n1538__19773267430, not_pi151_0);
  and g_20175 (new_n5714_, new_n5915_, new_n5968_);
  or g_20176 (new_n5233_, not_new_n4999__0, not_new_n5232_);
  or g_20177 (new_n7310_, not_new_n7023_, not_new_n741_);
  not g_20178 (not_new_n1585__6782230728490, new_n1585_);
  not g_20179 (not_new_n3529_, new_n3529_);
  not g_20180 (not_new_n3986__0, new_n3986_);
  not g_20181 (not_new_n9942_, new_n9942_);
  not g_20182 (not_new_n1047__3430, new_n1047_);
  or g_20183 (po154, not_new_n3534_, not_new_n3535_);
  or g_20184 (new_n6170_, not_new_n5777__0, not_new_n1604__490);
  not g_20185 (not_new_n3378_, new_n3378_);
  not g_20186 (not_new_n8108__0, new_n8108_);
  not g_20187 (not_new_n9408__0, new_n9408_);
  buf g_20188 (po042, pi222);
  not g_20189 (not_pi055_2, pi055);
  not g_20190 (not_new_n8163_, new_n8163_);
  not g_20191 (not_new_n2319_, new_n2319_);
  not g_20192 (new_n6978_, new_n738_);
  not g_20193 (not_new_n1580__8235430, new_n1580_);
  not g_20194 (not_new_n7447_, new_n7447_);
  not g_20195 (not_new_n1061__16284135979104490, new_n1061_);
  or g_20196 (new_n9639_, not_new_n9422_, not_new_n9638_);
  not g_20197 (not_new_n1594__4, new_n1594_);
  or g_20198 (new_n6901_, not_new_n6629_, not_new_n6758_);
  not g_20199 (not_new_n4755_, new_n4755_);
  not g_20200 (not_new_n8413_, new_n8413_);
  not g_20201 (not_new_n599__968890104070, new_n599_);
  not g_20202 (not_new_n5300_, new_n5300_);
  not g_20203 (not_new_n8422_, new_n8422_);
  or g_20204 (new_n4403_, not_new_n4284_, not_new_n682_);
  not g_20205 (new_n6245_, new_n621_);
  not g_20206 (not_new_n3097_, new_n3097_);
  not g_20207 (not_new_n6325_, new_n6325_);
  not g_20208 (not_pi122, pi122);
  or g_20209 (new_n1029_, not_new_n3389_, not_new_n3388_);
  not g_20210 (not_new_n1538__0, new_n1538_);
  or g_20211 (new_n7464_, not_new_n7263_, or_not_new_n7463__not_new_n7312_);
  not g_20212 (not_new_n4839_, new_n4839_);
  not g_20213 (not_new_n5006_, new_n5006_);
  not g_20214 (not_new_n646__24010, new_n646_);
  or g_20215 (or_not_new_n6782__not_new_n6621_, not_new_n6782_, not_new_n6621_);
  not g_20216 (not_pi254, pi254);
  not g_20217 (new_n7406_, new_n7045_);
  not g_20218 (new_n10043_, new_n10022_);
  or g_20219 (new_n3468_, not_new_n1594__490, not_new_n1016__1);
  or g_20220 (new_n9915_, not_new_n637__16284135979104490, not_new_n1065__5585458640832840070);
  or g_20221 (new_n3712_, not_pi242, not_new_n989__16284135979104490);
  not g_20222 (not_new_n9417_, new_n9417_);
  not g_20223 (not_new_n1019__5, new_n1019_);
  not g_20224 (not_new_n635__5, new_n635_);
  not g_20225 (not_new_n595__2326305139872070, new_n595_);
  not g_20226 (new_n4577_, new_n4451_);
  not g_20227 (new_n8636_, new_n1149_);
  not g_20228 (new_n9509_, new_n9356_);
  not g_20229 (not_new_n1611__19773267430, new_n1611_);
  or g_20230 (new_n5144_, new_n626_, new_n1053_);
  not g_20231 (not_new_n5742__0, new_n5742_);
  not g_20232 (not_new_n1790_, new_n1790_);
  not g_20233 (not_new_n7534_, new_n7534_);
  not g_20234 (not_new_n3938_, new_n3938_);
  or g_20235 (new_n3412_, not_new_n1536__168070, not_pi030_0);
  not g_20236 (not_new_n735_, new_n735_);
  not g_20237 (not_new_n1376_, new_n1376_);
  xnor g_20238 (key_gate_50, new_n1181_, key_50);
  or g_20239 (new_n1673_, not_new_n1631__490, not_pi046);
  or g_20240 (or_not_new_n1554__not_new_n2429_, not_new_n1554_, not_new_n2429_);
  or g_20241 (new_n4670_, not_pi177_3, not_new_n4446__0);
  not g_20242 (not_new_n10018_, new_n10018_);
  not g_20243 (not_new_n642__403536070, new_n642_);
  or g_20244 (new_n9134_, not_new_n8950_, not_new_n9133_);
  not g_20245 (not_pi091, pi091);
  not g_20246 (not_new_n6185_, new_n6185_);
  or g_20247 (new_n1041_, not_new_n3422_, not_new_n3423_);
  or g_20248 (new_n2006_, not_new_n6558_, not_new_n1580__490);
  or g_20249 (new_n6048_, not_new_n6047_, not_new_n5977_);
  not g_20250 (not_new_n618__968890104070, new_n618_);
  not g_20251 (not_new_n1031__9, new_n1031_);
  or g_20252 (new_n937_, or_not_new_n1024__0_not_new_n3384__2, not_new_n3387__0);
  not g_20253 (not_new_n7405_, new_n7405_);
  not g_20254 (not_new_n1611__3, new_n1611_);
  or g_20255 (new_n5636_, not_new_n5434_, not_pi131_2);
  not g_20256 (not_new_n8688_, new_n8688_);
  not g_20257 (not_new_n9833_, new_n9833_);
  not g_20258 (not_new_n633__57648010, new_n633_);
  not g_20259 (not_new_n759_, new_n759_);
  not g_20260 (not_new_n5405_, new_n5405_);
  not g_20261 (new_n8108_, new_n1041_);
  not g_20262 (not_new_n4190_, new_n4190_);
  not g_20263 (not_new_n6977__1, new_n6977_);
  or g_20264 (new_n2049_, not_new_n593__3430, not_new_n638_);
  or g_20265 (new_n2321_, not_new_n588__113988951853731430, not_pi127);
  or g_20266 (new_n6207_, not_new_n5789__0, not_new_n644__57648010);
  not g_20267 (not_new_n4422__0, new_n4422_);
  not g_20268 (not_new_n1319_, new_n1319_);
  not g_20269 (not_new_n638__3430, new_n638_);
  not g_20270 (not_new_n5438__0, new_n5438_);
  not g_20271 (not_new_n3172_, new_n3172_);
  or g_20272 (new_n9972_, not_new_n3897_, not_new_n3898_);
  not g_20273 (not_new_n5915_, new_n5915_);
  or g_20274 (new_n3788_, not_new_n1063__6, not_new_n638__10);
  not g_20275 (new_n6293_, new_n1065_);
  not g_20276 (not_new_n8368__1, new_n8368_);
  or g_20277 (new_n1659_, not_po296_8, not_pi023);
  not g_20278 (not_new_n1043__2326305139872070, new_n1043_);
  or g_20279 (new_n8169_, not_new_n621__968890104070, not_new_n8128_);
  not g_20280 (not_new_n581__367033682172941254412302110320336601888010, new_n581_);
  not g_20281 (not_new_n9313_, new_n9313_);
  not g_20282 (not_new_n5717_, new_n5717_);
  not g_20283 (not_new_n10293_, new_n10293_);
  or g_20284 (new_n4179_, not_new_n4077_, not_pi266_2);
  not g_20285 (not_new_n1944_, new_n1944_);
  not g_20286 (not_new_n3742_, new_n3742_);
  not g_20287 (not_new_n589__541169560379521116689596608490, new_n589_);
  not g_20288 (not_new_n723_, new_n723_);
  or g_20289 (new_n6198_, not_new_n5799__0, not_new_n1063__490);
  not g_20290 (not_new_n1035__5, new_n1035_);
  not g_20291 (not_new_n8917_, new_n8917_);
  or g_20292 (or_not_new_n6239__not_new_n6350_, not_new_n6350_, not_new_n6239_);
  not g_20293 (not_new_n1612__57648010, new_n1612_);
  not g_20294 (not_new_n1602__1176490, new_n1602_);
  not g_20295 (not_new_n3237_, new_n3237_);
  not g_20296 (new_n6661_, new_n6634_);
  not g_20297 (not_new_n4230_, new_n4230_);
  or g_20298 (or_not_new_n3140__not_new_n3139_, not_new_n3140_, not_new_n3139_);
  or g_20299 (new_n2541_, not_new_n606__2, not_new_n5486__0);
  or g_20300 (new_n6913_, not_new_n6633__1, not_new_n642__403536070);
  not g_20301 (new_n5463_, new_n1015_);
  or g_20302 (or_not_new_n934__not_new_n933__0, not_new_n933__0, not_new_n934_);
  or g_20303 (new_n944_, not_new_n1792_, or_or_not_new_n1231__not_new_n1229__not_new_n1793_);
  not g_20304 (not_new_n7931_, new_n7931_);
  not g_20305 (not_new_n4121__1, new_n4121_);
  or g_20306 (new_n3656_, not_new_n989__0, not_pi214);
  or g_20307 (or_not_new_n1562__not_new_n2469_, not_new_n1562_, not_new_n2469_);
  and g_20308 (new_n1307_, new_n2159_, and_new_n1306__new_n2160_);
  or g_20309 (new_n4223_, not_pi251_1, not_new_n4152_);
  not g_20310 (not_new_n5817_, new_n5817_);
  not g_20311 (not_new_n8869__0, new_n8869_);
  and g_20312 (new_n600_, new_n1587_, new_n1611_);
  and g_20313 (new_n5035_, new_n4906_, new_n4900_);
  not g_20314 (not_pi099, pi099);
  not g_20315 (not_new_n619__9, new_n619_);
  not g_20316 (not_new_n7097_, new_n7097_);
  not g_20317 (not_new_n8635_, new_n8635_);
  not g_20318 (not_new_n3573_, new_n3573_);
  or g_20319 (new_n5734_, not_new_n6078_, not_new_n5966_);
  or g_20320 (new_n1023_, not_new_n3371_, not_new_n3370_);
  and g_20321 (new_n1357_, and_new_n2379__new_n2378_, new_n2377_);
  not g_20322 (not_new_n8286_, new_n8286_);
  not g_20323 (new_n7912_, new_n7654_);
  not g_20324 (not_new_n1556_, new_n1556_);
  not g_20325 (not_new_n1063__6, new_n1063_);
  or g_20326 (new_n3411_, not_new_n1805_, not_new_n1613__0);
  or g_20327 (new_n7361_, not_new_n7107_, not_new_n775__8);
  not g_20328 (not_new_n8400_, new_n8400_);
  not g_20329 (new_n3419_, new_n1039_);
  not g_20330 (not_new_n8625_, new_n8625_);
  not g_20331 (new_n9637_, new_n9422_);
  not g_20332 (not_new_n6603_, new_n6603_);
  not g_20333 (not_new_n6479__1, new_n6479_);
  and g_20334 (new_n1565_, new_n3642_, new_n3643_);
  not g_20335 (not_new_n5494_, new_n5494_);
  and g_20336 (new_n1554_, new_n3620_, new_n3621_);
  not g_20337 (not_new_n1599__2824752490, new_n1599_);
  or g_20338 (new_n9206_, not_new_n9204_, not_new_n9205_);
  not g_20339 (not_new_n3318_, new_n3318_);
  not g_20340 (not_new_n684_, new_n684_);
  not g_20341 (not_new_n589__403536070, new_n589_);
  not g_20342 (not_new_n4770_, new_n4770_);
  or g_20343 (new_n3457_, not_pi021_0, not_new_n1536__6782230728490);
  not g_20344 (not_new_n6538__0, new_n6538_);
  not g_20345 (not_new_n1585__8, new_n1585_);
  not g_20346 (not_new_n4698_, new_n4698_);
  or g_20347 (new_n1999_, not_new_n585__490, not_new_n4134_);
  and g_20348 (new_n6339_, and_new_n6373__new_n6386_, new_n6262_);
  not g_20349 (not_new_n622__968890104070, new_n622_);
  not g_20350 (not_new_n635__2, new_n635_);
  or g_20351 (new_n6689_, not_new_n6473__1, not_new_n6656__0);
  not g_20352 (not_new_n640__490, new_n640_);
  not g_20353 (not_new_n3185__1, new_n3185_);
  or g_20354 (new_n7416_, not_new_n7120_, not_new_n775__24010);
  or g_20355 (new_n4047_, not_new_n3954_, not_pi043_3);
  and g_20356 (new_n1284_, and_and_new_n2048__new_n2051__new_n2049_, new_n2050_);
  or g_20357 (new_n10201_, not_new_n10080_, not_new_n9888__1);
  not g_20358 (not_new_n5496__0, new_n5496_);
  not g_20359 (not_new_n1067__2, new_n1067_);
  and g_20360 (new_n6228_, new_n6398_, new_n6399_);
  not g_20361 (not_new_n5593_, new_n5593_);
  not g_20362 (not_new_n7452_, new_n7452_);
  not g_20363 (not_po296_1, po296);
  not g_20364 (not_new_n4735_, new_n4735_);
  not g_20365 (not_new_n5694_, new_n5694_);
  or g_20366 (new_n8174_, not_new_n8424_, not_new_n8370_);
  or g_20367 (new_n651_, or_not_new_n3113__not_new_n3112_, not_new_n3111_);
  not g_20368 (not_new_n5891_, new_n5891_);
  not g_20369 (not_new_n7722_, new_n7722_);
  not g_20370 (not_new_n646__138412872010, new_n646_);
  or g_20371 (new_n2966_, not_new_n1616__6782230728490, not_new_n2963_);
  not g_20372 (not_new_n973_, new_n973_);
  or g_20373 (new_n1935_, not_new_n593__7, not_new_n647_);
  not g_20374 (not_new_n3670_, new_n3670_);
  or g_20375 (new_n9585_, new_n644_, new_n1059_);
  not g_20376 (not_new_n8937_, new_n8937_);
  not g_20377 (not_new_n594__7, new_n594_);
  or g_20378 (new_n7166_, not_new_n7027_, not_new_n7165_);
  or g_20379 (new_n1754_, not_new_n1728__138412872010, not_pi068);
  not g_20380 (not_new_n7753__0, new_n7753_);
  not g_20381 (not_new_n8553_, new_n8553_);
  not g_20382 (new_n8456_, new_n8266_);
  not g_20383 (not_new_n7041_, new_n7041_);
  or g_20384 (new_n7534_, not_new_n7424__1, not_new_n730__1);
  not g_20385 (not_new_n2890_, new_n2890_);
  not g_20386 (not_new_n9940_, new_n9940_);
  or g_20387 (new_n7184_, not_new_n6978__0, not_new_n6977_);
  not g_20388 (not_new_n3372__113988951853731430, new_n3372_);
  or g_20389 (new_n7049_, not_new_n7374_, not_new_n7375_);
  not g_20390 (not_new_n9958__0, new_n9958_);
  and g_20391 (new_n1381_, new_n2437_, new_n2438_);
  and g_20392 (new_n7697_, new_n7578_, new_n7577_);
  or g_20393 (new_n9890_, not_new_n1035__1176490, not_new_n642__16284135979104490);
  or g_20394 (new_n8235_, not_new_n8554_, not_new_n8553_);
  not g_20395 (not_new_n4214_, new_n4214_);
  or g_20396 (new_n4148_, not_new_n4174_, not_pi273_0);
  not g_20397 (not_new_n9742_, new_n9742_);
  or g_20398 (new_n6140_, not_new_n617__57648010, not_new_n5807__1);
  not g_20399 (not_new_n10032__0, new_n10032_);
  or g_20400 (new_n10066_, new_n1045_, new_n635_);
  not g_20401 (not_new_n2851_, new_n2851_);
  not g_20402 (not_new_n9566_, new_n9566_);
  not g_20403 (not_new_n7345__1, new_n7345_);
  or g_20404 (new_n6124_, not_new_n1607__7, not_new_n5885_);
  not g_20405 (not_new_n4134__0, new_n4134_);
  not g_20406 (not_new_n10017_, new_n10017_);
  not g_20407 (new_n9597_, new_n9412_);
  not g_20408 (not_new_n9957__0, new_n9957_);
  or g_20409 (new_n5188_, not_new_n5185_, not_new_n5187_);
  not g_20410 (not_new_n620__0, new_n620_);
  not g_20411 (not_new_n9345_, new_n9345_);
  not g_20412 (not_new_n4566_, new_n4566_);
  or g_20413 (new_n8038_, not_new_n1069__8235430, not_new_n7639__0);
  not g_20414 (not_new_n3446_, new_n3446_);
  or g_20415 (new_n9615_, new_n1603_, new_n639_);
  not g_20416 (not_new_n9880_, new_n9880_);
  and g_20417 (new_n8238_, new_n8282_, new_n8565_);
  not g_20418 (new_n4777_, new_n1602_);
  not g_20419 (not_pi194, pi194);
  and g_20420 (new_n8089_, new_n8359_, new_n8361_);
  not g_20421 (not_new_n5148_, new_n5148_);
  not g_20422 (not_new_n1702_, key_gate_24);
  not g_20423 (not_new_n610__3430, new_n610_);
  or g_20424 (new_n9959_, not_new_n10264_, not_new_n10263_);
  not g_20425 (not_new_n1599__490, new_n1599_);
  not g_20426 (not_new_n3814_, new_n3814_);
  not g_20427 (not_new_n1049__332329305696010, new_n1049_);
  not g_20428 (not_new_n3834_, new_n3834_);
  and g_20429 (new_n1372_, new_n2416_, new_n2415_);
  not g_20430 (not_new_n1039__6782230728490, new_n1039_);
  not g_20431 (not_new_n639__8235430, new_n639_);
  and g_20432 (new_n8231_, and_new_n8082__new_n8430_, new_n8387_);
  not g_20433 (not_new_n591__57648010, new_n591_);
  and g_20434 (new_n3975_, not_pi043_2, not_pi044_2);
  not g_20435 (not_new_n2286_, new_n2286_);
  or g_20436 (new_n5916_, not_new_n1063__70, not_new_n5799_);
  not g_20437 (new_n5760_, new_n647_);
  not g_20438 (not_new_n10216_, new_n10216_);
  or g_20439 (new_n8248_, not_new_n8202_, not_new_n8450_);
  or g_20440 (new_n7874_, not_new_n7771__0, not_new_n7662__1);
  or g_20441 (new_n6959_, not_new_n6643_, not_new_n6812__0);
  or g_20442 (new_n9616_, not_new_n9615_, not_new_n9613_);
  not g_20443 (not_new_n10205_, new_n10205_);
  or g_20444 (new_n9950_, not_new_n10164_, not_new_n9909_);
  not g_20445 (not_new_n3511_, new_n3511_);
  not g_20446 (not_pi060_2, pi060);
  not g_20447 (not_new_n1027__16284135979104490, new_n1027_);
  or g_20448 (new_n8337_, not_new_n8291_, not_new_n8077_);
  or g_20449 (new_n8476_, not_new_n631__5585458640832840070, not_new_n8106__2);
  not g_20450 (not_new_n1264_, new_n1264_);
  not g_20451 (not_new_n9708_, new_n9708_);
  or g_20452 (po271, not_new_n2768_, or_not_new_n2769__not_new_n1476_);
  or g_20453 (new_n4378_, not_new_n4309_, not_new_n4375_);
  and g_20454 (new_n9873_, new_n10087_, new_n10084_);
  not g_20455 (not_new_n9694_, new_n9694_);
  not g_20456 (not_new_n2963_, new_n2963_);
  or g_20457 (new_n2346_, not_new_n4756_, not_new_n591__5585458640832840070);
  not g_20458 (not_new_n8841_, new_n8841_);
  not g_20459 (not_new_n9333_, new_n9333_);
  not g_20460 (not_new_n634__1176490, new_n634_);
  not g_20461 (not_new_n3919_, new_n3919_);
  not g_20462 (not_new_n9195_, new_n9195_);
  not g_20463 (not_pi041, pi041);
  or g_20464 (new_n4108_, not_new_n4172_, not_pi262_0);
  not g_20465 (not_new_n1613__4, new_n1613_);
  and g_20466 (and_new_n2414__new_n2413_, new_n2413_, new_n2414_);
  not g_20467 (new_n5160_, new_n5077_);
  not g_20468 (not_new_n642__8, new_n642_);
  or g_20469 (new_n3437_, not_new_n1536__2824752490, not_pi025_0);
  or g_20470 (new_n770_, not_new_n3196_, not_new_n3197_);
  or g_20471 (or_or_not_new_n1335__not_new_n1333__not_new_n2287_, or_not_new_n1335__not_new_n1333_, not_new_n2287_);
  or g_20472 (new_n2749_, not_new_n3311__0, not_new_n1045__1);
  not g_20473 (not_new_n4201_, new_n4201_);
  not g_20474 (new_n4443_, pi176);
  not g_20475 (not_new_n1355_, new_n1355_);
  not g_20476 (not_new_n5816_, new_n5816_);
  or g_20477 (new_n4999_, or_not_new_n5276__not_new_n5277_, not_new_n5165_);
  not g_20478 (not_new_n627__1, new_n627_);
  and g_20479 (new_n3979_, new_n4051_, new_n4052_);
  not g_20480 (not_new_n5431__0, new_n5431_);
  not g_20481 (not_new_n8959__0, new_n8959_);
  not g_20482 (not_new_n3757_, new_n3757_);
  not g_20483 (not_new_n3443_, new_n3443_);
  or g_20484 (new_n1733_, not_pi077, not_new_n1728__1);
  not g_20485 (not_new_n1051__168070, new_n1051_);
  not g_20486 (not_new_n593__403536070, new_n593_);
  not g_20487 (not_new_n1260_, new_n1260_);
  not g_20488 (new_n4176_, new_n4146_);
  not g_20489 (not_new_n5092_, new_n5092_);
  or g_20490 (new_n2059_, not_new_n1583__24010, not_new_n7692_);
  or g_20491 (new_n5187_, new_n1603_, new_n639_);
  not g_20492 (not_new_n1599__1176490, new_n1599_);
  not g_20493 (not_new_n1581__9, new_n1581_);
  not g_20494 (not_new_n638__273687473400809163430, new_n638_);
  not g_20495 (not_new_n1579_, new_n1579_);
  not g_20496 (not_new_n6762_, new_n6762_);
  not g_20497 (not_new_n627__6782230728490, new_n627_);
  or g_20498 (new_n932_, not_new_n1027__1, not_new_n1024_);
  not g_20499 (not_new_n6979__1, new_n6979_);
  or g_20500 (new_n2223_, not_new_n2218_, not_new_n1320_);
  or g_20501 (new_n8559_, not_new_n8148__0, not_new_n633__968890104070);
  not g_20502 (not_new_n7553_, new_n7553_);
  not g_20503 (not_new_n9080_, new_n9080_);
  not g_20504 (not_new_n9744_, new_n9744_);
  not g_20505 (not_new_n4565_, new_n4565_);
  or g_20506 (new_n7684_, not_new_n7951_, not_new_n7950_);
  or g_20507 (new_n9255_, not_new_n9253_, not_new_n9096_);
  not g_20508 (not_new_n1599__3430, new_n1599_);
  or g_20509 (new_n4930_, not_new_n642__490, not_new_n1035__8);
  not g_20510 (not_new_n7053_, new_n7053_);
  not g_20511 (not_new_n1041__8235430, new_n1041_);
  not g_20512 (not_new_n3558_, new_n3558_);
  not g_20513 (not_new_n5045_, new_n5045_);
  not g_20514 (not_new_n6702_, new_n6702_);
  or g_20515 (new_n7333_, not_new_n6974_, not_new_n765_);
  not g_20516 (not_new_n9584__0, new_n9584_);
  not g_20517 (not_new_n4065_, new_n4065_);
  not g_20518 (new_n6502_, new_n1600_);
  or g_20519 (new_n1769_, not_new_n1583_, not_new_n7595_);
  and g_20520 (and_new_n6326__new_n6241_, new_n6326_, new_n6241_);
  not g_20521 (not_new_n2714_, new_n2714_);
  or g_20522 (new_n3312_, not_new_n3321_, not_new_n3318__0);
  not g_20523 (not_new_n3372__168070, new_n3372_);
  or g_20524 (new_n9948_, not_new_n10115_, not_new_n10116_);
  not g_20525 (not_new_n8039_, new_n8039_);
  not g_20526 (not_new_n6728_, new_n6728_);
  not g_20527 (new_n9922_, new_n1057_);
  not g_20528 (not_new_n7512_, new_n7512_);
  not g_20529 (not_new_n5009_, new_n5009_);
  or g_20530 (or_or_not_new_n1555__not_new_n2434__not_new_n1379_, or_not_new_n1555__not_new_n2434_, not_new_n1379_);
  not g_20531 (not_new_n3295_, new_n3295_);
  or g_20532 (new_n5182_, not_new_n5180_, not_new_n5181_);
  or g_20533 (new_n2264_, not_pi124, not_new_n588__332329305696010);
  or g_20534 (new_n5334_, not_new_n5333_, not_new_n5332_);
  or g_20535 (new_n5712_, not_pi129_3, not_new_n5429_);
  and g_20536 (new_n8270_, new_n8571_, new_n8570_);
  not g_20537 (new_n5472_, pi147);
  not g_20538 (not_new_n8472_, new_n8472_);
  or g_20539 (new_n6944_, not_new_n644__19773267430, not_new_n6522__0);
  not g_20540 (not_new_n6999_, new_n6999_);
  not g_20541 (not_new_n6297_, new_n6297_);
  and g_20542 (new_n5875_, new_n5715_, new_n6037_);
  or g_20543 (new_n2263_, not_pi156, not_new_n587__332329305696010);
  not g_20544 (not_new_n746_, new_n746_);
  or g_20545 (new_n5344_, not_new_n4951__0, not_new_n621__168070);
  or g_20546 (new_n2919_, not_new_n1596__1, not_new_n613__5);
  not g_20547 (not_new_n644__3430, new_n644_);
  not g_20548 (not_new_n637__8, new_n637_);
  not g_20549 (not_new_n9358_, new_n9358_);
  not g_20550 (not_new_n1976__0, new_n1976_);
  not g_20551 (not_new_n635__6, new_n635_);
  not g_20552 (not_new_n1561_, new_n1561_);
  not g_20553 (not_new_n7002__0, new_n7002_);
  not g_20554 (not_new_n2581_, new_n2581_);
  and g_20555 (new_n5512_, new_n5666_, new_n5667_);
  not g_20556 (not_new_n10105_, new_n10105_);
  not g_20557 (not_new_n6110_, new_n6110_);
  or g_20558 (new_n4524_, not_pi165_1, not_new_n1007__2);
  not g_20559 (not_new_n4116__1, new_n4116_);
  and g_20560 (new_n3972_, not_pi052_2, not_pi051_2);
  not g_20561 (not_new_n9947_, new_n9947_);
  xor g_20562 (key_gate_109, not_new_n1651_, key_109);
  or g_20563 (new_n5127_, not_new_n628__3430, not_new_n1039__8);
  not g_20564 (not_new_n7468_, new_n7468_);
  or g_20565 (new_n3431_, not_new_n1881_, not_new_n1613__4);
  or g_20566 (new_n5238_, new_n637_, new_n1065_);
  not g_20567 (not_new_n7879_, new_n7879_);
  or g_20568 (new_n6650_, not_new_n1053__24010, not_new_n6525_);
  not g_20569 (not_new_n2769_, new_n2769_);
  or g_20570 (new_n5106_, not_new_n4938_, not_new_n4937_);
  or g_20571 (new_n10281_, not_new_n617__93874803376477543056490, not_new_n9943_);
  not g_20572 (not_new_n6992__1, new_n6992_);
  not g_20573 (not_new_n597__168070, new_n597_);
  buf g_20574 (po035, pi229);
  or g_20575 (new_n8471_, not_new_n8308__0, not_new_n8245_);
  not g_20576 (not_new_n5682_, new_n5682_);
  or g_20577 (new_n2052_, not_new_n2047_, not_new_n1284_);
  or g_20578 (new_n4575_, not_new_n4494_, not_new_n4574_);
  or g_20579 (new_n7691_, not_new_n8022_, not_new_n8021_);
  not g_20580 (not_new_n588__6, new_n588_);
  not g_20581 (not_new_n5848_, new_n5848_);
  not g_20582 (not_new_n637__2824752490, new_n637_);
  not g_20583 (not_new_n7538_, new_n7538_);
  not g_20584 (not_new_n2880_, new_n2880_);
  not g_20585 (not_new_n7352_, new_n7352_);
  or g_20586 (new_n6877_, not_new_n617__138412872010, not_new_n6498__1);
  or g_20587 (new_n8744_, not_new_n1153__0, not_new_n8605_);
  and g_20588 (new_n6638_, new_n6936_, new_n6935_);
  not g_20589 (not_new_n5649_, new_n5649_);
  or g_20590 (new_n7137_, not_new_n7261_, not_new_n7260_);
  not g_20591 (not_new_n1057__24010, new_n1057_);
  not g_20592 (not_new_n7824_, new_n7824_);
  or g_20593 (new_n6764_, not_new_n6763_, not_new_n6607_);
  or g_20594 (new_n3054_, not_new_n1170_, not_new_n1027__6782230728490);
  not g_20595 (new_n9904_, new_n645_);
  or g_20596 (new_n4061_, not_new_n3989_, not_pi056_2);
  not g_20597 (not_new_n1538__6, new_n1538_);
  not g_20598 (new_n8425_, new_n8174_);
  not g_20599 (not_new_n7925_, new_n7925_);
  or g_20600 (po214, not_new_n1415_, not_new_n1413_);
  not g_20601 (not_new_n1069__5, new_n1069_);
  or g_20602 (new_n7686_, not_new_n7967_, not_new_n7966_);
  not g_20603 (not_new_n10024__0, new_n10024_);
  not g_20604 (not_pi152_0, pi152);
  not g_20605 (not_new_n3126_, new_n3126_);
  not g_20606 (not_new_n6373__3, new_n6373_);
  not g_20607 (not_new_n1941_, new_n1941_);
  or g_20608 (new_n1949_, not_new_n6559_, not_new_n1580__9);
  not g_20609 (not_new_n5641_, new_n5641_);
  or g_20610 (new_n10250_, not_new_n10248_, not_new_n10249_);
  and g_20611 (new_n1477_, new_n2771_, new_n2770_);
  or g_20612 (new_n3282_, not_new_n646__8, not_new_n3184__8235430);
  not g_20613 (not_new_n1602__4, new_n1602_);
  or g_20614 (new_n9592_, new_n1063_, new_n638_);
  or g_20615 (new_n6833_, not_new_n6479__0, not_new_n648__2824752490);
  or g_20616 (new_n5599_, not_new_n5597__0, not_new_n5598_);
  and g_20617 (new_n7575_, new_n7850_, new_n7770_);
  or g_20618 (new_n2631_, not_new_n606__70, not_new_n5478__0);
  not g_20619 (new_n9891_, new_n1031_);
  not g_20620 (not_pi161_1, pi161);
  not g_20621 (not_pi218, pi218);
  not g_20622 (not_pi019, pi019);
  not g_20623 (not_new_n8411_, new_n8411_);
  or g_20624 (new_n7878_, not_new_n7876_, not_new_n7877_);
  not g_20625 (not_new_n1611__3430, new_n1611_);
  not g_20626 (not_pi055, pi055);
  not g_20627 (not_new_n632__6, new_n632_);
  not g_20628 (not_new_n10136_, new_n10136_);
  not g_20629 (not_new_n6873_, new_n6873_);
  not g_20630 (not_new_n3538_, new_n3538_);
  not g_20631 (not_new_n7598__0, new_n7598_);
  not g_20632 (not_new_n2040_, new_n2040_);
  not g_20633 (not_new_n8154_, new_n8154_);
  not g_20634 (not_new_n6449_, new_n6449_);
  or g_20635 (new_n1009_, not_new_n3340_, not_new_n3339_);
  not g_20636 (new_n6950_, new_n6609_);
  not g_20637 (not_new_n8721_, new_n8721_);
  not g_20638 (not_new_n7043_, new_n7043_);
  or g_20639 (new_n8534_, not_new_n1603__403536070, not_new_n8136__0);
  not g_20640 (not_new_n2204_, new_n2204_);
  not g_20641 (new_n1589_, new_n938_);
  not g_20642 (not_new_n7153_, new_n7153_);
  not g_20643 (not_new_n1605__4, new_n1605_);
  not g_20644 (not_new_n1071_, new_n1071_);
  not g_20645 (not_new_n8248__0, new_n8248_);
  not g_20646 (not_new_n4113__2, new_n4113_);
  not g_20647 (not_new_n6131_, new_n6131_);
  not g_20648 (not_new_n8176_, new_n8176_);
  not g_20649 (not_new_n8085_, new_n8085_);
  not g_20650 (not_new_n6226_, new_n6226_);
  and g_20651 (new_n7112_, new_n7384_, new_n7383_);
  not g_20652 (not_new_n625__16284135979104490, new_n625_);
  not g_20653 (not_new_n4933__0, new_n4933_);
  not g_20654 (not_new_n1596__6, new_n1596_);
  or g_20655 (new_n6778_, not_new_n6650__0, not_new_n6777_);
  not g_20656 (not_new_n8205_, new_n8205_);
  not g_20657 (not_new_n2207_, new_n2207_);
  not g_20658 (not_new_n1309_, new_n1309_);
  or g_20659 (new_n5979_, not_new_n1065__10, not_new_n5798_);
  not g_20660 (not_new_n4114__1, new_n4114_);
  not g_20661 (not_new_n2792_, new_n2792_);
  or g_20662 (new_n6753_, not_new_n6538__0, not_new_n6653_);
  not g_20663 (not_new_n8188_, new_n8188_);
  not g_20664 (not_new_n627__70, new_n627_);
  not g_20665 (not_new_n593__8235430, new_n593_);
  not g_20666 (not_new_n5431__1, new_n5431_);
  not g_20667 (not_new_n6483__0, new_n6483_);
  not g_20668 (not_new_n6967_, new_n6967_);
  and g_20669 (new_n608_, new_n592_, new_n3366_);
  not g_20670 (not_new_n7155__0, new_n7155_);
  not g_20671 (new_n4112_, pi273);
  or g_20672 (new_n4326_, not_new_n4289_, not_new_n4288_);
  or g_20673 (new_n5329_, not_new_n5327_, not_new_n5207_);
  or g_20674 (new_n5181_, not_new_n4975_, not_new_n4974_);
  not g_20675 (new_n1582_, new_n935_);
  not g_20676 (not_new_n8366_, new_n8366_);
  not g_20677 (not_new_n7462_, new_n7462_);
  not g_20678 (not_new_n3405_, new_n3405_);
  or g_20679 (new_n4451_, not_new_n4576_, not_new_n4575_);
  and g_20680 (and_and_and_new_n6227__new_n6232__new_n6229__new_n6317_, new_n6317_, and_and_new_n6227__new_n6232__new_n6229_);
  not g_20681 (not_new_n8265__1, new_n8265_);
  not g_20682 (not_new_n9549_, new_n9549_);
  or g_20683 (new_n4027_, not_new_n3945_, not_pi059_2);
  or g_20684 (new_n6927_, not_new_n6516__0, not_new_n1067__24010);
  not g_20685 (not_new_n6649_, new_n6649_);
  not g_20686 (not_new_n4841_, new_n4841_);
  not g_20687 (not_new_n591_, new_n591_);
  or g_20688 (or_or_not_new_n2587__not_new_n2591__not_new_n1433_, or_not_new_n2587__not_new_n2591_, not_new_n1433_);
  not g_20689 (not_new_n3372__490, new_n3372_);
  not g_20690 (not_new_n3841_, new_n3841_);
  not g_20691 (not_new_n630__39098210485829880490, new_n630_);
  or g_20692 (new_n8572_, not_new_n8271__2, not_new_n8401_);
  not g_20693 (not_new_n1031__5, new_n1031_);
  not g_20694 (not_new_n5399_, new_n5399_);
  not g_20695 (not_new_n4969_, new_n4969_);
  or g_20696 (new_n8364_, not_new_n8137_, not_new_n630__138412872010);
  not g_20697 (not_new_n4494_, new_n4494_);
  not g_20698 (not_new_n5451__0, new_n5451_);
  not g_20699 (not_pi124_0, pi124);
  not g_20700 (not_new_n2498_, new_n2498_);
  not g_20701 (not_new_n6739_, new_n6739_);
  not g_20702 (not_pi054_1, pi054);
  not g_20703 (not_new_n1071__70, new_n1071_);
  not g_20704 (new_n10008_, new_n619_);
  not g_20705 (not_new_n2028_, new_n2028_);
  not g_20706 (not_new_n8860_, new_n8860_);
  xor g_20707 (key_gate_78, not_new_n596_, key_78);
  not g_20708 (not_new_n4433__0, new_n4433_);
  not g_20709 (not_new_n5785_, new_n5785_);
  or g_20710 (new_n3347_, not_pi049_0, not_new_n1534__168070);
  not g_20711 (not_new_n760_, new_n760_);
  not g_20712 (new_n9937_, new_n622_);
  not g_20713 (not_new_n5558_, new_n5558_);
  or g_20714 (or_not_new_n5917__not_new_n5719__0, not_new_n5917_, not_new_n5719__0);
  or g_20715 (new_n1022_, not_new_n3367_, not_new_n3368_);
  not g_20716 (not_new_n10115_, new_n10115_);
  not g_20717 (not_new_n624__5, new_n624_);
  or g_20718 (new_n3247_, not_new_n1049__5, not_new_n589__113988951853731430);
  not g_20719 (not_new_n6519__1, new_n6519_);
  not g_20720 (new_n6505_, new_n639_);
  not g_20721 (not_new_n2955_, new_n2955_);
  not g_20722 (new_n4521_, new_n4483_);
  or g_20723 (po145, not_new_n3517_, not_new_n3516_);
  or g_20724 (new_n4385_, not_new_n4272_, not_new_n688_);
  or g_20725 (new_n2187_, not_pi152, not_new_n587__138412872010);
  not g_20726 (not_new_n6531__2, new_n6531_);
  or g_20727 (new_n8001_, not_new_n7932__0, not_new_n7745_);
  not g_20728 (not_new_n3855_, new_n3855_);
  not g_20729 (not_new_n6984__1, new_n6984_);
  or g_20730 (new_n9021_, new_n1045_, new_n635_);
  or g_20731 (new_n2602_, not_pi202, not_new_n2509__8);
  and g_20732 (new_n9348_, new_n9545_, new_n9548_);
  or g_20733 (new_n4324_, not_new_n679_, not_new_n4321__0);
  not g_20734 (not_new_n10008_, new_n10008_);
  not g_20735 (not_new_n1047__19773267430, new_n1047_);
  or g_20736 (new_n3220_, not_new_n1071__4, not_new_n3185__1176490);
  not g_20737 (not_new_n9139_, new_n9139_);
  and g_20738 (new_n9337_, new_n9589_, new_n9335_);
  and g_20739 (new_n7737_, new_n7964_, new_n7965_);
  or g_20740 (new_n8417_, not_new_n8342_, not_new_n8340__0);
  not g_20741 (not_new_n2791_, new_n2791_);
  or g_20742 (new_n3056_, not_new_n581__138412872010, not_new_n1067__2);
  not g_20743 (not_new_n2454_, new_n2454_);
  not g_20744 (not_new_n628_, new_n628_);
  or g_20745 (new_n5244_, not_new_n5240_, not_new_n5083_);
  or g_20746 (new_n3047_, not_new_n1037__2, not_new_n581__403536070);
  or g_20747 (new_n2978_, not_new_n604__332329305696010, not_new_n635__3);
  or g_20748 (new_n7780_, not_new_n7753__1, not_new_n642__2824752490);
  not g_20749 (not_new_n1580__6, new_n1580_);
  not g_20750 (not_new_n606__57648010, new_n606_);
  not g_20751 (not_new_n1602__70, new_n1602_);
  not g_20752 (not_new_n600__1176490, new_n600_);
  or g_20753 (new_n6473_, not_new_n634__403536070, not_new_n6478_);
  not g_20754 (not_new_n989__1176490, new_n989_);
  and g_20755 (new_n9864_, new_n10100_, new_n9858_);
  not g_20756 (not_new_n9207_, new_n9207_);
  not g_20757 (not_new_n8393_, new_n8393_);
  not g_20758 (not_new_n3434_, new_n3434_);
  not g_20759 (not_new_n9470_, new_n9470_);
  not g_20760 (not_pi249, pi249);
  not g_20761 (not_new_n3185__2824752490, new_n3185_);
  not g_20762 (not_new_n3372__138412872010, new_n3372_);
  not g_20763 (not_new_n3391_, new_n3391_);
  not g_20764 (not_new_n9622_, new_n9622_);
  not g_20765 (not_new_n1602_, new_n1602_);
  not g_20766 (new_n4935_, new_n635_);
  not g_20767 (not_new_n4469__0, new_n4469_);
  not g_20768 (not_new_n1024__2, new_n1024_);
  not g_20769 (not_new_n7414_, new_n7414_);
  and g_20770 (and_new_n1254__new_n1913_, new_n1254_, new_n1913_);
  not g_20771 (not_new_n7151_, new_n7151_);
  or g_20772 (new_n9004_, new_n1045_, new_n635_);
  not g_20773 (not_new_n644__6782230728490, new_n644_);
  not g_20774 (not_new_n3315__8, new_n3315_);
  or g_20775 (new_n6464_, not_new_n6764_, not_new_n6767_);
  not g_20776 (new_n4818_, new_n4732_);
  or g_20777 (new_n7281_, not_new_n7277_, not_new_n7160_);
  not g_20778 (not_new_n648__24010, new_n648_);
  or g_20779 (new_n5708_, not_new_n5706__0, not_new_n5707_);
  not g_20780 (new_n9140_, new_n8900_);
  not g_20781 (not_new_n4014_, new_n4014_);
  not g_20782 (not_new_n7406_, new_n7406_);
  not g_20783 (not_new_n3999_, new_n3999_);
  or g_20784 (new_n9846_, not_new_n1055__5585458640832840070, not_new_n9393_);
  not g_20785 (not_new_n9511__0, new_n9511_);
  or g_20786 (new_n1171_, not_new_n3872_, not_new_n3871_);
  not g_20787 (not_new_n1011__8, new_n1011_);
  xor g_20788 (key_gate_10, new_n1717_, key_10);
  not g_20789 (not_new_n9590_, new_n9590_);
  not g_20790 (not_pi137_0, pi137);
  or g_20791 (new_n6376_, not_new_n1600__490, not_new_n6280_);
  or g_20792 (new_n2206_, not_new_n587__968890104070, not_pi153);
  not g_20793 (not_new_n4003_, new_n4003_);
  buf g_20794 (po000, pi193);
  not g_20795 (not_new_n1065__968890104070, new_n1065_);
  not g_20796 (not_new_n6951_, new_n6951_);
  and g_20797 (new_n4139_, pi270, pi251);
  or g_20798 (new_n10182_, new_n637_, new_n1065_);
  or g_20799 (new_n10290_, not_new_n9936_, not_new_n622__113988951853731430);
  or g_20800 (new_n9582_, not_new_n644__113988951853731430, not_new_n1059__47475615099430);
  or g_20801 (new_n2588_, not_new_n4468__0, not_new_n610__7);
  or g_20802 (new_n6107_, not_new_n1043__490, not_new_n5755__0);
  not g_20803 (not_new_n8265__0, new_n8265_);
  not g_20804 (not_new_n4081_, new_n4081_);
  not g_20805 (not_new_n588__968890104070, new_n588_);
  or g_20806 (new_n2188_, not_new_n588__138412872010, not_pi120);
  not g_20807 (not_new_n591__2326305139872070, new_n591_);
  not g_20808 (new_n9925_, new_n627_);
  or g_20809 (new_n2736_, not_new_n1588__39098210485829880490, not_new_n994__2);
  not g_20810 (not_new_n637__10, new_n637_);
  not g_20811 (not_new_n7792_, new_n7792_);
  not g_20812 (not_new_n5507__0, new_n5507_);
  not g_20813 (not_new_n6191_, new_n6191_);
  not g_20814 (not_new_n8134__1, new_n8134_);
  or g_20815 (new_n4477_, not_new_n4532_, not_new_n4531_);
  not g_20816 (new_n9397_, new_n1061_);
  not g_20817 (not_new_n7603__1, new_n7603_);
  or g_20818 (new_n7400_, not_new_n7024__0, not_new_n6982__2);
  or g_20819 (new_n8439_, not_new_n8230_, not_new_n8266__3);
  not g_20820 (not_new_n7626_, new_n7626_);
  not g_20821 (not_new_n7008_, new_n7008_);
  or g_20822 (or_or_not_new_n2597__not_new_n2601__not_new_n1435_, not_new_n1435_, or_not_new_n2597__not_new_n2601_);
  not g_20823 (not_new_n3184__2824752490, new_n3184_);
  and g_20824 (new_n4900_, new_n5103_, new_n5104_);
  not g_20825 (not_new_n6459_, new_n6459_);
  not g_20826 (not_new_n5523_, new_n5523_);
  not g_20827 (not_new_n7325_, new_n7325_);
  or g_20828 (new_n8176_, not_new_n8135_, not_new_n1602__57648010);
  or g_20829 (new_n2105_, not_new_n9869_, not_new_n594__1176490);
  or g_20830 (new_n5413_, not_new_n1057__10, not_new_n4963_);
  not g_20831 (not_new_n7950_, new_n7950_);
  or g_20832 (new_n6766_, not_new_n6531__1, not_new_n1065__1176490);
  or g_20833 (or_or_not_new_n2919__not_new_n2922__not_new_n2921_, not_new_n2921_, or_not_new_n2919__not_new_n2922_);
  or g_20834 (new_n9618_, new_n625_, new_n1602_);
  or g_20835 (new_n5348_, not_new_n5346_, not_new_n5347_);
  or g_20836 (new_n6664_, not_new_n1039__168070, not_new_n6482_);
  or g_20837 (new_n6840_, not_new_n6677__0, not_new_n6614_);
  or g_20838 (new_n623_, or_not_new_n2319__not_new_n2320_, not_new_n2321_);
  or g_20839 (new_n3673_, not_new_n647__9, not_po298_9);
  not g_20840 (not_new_n3093_, new_n3093_);
  not g_20841 (not_pi052_0, pi052);
  or g_20842 (new_n5899_, not_new_n5815_, not_new_n1031__3430);
  not g_20843 (not_new_n3254_, new_n3254_);
  or g_20844 (new_n5833_, not_new_n6169_, not_new_n6168_);
  not g_20845 (not_new_n642__7, new_n642_);
  not g_20846 (not_new_n6986_, new_n6986_);
  not g_20847 (not_new_n7706_, new_n7706_);
  not g_20848 (new_n3995_, pi049);
  not g_20849 (not_po298_1176490, po298);
  or g_20850 (new_n9694_, not_new_n618__1915812313805664144010, not_new_n1596__113988951853731430);
  not g_20851 (not_new_n9229_, new_n9229_);
  not g_20852 (not_new_n8142_, new_n8142_);
  not g_20853 (not_new_n598__9, new_n598_);
  or g_20854 (new_n4092_, not_new_n4142_, not_new_n4163_);
  not g_20855 (not_new_n3525_, new_n3525_);
  or g_20856 (new_n1702_, key_gate_104, not_new_n596__138412872010);
  and g_20857 (and_new_n2124__new_n2127_, new_n2124_, new_n2127_);
  not g_20858 (not_new_n1067__2824752490, new_n1067_);
  not g_20859 (not_new_n9336_, new_n9336_);
  not g_20860 (not_new_n635__490, new_n635_);
  not g_20861 (new_n1598_, new_n975_);
  and g_20862 (and_new_n2642__new_n2641_, new_n2641_, new_n2642_);
  not g_20863 (not_new_n598__1176490, new_n598_);
  not g_20864 (not_new_n5068_, new_n5068_);
  not g_20865 (new_n9594_, new_n9427_);
  not g_20866 (not_pi145, pi145);
  or g_20867 (new_n10130_, not_new_n10129_, not_new_n10127_);
  not g_20868 (not_new_n5819_, new_n5819_);
  or g_20869 (new_n1909_, not_new_n1584__6, not_new_n9348_);
  or g_20870 (new_n1770_, not_new_n1585_, not_new_n5737_);
  or g_20871 (new_n969_, not_pi009, not_new_n1536__2);
  not g_20872 (new_n7222_, new_n7016_);
  not g_20873 (not_new_n3197_, new_n3197_);
  not g_20874 (not_new_n1919_, new_n1919_);
  not g_20875 (not_new_n9893__0, new_n9893_);
  not g_20876 (not_new_n7723_, new_n7723_);
  or g_20877 (new_n7513_, not_new_n7442__0, not_new_n726__0);
  not g_20878 (not_new_n9235_, new_n9235_);
  not g_20879 (not_new_n3962_, new_n3962_);
  not g_20880 (not_new_n1598__968890104070, new_n1598_);
  or g_20881 (new_n722_, not_new_n3270_, not_new_n3269_);
  not g_20882 (not_new_n9690_, new_n9690_);
  or g_20883 (new_n6116_, not_new_n5753__0, not_new_n628__8235430);
  or g_20884 (new_n3210_, not_new_n1601__4, not_new_n3185__70);
  or g_20885 (new_n5974_, not_new_n5972_, not_new_n5973_);
  not g_20886 (not_new_n2242_, new_n2242_);
  or g_20887 (new_n1655_, not_new_n1631__6, not_pi040);
  not g_20888 (new_n3429_, new_n1043_);
  not g_20889 (not_new_n10124_, new_n10124_);
  not g_20890 (not_new_n5202_, new_n5202_);
  or g_20891 (or_not_new_n2284__not_new_n2281_, not_new_n2281_, not_new_n2284_);
  not g_20892 (not_new_n3044_, new_n3044_);
  not g_20893 (not_new_n9602_, new_n9602_);
  not g_20894 (not_new_n736_, new_n736_);
  not g_20895 (not_new_n6974__4, new_n6974_);
  not g_20896 (not_new_n3806_, new_n3806_);
  or g_20897 (new_n7510_, not_new_n7508_, not_new_n7509_);
  or g_20898 (new_n4669_, not_new_n1013__4, not_new_n4445__0);
  or g_20899 (new_n1842_, not_new_n1588__3, not_new_n1039_);
  not g_20900 (not_new_n1297_, new_n1297_);
  not g_20901 (not_new_n10306_, new_n10306_);
  or g_20902 (new_n3036_, not_new_n581__168070, not_new_n1601__2);
  not g_20903 (not_new_n2185_, new_n2185_);
  not g_20904 (not_new_n7331_, new_n7331_);
  not g_20905 (not_new_n7585_, new_n7585_);
  not g_20906 (not_new_n6479__0, new_n6479_);
  not g_20907 (not_new_n9380_, new_n9380_);
  not g_20908 (not_new_n10327_, new_n10327_);
  or g_20909 (new_n2895_, not_new_n6970_, not_new_n595__8235430);
  not g_20910 (not_new_n928__47475615099430, new_n928_);
  not g_20911 (not_new_n6298_, new_n6298_);
  or g_20912 (new_n9318_, not_new_n1055__113988951853731430, not_new_n8865_);
  not g_20913 (not_new_n1580__2326305139872070, new_n1580_);
  not g_20914 (not_new_n8266__4, new_n8266_);
  not g_20915 (not_new_n10101_, new_n10101_);
  not g_20916 (not_new_n8803_, new_n8803_);
  or g_20917 (new_n8513_, not_new_n8384_, not_new_n8256__1);
  or g_20918 (new_n6942_, not_new_n6639_, not_new_n6818_);
  and g_20919 (new_n6615_, new_n6844_, new_n6845_);
  and g_20920 (new_n9462_, new_n9574_, new_n9510_);
  not g_20921 (not_new_n8248_, new_n8248_);
  or g_20922 (new_n7393_, not_new_n6981__1, not_new_n7023__1);
  or g_20923 (new_n5638_, not_new_n5434__0, not_pi131_3);
  not g_20924 (new_n3434_, new_n1045_);
  not g_20925 (not_new_n3927__0, new_n3927_);
  not g_20926 (not_new_n1039__490, new_n1039_);
  not g_20927 (not_new_n1027__4, new_n1027_);
  not g_20928 (not_new_n634__1, new_n634_);
  not g_20929 (not_new_n1008__3, new_n1008_);
  or g_20930 (new_n9445_, not_new_n9822_, not_new_n9823_);
  not g_20931 (not_new_n2109__0, new_n2109_);
  or g_20932 (new_n2314_, not_new_n594__2326305139872070, not_new_n9961_);
  not g_20933 (not_new_n7257_, new_n7257_);
  not g_20934 (not_new_n4071__3, new_n4071_);
  or g_20935 (new_n10285_, not_new_n10283_, not_new_n10284_);
  not g_20936 (not_new_n4117__0, new_n4117_);
  not g_20937 (not_new_n588__19773267430, new_n588_);
  not g_20938 (not_new_n1768__1, new_n1768_);
  not g_20939 (not_new_n599__47475615099430, new_n599_);
  not g_20940 (not_new_n8417_, new_n8417_);
  not g_20941 (not_new_n6242__4, new_n6242_);
  or g_20942 (new_n2921_, not_new_n1616__403536070, not_new_n2918_);
  not g_20943 (new_n943_, pi161);
  or g_20944 (new_n2782_, not_new_n630__2, not_new_n602__5);
  or g_20945 (new_n2920_, not_new_n612__5, not_new_n4119__2);
  or g_20946 (or_not_new_n1557__not_new_n2444_, not_new_n1557_, not_new_n2444_);
  or g_20947 (new_n9271_, not_new_n8880_, not_new_n1603__138412872010);
  not g_20948 (not_new_n6993_, new_n6993_);
  not g_20949 (not_new_n622__57648010, new_n622_);
  or g_20950 (new_n673_, not_new_n3092_, or_not_new_n3094__not_new_n3093_);
  not g_20951 (not_new_n6959_, new_n6959_);
  xnor g_20952 (key_gate_14, new_n1690_, key_14);
  or g_20953 (new_n1917_, not_new_n591__7, not_new_n4728_);
  or g_20954 (new_n1991_, not_new_n594__10, not_new_n9973_);
  or g_20955 (new_n9804_, not_new_n9425__0, not_new_n1604__332329305696010);
  not g_20956 (not_new_n3515_, new_n3515_);
  or g_20957 (new_n10276_, not_new_n618__225393402906922580878632490, not_new_n9946__0);
  and g_20958 (new_n1532_, new_n3244_, new_n3243_);
  not g_20959 (not_new_n9901__0, new_n9901_);
  not g_20960 (not_new_n984__3430, new_n984_);
  not g_20961 (not_new_n6349_, new_n6349_);
  not g_20962 (new_n5914_, new_n5740_);
  or g_20963 (new_n5258_, not_new_n5138_, not_new_n5091__0);
  not g_20964 (not_new_n5690_, new_n5690_);
  or g_20965 (new_n4119_, not_new_n4189_, not_new_n4190_);
  not g_20966 (not_new_n5031_, new_n5031_);
  not g_20967 (not_new_n9917__0, new_n9917_);
  not g_20968 (not_new_n6477__0, new_n6477_);
  not g_20969 (not_new_n3541_, new_n3541_);
  or g_20970 (new_n8450_, not_new_n8127_, not_new_n8201_);
  or g_20971 (new_n5176_, new_n645_, new_n1071_);
  not g_20972 (new_n4111_, pi267);
  not g_20973 (not_new_n1588__70, new_n1588_);
  not g_20974 (not_new_n8644_, new_n8644_);
  not g_20975 (new_n4248_, new_n699_);
  not g_20976 (not_new_n4177_, new_n4177_);
  not g_20977 (not_new_n1485_, new_n1485_);
  or g_20978 (new_n1828_, not_new_n585__3, not_new_n4118_);
  or g_20979 (or_not_new_n5448__not_new_n5597__1, not_new_n5448_, not_new_n5597__1);
  not g_20980 (not_new_n1007__4, new_n1007_);
  not g_20981 (not_new_n6358_, new_n6358_);
  not g_20982 (new_n4427_, pi168);
  or g_20983 (new_n7390_, not_new_n7342__0, not_new_n741__0);
  not g_20984 (not_new_n1614__0, new_n1614_);
  not g_20985 (not_new_n5912_, new_n5912_);
  not g_20986 (not_new_n1591__57648010, new_n1591_);
  or g_20987 (new_n6090_, not_new_n5865_, not_new_n6064_);
  not g_20988 (not_new_n594__968890104070, new_n594_);
  not g_20989 (not_pi033_0, pi033);
  not g_20990 (not_new_n6490_, new_n6490_);
  not g_20991 (not_new_n3724_, new_n3724_);
  or g_20992 (new_n1037_, not_new_n3412_, not_new_n3413_);
  not g_20993 (not_new_n7242_, new_n7242_);
  not g_20994 (new_n3409_, new_n1035_);
  not g_20995 (not_pi250, pi250);
  and g_20996 (and_and_new_n2257__new_n2260__new_n2258_, new_n2258_, and_new_n2257__new_n2260_);
  not g_20997 (not_new_n6464_, new_n6464_);
  not g_20998 (new_n6914_, new_n6602_);
  or g_20999 (new_n7952_, not_new_n1049__57648010, not_new_n7598__1);
  not g_21000 (not_new_n10063_, new_n10063_);
  not g_21001 (not_new_n3912_, new_n3912_);
  not g_21002 (not_new_n1848_, new_n1848_);
  not g_21003 (not_new_n5379_, new_n5379_);
  not g_21004 (not_new_n6170_, new_n6170_);
  not g_21005 (not_new_n9414_, new_n9414_);
  not g_21006 (not_pi026, pi026);
  not g_21007 (not_new_n591__5585458640832840070, new_n591_);
  not g_21008 (not_new_n2534_, new_n2534_);
  not g_21009 (not_new_n9910__0, new_n9910_);
  or g_21010 (new_n3501_, not_new_n2147_, not_new_n1613__57648010);
  not g_21011 (not_new_n608__490, new_n608_);
  not g_21012 (not_new_n5958_, new_n5958_);
  not g_21013 (not_new_n9412_, new_n9412_);
  or g_21014 (or_not_pi257_3_not_pi260_3, not_pi257_3, not_pi260_3);
  not g_21015 (not_pi014, pi014);
  not g_21016 (not_new_n5787_, new_n5787_);
  and g_21017 (new_n5721_, new_n5920_, and_new_n5938__new_n5933_);
  or g_21018 (new_n6051_, not_new_n5995_, not_new_n5994_);
  not g_21019 (not_new_n6240_, new_n6240_);
  not g_21020 (not_new_n979_, new_n979_);
  or g_21021 (new_n10020_, not_new_n10234_, not_new_n9992_);
  or g_21022 (new_n3911_, not_new_n10107_, not_new_n10344_);
  or g_21023 (or_not_new_n1024__0_not_new_n3384__2, not_new_n3384__2, not_new_n1024__0);
  not g_21024 (not_new_n1793_, new_n1793_);
  or g_21025 (new_n6055_, not_new_n6005_, not_new_n5810_);
  not g_21026 (not_new_n1546_, new_n1546_);
  not g_21027 (new_n4254_, new_n697_);
  not g_21028 (not_new_n6583_, new_n6583_);
  not g_21029 (not_new_n8144_, new_n8144_);
  not g_21030 (not_new_n8162__1, new_n8162_);
  and g_21031 (new_n5864_, new_n5775_, new_n6056_);
  not g_21032 (not_new_n8713__2, new_n8713_);
  not g_21033 (not_new_n594_, new_n594_);
  or g_21034 (or_or_not_new_n1557__not_new_n2444__not_new_n1383_, not_new_n1383_, or_not_new_n1557__not_new_n2444_);
  not g_21035 (not_new_n3684_, new_n3684_);
  not g_21036 (new_n8600_, new_n1053_);
  not g_21037 (new_n6729_, new_n6513_);
  not g_21038 (not_new_n2320_, new_n2320_);
  not g_21039 (not_new_n8208_, new_n8208_);
  not g_21040 (not_new_n1537__2, new_n1537_);
  not g_21041 (not_new_n3517_, new_n3517_);
  not g_21042 (not_new_n5805__0, new_n5805_);
  or g_21043 (new_n7750_, not_new_n7925_, not_new_n7917_);
  not g_21044 (not_new_n2917_, new_n2917_);
  not g_21045 (not_new_n4217_, new_n4217_);
  not g_21046 (not_new_n3500_, new_n3500_);
  not g_21047 (not_pi173_2, pi173);
  not g_21048 (not_new_n1045__16284135979104490, new_n1045_);
  or g_21049 (or_not_new_n5893__0_not_new_n6159__0, not_new_n6159__0, not_new_n5893__0);
  not g_21050 (not_new_n581__881247870897231951843937366879128181133112010, new_n581_);
  or g_21051 (new_n8588_, not_new_n8158__2, not_new_n626__273687473400809163430);
  not g_21052 (new_n6476_, new_n1045_);
  not g_21053 (not_new_n738__0, new_n738_);
  or g_21054 (new_n9768_, not_new_n1597__113988951853731430, not_new_n9377__0);
  or g_21055 (new_n3215_, not_new_n589__3430, not_new_n639__7);
  not g_21056 (not_new_n5594_, new_n5594_);
  or g_21057 (new_n4041_, not_pi050_3, not_new_n4040_);
  not g_21058 (not_new_n609__3430, new_n609_);
  not g_21059 (new_n4243_, new_n704_);
  not g_21060 (not_new_n5793__0, new_n5793_);
  not g_21061 (not_new_n6999__1, new_n6999_);
  not g_21062 (not_new_n5737_, new_n5737_);
  or g_21063 (new_n8112_, not_new_n632__968890104070, not_new_n8114_);
  or g_21064 (or_or_not_new_n6349__not_new_n6373__7_not_new_n1041__490, or_not_new_n6349__not_new_n6373__7, not_new_n1041__490);
  or g_21065 (new_n2741_, not_new_n612_, not_new_n4121__2);
  not g_21066 (not_new_n1596__2, new_n1596_);
  not g_21067 (not_new_n3311_, new_n3311_);
  not g_21068 (not_po296_93874803376477543056490, po296);
  not g_21069 (not_pi260_4, pi260);
  not g_21070 (not_new_n4473__0, new_n4473_);
  not g_21071 (not_new_n9519_, new_n9519_);
  or g_21072 (new_n9227_, not_new_n9226_, not_new_n9225_);
  not g_21073 (not_new_n6694_, new_n6694_);
  not g_21074 (not_new_n7189_, new_n7189_);
  not g_21075 (not_new_n9679_, new_n9679_);
  or g_21076 (new_n3589_, not_new_n1612__797922662976120010, not_new_n2348__0);
  or g_21077 (new_n4872_, not_new_n1603__7, not_new_n4743_);
  not g_21078 (not_new_n10016_, new_n10016_);
  not g_21079 (not_new_n604__1, new_n604_);
  or g_21080 (new_n4658_, not_new_n4492_, not_new_n4451__0);
  not g_21081 (not_new_n631__4, new_n631_);
  not g_21082 (new_n8142_, new_n645_);
  not g_21083 (not_new_n6168_, new_n6168_);
  not g_21084 (not_new_n1907_, new_n1907_);
  and g_21085 (and_new_n2995__new_n998_, new_n998_, new_n2995_);
  not g_21086 (not_new_n5579_, new_n5579_);
  not g_21087 (not_new_n2808_, new_n2808_);
  not g_21088 (not_new_n4786_, new_n4786_);
  not g_21089 (not_new_n2096_, new_n2096_);
  not g_21090 (new_n6257_, new_n1601_);
  not g_21091 (not_new_n7272_, new_n7272_);
  not g_21092 (not_new_n1065__3, new_n1065_);
  and g_21093 (po095, pi074, key_gate_101);
  not g_21094 (not_new_n7732_, new_n7732_);
  not g_21095 (new_n9404_, new_n1069_);
  or g_21096 (new_n2989_, or_not_new_n7047__0_not_new_n3369__0, not_new_n1021__0);
  not g_21097 (not_new_n8293_, new_n8293_);
  or g_21098 (or_not_new_n1342__not_new_n1343_, not_new_n1342_, not_new_n1343_);
  or g_21099 (or_not_new_n2926__not_new_n2925_, not_new_n2926_, not_new_n2925_);
  not g_21100 (new_n7098_, new_n765_);
  not g_21101 (not_new_n3734_, new_n3734_);
  not g_21102 (not_new_n8799__0, new_n8799_);
  or g_21103 (new_n4697_, not_new_n4437__0, not_new_n1017__4);
  not g_21104 (not_new_n5749__0, new_n5749_);
  not g_21105 (not_new_n680_, new_n680_);
  not g_21106 (new_n8119_, new_n631_);
  or g_21107 (new_n7548_, not_new_n733__0, not_new_n7415__2);
  or g_21108 (new_n9014_, new_n1051_, new_n647_);
  or g_21109 (new_n2292_, not_new_n1591__332329305696010, not_new_n8910_);
  not g_21110 (not_new_n2923_, new_n2923_);
  not g_21111 (not_new_n6665_, new_n6665_);
  or g_21112 (new_n6377_, not_new_n6376_, not_new_n6308_);
  or g_21113 (new_n9601_, not_new_n9331_, not_new_n9427_);
  not g_21114 (not_new_n4133__2, new_n4133_);
  not g_21115 (not_new_n7974_, new_n7974_);
  not g_21116 (not_new_n3778_, new_n3778_);
  or g_21117 (new_n3348_, not_new_n3996__0, not_pi064_168070);
  or g_21118 (new_n994_, not_new_n1472_, not_new_n584_);
  or g_21119 (new_n8910_, not_new_n9242_, not_new_n9243_);
  and g_21120 (new_n1446_, new_n1620_, new_n2657_);
  or g_21121 (new_n2331_, not_new_n6467_, not_new_n1580__113988951853731430);
  not g_21122 (not_new_n4253_, new_n4253_);
  and g_21123 (new_n6449_, new_n6716_, new_n6715_);
  and g_21124 (new_n9492_, new_n9766_, new_n9765_);
  or g_21125 (new_n2857_, not_new_n3310__8, not_new_n4117__2);
  or g_21126 (new_n8759_, not_new_n8613_, not_new_n1059__19773267430);
  not g_21127 (new_n8709_, new_n1162_);
  or g_21128 (new_n5312_, not_new_n1041__9, not_new_n4926_);
  not g_21129 (not_new_n1057__3430, new_n1057_);
  or g_21130 (new_n3527_, not_new_n1612_, not_new_n1781__0);
  not g_21131 (not_new_n5060_, new_n5060_);
  not g_21132 (not_new_n586__1, new_n586_);
  not g_21133 (not_new_n622__0, new_n622_);
  or g_21134 (new_n4483_, not_new_n4520_, not_new_n4519_);
  not g_21135 (not_new_n603__1176490, new_n603_);
  or g_21136 (new_n6849_, not_new_n624__403536070, not_new_n6477__0);
  xnor g_21137 (key_gate_79, key_79, new_n1639_);
  and g_21138 (po090, key_gate_101, pi069);
  and g_21139 (new_n599_, new_n1579_, new_n1611_);
  not g_21140 (new_n6619_, new_n1607_);
  or g_21141 (new_n2448_, not_new_n4128__0, not_new_n600__57648010);
  not g_21142 (not_new_n1588__4, new_n1588_);
  not g_21143 (not_new_n8532_, new_n8532_);
  or g_21144 (new_n6470_, not_new_n6686_, not_new_n6688_);
  or g_21145 (new_n8563_, not_new_n1065__47475615099430, not_new_n8162__2);
  not g_21146 (not_new_n643__332329305696010, new_n643_);
  not g_21147 (not_new_n7650__0, new_n7650_);
  not g_21148 (not_new_n634__490, new_n634_);
  or g_21149 (or_not_new_n6508__1_not_new_n6600_, not_new_n6508__1, not_new_n6600_);
  or g_21150 (new_n1021_, not_new_n3365_, not_new_n3364_);
  not g_21151 (not_new_n8574_, new_n8574_);
  or g_21152 (new_n5671_, not_new_n5512_, not_new_n5513__0);
  or g_21153 (new_n2651_, not_new_n606__3430, not_new_n5480__0);
  not g_21154 (not_new_n8219_, new_n8219_);
  or g_21155 (new_n9012_, not_new_n8956_, not_new_n9011_);
  not g_21156 (not_new_n3669_, new_n3669_);
  not g_21157 (not_new_n7747_, new_n7747_);
  and g_21158 (new_n1202_, new_n1695_, new_n1697_);
  not g_21159 (new_n6493_, new_n647_);
  or g_21160 (new_n1925_, not_new_n634__0, not_new_n601__6);
  not g_21161 (not_new_n7781_, new_n7781_);
  not g_21162 (not_new_n10107_, new_n10107_);
  not g_21163 (not_new_n5078__3, new_n5078_);
  not g_21164 (new_n8129_, new_n1597_);
  not g_21165 (not_new_n6780_, new_n6780_);
  not g_21166 (not_new_n2509__1176490, new_n2509_);
  or g_21167 (new_n4614_, not_new_n4529_, not_new_n4612_);
  not g_21168 (not_new_n640__2326305139872070, new_n640_);
  or g_21169 (po058, key_gate_97, not_new_n1185_);
  not g_21170 (new_n3384_, new_n1028_);
  not g_21171 (not_new_n5275_, new_n5275_);
  not g_21172 (not_pi051_0, pi051);
  not g_21173 (not_new_n1069__6, new_n1069_);
  not g_21174 (not_new_n6723_, new_n6723_);
  not g_21175 (not_new_n1534__490, key_gate_5);
  not g_21176 (not_new_n4113__0, new_n4113_);
  not g_21177 (not_new_n8108_, new_n8108_);
  not g_21178 (not_new_n1053__8, new_n1053_);
  not g_21179 (not_new_n1766_, new_n1766_);
  not g_21180 (not_new_n4809_, new_n4809_);
  and g_21181 (and_new_n1972__new_n1975_, new_n1972_, new_n1975_);
  or g_21182 (new_n9600_, not_new_n9597_, not_new_n1067__138412872010);
  not g_21183 (not_new_n9011_, new_n9011_);
  or g_21184 (new_n2286_, not_new_n601__47475615099430, not_new_n621__0);
  or g_21185 (new_n7791_, not_new_n1041__168070, not_new_n7613_);
  or g_21186 (new_n9837_, not_new_n9835_, not_new_n9588_);
  or g_21187 (new_n2576_, not_new_n2573_, or_not_new_n2575__not_new_n2574_);
  not g_21188 (not_new_n751_, new_n751_);
  not g_21189 (not_new_n8369_, new_n8369_);
  not g_21190 (not_new_n9587_, new_n9587_);
  not g_21191 (not_new_n6124_, new_n6124_);
  not g_21192 (not_new_n5492__0, new_n5492_);
  not g_21193 (not_pi265_1, pi265);
  not g_21194 (not_new_n4233_, new_n4233_);
  and g_21195 (po109, key_gate_101, pi088);
  not g_21196 (not_new_n4726_, new_n4726_);
  not g_21197 (not_new_n6526__0, new_n6526_);
  not g_21198 (not_new_n10309_, new_n10309_);
  or g_21199 (new_n5374_, not_new_n5373_, not_new_n5372_);
  not g_21200 (not_new_n591__2, new_n591_);
  not g_21201 (not_new_n4515_, new_n4515_);
  not g_21202 (not_new_n6478_, new_n6478_);
  not g_21203 (not_new_n644__47475615099430, new_n644_);
  or g_21204 (new_n5330_, not_new_n4993_, not_new_n618__24010);
  not g_21205 (not_new_n5496_, new_n5496_);
  not g_21206 (not_new_n4691_, new_n4691_);
  not g_21207 (not_new_n1607__24010, new_n1607_);
  not g_21208 (not_new_n1039__1, new_n1039_);
  not g_21209 (not_new_n7635__0, new_n7635_);
  not g_21210 (not_new_n622__47475615099430, new_n622_);
  not g_21211 (not_new_n6487__2, new_n6487_);
  not g_21212 (not_new_n1374_, new_n1374_);
  or g_21213 (new_n7344_, not_new_n6974__1, not_new_n773_);
  or g_21214 (new_n7589_, not_new_n7879_, not_new_n7882_);
  not g_21215 (not_new_n8098_, new_n8098_);
  not g_21216 (not_new_n1053__403536070, new_n1053_);
  not g_21217 (not_new_n4025_, new_n4025_);
  or g_21218 (new_n6069_, not_new_n5878__0, not_new_n5723_);
  and g_21219 (and_new_n6373__new_n6389_, new_n6373_, new_n6389_);
  not g_21220 (not_new_n600__0, new_n600_);
  and g_21221 (and_new_n6451__new_n6799_, new_n6799_, new_n6451_);
  or g_21222 (new_n5640_, not_new_n5503_, not_new_n5504__0);
  not g_21223 (not_new_n1538__403536070, new_n1538_);
  or g_21224 (new_n5016_, not_new_n5387_, not_new_n5388_);
  not g_21225 (new_n7649_, new_n626_);
  or g_21226 (new_n3615_, not_new_n955_, not_new_n1611__70);
  or g_21227 (new_n3830_, not_new_n1576__0, not_new_n648__490);
  not g_21228 (not_new_n9539__0, new_n9539_);
  or g_21229 (new_n2822_, not_new_n1616__8, not_new_n2819_);
  or g_21230 (new_n3677_, not_new_n627__9, not_po298_70);
  or g_21231 (new_n9231_, not_new_n1596__332329305696010, not_new_n8892_);
  not g_21232 (not_new_n4664_, new_n4664_);
  not g_21233 (not_new_n10141_, new_n10141_);
  or g_21234 (new_n9054_, not_new_n644__332329305696010, not_new_n1059__138412872010);
  not g_21235 (not_new_n3096_, new_n3096_);
  not g_21236 (not_new_n8041_, new_n8041_);
  not g_21237 (not_new_n8788_, new_n8788_);
  not g_21238 (not_new_n6179_, new_n6179_);
  and g_21239 (new_n1414_, new_n2514_, new_n2511_);
  not g_21240 (not_new_n1228_, new_n1228_);
  or g_21241 (new_n3059_, not_new_n581__968890104070, not_new_n1065__2);
  not g_21242 (not_new_n600__403536070, new_n600_);
  not g_21243 (not_new_n5012_, new_n5012_);
  or g_21244 (new_n2456_, not_new_n4784__0, not_new_n597__403536070);
  or g_21245 (new_n3410_, not_new_n1537__0, not_pi098_0);
  not g_21246 (not_new_n2899_, new_n2899_);
  not g_21247 (new_n5281_, new_n4991_);
  and g_21248 (new_n6579_, and_new_n6481__new_n6853_, new_n6852_);
  or g_21249 (new_n5170_, not_new_n4985_, not_new_n4984_);
  or g_21250 (new_n5686_, not_new_n5562_, not_new_n5461_);
  not g_21251 (new_n4447_, pi178);
  not g_21252 (not_new_n7611__2, new_n7611_);
  not g_21253 (not_new_n9365_, new_n9365_);
  not g_21254 (not_new_n5982_, new_n5982_);
  not g_21255 (not_new_n1576__24010, new_n1576_);
  not g_21256 (not_new_n5395_, new_n5395_);
  and g_21257 (new_n9995_, new_n10288_, and_new_n10034__new_n10289_);
  not g_21258 (not_new_n595__6, new_n595_);
  not g_21259 (not_new_n603__47475615099430, new_n603_);
  or g_21260 (new_n9382_, not_new_n1600__968890104070, not_new_n629__332329305696010);
  or g_21261 (new_n1854_, not_new_n6562_, not_new_n1580__4);
  not g_21262 (not_new_n3194_, new_n3194_);
  not g_21263 (not_new_n1693_, key_gate_52);
  or g_21264 (new_n2584_, not_new_n1018_, not_new_n607__5);
  or g_21265 (new_n4668_, not_pi177_2, not_new_n4446_);
  or g_21266 (new_n3399_, not_new_n1728__113988951853731430, not_pi066_0);
  or g_21267 (new_n8574_, not_new_n8152__0, not_new_n1059__2824752490);
  or g_21268 (new_n3279_, not_new_n1071__5, not_new_n589__3788186922656647816827176259430);
  or g_21269 (new_n2259_, not_new_n591__47475615099430, not_new_n4771_);
  not g_21270 (not_new_n2115_, new_n2115_);
  not g_21271 (not_new_n7572_, new_n7572_);
  not g_21272 (not_new_n606__1, new_n606_);
  or g_21273 (new_n6823_, not_new_n6481__1, not_new_n6663_);
  or g_21274 (new_n3273_, not_new_n589__11044276742439206463052992010, not_new_n1603__5);
  not g_21275 (not_new_n1585__1176490, new_n1585_);
  not g_21276 (not_new_n9335_, new_n9335_);
  not g_21277 (not_new_n7917_, new_n7917_);
  or g_21278 (new_n7786_, not_new_n7611_, not_new_n1045__403536070);
  not g_21279 (not_new_n4459_, new_n4459_);
  not g_21280 (not_new_n4604_, new_n4604_);
  not g_21281 (not_pi147_2, pi147);
  not g_21282 (not_new_n5435__1, new_n5435_);
  not g_21283 (not_new_n2985_, new_n2985_);
  not g_21284 (not_new_n9633_, new_n9633_);
  not g_21285 (new_n4964_, new_n1055_);
  not g_21286 (not_new_n2726_, new_n2726_);
  or g_21287 (new_n9313_, not_new_n1057__138412872010, not_new_n8863_);
  not g_21288 (not_new_n6564_, new_n6564_);
  not g_21289 (not_new_n7648_, new_n7648_);
  and g_21290 (new_n1208_, new_n1715_, new_n1713_);
  not g_21291 (not_new_n9036_, new_n9036_);
  or g_21292 (new_n2050_, not_new_n4801_, not_new_n591__24010);
  or g_21293 (new_n8570_, not_new_n1061__2824752490, not_new_n8164__0);
  not g_21294 (not_new_n8249_, new_n8249_);
  not g_21295 (not_new_n611__7, new_n611_);
  not g_21296 (new_n7118_, new_n761_);
  or g_21297 (new_n5818_, not_new_n6156_, not_new_n6155_);
  not g_21298 (new_n10224_, new_n10006_);
  not g_21299 (not_new_n3432_, new_n3432_);
  not g_21300 (not_new_n1536__2, new_n1536_);
  and g_21301 (new_n8690_, and_and_new_n8753__new_n8754__new_n8761_, new_n8755_);
  not g_21302 (not_new_n1558_, new_n1558_);
  or g_21303 (new_n7428_, not_new_n7124_, not_new_n775__57648010);
  and g_21304 (new_n1299_, new_n2121_, and_new_n1298__new_n2122_);
  not g_21305 (not_new_n640__70, new_n640_);
  and g_21306 (new_n4476_, new_n4602_, new_n4601_);
  not g_21307 (not_pi257_5, pi257);
  not g_21308 (not_new_n9720_, new_n9720_);
  not g_21309 (not_new_n581__968890104070, new_n581_);
  or g_21310 (new_n2711_, not_new_n998_, not_new_n2709_);
  not g_21311 (not_new_n7284_, new_n7284_);
  and g_21312 (new_n6573_, new_n6681_, new_n6680_);
  or g_21313 (new_n7371_, not_new_n7357__1, not_new_n737__1);
  not g_21314 (new_n9170_, new_n8896_);
  not g_21315 (not_new_n1013__0, new_n1013_);
  not g_21316 (not_new_n4779_, new_n4779_);
  not g_21317 (not_new_n7624__0, new_n7624_);
  not g_21318 (not_new_n1607__2, new_n1607_);
  or g_21319 (new_n2519_, not_pi249, not_po296_39098210485829880490);
  or g_21320 (new_n749_, not_new_n3206_, not_new_n3207_);
  not g_21321 (not_new_n6643_, new_n6643_);
  not g_21322 (not_new_n1594__2, new_n1594_);
  or g_21323 (new_n687_, not_new_n3029_, not_new_n1504_);
  not g_21324 (not_new_n2294_, new_n2294_);
  or g_21325 (new_n7239_, not_new_n7237_, not_new_n7083_);
  or g_21326 (new_n3134_, not_new_n639__5, not_new_n3315__1176490);
  or g_21327 (po285, not_new_n2893_, or_or_or_not_new_n2892__not_new_n2895__not_new_n2894__not_new_n2896_);
  not g_21328 (not_new_n6576_, new_n6576_);
  not g_21329 (not_new_n7343_, new_n7343_);
  not g_21330 (new_n4430_, new_n1003_);
  not g_21331 (not_new_n8164_, new_n8164_);
  not g_21332 (not_new_n1069__24010, new_n1069_);
  or g_21333 (new_n2752_, not_new_n595__1, not_new_n7050_);
  not g_21334 (not_new_n4538_, new_n4538_);
  not g_21335 (not_new_n7840_, new_n7840_);
  not g_21336 (not_new_n8833__0, new_n8833_);
  not g_21337 (not_new_n3342_, new_n3342_);
  not g_21338 (new_n5987_, new_n5802_);
  not g_21339 (not_new_n9078_, new_n9078_);
  not g_21340 (not_pi083, pi083);
  or g_21341 (new_n3751_, not_new_n1602__6, not_new_n625__10);
  not g_21342 (not_new_n8805_, new_n8805_);
  or g_21343 (new_n10320_, not_new_n9949__0, not_new_n1604__113988951853731430);
  not g_21344 (not_new_n1607__7, new_n1607_);
  and g_21345 (new_n1197_, new_n1682_, new_n1680_);
  or g_21346 (new_n4151_, not_pi263_1, not_new_n4159__0);
  not g_21347 (not_new_n6635__2, new_n6635_);
  not g_21348 (not_new_n1028_, new_n1028_);
  not g_21349 (not_new_n6712_, new_n6712_);
  not g_21350 (new_n4836_, new_n4778_);
  not g_21351 (not_new_n2796_, new_n2796_);
  not g_21352 (not_new_n1583__57648010, new_n1583_);
  not g_21353 (not_new_n1045__7, new_n1045_);
  not g_21354 (not_new_n597__332329305696010, new_n597_);
  not g_21355 (new_n9102_, new_n8965_);
  not g_21356 (not_new_n2149_, new_n2149_);
  or g_21357 (new_n2649_, not_po296_3788186922656647816827176259430, not_pi260);
  or g_21358 (new_n2098_, not_new_n1585__1176490, not_new_n5823_);
  not g_21359 (not_new_n2777_, new_n2777_);
  not g_21360 (not_new_n928__5, new_n928_);
  not g_21361 (not_new_n1631__3430, key_gate_76);
  buf g_21362 (po014, pi207);
  not g_21363 (not_new_n6898_, new_n6898_);
  not g_21364 (not_new_n8088_, new_n8088_);
  or g_21365 (new_n8017_, not_new_n7670__0, not_new_n7884_);
  and g_21366 (and_new_n10033__new_n3902_, new_n3902_, new_n10033_);
  not g_21367 (not_new_n1589__3, new_n1589_);
  not g_21368 (not_new_n1612__4, new_n1612_);
  not g_21369 (not_new_n3372__1915812313805664144010, new_n3372_);
  not g_21370 (not_new_n2709_, new_n2709_);
  or g_21371 (new_n4029_, not_pi058_3, not_new_n4028_);
  or g_21372 (new_n9049_, not_new_n9047_, not_new_n9048_);
  not g_21373 (not_new_n7277_, new_n7277_);
  or g_21374 (new_n5369_, not_new_n5189_, not_new_n5367_);
  not g_21375 (not_new_n1043__24010, new_n1043_);
  and g_21376 (new_n8928_, and_new_n8837__new_n9203_, new_n9202_);
  not g_21377 (not_new_n7293_, new_n7293_);
  or g_21378 (new_n4629_, not_new_n1008__3, not_new_n4419_);
  not g_21379 (not_new_n2979_, new_n2979_);
  not g_21380 (not_new_n8113__2, new_n8113_);
  or g_21381 (new_n2620_, not_new_n608__10, not_new_n1003__0);
  not g_21382 (not_new_n8223_, new_n8223_);
  or g_21383 (or_not_new_n2072__not_new_n2073_, not_new_n2072_, not_new_n2073_);
  not g_21384 (not_new_n6488__0, new_n6488_);
  not g_21385 (not_new_n9589_, new_n9589_);
  or g_21386 (new_n7493_, not_new_n7008__0, not_new_n7040__0);
  or g_21387 (or_not_new_n2208__not_new_n2205_, not_new_n2205_, not_new_n2208_);
  not g_21388 (new_n4436_, new_n1018_);
  not g_21389 (not_new_n9523__1, new_n9523_);
  not g_21390 (not_new_n9097_, new_n9097_);
  not g_21391 (not_new_n1059__7, new_n1059_);
  not g_21392 (not_new_n7739__1, new_n7739_);
  or g_21393 (new_n10098_, not_new_n644__39098210485829880490, not_new_n1059__16284135979104490);
  not g_21394 (new_n6522_, new_n1059_);
  or g_21395 (new_n2476_, not_new_n4774__0, not_new_n597__968890104070);
  not g_21396 (not_new_n1594__3430, new_n1594_);
  not g_21397 (not_new_n596__968890104070, key_gate_88);
  not g_21398 (not_new_n618__332329305696010, new_n618_);
  not g_21399 (not_new_n7192_, new_n7192_);
  not g_21400 (not_new_n634__8235430, new_n634_);
  not g_21401 (not_new_n5928_, new_n5928_);
  or g_21402 (new_n3012_, not_new_n581__7, not_new_n1606__1);
  or g_21403 (new_n7275_, not_new_n7454__1, not_new_n7010__1);
  or g_21404 (new_n2073_, not_pi146, not_new_n587__1176490);
  not g_21405 (not_new_n1601__5, new_n1601_);
  not g_21406 (not_new_n1170_, new_n1170_);
  not g_21407 (not_new_n3315__57648010, new_n3315_);
  not g_21408 (not_new_n4239_, new_n4239_);
  not g_21409 (not_pi011_0, pi011);
  not g_21410 (not_new_n1039__968890104070, new_n1039_);
  or g_21411 (new_n6421_, or_or_or_not_new_n6240__not_new_n6330__not_new_n6331__not_new_n6242__1, not_new_n6227_);
  not g_21412 (not_new_n5795_, new_n5795_);
  not g_21413 (not_pi119, pi119);
  not g_21414 (not_new_n1537__10, new_n1537_);
  not g_21415 (not_new_n2497_, new_n2497_);
  not g_21416 (not_new_n8132_, new_n8132_);
  or g_21417 (new_n5303_, not_new_n4936_, not_new_n1047__10);
  not g_21418 (not_new_n7458_, new_n7458_);
  not g_21419 (not_new_n1067__2326305139872070, new_n1067_);
  or g_21420 (new_n9686_, not_new_n9519__0, not_new_n9566_);
  not g_21421 (not_new_n1945_, new_n1945_);
  not g_21422 (not_new_n587__16284135979104490, new_n587_);
  or g_21423 (new_n9610_, not_new_n9608_, not_new_n9609_);
  xnor g_21424 (key_gate_96, not_new_n1708_, key_96);
  not g_21425 (not_new_n9410_, new_n9410_);
  or g_21426 (po069, key_gate_92, not_new_n1196_);
  and g_21427 (new_n3927_, new_n4024_, new_n4018_);
  not g_21428 (not_new_n4411__0, new_n4411_);
  or g_21429 (or_or_not_new_n1559__not_new_n2454__not_new_n1387_, or_not_new_n1559__not_new_n2454_, not_new_n1387_);
  or g_21430 (new_n7970_, not_new_n7739__2, not_new_n7818_);
  not g_21431 (not_new_n1720_, key_gate_83);
  not g_21432 (new_n8635_, new_n1150_);
  not g_21433 (not_new_n953_, new_n953_);
  not g_21434 (not_new_n680__0, new_n680_);
  or g_21435 (new_n2496_, not_new_n597__2326305139872070, not_new_n4764__0);
  not g_21436 (not_new_n7597__1, new_n7597_);
  not g_21437 (not_new_n5629_, new_n5629_);
  not g_21438 (not_new_n1049__2, new_n1049_);
  or g_21439 (new_n2794_, not_new_n1059__1, not_new_n3311__4);
  not g_21440 (not_new_n2966_, new_n2966_);
  not g_21441 (not_new_n7680_, new_n7680_);
  not g_21442 (not_new_n9867__0, new_n9867_);
  or g_21443 (new_n2881_, not_new_n4135__1, not_new_n994__57648010);
  or g_21444 (new_n1153_, not_new_n3836_, not_new_n3835_);
  not g_21445 (not_new_n4115__1, new_n4115_);
  not g_21446 (not_new_n1067__168070, new_n1067_);
  or g_21447 (new_n5823_, not_new_n6194_, not_new_n6193_);
  or g_21448 (new_n5821_, not_new_n6183_, not_new_n6184_);
  or g_21449 (new_n5557_, not_pi140_1, not_new_n1018__5);
  not g_21450 (not_new_n7170_, new_n7170_);
  or g_21451 (new_n2834_, not_new_n604__10, not_new_n630__3);
  not g_21452 (not_new_n5790_, new_n5790_);
  not g_21453 (not_new_n6083_, new_n6083_);
  not g_21454 (not_new_n1596__13410686196639649008070, new_n1596_);
  or g_21455 (new_n3493_, not_new_n1594__8235430, not_new_n1011__0);
  or g_21456 (new_n3707_, not_po298_332329305696010, not_new_n621__9);
  not g_21457 (new_n7765_, new_n7662_);
  not g_21458 (not_new_n6709__0, new_n6709_);
  or g_21459 (new_n9291_, not_new_n8881_, not_new_n637__47475615099430);
  not g_21460 (not_new_n9056_, new_n9056_);
  not g_21461 (not_new_n3927_, new_n3927_);
  not g_21462 (not_new_n4001__1, new_n4001_);
  not g_21463 (not_new_n3827_, new_n3827_);
  or g_21464 (new_n10056_, not_new_n9879_, not_new_n9880_);
  or g_21465 (or_not_new_n2577__not_new_n2581_, not_new_n2581_, not_new_n2577_);
  or g_21466 (new_n2308_, not_new_n1584__2326305139872070, not_new_n9437_);
  or g_21467 (or_not_new_n1763__not_new_n1764_, not_new_n1763_, not_new_n1764_);
  or g_21468 (new_n7896_, not_new_n7837__0, not_new_n7658__0);
  or g_21469 (new_n7948_, not_new_n1051__1176490, not_new_n7617__0);
  not g_21470 (not_new_n611__4, new_n611_);
  or g_21471 (new_n9163_, not_new_n9138_, not_new_n8884__1);
  not g_21472 (not_new_n2479_, new_n2479_);
  not g_21473 (not_new_n2719_, new_n2719_);
  not g_21474 (not_new_n626__8235430, new_n626_);
  or g_21475 (new_n4365_, not_new_n4261_, not_new_n662_);
  not g_21476 (not_new_n8046_, new_n8046_);
  not g_21477 (not_new_n5984__0, new_n5984_);
  or g_21478 (new_n2215_, not_new_n6465_, not_new_n1580__968890104070);
  not g_21479 (not_new_n4154_, new_n4154_);
  or g_21480 (new_n3574_, not_new_n1538__968890104070, not_pi153_0);
  or g_21481 (new_n10255_, not_new_n624__113988951853731430, not_new_n9885_);
  or g_21482 (new_n2116_, not_new_n7680_, not_new_n1583__8235430);
  or g_21483 (or_not_new_n9694__not_new_n9634_, not_new_n9694_, not_new_n9634_);
  not g_21484 (not_new_n2078_, new_n2078_);
  not g_21485 (not_new_n642__2326305139872070, new_n642_);
  not g_21486 (not_new_n6731_, new_n6731_);
  not g_21487 (not_new_n588__797922662976120010, new_n588_);
  buf g_21488 (po049, pi215);
  or g_21489 (new_n10109_, not_new_n638__32199057558131797268376070, not_new_n1063__332329305696010);
  not g_21490 (not_new_n10109_, new_n10109_);
  not g_21491 (not_new_n6161_, new_n6161_);
  not g_21492 (not_pi044_1, pi044);
  not g_21493 (not_new_n4950__0, new_n4950_);
  not g_21494 (not_new_n7388_, new_n7388_);
  not g_21495 (not_new_n646__490, new_n646_);
  or g_21496 (new_n8729_, not_new_n1045__2326305139872070, not_new_n8633_);
  not g_21497 (new_n9883_, new_n1039_);
  not g_21498 (not_new_n1576__7, new_n1576_);
  not g_21499 (not_new_n640__168070, new_n640_);
  or g_21500 (new_n3304_, not_new_n6467__0, not_new_n1580__797922662976120010);
  not g_21501 (not_new_n4470_, new_n4470_);
  not g_21502 (not_new_n5739__0, new_n5739_);
  or g_21503 (new_n3958_, not_new_n4053_, not_new_n4054_);
  not g_21504 (not_new_n4974__0, new_n4974_);
  not g_21505 (not_new_n1265_, new_n1265_);
  or g_21506 (or_not_new_n2605__not_new_n2604_, not_new_n2604_, not_new_n2605_);
  and g_21507 (new_n1374_, new_n2420_, new_n2421_);
  or g_21508 (new_n3293_, not_new_n1057__5, not_new_n589__3119734822845423713013303218219760490);
  or g_21509 (new_n7087_, not_new_n7459_, not_new_n7458_);
  or g_21510 (new_n3684_, not_pi228, not_new_n989__24010);
  not g_21511 (not_new_n1537__332329305696010, new_n1537_);
  or g_21512 (new_n4747_, or_not_new_n4841__not_new_n4762_, not_new_n4765_);
  or g_21513 (new_n9372_, not_new_n9387_, not_new_n9540_);
  not g_21514 (not_new_n638__1915812313805664144010, new_n638_);
  not g_21515 (not_new_n7179_, new_n7179_);
  or g_21516 (new_n6926_, not_new_n6604_, not_new_n6636__0);
  or g_21517 (new_n2449_, not_new_n599__57648010, not_new_n9967__0);
  or g_21518 (new_n7257_, not_new_n7085_, not_new_n7255_);
  not g_21519 (not_new_n4757__0, new_n4757_);
  not g_21520 (not_new_n640__968890104070, new_n640_);
  not g_21521 (not_new_n2740_, new_n2740_);
  and g_21522 (new_n1302_, new_n2139_, new_n2138_);
  not g_21523 (not_new_n689_, new_n689_);
  and g_21524 (new_n8803_, new_n9068_, new_n9067_);
  not g_21525 (not_pi061_1, pi061);
  or g_21526 (new_n10306_, not_new_n10134_, not_new_n10304_);
  or g_21527 (new_n3130_, not_new_n581__185621159210175743024531636712070, not_new_n630__6);
  and g_21528 (new_n1353_, and_new_n2369__new_n2368_, new_n2367_);
  or g_21529 (new_n7871_, not_new_n7870_, not_new_n7718_);
  not g_21530 (not_new_n3311__168070, new_n3311_);
  not g_21531 (not_new_n5710_, new_n5710_);
  not g_21532 (not_new_n9624_, new_n9624_);
  not g_21533 (not_new_n7252_, new_n7252_);
  not g_21534 (not_new_n4072_, new_n4072_);
  not g_21535 (not_new_n1329_, new_n1329_);
  or g_21536 (new_n9367_, not_new_n9535_, not_new_n9536_);
  not g_21537 (not_new_n4204_, new_n4204_);
  or g_21538 (new_n8854_, not_new_n1600__19773267430, not_new_n629__6782230728490);
  or g_21539 (new_n2916_, not_new_n602__2824752490, not_new_n619__1);
  not g_21540 (not_new_n2710_, new_n2710_);
  not g_21541 (not_new_n7716_, new_n7716_);
  not g_21542 (not_new_n3480_, new_n3480_);
  not g_21543 (not_new_n2054_, new_n2054_);
  not g_21544 (not_new_n6233__0, new_n6233_);
  not g_21545 (not_new_n1612__2, new_n1612_);
  not g_21546 (not_new_n5833_, new_n5833_);
  and g_21547 (new_n7086_, new_n7261_, new_n7264_);
  or g_21548 (new_n6173_, not_new_n6172_, not_new_n6058_);
  and g_21549 (new_n10012_, new_n10274_, new_n10275_);
  or g_21550 (po138, not_new_n3502_, not_new_n3503_);
  and g_21551 (new_n9327_, new_n9520_, new_n9519_);
  not g_21552 (not_new_n6443__403536070, new_n6443_);
  or g_21553 (new_n3017_, not_new_n1027__490, not_new_n1158_);
  or g_21554 (new_n7191_, not_new_n7190_, not_new_n7074_);
  or g_21555 (new_n8489_, not_new_n8114__0, not_new_n632__6782230728490);
  not g_21556 (new_n4545_, new_n4508_);
  or g_21557 (new_n708_, not_new_n3006_, not_new_n1492_);
  not g_21558 (not_new_n1597__403536070, new_n1597_);
  not g_21559 (new_n4831_, new_n4741_);
  or g_21560 (new_n7772_, not_new_n7604_, not_new_n1037__1176490);
  not g_21561 (not_pi170_1, pi170);
  not g_21562 (not_new_n7216_, new_n7216_);
  not g_21563 (not_new_n5823_, new_n5823_);
  not g_21564 (new_n7321_, new_n6990_);
  not g_21565 (not_new_n6104_, new_n6104_);
  or g_21566 (new_n3357_, not_new_n1534__2824752490, not_pi044_0);
  or g_21567 (new_n5687_, not_new_n5459__1, not_pi142_3);
  or g_21568 (new_n9250_, not_new_n9248_, not_new_n9109__0);
  or g_21569 (new_n10296_, not_new_n1600__332329305696010, not_new_n9939_);
  not g_21570 (not_new_n8271__0, new_n8271_);
  not g_21571 (not_new_n8230_, new_n8230_);
  not g_21572 (not_new_n5514_, new_n5514_);
  not g_21573 (not_new_n7543_, new_n7543_);
  or g_21574 (new_n2473_, not_new_n4123__0, not_new_n600__968890104070);
  or g_21575 (new_n5660_, not_new_n5471_, not_pi146_2);
  and g_21576 (new_n9999_, new_n9860_, new_n10174_);
  not g_21577 (not_new_n3327_, new_n3327_);
  and g_21578 (new_n5886_, new_n6130_, new_n6129_);
  not g_21579 (not_new_n4305_, new_n4305_);
  or g_21580 (new_n1691_, not_pi052, not_new_n1631__57648010);
  not g_21581 (not_new_n1847_, new_n1847_);
  not g_21582 (not_new_n1611__6782230728490, new_n1611_);
  or g_21583 (new_n3954_, not_new_n3961_, not_new_n4001__0);
  not g_21584 (not_new_n4928_, new_n4928_);
  or g_21585 (new_n2097_, not_new_n7681_, not_new_n1583__1176490);
  not g_21586 (new_n4246_, new_n701_);
  not g_21587 (not_new_n9637_, new_n9637_);
  or g_21588 (new_n3014_, not_new_n581__8, not_new_n1039__2);
  not g_21589 (not_new_n2717_, new_n2717_);
  not g_21590 (not_new_n3287_, new_n3287_);
  not g_21591 (not_new_n589__77309937197074445241370944070, new_n589_);
  not g_21592 (not_new_n1455_, new_n1455_);
  and g_21593 (new_n9983_, and_new_n9888__new_n10254_, new_n10253_);
  or g_21594 (new_n2915_, not_new_n617__3, not_new_n604__403536070);
  not g_21595 (not_new_n1425_, new_n1425_);
  not g_21596 (new_n8873_, new_n645_);
  not g_21597 (not_pi230, pi230);
  not g_21598 (not_new_n603_, new_n603_);
  or g_21599 (new_n5827_, not_new_n6103_, not_new_n6102_);
  and g_21600 (and_new_n5938__new_n5933_, new_n5933_, new_n5938_);
  not g_21601 (not_new_n632__16284135979104490, new_n632_);
  not g_21602 (not_new_n8287__0, new_n8287_);
  not g_21603 (not_new_n6008_, new_n6008_);
  not g_21604 (new_n6810_, new_n6625_);
  not g_21605 (not_new_n3384__3, new_n3384_);
  not g_21606 (not_new_n5063__1, new_n5063_);
  not g_21607 (new_n5941_, new_n5758_);
  not g_21608 (not_new_n1728__16284135979104490, new_n1728_);
  not g_21609 (not_new_n596__168070, key_gate_88);
  or g_21610 (new_n5874_, not_new_n6212_, not_new_n6211_);
  not g_21611 (not_new_n2765_, new_n2765_);
  not g_21612 (not_new_n645__1176490, new_n645_);
  not g_21613 (not_new_n4292_, new_n4292_);
  not g_21614 (not_new_n4775__0, new_n4775_);
  not g_21615 (not_new_n7321_, new_n7321_);
  not g_21616 (not_new_n8316_, new_n8316_);
  not g_21617 (not_new_n6620_, new_n6620_);
  not g_21618 (new_n1603_, new_n965_);
  not g_21619 (new_n5230_, new_n5072_);
  and g_21620 (new_n5903_, new_n6199_, new_n6198_);
  and g_21621 (new_n9329_, new_n9572_, new_n9571_);
  not g_21622 (new_n5741_, new_n648_);
  or g_21623 (new_n3798_, not_new_n3796_, not_new_n3797_);
  or g_21624 (new_n7530_, not_new_n7016__1, not_new_n7307_);
  or g_21625 (new_n3820_, not_new_n992_, or_not_new_n1028__8_not_new_n1622__1);
  or g_21626 (new_n10314_, not_new_n639__39098210485829880490, not_new_n9910_);
  not g_21627 (not_pi270_0, pi270);
  not g_21628 (not_new_n610__6, new_n610_);
  or g_21629 (new_n2831_, not_new_n1616__9, not_new_n2828_);
  not g_21630 (new_n4283_, new_n651_);
  not g_21631 (not_new_n604__6, new_n604_);
  or g_21632 (new_n4597_, not_pi169_3, not_new_n4430__0);
  not g_21633 (not_new_n6486__0, new_n6486_);
  not g_21634 (not_new_n4928__0, new_n4928_);
  or g_21635 (new_n10266_, not_new_n1037__113988951853731430, not_new_n9882_);
  not g_21636 (not_new_n1583__5, new_n1583_);
  not g_21637 (not_new_n603__2824752490, new_n603_);
  not g_21638 (not_new_n6114_, new_n6114_);
  or g_21639 (po255, not_new_n3696_, not_new_n3697_);
  not g_21640 (not_new_n8196_, new_n8196_);
  and g_21641 (and_new_n9412__new_n9818_, new_n9412_, new_n9818_);
  not g_21642 (not_new_n1018__3, new_n1018_);
  not g_21643 (not_new_n2969_, new_n2969_);
  not g_21644 (not_new_n3931_, key_gate_6);
  not g_21645 (not_new_n601__7, new_n601_);
  not g_21646 (not_new_n3913__0, new_n3913_);
  or g_21647 (new_n7299_, not_new_n7297_, not_new_n7096_);
  or g_21648 (new_n5549_, not_new_n5496_, not_new_n5548_);
  or g_21649 (new_n8394_, not_new_n8393_, not_new_n8392_);
  or g_21650 (new_n9678_, not_new_n9677_, not_new_n9482_);
  or g_21651 (new_n9247_, not_new_n8890_, not_new_n1599__19773267430);
  not g_21652 (not_new_n589__1176490, new_n589_);
  not g_21653 (not_new_n1049__138412872010, new_n1049_);
  or g_21654 (or_not_new_n2847__not_new_n2850_, not_new_n2850_, not_new_n2847_);
  not g_21655 (not_new_n2190_, new_n2190_);
  not g_21656 (not_new_n5644_, new_n5644_);
  not g_21657 (not_new_n2509__2, new_n2509_);
  not g_21658 (not_new_n1272_, new_n1272_);
  not g_21659 (not_new_n8150__1, new_n8150_);
  not g_21660 (not_new_n591__6, new_n591_);
  not g_21661 (not_new_n6631__0, new_n6631_);
  not g_21662 (not_new_n3184__8, new_n3184_);
  not g_21663 (not_new_n4157__0, new_n4157_);
  not g_21664 (not_new_n6373_, new_n6373_);
  not g_21665 (not_new_n1596__797922662976120010, new_n1596_);
  not g_21666 (not_new_n2957_, new_n2957_);
  not g_21667 (not_pi023, pi023);
  not g_21668 (new_n7363_, new_n7021_);
  not g_21669 (not_pi260_0, pi260);
  or g_21670 (new_n5498_, not_new_n5539_, not_new_n5538_);
  not g_21671 (not_new_n3675_, new_n3675_);
  not g_21672 (not_new_n5687_, new_n5687_);
  not g_21673 (not_new_n3310__7, new_n3310_);
  not g_21674 (not_new_n1011__3, new_n1011_);
  or g_21675 (new_n2628_, not_new_n610__70, not_new_n4455__0);
  or g_21676 (new_n4544_, not_new_n1002__2, not_pi170_1);
  not g_21677 (not_new_n3184__57648010, new_n3184_);
  not g_21678 (not_new_n4293_, new_n4293_);
  or g_21679 (new_n4012_, not_new_n3956_, not_new_n4004__0);
  not g_21680 (new_n6290_, new_n1059_);
  or g_21681 (new_n8430_, not_new_n8368__1, not_new_n8175__0);
  not g_21682 (not_new_n8231_, new_n8231_);
  or g_21683 (new_n5523_, new_n1009_, pi131);
  not g_21684 (not_new_n2037_, new_n2037_);
  not g_21685 (not_new_n7618__0, new_n7618_);
  or g_21686 (new_n9168_, or_not_new_n8995__1_not_new_n8799__1, not_new_n8798__2);
  not g_21687 (not_new_n591__168070, new_n591_);
  not g_21688 (not_new_n948_, new_n948_);
  not g_21689 (not_new_n4984_, new_n4984_);
  not g_21690 (not_new_n4441_, new_n4441_);
  not g_21691 (not_new_n8871_, new_n8871_);
  not g_21692 (not_new_n6443__24010, new_n6443_);
  or g_21693 (new_n5420_, not_new_n5078__3, not_new_n5265_);
  or g_21694 (new_n1950_, not_new_n1591__8, not_new_n8903_);
  not g_21695 (not_new_n3932_, key_gate_15);
  not g_21696 (not_new_n9814_, new_n9814_);
  not g_21697 (not_new_n994__1, new_n994_);
  or g_21698 (new_n3792_, not_new_n3790_, not_new_n3791_);
  not g_21699 (not_new_n10073_, new_n10073_);
  not g_21700 (not_new_n5733_, new_n5733_);
  not g_21701 (not_new_n8490_, new_n8490_);
  not g_21702 (not_new_n1004__2, new_n1004_);
  not g_21703 (not_new_n1589__70, new_n1589_);
  or g_21704 (new_n6684_, not_new_n6683_, not_new_n6528__0);
  not g_21705 (new_n6909_, new_n6601_);
  not g_21706 (not_new_n7436_, new_n7436_);
  or g_21707 (new_n666_, or_not_new_n3161__not_new_n3160_, not_new_n3159_);
  not g_21708 (not_new_n625__5, new_n625_);
  not g_21709 (not_new_n591__70, new_n591_);
  or g_21710 (new_n7295_, not_new_n7294_, not_new_n7017_);
  not g_21711 (not_new_n5458_, new_n5458_);
  not g_21712 (not_new_n4793__0, new_n4793_);
  not g_21713 (not_pi048_4, pi048);
  not g_21714 (not_new_n600__57648010, new_n600_);
  not g_21715 (not_pi258, pi258);
  not g_21716 (not_new_n6651_, new_n6651_);
  not g_21717 (not_new_n9447_, new_n9447_);
  not g_21718 (not_new_n4261_, new_n4261_);
  not g_21719 (not_new_n9900__2, new_n9900_);
  or g_21720 (new_n2110_, not_pi180, not_new_n586__57648010);
  not g_21721 (not_new_n2225_, new_n2225_);
  not g_21722 (not_new_n7943_, new_n7943_);
  not g_21723 (not_new_n8991__0, new_n8991_);
  not g_21724 (not_new_n2536_, new_n2536_);
  or g_21725 (new_n2936_, not_new_n2933_, or_not_new_n2935__not_new_n2934_);
  not g_21726 (not_new_n1588__403536070, new_n1588_);
  not g_21727 (not_pi142, pi142);
  not g_21728 (not_new_n1920_, new_n1920_);
  not g_21729 (not_new_n9374_, new_n9374_);
  not g_21730 (not_pi132_1, pi132);
  and g_21731 (new_n1410_, new_n985_, new_n920_);
  or g_21732 (new_n9644_, new_n1599_, new_n622_);
  or g_21733 (new_n8571_, not_new_n643__332329305696010, not_new_n8151__0);
  not g_21734 (not_new_n3384__6, new_n3384_);
  not g_21735 (not_new_n6974__70, new_n6974_);
  not g_21736 (not_pi143_1, pi143);
  and g_21737 (new_n1340_, new_n2316_, and_and_new_n2314__new_n2317__new_n2315_);
  not g_21738 (not_new_n7735_, new_n7735_);
  not g_21739 (not_new_n7713_, new_n7713_);
  or g_21740 (new_n8381_, not_new_n1596__19773267430, not_new_n8172_);
  and g_21741 (po104, key_gate_101, pi083);
  not g_21742 (not_new_n1059__0, new_n1059_);
  and g_21743 (and_new_n7662__new_n7994_, new_n7662_, new_n7994_);
  not g_21744 (not_new_n8546_, new_n8546_);
  not g_21745 (not_new_n7064_, new_n7064_);
  not g_21746 (not_new_n8596__1, new_n8596_);
  not g_21747 (new_n4814_, new_n4730_);
  or g_21748 (new_n8194_, not_new_n8490_, not_new_n8491_);
  not g_21749 (not_new_n1728__3430, new_n1728_);
  not g_21750 (not_pi164_2, pi164);
  and g_21751 (new_n8813_, new_n9143_, new_n9146_);
  or g_21752 (or_or_not_new_n4240__not_new_n4343__not_new_n704_, not_new_n704_, or_not_new_n4240__not_new_n4343_);
  or g_21753 (new_n4206_, not_new_n4167__0, not_new_n4097_);
  not g_21754 (not_new_n1584__3, new_n1584_);
  not g_21755 (not_new_n626__39098210485829880490, new_n626_);
  not g_21756 (not_new_n4825_, new_n4825_);
  not g_21757 (not_new_n7849_, new_n7849_);
  or g_21758 (new_n2868_, not_new_n595__24010, not_new_n7064_);
  not g_21759 (new_n4105_, pi258);
  not g_21760 (not_new_n1051__7, new_n1051_);
  not g_21761 (not_new_n587__3, new_n587_);
  or g_21762 (new_n714_, not_new_n3375_, not_new_n939_);
  or g_21763 (new_n10344_, not_new_n10343_, not_new_n10342_);
  not g_21764 (not_new_n1008__1, new_n1008_);
  not g_21765 (not_new_n4572_, new_n4572_);
  not g_21766 (not_new_n1611__7, new_n1611_);
  and g_21767 (new_n1199_, new_n1688_, new_n1686_);
  or g_21768 (new_n9526_, not_new_n9452_, not_new_n9326__0);
  not g_21769 (new_n9066_, new_n8899_);
  not g_21770 (not_new_n8279_, new_n8279_);
  not g_21771 (not_new_n1018__0, new_n1018_);
  not g_21772 (not_pi118, pi118);
  or g_21773 (new_n8395_, not_new_n8238_, not_new_n8394_);
  not g_21774 (not_new_n2855_, new_n2855_);
  not g_21775 (not_new_n6154_, new_n6154_);
  or g_21776 (new_n4356_, not_new_n697_, not_new_n4255_);
  or g_21777 (new_n1787_, not_pi097, not_new_n588__1);
  not g_21778 (not_new_n2755_, new_n2755_);
  not g_21779 (not_new_n8129__0, new_n8129_);
  not g_21780 (not_new_n1690_, key_gate_14);
  not g_21781 (not_new_n7947_, new_n7947_);
  not g_21782 (not_new_n4174__0, new_n4174_);
  and g_21783 (new_n8203_, new_n8084_, new_n8083_);
  or g_21784 (new_n7043_, not_new_n7450_, not_new_n7449_);
  or g_21785 (new_n8528_, not_new_n8439_, or_not_new_n8139__1_not_new_n8231_);
  not g_21786 (not_new_n8630_, new_n8630_);
  not g_21787 (not_new_n4017__0, new_n4017_);
  or g_21788 (new_n2800_, not_new_n602__7, not_new_n639__3);
  not g_21789 (not_new_n744__0, new_n744_);
  or g_21790 (new_n1809_, not_new_n585__2, not_new_n4071_);
  not g_21791 (not_new_n652_, new_n652_);
  not g_21792 (not_new_n8899__3, new_n8899_);
  or g_21793 (new_n3483_, not_new_n1013__1, not_new_n1594__168070);
  or g_21794 (new_n2735_, or_not_new_n2734__not_new_n2733_, not_new_n2732_);
  or g_21795 (new_n2796_, not_new_n2793_, not_new_n1616__6);
  not g_21796 (not_new_n8599_, new_n8599_);
  not g_21797 (not_new_n8098__0, new_n8098_);
  not g_21798 (not_new_n9133_, new_n9133_);
  or g_21799 (new_n6079_, not_new_n5748__1, not_new_n5928_);
  not g_21800 (not_new_n1037__57648010, new_n1037_);
  not g_21801 (not_new_n1584__4, new_n1584_);
  or g_21802 (new_n9304_, not_new_n8870_, not_new_n1061__968890104070);
  or g_21803 (new_n8409_, not_new_n8281__0, not_new_n8408_);
  not g_21804 (not_new_n1470_, new_n1470_);
  not g_21805 (not_new_n5445_, new_n5445_);
  not g_21806 (not_new_n6974__8235430, new_n6974_);
  or g_21807 (new_n3269_, not_new_n589__225393402906922580878632490, not_new_n1601__5);
  not g_21808 (new_n9408_, new_n639_);
  not g_21809 (not_new_n3926_, new_n3926_);
  or g_21810 (new_n7362_, not_new_n6974__7, not_new_n767_);
  not g_21811 (not_new_n8109_, new_n8109_);
  not g_21812 (not_new_n8092_, new_n8092_);
  or g_21813 (new_n1931_, not_new_n8904_, not_new_n1591__7);
  or g_21814 (new_n7286_, not_new_n7285_, not_new_n7016__0);
  and g_21815 (new_n1264_, and_and_new_n1953__new_n1956__new_n1954_, new_n1955_);
  not g_21816 (not_new_n1063__2326305139872070, new_n1063_);
  not g_21817 (not_new_n1530_, new_n1530_);
  not g_21818 (not_pi086, pi086);
  and g_21819 (new_n4788_, new_n4879_, new_n4878_);
  not g_21820 (not_new_n604__138412872010, new_n604_);
  not g_21821 (not_new_n690_, new_n690_);
  or g_21822 (new_n3477_, not_new_n1536__16284135979104490, not_pi017_0);
  not g_21823 (new_n10134_, new_n10018_);
  not g_21824 (not_new_n1161_, new_n1161_);
  or g_21825 (new_n5944_, not_new_n5740_, not_new_n5741__0);
  or g_21826 (new_n8455_, not_new_n8358_, not_new_n8267_);
  not g_21827 (not_new_n4366_, new_n4366_);
  not g_21828 (not_new_n599__168070, new_n599_);
  not g_21829 (not_new_n4583_, new_n4583_);
  not g_21830 (not_pi175_2, pi175);
  or g_21831 (new_n9000_, not_new_n8999_, not_new_n631__39098210485829880490);
  or g_21832 (new_n1960_, not_pi108, not_new_n588__10);
  not g_21833 (not_new_n9892_, new_n9892_);
  not g_21834 (new_n6300_, new_n1602_);
  not g_21835 (not_new_n1047__70, new_n1047_);
  not g_21836 (not_new_n10183_, new_n10183_);
  or g_21837 (new_n4516_, not_pi163_1, not_new_n1009__2);
  not g_21838 (not_new_n594__19773267430, new_n594_);
  not g_21839 (not_new_n4935_, new_n4935_);
  or g_21840 (new_n4200_, not_new_n4170__0, not_new_n4103_);
  or g_21841 (new_n3250_, not_new_n3184__1, not_new_n634__8);
  not g_21842 (not_new_n5774_, new_n5774_);
  not g_21843 (not_new_n6171_, new_n6171_);
  or g_21844 (new_n10100_, new_n627_, new_n1055_);
  not g_21845 (new_n8438_, new_n8257_);
  or g_21846 (new_n9319_, not_new_n9317_, not_new_n9318_);
  or g_21847 (new_n9971_, not_new_n3905_, not_new_n3904_);
  not g_21848 (not_new_n6525_, new_n6525_);
  and g_21849 (and_new_n6016__new_n5855_, new_n6016_, new_n5855_);
  not g_21850 (not_new_n3362_, new_n3362_);
  not g_21851 (not_new_n1039__5, new_n1039_);
  or g_21852 (new_n7307_, not_new_n6993__1, not_new_n7291_);
  not g_21853 (not_new_n633__168070, new_n633_);
  not g_21854 (not_new_n1287_, new_n1287_);
  not g_21855 (not_new_n10235_, new_n10235_);
  not g_21856 (not_new_n619__403536070, new_n619_);
  or g_21857 (new_n9108_, not_new_n8966_, not_new_n9099_);
  not g_21858 (not_new_n1537__7, new_n1537_);
  not g_21859 (not_new_n627__0, new_n627_);
  not g_21860 (new_n4425_, pi167);
  or g_21861 (new_n9811_, not_new_n9646__0, not_new_n9809_);
  not g_21862 (not_new_n2109_, new_n2109_);
  not g_21863 (not_new_n626__10, new_n626_);
  not g_21864 (not_new_n588__490, new_n588_);
  not g_21865 (new_n6825_, new_n6635_);
  not g_21866 (not_new_n5162_, new_n5162_);
  not g_21867 (not_new_n5686_, new_n5686_);
  not g_21868 (new_n6820_, new_n6617_);
  or g_21869 (new_n8994_, new_n642_, new_n1035_);
  not g_21870 (not_new_n1051__1, new_n1051_);
  not g_21871 (not_new_n7646_, new_n7646_);
  not g_21872 (not_new_n2902_, new_n2902_);
  or g_21873 (new_n3140_, not_new_n645__5, not_new_n3315__57648010);
  not g_21874 (not_new_n1057__8235430, new_n1057_);
  not g_21875 (not_pi134_0, pi134);
  not g_21876 (not_new_n928__3, new_n928_);
  or g_21877 (new_n9799_, not_new_n1603__47475615099430, not_new_n9408_);
  not g_21878 (not_new_n627__9, new_n627_);
  not g_21879 (not_new_n5696_, new_n5696_);
  not g_21880 (not_new_n3709_, new_n3709_);
  not g_21881 (not_new_n928__403536070, new_n928_);
  or g_21882 (new_n10118_, new_n645_, new_n1071_);
  or g_21883 (new_n2852_, not_new_n604__490, not_new_n624__2);
  or g_21884 (new_n7232_, not_new_n7231_, not_new_n7148_);
  or g_21885 (new_n5939_, not_new_n1045__70, not_new_n5754__0);
  or g_21886 (new_n5613_, not_new_n5612_, not_new_n5611_);
  not g_21887 (not_new_n617__273687473400809163430, new_n617_);
  not g_21888 (new_n5988_, new_n5902_);
  or g_21889 (new_n9702_, not_new_n9587__0, not_new_n9590_);
  not g_21890 (not_new_n5199__0, new_n5199_);
  not g_21891 (not_new_n635__6782230728490, new_n635_);
  not g_21892 (not_new_n10026_, new_n10026_);
  or g_21893 (or_or_not_new_n4933__not_new_n4930__0_not_new_n5322_, not_new_n5322_, or_not_new_n4933__not_new_n4930__0);
  not g_21894 (new_n6292_, new_n1604_);
  not g_21895 (not_new_n5978_, new_n5978_);
  or g_21896 (new_n3683_, not_new_n643__9, not_po298_24010);
  not g_21897 (not_new_n1583__19773267430, new_n1583_);
  not g_21898 (not_new_n10199_, new_n10199_);
  not g_21899 (not_new_n6893_, new_n6893_);
  or g_21900 (new_n5362_, not_new_n5360_, not_new_n5192__0);
  not g_21901 (not_new_n601__2, new_n601_);
  or g_21902 (new_n3153_, not_new_n1065__3, not_new_n928__138412872010);
  not g_21903 (not_new_n4159__1, new_n4159_);
  not g_21904 (not_new_n630__7, new_n630_);
  or g_21905 (new_n3180_, not_new_n986__0, not_new_n937_);
  not g_21906 (not_new_n4457_, new_n4457_);
  or g_21907 (or_not_new_n2607__not_new_n2611_, not_new_n2611_, not_new_n2607_);
  or g_21908 (new_n1788_, not_pi129, not_new_n587__1);
  and g_21909 (new_n9994_, new_n10142_, new_n10034_);
  not g_21910 (not_new_n7446_, new_n7446_);
  and g_21911 (new_n1482_, new_n2859_, new_n2860_);
  not g_21912 (not_new_n8370_, new_n8370_);
  or g_21913 (new_n6925_, not_new_n6924_, not_new_n6726_);
  not g_21914 (not_new_n1601__168070, new_n1601_);
  or g_21915 (new_n9179_, not_new_n8808_, not_new_n8896_);
  or g_21916 (new_n9691_, not_new_n9666_, not_new_n9412__1);
  or g_21917 (new_n3504_, not_new_n1537__2824752490, not_pi118_0);
  or g_21918 (new_n758_, not_new_n3227_, not_new_n3226_);
  and g_21919 (new_n5068_, new_n5364_, new_n5363_);
  not g_21920 (not_new_n1536__2326305139872070, new_n1536_);
  not g_21921 (not_new_n3572_, new_n3572_);
  not g_21922 (not_new_n4455__0, new_n4455_);
  and g_21923 (new_n1484_, new_n2904_, new_n2905_);
  not g_21924 (not_new_n596__1, key_gate_88);
  not g_21925 (new_n7439_, new_n7039_);
  not g_21926 (not_new_n630__1176490, new_n630_);
  not g_21927 (not_new_n5654_, new_n5654_);
  not g_21928 (new_n5429_, new_n1020_);
  not g_21929 (new_n9417_, new_n1599_);
  not g_21930 (not_new_n8137__0, new_n8137_);
  not g_21931 (not_new_n6018_, new_n6018_);
  or g_21932 (new_n6186_, not_new_n5803__0, not_new_n646__1176490);
  not g_21933 (not_new_n8202_, new_n8202_);
  not g_21934 (not_new_n4438_, new_n4438_);
  not g_21935 (not_new_n6328_, new_n6328_);
  not g_21936 (not_pi168, pi168);
  or g_21937 (new_n8762_, not_new_n8596__0, not_new_n8683_);
  xnor g_21938 (key_gate_63, key_63, not_pi033);
  not g_21939 (not_new_n8595__5, new_n8595_);
  not g_21940 (not_new_n670_, new_n670_);
  or g_21941 (or_or_not_new_n6363__not_new_n6358__not_new_n6361_, or_not_new_n6363__not_new_n6358_, not_new_n6361_);
  not g_21942 (new_n4719_, new_n620_);
  not g_21943 (not_new_n9491_, new_n9491_);
  not g_21944 (not_new_n7748_, new_n7748_);
  or g_21945 (or_not_new_n6318__not_new_n6373__0, not_new_n6373__0, not_new_n6318_);
  not g_21946 (not_new_n631__332329305696010, new_n631_);
  not g_21947 (not_new_n641__9, new_n641_);
  not g_21948 (not_new_n1590_, new_n1590_);
  not g_21949 (not_new_n642__968890104070, new_n642_);
  not g_21950 (not_new_n3280_, new_n3280_);
  not g_21951 (not_new_n8875__0, new_n8875_);
  not g_21952 (not_new_n3310__5, new_n3310_);
  or g_21953 (new_n4388_, not_new_n4274_, not_new_n655_);
  and g_21954 (new_n1406_, and_new_n934__new_n986_, new_n937_);
  or g_21955 (new_n2841_, not_new_n7057_, not_new_n595__70);
  or g_21956 (new_n4700_, not_new_n4503_, not_new_n4504__0);
  not g_21957 (not_new_n7735__0, new_n7735_);
  not g_21958 (not_new_n5084__0, new_n5084_);
  or g_21959 (new_n6748_, not_new_n6647_, not_new_n617__2824752490);
  not g_21960 (not_new_n4082_, new_n4082_);
  or g_21961 (new_n6390_, not_new_n6264_, not_new_n646__8235430);
  not g_21962 (not_new_n4534_, new_n4534_);
  not g_21963 (not_new_n1666_, key_gate_115);
  or g_21964 (new_n9316_, not_new_n9314_, not_new_n9140__0);
  not g_21965 (not_new_n5719__0, new_n5719_);
  not g_21966 (not_new_n1708_, key_gate_111);
  not g_21967 (not_new_n4797__1, new_n4797_);
  or g_21968 (new_n7820_, not_new_n7605__0, not_new_n7772_);
  not g_21969 (not_new_n3176_, new_n3176_);
  or g_21970 (new_n9730_, not_new_n9366__0, not_new_n634__797922662976120010);
  or g_21971 (new_n4207_, not_pi268_2, not_new_n4094_);
  and g_21972 (and_new_n8984__new_n9245_, new_n9245_, new_n8984_);
  or g_21973 (new_n9307_, not_new_n9306_, not_new_n9305_);
  and g_21974 (new_n6354_, new_n6232_, new_n6265_);
  not g_21975 (not_new_n8158__2, new_n8158_);
  not g_21976 (not_new_n989__332329305696010, new_n989_);
  not g_21977 (new_n4826_, new_n4805_);
  not g_21978 (not_new_n4136_, new_n4136_);
  not g_21979 (not_new_n1059__57648010, new_n1059_);
  or g_21980 (po189, or_not_new_n1546__not_new_n1362_, not_new_n1361_);
  or g_21981 (new_n776_, not_new_n3825_, or_not_new_n2989__not_new_n3826_);
  not g_21982 (not_new_n5374_, new_n5374_);
  and g_21983 (new_n7578_, new_n7796_, new_n7774_);
  not g_21984 (not_new_n5534_, new_n5534_);
  not g_21985 (not_new_n3466_, new_n3466_);
  not g_21986 (not_new_n8134__0, new_n8134_);
  not g_21987 (not_new_n7874_, new_n7874_);
  not g_21988 (new_n8632_, new_n1153_);
  and g_21989 (new_n8077_, new_n8281_, new_n8334_);
  not g_21990 (not_new_n3426_, new_n3426_);
  not g_21991 (not_new_n1783_, new_n1783_);
  not g_21992 (not_new_n598__10, new_n598_);
  not g_21993 (not_pi151, pi151);
  not g_21994 (not_new_n588_, new_n588_);
  not g_21995 (not_new_n4921_, new_n4921_);
  not g_21996 (not_new_n5424_, new_n5424_);
  not g_21997 (not_new_n628__70, new_n628_);
  or g_21998 (new_n958_, or_or_not_new_n1287__not_new_n1285__not_new_n2059_, not_new_n2058_);
  or g_21999 (new_n10207_, not_new_n10182_, not_new_n9915__0);
  or g_22000 (new_n2810_, not_new_n2809_, not_new_n1617_);
  not g_22001 (not_new_n4544_, new_n4544_);
  not g_22002 (not_new_n1594__70, new_n1594_);
  or g_22003 (new_n9820_, not_new_n9410_, not_new_n1065__797922662976120010);
  or g_22004 (new_n9387_, not_new_n1049__332329305696010, not_new_n648__797922662976120010);
  or g_22005 (new_n6411_, not_new_n6375_, not_new_n6307_);
  or g_22006 (po250, not_new_n3686_, not_new_n3687_);
  not g_22007 (not_new_n3020_, new_n3020_);
  or g_22008 (or_not_new_n3965__not_new_n3966_, not_new_n3966_, not_new_n3965_);
  not g_22009 (not_new_n4455_, new_n4455_);
  not g_22010 (not_new_n3177_, new_n3177_);
  not g_22011 (not_new_n6769_, new_n6769_);
  not g_22012 (not_new_n9946__0, new_n9946_);
  or g_22013 (new_n10176_, new_n642_, new_n1035_);
  or g_22014 (new_n9441_, not_new_n9790_, not_new_n9789_);
  not g_22015 (not_new_n6635_, new_n6635_);
  and g_22016 (new_n1341_, new_n2324_, new_n1609_);
  not g_22017 (new_n7940_, new_n7759_);
  or g_22018 (or_not_new_n2903__not_new_n1483_, not_new_n2903_, not_new_n1483_);
  or g_22019 (new_n3195_, not_new_n631__7, not_new_n589__3);
  or g_22020 (new_n4632_, not_pi164_3, not_new_n4420__0);
  or g_22021 (po120, not_new_n3415_, not_new_n3416_);
  or g_22022 (new_n4526_, new_n1006_, pi166);
  and g_22023 (and_new_n1915__new_n1918_, new_n1915_, new_n1918_);
  not g_22024 (not_new_n6040_, new_n6040_);
  or g_22025 (or_not_new_n2872__not_new_n2871_, not_new_n2871_, not_new_n2872_);
  and g_22026 (new_n9468_, new_n9711_, new_n9619_);
  or g_22027 (new_n2912_, not_new_n2909_, not_new_n1616__57648010);
  or g_22028 (new_n735_, not_new_n3297_, not_new_n3298_);
  not g_22029 (not_new_n6964_, new_n6964_);
  or g_22030 (new_n3511_, not_new_n1613__968890104070, not_new_n2242_);
  or g_22031 (new_n9569_, not_new_n1037__47475615099430, not_new_n632__113988951853731430);
  xnor g_22032 (key_gate_62, key_62, not_new_n1669_);
  not g_22033 (not_new_n8538_, new_n8538_);
  or g_22034 (new_n9311_, not_new_n8868_, not_new_n1059__6782230728490);
  not g_22035 (not_new_n9337_, new_n9337_);
  not g_22036 (not_new_n4310_, new_n4310_);
  not g_22037 (not_new_n4117_, new_n4117_);
  not g_22038 (not_new_n4414__0, new_n4414_);
  or g_22039 (new_n5948_, not_new_n1051__10, not_new_n5760_);
  not g_22040 (new_n4235_, new_n706_);
  or g_22041 (new_n5216_, new_n1599_, new_n622_);
  not g_22042 (not_new_n5238_, new_n5238_);
  not g_22043 (not_new_n6974__168070, new_n6974_);
  not g_22044 (not_new_n9173_, new_n9173_);
  or g_22045 (new_n8393_, not_new_n638__797922662976120010, not_new_n8150__0);
  not g_22046 (not_new_n6465_, new_n6465_);
  not g_22047 (not_pi172_2, pi172);
  not g_22048 (not_new_n648__2, new_n648_);
  not g_22049 (not_new_n4765__0, new_n4765_);
  or g_22050 (new_n5383_, not_new_n5381_, not_new_n5218__0);
  and g_22051 (new_n5853_, new_n6013_, new_n6014_);
  not g_22052 (not_new_n1067__6782230728490, new_n1067_);
  or g_22053 (new_n2805_, not_new_n1616__7, not_new_n2802_);
  or g_22054 (new_n2693_, not_new_n4452_, not_new_n609__57648010);
  not g_22055 (not_new_n1600__7, new_n1600_);
  and g_22056 (new_n8818_, new_n9042_, new_n9039_);
  or g_22057 (new_n2053_, not_new_n586__168070, not_pi177);
  not g_22058 (new_n4259_, new_n663_);
  or g_22059 (new_n5980_, not_new_n5785_, not_new_n637__168070);
  not g_22060 (not_new_n646__57648010, new_n646_);
  or g_22061 (new_n9505_, not_new_n9586_, not_new_n9587_);
  not g_22062 (not_new_n636__3, new_n636_);
  not g_22063 (not_new_n5229_, new_n5229_);
  or g_22064 (new_n2389_, not_new_n9875__0, not_new_n599__6);
  not g_22065 (not_new_n4464_, new_n4464_);
  or g_22066 (new_n7064_, not_new_n7531_, not_new_n7530_);
  or g_22067 (new_n5953_, not_new_n5952_, not_new_n5842_);
  not g_22068 (not_new_n587__138412872010, new_n587_);
  or g_22069 (new_n10343_, not_new_n1063__16284135979104490, not_new_n9918__0);
  or g_22070 (new_n8772_, not_new_n8645__0, not_new_n1602__19773267430);
  not g_22071 (not_new_n1631__797922662976120010, key_gate_76);
  not g_22072 (not_new_n647__7, new_n647_);
  not g_22073 (not_new_n5631_, new_n5631_);
  or g_22074 (new_n7288_, not_new_n6993__0, not_new_n7222_);
  not g_22075 (new_n8149_, new_n1065_);
  not g_22076 (new_n7741_, new_n1607_);
  or g_22077 (new_n10029_, not_new_n10227_, not_new_n9988_);
  not g_22078 (not_new_n9845_, new_n9845_);
  not g_22079 (not_new_n8984__0, new_n8984_);
  not g_22080 (not_new_n1049_, new_n1049_);
  not g_22081 (not_new_n616_, new_n616_);
  not g_22082 (not_new_n1529_, new_n1529_);
  or g_22083 (new_n3668_, not_new_n989__6, not_pi220);
  not g_22084 (not_new_n619__6, new_n619_);
  not g_22085 (not_new_n1063__24010, new_n1063_);
  or g_22086 (new_n2196_, not_new_n1580__138412872010, not_new_n6565_);
  not g_22087 (not_new_n4951__0, new_n4951_);
  or g_22088 (new_n6544_, not_new_n6791_, not_new_n6731_);
  not g_22089 (not_new_n5083__0, new_n5083_);
  not g_22090 (not_new_n5868_, new_n5868_);
  or g_22091 (new_n5161_, new_n643_, new_n1061_);
  not g_22092 (not_new_n1607__3430, new_n1607_);
  or g_22093 (new_n5527_, not_new_n5630_, not_new_n1008__5);
  not g_22094 (new_n9383_, new_n1602_);
  not g_22095 (not_new_n644__19773267430, new_n644_);
  or g_22096 (new_n10160_, not_new_n10156_, not_new_n10034_);
  not g_22097 (not_new_n3799_, new_n3799_);
  or g_22098 (new_n8095_, not_new_n8395_, not_new_n8398_);
  not g_22099 (not_new_n4898_, new_n4898_);
  not g_22100 (new_n3983_, pi060);
  not g_22101 (not_new_n6290_, new_n6290_);
  or g_22102 (new_n7619_, not_new_n7614_, not_new_n7808_);
  and g_22103 (new_n8087_, new_n8368_, new_n8081_);
  or g_22104 (new_n7335_, not_new_n736__1, not_new_n7334_);
  and g_22105 (new_n5023_, new_n1037_, new_n632_);
  not g_22106 (not_pi033_4, pi033);
  not g_22107 (not_new_n1011__4, new_n1011_);
  and g_22108 (new_n8237_, new_n8397_, new_n8080_);
  not g_22109 (not_new_n4964_, new_n4964_);
  not g_22110 (not_new_n7360_, new_n7360_);
  or g_22111 (new_n1834_, not_new_n1581__2, not_new_n8099_);
  or g_22112 (new_n7500_, not_new_n7007__1, not_new_n7038__1);
  not g_22113 (not_new_n7932__0, new_n7932_);
  not g_22114 (not_new_n2345__0, new_n2345_);
  xor g_22115 (key_gate_19, not_new_n3931_, key_19);
  or g_22116 (new_n4574_, new_n1012_, pi178);
  or g_22117 (or_not_new_n4843__not_new_n4757_, not_new_n4757_, not_new_n4843_);
  not g_22118 (not_new_n5285_, new_n5285_);
  not g_22119 (not_new_n5803__0, new_n5803_);
  not g_22120 (not_new_n1534__0, key_gate_5);
  not g_22121 (not_new_n4723__0, new_n4723_);
  not g_22122 (not_new_n6337_, new_n6337_);
  or g_22123 (new_n9094_, not_new_n9093_, not_new_n8888_);
  not g_22124 (not_pi162_1, pi162);
  or g_22125 (new_n3326_, not_pi064_4, not_new_n3934__0);
  not g_22126 (new_n5059_, new_n1607_);
  or g_22127 (new_n4187_, not_new_n4071__3, not_pi257_5);
  or g_22128 (new_n7875_, not_new_n7855_, not_new_n7750_);
  not g_22129 (not_new_n7240_, new_n7240_);
  or g_22130 (new_n9195_, not_new_n9154_, not_new_n8844__0);
  not g_22131 (not_new_n7056_, new_n7056_);
  not g_22132 (not_pi106_0, pi106);
  not g_22133 (not_new_n8564_, new_n8564_);
  or g_22134 (new_n1683_, not_pi015, not_po296_1176490);
  and g_22135 (new_n1555_, new_n3623_, new_n3622_);
  and g_22136 (new_n4314_, new_n4391_, new_n4392_);
  not g_22137 (new_n9602_, new_n9501_);
  or g_22138 (new_n7326_, not_new_n7178_, not_new_n7115_);
  or g_22139 (new_n7541_, not_new_n731__1, not_new_n7421__1);
  not g_22140 (not_new_n3413_, new_n3413_);
  and g_22141 (new_n8218_, new_n8379_, new_n8378_);
  or g_22142 (new_n8590_, not_new_n8274_, not_new_n8443__0);
  not g_22143 (not_new_n4427_, new_n4427_);
  not g_22144 (not_new_n1595__0, new_n1595_);
  not g_22145 (not_new_n1612__47475615099430, new_n1612_);
  or g_22146 (new_n5371_, not_new_n1603__9, not_new_n4980_);
  not g_22147 (not_new_n617__6782230728490, new_n617_);
  not g_22148 (new_n6054_, new_n5810_);
  or g_22149 (new_n3109_, not_new_n581__225393402906922580878632490, not_new_n628__6);
  or g_22150 (new_n1860_, not_new_n4725_, not_new_n591__4);
  not g_22151 (new_n4244_, new_n703_);
  not g_22152 (not_new_n624__4, new_n624_);
  not g_22153 (not_new_n587__57648010, new_n587_);
  not g_22154 (not_new_n9967_, new_n9967_);
  or g_22155 (new_n9188_, or_not_new_n8941__not_new_n8811_, not_new_n9186__0);
  or g_22156 (new_n762_, not_new_n3234_, not_new_n3235_);
  or g_22157 (new_n3644_, not_new_n984__332329305696010, not_pi188_0);
  or g_22158 (new_n1149_, not_new_n3828_, not_new_n3827_);
  not g_22159 (not_new_n6840_, new_n6840_);
  not g_22160 (not_pi065_0, pi065);
  not g_22161 (not_pi249_1, pi249);
  not g_22162 (not_new_n8321_, new_n8321_);
  or g_22163 (new_n2754_, not_new_n604__2, not_new_n633__2);
  not g_22164 (not_new_n775__168070, new_n775_);
  not g_22165 (not_new_n1603__2, new_n1603_);
  not g_22166 (not_new_n643__1, new_n643_);
  not g_22167 (not_new_n6896_, new_n6896_);
  or g_22168 (new_n3602_, not_new_n984__5, not_pi167_0);
  not g_22169 (not_new_n1728__57648010, new_n1728_);
  not g_22170 (not_pi165_2, pi165);
  not g_22171 (not_new_n631__3430, new_n631_);
  or g_22172 (new_n6876_, not_new_n1597__1176490, not_new_n6539__2);
  not g_22173 (not_new_n4994__0, new_n4994_);
  or g_22174 (or_not_new_n6817__not_new_n6788_, not_new_n6817_, not_new_n6788_);
  or g_22175 (new_n4703_, not_pi172_2, not_new_n4436_);
  not g_22176 (not_new_n1027_, new_n1027_);
  and g_22177 (po093, key_gate_101, pi072);
  not g_22178 (not_new_n643__797922662976120010, new_n643_);
  not g_22179 (not_new_n601__403536070, new_n601_);
  not g_22180 (not_new_n4680_, new_n4680_);
  or g_22181 (new_n9234_, not_new_n9233_, not_new_n9232_);
  or g_22182 (new_n5071_, not_new_n1031__70, not_new_n641__70);
  not g_22183 (not_new_n1057__490, new_n1057_);
  and g_22184 (new_n1424_, new_n2549_, new_n2548_);
  or g_22185 (new_n4396_, not_new_n4393_, not_new_n4315_);
  or g_22186 (new_n2479_, not_new_n599__6782230728490, not_new_n9963__0);
  not g_22187 (not_new_n604_, new_n604_);
  or g_22188 (new_n3002_, not_new_n1043__2, not_new_n581__4);
  not g_22189 (new_n5928_, new_n5763_);
  or g_22190 (or_not_new_n1255__not_new_n1253_, not_new_n1255_, not_new_n1253_);
  not g_22191 (not_new_n6555_, new_n6555_);
  or g_22192 (new_n1863_, not_new_n586__5, not_pi167);
  or g_22193 (new_n3542_, not_pi137_0, not_new_n1538__7);
  not g_22194 (new_n7641_, new_n1067_);
  buf g_22195 (po030, pi234);
  not g_22196 (not_pi173_3, pi173);
  not g_22197 (not_new_n691_, new_n691_);
  or g_22198 (new_n7527_, not_new_n7430__2, not_new_n729__0);
  not g_22199 (not_new_n6541__0, new_n6541_);
  and g_22200 (new_n5718_, new_n5893_, new_n5997_);
  xor g_22201 (key_gate_77, key_77, new_n924_);
  not g_22202 (not_new_n5447__0, new_n5447_);
  not g_22203 (not_new_n8528_, new_n8528_);
  not g_22204 (not_new_n1053__16284135979104490, new_n1053_);
  not g_22205 (not_new_n5807__1, new_n5807_);
  not g_22206 (new_n7612_, new_n631_);
  or g_22207 (new_n9793_, not_new_n9383__0, not_new_n625__13410686196639649008070);
  not g_22208 (not_new_n3310__3, new_n3310_);
  not g_22209 (not_new_n4166_, new_n4166_);
  and g_22210 (new_n6452_, and_new_n6673__new_n6668_, new_n6655_);
  not g_22211 (not_new_n633__6, new_n633_);
  not g_22212 (new_n9533_, new_n9365_);
  or g_22213 (new_n8048_, not_new_n1065__19773267430, not_new_n7655__2);
  or g_22214 (new_n8296_, not_new_n8113__0, not_new_n8112_);
  not g_22215 (not_new_n1051__2, new_n1051_);
  not g_22216 (new_n7627_, new_n630_);
  or g_22217 (new_n9432_, not_new_n9728_, not_new_n9729_);
  and g_22218 (new_n4308_, new_n4374_, new_n4373_);
  not g_22219 (not_new_n5456_, new_n5456_);
  or g_22220 (or_or_not_new_n2785__not_new_n2788__not_new_n2787_, or_not_new_n2785__not_new_n2788_, not_new_n2787_);
  or g_22221 (new_n2957_, not_new_n2954_, not_new_n1616__968890104070);
  or g_22222 (new_n7172_, not_new_n7354_, not_new_n6982_);
  or g_22223 (new_n3473_, not_new_n1015__1, not_new_n1594__3430);
  not g_22224 (not_new_n6923_, new_n6923_);
  not g_22225 (not_new_n6636_, new_n6636_);
  and g_22226 (new_n613_, new_n590_, new_n2739_);
  not g_22227 (not_new_n1601__138412872010, new_n1601_);
  not g_22228 (not_new_n2861_, new_n2861_);
  or g_22229 (new_n7564_, not_new_n7204_, not_new_n7562_);
  not g_22230 (not_new_n4824_, new_n4824_);
  not g_22231 (not_new_n1300_, new_n1300_);
  not g_22232 (not_new_n585__968890104070, new_n585_);
  not g_22233 (not_new_n8086_, new_n8086_);
  or g_22234 (new_n8477_, not_new_n8126__0, not_new_n8330_);
  not g_22235 (not_new_n588__2824752490, new_n588_);
  and g_22236 (and_new_n3055__new_n998_, new_n3055_, new_n998_);
  not g_22237 (not_new_n3240_, new_n3240_);
  not g_22238 (not_new_n3121_, new_n3121_);
  not g_22239 (not_new_n9201_, new_n9201_);
  or g_22240 (new_n1866_, not_new_n585__5, not_new_n4116_);
  or g_22241 (new_n2309_, not_new_n1581__2326305139872070, not_new_n8180_);
  or g_22242 (new_n5486_, not_new_n5672_, not_new_n5671_);
  not g_22243 (not_new_n624__2, new_n624_);
  or g_22244 (new_n10034_, not_new_n1599__6782230728490, not_new_n622__16284135979104490);
  not g_22245 (not_new_n1041__138412872010, new_n1041_);
  and g_22246 (new_n6972_, new_n7198_, new_n7201_);
  not g_22247 (not_new_n3398_, new_n3398_);
  and g_22248 (and_new_n2394__new_n2393_, new_n2393_, new_n2394_);
  not g_22249 (not_new_n3425_, new_n3425_);
  or g_22250 (new_n652_, or_not_new_n3116__not_new_n3115_, not_new_n3114_);
  or g_22251 (new_n6838_, not_new_n6478__0, not_new_n634__2824752490);
  not g_22252 (not_new_n1537__47475615099430, new_n1537_);
  not g_22253 (not_new_n1257_, new_n1257_);
  or g_22254 (new_n2460_, not_new_n1603__0, not_new_n598__2824752490);
  not g_22255 (not_new_n9968__0, new_n9968_);
  not g_22256 (not_pi058_1, pi058);
  not g_22257 (not_new_n8289__0, new_n8289_);
  not g_22258 (not_new_n726_, new_n726_);
  or g_22259 (new_n1927_, not_new_n1585__7, not_new_n5736_);
  not g_22260 (not_new_n6850_, new_n6850_);
  not g_22261 (not_new_n612__4, new_n612_);
  or g_22262 (new_n3065_, not_new_n1061__2, not_new_n581__47475615099430);
  not g_22263 (not_new_n1071__2824752490, new_n1071_);
  or g_22264 (new_n1651_, key_gate_86, not_new_n596__5);
  or g_22265 (new_n10172_, not_new_n9998_, not_new_n10171_);
  not g_22266 (not_new_n984__138412872010, new_n984_);
  not g_22267 (not_new_n631__4599865365447399609768010, new_n631_);
  not g_22268 (not_new_n3185__3430, new_n3185_);
  not g_22269 (not_new_n6054_, new_n6054_);
  and g_22270 (new_n5055_, new_n5252_, new_n4901_);
  or g_22271 (new_n6907_, not_new_n1604__168070, not_new_n6510__0);
  or g_22272 (new_n5197_, new_n1599_, new_n622_);
  not g_22273 (not_new_n3103_, new_n3103_);
  not g_22274 (not_new_n4413_, new_n4413_);
  or g_22275 (new_n9652_, not_new_n9651_, not_new_n9426__0);
  not g_22276 (new_n4172_, new_n4106_);
  not g_22277 (not_new_n6021_, new_n6021_);
  or g_22278 (new_n3502_, not_pi117_0, not_new_n1537__403536070);
  not g_22279 (not_new_n5775_, new_n5775_);
  not g_22280 (not_new_n7450_, new_n7450_);
  not g_22281 (not_new_n1585__5, new_n1585_);
  not g_22282 (not_new_n2575_, new_n2575_);
  not g_22283 (not_new_n4754_, new_n4754_);
  not g_22284 (not_new_n9072_, new_n9072_);
  not g_22285 (not_new_n1160__0, new_n1160_);
  not g_22286 (not_new_n1589__2326305139872070, new_n1589_);
  or g_22287 (new_n9128_, not_new_n9126_, not_new_n8949_);
  not g_22288 (not_new_n628__13410686196639649008070, new_n628_);
  or g_22289 (or_not_new_n1561__not_new_n2464_, not_new_n1561_, not_new_n2464_);
  or g_22290 (new_n1015_, not_new_n3351_, not_new_n3352_);
  not g_22291 (not_new_n9587__0, new_n9587_);
  not g_22292 (not_new_n1035__7, new_n1035_);
  or g_22293 (new_n1932_, not_new_n1589__7, not_new_n5004_);
  and g_22294 (po100, pi079, key_gate_101);
  or g_22295 (new_n5545_, not_new_n5597_, not_new_n1003__5);
  not g_22296 (not_new_n3230_, new_n3230_);
  not g_22297 (not_pi252_1, pi252);
  not g_22298 (not_po298_1, po298);
  or g_22299 (new_n718_, not_new_n3261_, not_new_n3262_);
  not g_22300 (not_new_n8639_, new_n8639_);
  not g_22301 (not_new_n6443_, new_n6443_);
  not g_22302 (new_n3369_, new_n1022_);
  or g_22303 (new_n6765_, not_new_n6546_, not_new_n6651_);
  not g_22304 (not_new_n7841_, new_n7841_);
  or g_22305 (new_n4810_, not_new_n4749__0, not_new_n4818__0);
  not g_22306 (new_n4091_, pi261);
  or g_22307 (or_or_not_new_n2034__not_new_n2035__not_new_n2037_, or_not_new_n2034__not_new_n2035_, not_new_n2037_);
  not g_22308 (not_new_n8737_, new_n8737_);
  or g_22309 (new_n4586_, not_new_n4645_, not_new_n4416__0);
  or g_22310 (new_n9741_, not_new_n9739_, not_new_n9740_);
  or g_22311 (new_n1156_, not_new_n3842_, not_new_n3841_);
  and g_22312 (new_n8666_, new_n8757_, new_n8665_);
  and g_22313 (new_n5881_, new_n6112_, new_n6111_);
  not g_22314 (not_new_n598__4, new_n598_);
  not g_22315 (not_new_n4148_, new_n4148_);
  or g_22316 (new_n2608_, not_new_n4453__0, not_new_n610__9);
  not g_22317 (not_new_n7366__0, new_n7366_);
  not g_22318 (not_new_n9599_, new_n9599_);
  or g_22319 (new_n8778_, not_new_n1600__2824752490, not_new_n8599_);
  not g_22320 (new_n3372_, new_n1023_);
  and g_22321 (new_n5908_, new_n6220_, new_n6219_);
  not g_22322 (not_new_n5447__1, new_n5447_);
  not g_22323 (not_pi048_3, pi048);
  not g_22324 (not_pi135_0, pi135);
  not g_22325 (not_new_n8873_, new_n8873_);
  not g_22326 (not_new_n1583__8235430, new_n1583_);
  and g_22327 (and_and_new_n8692__new_n8691__new_n8695_, new_n8695_, and_new_n8692__new_n8691_);
  or g_22328 (new_n2685_, not_new_n605__8235430, not_new_n5427_);
  not g_22329 (not_new_n951_, new_n951_);
  not g_22330 (not_new_n3239_, new_n3239_);
  not g_22331 (new_n5461_, pi142);
  or g_22332 (new_n2269_, not_new_n5831_, not_new_n1585__47475615099430);
  not g_22333 (not_new_n657_, new_n657_);
  or g_22334 (new_n10062_, new_n1051_, new_n647_);
  not g_22335 (not_new_n5484_, new_n5484_);
  not g_22336 (not_new_n7763_, new_n7763_);
  not g_22337 (not_new_n9312_, new_n9312_);
  not g_22338 (not_new_n10303_, new_n10303_);
  not g_22339 (not_new_n8004_, new_n8004_);
  or g_22340 (new_n1795_, not_new_n9429_, not_new_n1584__0);
  not g_22341 (not_new_n1601__6782230728490, new_n1601_);
  and g_22342 (new_n1360_, new_n2385_, new_n2386_);
  not g_22343 (not_new_n591__113988951853731430, new_n591_);
  not g_22344 (not_new_n10029_, new_n10029_);
  not g_22345 (not_new_n3333_, new_n3333_);
  not g_22346 (not_new_n1616__3430, new_n1616_);
  and g_22347 (new_n1324_, new_n2240_, and_and_new_n2238__new_n2241__new_n2239_);
  or g_22348 (new_n3811_, not_new_n1810_, not_new_n3419_);
  not g_22349 (new_n9939_, new_n629_);
  not g_22350 (not_new_n604__2, new_n604_);
  not g_22351 (not_new_n1600__24010, new_n1600_);
  not g_22352 (not_new_n1584__10, new_n1584_);
  not g_22353 (new_n7360_, new_n7022_);
  or g_22354 (new_n7987_, or_not_new_n1596__403536070_not_new_n7586_, not_new_n7665__0);
  not g_22355 (not_new_n1362_, new_n1362_);
  not g_22356 (not_new_n10342_, new_n10342_);
  not g_22357 (not_new_n8337_, new_n8337_);
  not g_22358 (not_pi056_0, pi056);
  or g_22359 (new_n2765_, not_new_n994__5, not_pi250_2);
  or g_22360 (new_n7802_, not_new_n7801_, not_new_n7652__0);
  not g_22361 (not_new_n4579_, new_n4579_);
  not g_22362 (new_n10104_, new_n10028_);
  not g_22363 (not_new_n1589__1, new_n1589_);
  not g_22364 (not_pi039_2, pi039);
  not g_22365 (not_new_n5221_, new_n5221_);
  not g_22366 (not_new_n1009__7, new_n1009_);
  or g_22367 (new_n7677_, not_new_n8026_, not_new_n8027_);
  not g_22368 (not_new_n8529_, new_n8529_);
  not g_22369 (not_new_n3281_, new_n3281_);
  or g_22370 (new_n10229_, not_new_n9915__1, not_new_n10110_);
  not g_22371 (not_new_n5776__0, new_n5776_);
  or g_22372 (new_n9598_, not_new_n9413_, not_new_n9412_);
  not g_22373 (not_new_n9367_, new_n9367_);
  not g_22374 (not_new_n9285_, new_n9285_);
  not g_22375 (not_new_n7570_, new_n7570_);
  or g_22376 (new_n10175_, not_new_n9999_, not_new_n10173_);
  not g_22377 (not_new_n9950__0, new_n9950_);
  and g_22378 (new_n6459_, new_n6458_, new_n6456_);
  not g_22379 (not_new_n5791__0, new_n5791_);
  not g_22380 (not_new_n8149_, new_n8149_);
  and g_22381 (new_n4725_, new_n4822_, new_n4730_);
  and g_22382 (and_new_n5097__new_n5098_, new_n5097_, new_n5098_);
  not g_22383 (not_new_n7820_, new_n7820_);
  buf g_22384 (po053, pi277);
  and g_22385 (and_new_n1541__new_n2366_, new_n1541_, new_n2366_);
  not g_22386 (not_new_n3338_, new_n3338_);
  not g_22387 (not_new_n2621_, new_n2621_);
  not g_22388 (not_new_n5871_, new_n5871_);
  or g_22389 (new_n1839_, not_new_n594__2, not_new_n9959_);
  or g_22390 (or_not_new_n1279__not_new_n1277_, not_new_n1277_, not_new_n1279_);
  or g_22391 (new_n8961_, not_new_n8980_, or_not_new_n9166__not_new_n9106_);
  not g_22392 (not_new_n6822_, new_n6822_);
  not g_22393 (not_new_n608__7, new_n608_);
  or g_22394 (new_n2644_, not_new_n607__70, not_new_n1006_);
  not g_22395 (not_new_n6351_, new_n6351_);
  not g_22396 (not_new_n1375_, new_n1375_);
  not g_22397 (not_pi043_0, pi043);
  and g_22398 (new_n5716_, new_n5916_, new_n5979_);
  or g_22399 (new_n5263_, not_new_n5238_, not_new_n4984__1);
  not g_22400 (not_new_n9261_, new_n9261_);
  not g_22401 (not_new_n7521_, new_n7521_);
  and g_22402 (new_n1230_, new_n1796_, new_n1797_);
  not g_22403 (not_new_n4700_, new_n4700_);
  not g_22404 (not_new_n6064_, new_n6064_);
  not g_22405 (not_new_n5678_, new_n5678_);
  not g_22406 (not_new_n9107_, new_n9107_);
  or g_22407 (new_n5061_, or_not_new_n5266__not_new_n5206_, not_new_n5080_);
  or g_22408 (new_n1887_, not_new_n601__4, not_new_n631__0);
  not g_22409 (not_new_n623__6, new_n623_);
  xnor g_22410 (key_gate_29, key_29, not_new_n3998_);
  not g_22411 (not_new_n9464_, new_n9464_);
  not g_22412 (not_new_n3504_, new_n3504_);
  not g_22413 (not_new_n3545_, new_n3545_);
  or g_22414 (new_n7264_, not_new_n7045_, not_new_n718_);
  not g_22415 (not_pi043, pi043);
  not g_22416 (not_new_n9437_, new_n9437_);
  or g_22417 (new_n3740_, not_new_n645__10, not_new_n1071__6);
  not g_22418 (not_new_n5800__0, new_n5800_);
  or g_22419 (new_n3533_, not_new_n1843__0, not_new_n1612__2);
  not g_22420 (not_pi060_1, pi060);
  not g_22421 (not_new_n9022_, new_n9022_);
  or g_22422 (new_n2689_, not_po296_9095436801298611408202050198891430, not_pi265_1);
  not g_22423 (not_new_n4899__0, new_n4899_);
  not g_22424 (not_new_n5693_, new_n5693_);
  not g_22425 (not_new_n1017__0, new_n1017_);
  or g_22426 (new_n3608_, not_pi170_0, not_new_n984__8);
  not g_22427 (not_new_n8991_, new_n8991_);
  not g_22428 (not_new_n3532_, new_n3532_);
  not g_22429 (not_new_n618__8235430, new_n618_);
  not g_22430 (not_new_n6492_, new_n6492_);
  not g_22431 (not_new_n3265_, new_n3265_);
  not g_22432 (not_new_n1027__5, new_n1027_);
  or g_22433 (new_n6836_, not_new_n6835_, not_new_n6834_);
  or g_22434 (new_n1176_, not_new_n3882_, not_new_n3881_);
  or g_22435 (new_n2240_, not_new_n4774_, not_new_n591__6782230728490);
  not g_22436 (new_n8432_, new_n8263_);
  not g_22437 (not_new_n5893__0, new_n5893_);
  not g_22438 (not_new_n1651_, key_gate_47);
  or g_22439 (new_n3517_, not_new_n2299_, not_new_n1613__332329305696010);
  not g_22440 (not_new_n3038_, new_n3038_);
  or g_22441 (new_n1732_, not_new_n1728__0, not_pi076);
  not g_22442 (new_n2038_, new_n638_);
  not g_22443 (new_n7917_, new_n7669_);
  not g_22444 (not_new_n8868_, new_n8868_);
  not g_22445 (not_new_n1527_, new_n1527_);
  or g_22446 (new_n1849_, not_new_n601__2, not_new_n628__0);
  not g_22447 (not_new_n6938_, new_n6938_);
  xor g_22448 (key_gate_60, key_60, not_new_n3957_);
  not g_22449 (not_new_n1019__2, new_n1019_);
  and g_22450 (new_n1344_, new_n2324_, new_n1609_);
  not g_22451 (not_new_n1204_, new_n1204_);
  not g_22452 (not_new_n618__5585458640832840070, new_n618_);
  not g_22453 (not_new_n7285_, new_n7285_);
  not g_22454 (not_new_n676_, new_n676_);
  or g_22455 (new_n5162_, not_new_n1061__10, not_new_n643__168070);
  or g_22456 (new_n9772_, not_new_n621__797922662976120010, not_new_n9379__0);
  and g_22457 (new_n5849_, new_n5724_, new_n5989_);
  and g_22458 (new_n6585_, new_n6743_, new_n6797_);
  or g_22459 (new_n7494_, not_new_n7445__1, not_new_n723__1);
  not g_22460 (not_new_n8118__1, new_n8118_);
  or g_22461 (new_n6692_, not_new_n6475__0, not_new_n631__19773267430);
  or g_22462 (new_n10256_, not_new_n1041__47475615099430, not_new_n9886_);
  not g_22463 (not_new_n3479_, new_n3479_);
  or g_22464 (new_n9280_, not_new_n1071__19773267430, not_new_n8873_);
  not g_22465 (not_new_n586__138412872010, new_n586_);
  or g_22466 (new_n656_, not_new_n3126_, or_not_new_n3128__not_new_n3127_);
  not g_22467 (not_new_n5905__0, new_n5905_);
  not g_22468 (not_new_n8147__0, new_n8147_);
  not g_22469 (not_new_n597__8235430, new_n597_);
  not g_22470 (not_new_n608__2, new_n608_);
  not g_22471 (new_n9934_, new_n1601_);
  and g_22472 (new_n10019_, new_n10308_, new_n10307_);
  or g_22473 (new_n4457_, not_new_n4620_, not_new_n4621_);
  not g_22474 (not_new_n645__57648010, new_n645_);
  not g_22475 (not_new_n1601__968890104070, new_n1601_);
  or g_22476 (new_n3786_, not_new_n3785_, not_new_n3784_);
  not g_22477 (not_new_n587__6, new_n587_);
  not g_22478 (not_new_n6525__0, new_n6525_);
  or g_22479 (new_n5878_, not_new_n5841_, not_new_n6044_);
  and g_22480 (and_and_new_n1839__new_n1842__new_n1840_, and_new_n1839__new_n1842_, new_n1840_);
  or g_22481 (new_n7590_, not_new_n7873_, not_new_n7871_);
  not g_22482 (not_new_n9249_, new_n9249_);
  not g_22483 (not_new_n6043_, new_n6043_);
  not g_22484 (not_new_n7709_, new_n7709_);
  not g_22485 (new_n8136_, new_n639_);
  not g_22486 (not_new_n5351_, new_n5351_);
  and g_22487 (new_n1401_, new_n2488_, new_n2487_);
  or g_22488 (new_n5541_, new_n1004_, pi136);
  not g_22489 (not_new_n10067_, new_n10067_);
  not g_22490 (not_new_n6510__0, new_n6510_);
  not g_22491 (not_new_n609__168070, new_n609_);
  not g_22492 (not_new_n2656_, new_n2656_);
  not g_22493 (not_new_n6600_, new_n6600_);
  not g_22494 (not_new_n3302_, new_n3302_);
  or g_22495 (new_n3371_, not_pi064_47475615099430, not_new_n3924__0);
  not g_22496 (not_new_n5900__1, new_n5900_);
  not g_22497 (not_new_n8211_, new_n8211_);
  not g_22498 (new_n4154_, new_n4145_);
  or g_22499 (new_n9152_, not_new_n1053__138412872010, not_new_n626__13410686196639649008070);
  or g_22500 (new_n1792_, not_new_n641__0, not_new_n601_);
  not g_22501 (not_new_n4687_, new_n4687_);
  or g_22502 (new_n5239_, not_new_n5156_, not_new_n5078__0);
  not g_22503 (not_new_n8973__0, new_n8973_);
  not g_22504 (not_new_n10114_, new_n10114_);
  not g_22505 (not_new_n1580__168070, new_n1580_);
  or g_22506 (new_n1972_, not_new_n9867_, not_new_n594__9);
  not g_22507 (new_n8040_, new_n7726_);
  not g_22508 (not_new_n5780_, new_n5780_);
  not g_22509 (not_new_n970_, new_n970_);
  not g_22510 (not_new_n4461_, new_n4461_);
  not g_22511 (not_pi154_0, pi154);
  not g_22512 (not_pi034_0, pi034);
  or g_22513 (new_n6997_, not_new_n734_, not_new_n7032_);
  or g_22514 (new_n7569_, not_new_n7097_, not_new_n7348_);
  not g_22515 (not_new_n607__490, new_n607_);
  not g_22516 (not_new_n8496_, new_n8496_);
  not g_22517 (not_new_n1925_, new_n1925_);
  or g_22518 (new_n8500_, not_new_n618__16284135979104490, not_new_n8171__1);
  or g_22519 (new_n3163_, not_new_n581__367033682172941254412302110320336601888010, not_new_n644__6);
  and g_22520 (new_n6315_, new_n6393_, new_n6383_);
  or g_22521 (new_n7818_, not_new_n7791__0, not_new_n7614__0);
  or g_22522 (new_n5236_, not_new_n633__24010, not_new_n1067__9);
  and g_22523 (new_n7729_, new_n8050_, new_n7769_);
  not g_22524 (not_new_n1061__3430, new_n1061_);
  or g_22525 (new_n7284_, not_new_n7439__1, not_new_n7004__1);
  not g_22526 (not_new_n621__16284135979104490, new_n621_);
  or g_22527 (new_n8398_, not_new_n8237_, not_new_n8396_);
  not g_22528 (not_new_n625__39098210485829880490, new_n625_);
  not g_22529 (not_new_n8743_, new_n8743_);
  and g_22530 (new_n1528_, new_n3083_, and_new_n3085__new_n998_);
  or g_22531 (new_n7432_, not_new_n6974__57648010, not_new_n756_);
  not g_22532 (not_new_n2527_, new_n2527_);
  not g_22533 (not_new_n3026_, new_n3026_);
  or g_22534 (new_n9822_, not_new_n9427__3, not_new_n9691_);
  or g_22535 (new_n9542_, new_n1051_, new_n647_);
  or g_22536 (new_n6418_, not_new_n6236_, or_or_or_not_new_n1055__168070_not_new_n6325__not_new_n6373__1_not_new_n6317_);
  not g_22537 (new_n4961_, new_n626_);
  not g_22538 (not_new_n928__168070, new_n928_);
  or g_22539 (or_or_not_new_n1782__not_new_n1783__not_new_n1785_, not_new_n1785_, or_not_new_n1782__not_new_n1783_);
  not g_22540 (not_new_n1596__403536070, new_n1596_);
  and g_22541 (new_n7094_, new_n7289_, new_n6963_);
  or g_22542 (new_n9776_, not_new_n9774_, not_new_n9775_);
  not g_22543 (not_new_n1599__7, new_n1599_);
  not g_22544 (not_new_n5767_, new_n5767_);
  not g_22545 (not_new_n665_, new_n665_);
  not g_22546 (not_new_n3000_, new_n3000_);
  not g_22547 (not_new_n6103_, new_n6103_);
  not g_22548 (not_new_n7361_, new_n7361_);
  or g_22549 (new_n2642_, not_new_n2509__490, not_pi206);
  not g_22550 (new_n4950_, new_n621_);
  or g_22551 (new_n5319_, not_new_n5057_, not_new_n5258_);
  not g_22552 (not_new_n2322_, new_n2322_);
  not g_22553 (not_new_n1598__9, new_n1598_);
  not g_22554 (not_new_n5385_, new_n5385_);
  not g_22555 (not_new_n647__8, new_n647_);
  and g_22556 (new_n6964_, new_n7235_, new_n7236_);
  not g_22557 (not_new_n9372__0, new_n9372_);
  and g_22558 (and_new_n1266__new_n1970_, new_n1970_, new_n1266_);
  not g_22559 (not_new_n7627__1, new_n7627_);
  not g_22560 (not_new_n2571_, new_n2571_);
  not g_22561 (not_new_n5099_, new_n5099_);
  or g_22562 (new_n5078_, not_new_n5271_, not_new_n5036_);
  not g_22563 (not_new_n644__5585458640832840070, new_n644_);
  not g_22564 (not_new_n6077_, new_n6077_);
  not g_22565 (not_new_n5092__0, new_n5092_);
  or g_22566 (new_n3308_, not_new_n994__797922662976120010, not_new_n1619_);
  and g_22567 (new_n8696_, and_and_new_n8692__new_n8691__new_n8695_, new_n8792_);
  and g_22568 (and_new_n4403__new_n4407_, new_n4403_, new_n4407_);
  not g_22569 (not_new_n601__490, new_n601_);
  not g_22570 (not_new_n8165__0, new_n8165_);
  and g_22571 (new_n9856_, new_n10053_, new_n10054_);
  or g_22572 (new_n2762_, not_pi249_0, not_po296_152867006319425761937651857692768264010);
  not g_22573 (not_new_n6321_, new_n6321_);
  not g_22574 (not_new_n1012__3, new_n1012_);
  or g_22575 (new_n1978_, not_pi141, not_new_n587__70);
  not g_22576 (not_new_n4417_, new_n4417_);
  or g_22577 (new_n3299_, not_new_n589__1070069044235980333563563003849377848070, not_new_n1035__5);
  not g_22578 (not_new_n4724__0, new_n4724_);
  or g_22579 (new_n617_, or_or_not_new_n2265__not_new_n2262__not_new_n2263_, not_new_n2264_);
  or g_22580 (new_n5490_, not_new_n5697_, not_new_n5696_);
  not g_22581 (new_n8838_, new_n1047_);
  not g_22582 (not_new_n9787_, new_n9787_);
  not g_22583 (not_new_n714_, new_n714_);
  buf g_22584 (po031, pi233);
  not g_22585 (not_new_n1534__24010, key_gate_5);
  not g_22586 (not_new_n5373_, new_n5373_);
  not g_22587 (not_new_n5554_, new_n5554_);
  not g_22588 (not_new_n648__8235430, new_n648_);
  or g_22589 (new_n9144_, not_new_n8983_, not_new_n9140_);
  or g_22590 (new_n9091_, not_new_n1602__138412872010, not_new_n625__797922662976120010);
  not g_22591 (not_new_n8523_, new_n8523_);
  or g_22592 (new_n3879_, not_new_n644__70, not_new_n6443__47475615099430);
  not g_22593 (new_n4255_, new_n665_);
  not g_22594 (not_new_n8425_, new_n8425_);
  not g_22595 (not_new_n8893_, new_n8893_);
  not g_22596 (not_new_n9357__0, new_n9357_);
  not g_22597 (not_new_n7428_, new_n7428_);
  not g_22598 (not_new_n6527__0, new_n6527_);
  or g_22599 (new_n7488_, not_new_n7041__1, not_new_n7009__1);
  not g_22600 (not_new_n5738_, new_n5738_);
  not g_22601 (not_new_n1761_, new_n1761_);
  not g_22602 (not_new_n1016_, new_n1016_);
  not g_22603 (not_new_n1063__138412872010, new_n1063_);
  xor g_22604 (key_gate_45, not_new_n3923_, key_45);
  not g_22605 (not_new_n583__0, new_n583_);
  not g_22606 (not_new_n8870__0, new_n8870_);
  or g_22607 (new_n6120_, not_new_n1037__490, not_new_n5747__0);
  or g_22608 (new_n8780_, not_new_n1599__403536070, not_new_n8709_);
  not g_22609 (new_n7454_, new_n7044_);
  or g_22610 (new_n9019_, not_new_n634__332329305696010, not_new_n1047__19773267430);
  not g_22611 (not_new_n3900_, new_n3900_);
  not g_22612 (not_new_n3754_, new_n3754_);
  and g_22613 (new_n6241_, new_n6377_, and_new_n6378__new_n6379_);
  or g_22614 (new_n5343_, not_new_n5341_, not_new_n5202_);
  or g_22615 (new_n1967_, not_new_n1581__9, not_new_n8200_);
  or g_22616 (new_n2751_, not_new_n1616__1, not_new_n2748_);
  or g_22617 (new_n9649_, not_new_n9610__0, not_new_n9647__0);
  or g_22618 (or_not_new_n9523__1_not_new_n9327__1, not_new_n9327__1, not_new_n9523__1);
  not g_22619 (not_new_n9746_, new_n9746_);
  not g_22620 (new_n6265_, new_n633_);
  not g_22621 (not_new_n8252_, new_n8252_);
  not g_22622 (not_new_n5165_, new_n5165_);
  or g_22623 (po181, not_new_n3589_, not_new_n3588_);
  xor g_22624 (key_gate_65, key_65, not_new_n3958_);
  or g_22625 (new_n1669_, not_new_n596__70, key_gate_29);
  not g_22626 (not_new_n8105__1, new_n8105_);
  not g_22627 (not_new_n1585__968890104070, new_n1585_);
  not g_22628 (not_new_n1617__0, new_n1617_);
  not g_22629 (not_new_n626__1577753820348458066150427430, new_n626_);
  or g_22630 (new_n4050_, not_new_n3976__0, not_new_n4003__0);
  not g_22631 (not_new_n3933_, new_n3933_);
  not g_22632 (not_new_n589__3430, new_n589_);
  not g_22633 (not_new_n4767_, new_n4767_);
  not g_22634 (not_new_n4782__0, new_n4782_);
  or g_22635 (or_or_not_pi269_2_not_pi248_2_not_pi257_2, not_pi257_2, or_not_pi269_2_not_pi248_2);
  and g_22636 (new_n8703_, new_n8797_, new_n8705_);
  or g_22637 (new_n5306_, not_new_n5305_, not_new_n5304_);
  not g_22638 (not_new_n1606__2, new_n1606_);
  or g_22639 (new_n7883_, not_new_n625__47475615099430, not_new_n7631__1);
  not g_22640 (not_new_n1584__168070, new_n1584_);
  not g_22641 (new_n4952_, new_n1600_);
  or g_22642 (new_n9788_, not_new_n9786_, not_new_n9787_);
  not g_22643 (not_pi117_0, pi117);
  or g_22644 (new_n3075_, not_new_n1027__5585458640832840070, not_new_n1177_);
  or g_22645 (new_n9761_, not_new_n1596__5585458640832840070, not_new_n9420__0);
  not g_22646 (not_new_n4798__0, new_n4798_);
  not g_22647 (not_new_n719__1, new_n719_);
  not g_22648 (not_new_n1728__6782230728490, new_n1728_);
  or g_22649 (new_n2934_, not_new_n602__138412872010, not_new_n624__3);
  or g_22650 (new_n3144_, not_new_n1071__3, not_new_n928__403536070);
  not g_22651 (not_new_n928__9, new_n928_);
  or g_22652 (new_n1855_, not_new_n8906_, not_new_n1591__3);
  not g_22653 (not_new_n2210_, new_n2210_);
  or g_22654 (new_n2977_, not_po296_29286449308136415160327158440136953416342323212091034008010, not_pi273);
  not g_22655 (not_new_n1006__0, new_n1006_);
  not g_22656 (not_new_n6912_, new_n6912_);
  or g_22657 (new_n5957_, not_new_n631__8235430, not_new_n5742__0);
  not g_22658 (not_new_n5741_, new_n5741_);
  not g_22659 (not_new_n6517__0, new_n6517_);
  or g_22660 (new_n9043_, new_n1051_, new_n647_);
  not g_22661 (not_new_n3858_, new_n3858_);
  not g_22662 (new_n8441_, new_n8256_);
  not g_22663 (new_n7990_, new_n7716_);
  not g_22664 (not_new_n1055__403536070, new_n1055_);
  not g_22665 (not_new_n1807_, new_n1807_);
  and g_22666 (new_n1335_, and_new_n1334__new_n2293_, new_n2292_);
  not g_22667 (not_new_n6520_, new_n6520_);
  or g_22668 (new_n7466_, not_new_n7406__1, not_new_n718__1);
  or g_22669 (new_n2510_, not_new_n4410__0, not_new_n610_);
  not g_22670 (not_new_n613_, new_n613_);
  not g_22671 (not_new_n9109_, new_n9109_);
  or g_22672 (new_n2941_, not_pi269_0, not_po296_12197604876358357001385738625629718207556152941312384010);
  or g_22673 (new_n9607_, not_new_n9606_, not_new_n1604__6782230728490);
  not g_22674 (not_pi174, pi174);
  or g_22675 (new_n5666_, not_new_n1013__6, not_new_n5468_);
  not g_22676 (not_new_n9933__0, new_n9933_);
  not g_22677 (not_new_n1069__70, new_n1069_);
  not g_22678 (not_new_n2349_, new_n2349_);
  or g_22679 (new_n9204_, not_new_n8834_, not_new_n635__47475615099430);
  and g_22680 (new_n6969_, new_n7287_, new_n7290_);
  not g_22681 (not_new_n2774_, new_n2774_);
  not g_22682 (not_new_n8874__1, new_n8874_);
  not g_22683 (not_new_n2509__3430, new_n2509_);
  not g_22684 (not_new_n597_, new_n597_);
  or g_22685 (new_n1647_, not_po296_4, not_pi027);
  or g_22686 (new_n3038_, not_new_n1027__403536070, not_new_n1165_);
  or g_22687 (new_n5231_, new_n645_, new_n1071_);
  or g_22688 (new_n6222_, not_new_n6068__0, not_new_n5908_);
  or g_22689 (new_n7908_, or_not_new_n7715__not_new_n7714_, not_new_n7863__0);
  or g_22690 (new_n10239_, not_new_n10198_, not_new_n9899__0);
  not g_22691 (not_new_n1612__3430, new_n1612_);
  not g_22692 (not_new_n642__16284135979104490, new_n642_);
  or g_22693 (new_n955_, not_new_n2001_, or_or_not_new_n1275__not_new_n1273__not_new_n2002_);
  not g_22694 (not_new_n9668_, new_n9668_);
  or g_22695 (new_n1689_, not_po296_57648010, not_pi013);
  or g_22696 (new_n2684_, not_new_n1010_, not_new_n607__168070);
  not g_22697 (not_new_n752_, new_n752_);
  and g_22698 (and_new_n6673__new_n6668_, new_n6668_, new_n6673_);
  not g_22699 (not_new_n1996_, new_n1996_);
  not g_22700 (not_new_n4114__0, new_n4114_);
  not g_22701 (not_new_n3459_, new_n3459_);
  not g_22702 (not_new_n581__6, new_n581_);
  not g_22703 (not_new_n596__3430, key_gate_88);
  not g_22704 (new_n7661_, new_n621_);
  not g_22705 (not_new_n591__403536070, new_n591_);
  not g_22706 (new_n7433_, new_n7036_);
  not g_22707 (not_pi063_0, pi063);
  not g_22708 (not_new_n2299__0, new_n2299_);
  not g_22709 (not_new_n1045__70, new_n1045_);
  not g_22710 (not_new_n7677_, new_n7677_);
  xnor g_22711 (key_gate_13, new_n1669_, key_13);
  not g_22712 (new_n7009_, new_n722_);
  not g_22713 (not_new_n9429_, new_n9429_);
  or g_22714 (new_n2343_, not_new_n591__797922662976120010, not_new_n4759_);
  not g_22715 (not_new_n1583__113988951853731430, new_n1583_);
  and g_22716 (new_n6970_, new_n7283_, new_n7280_);
  not g_22717 (not_new_n6317_, new_n6317_);
  and g_22718 (new_n8665_, new_n8719_, new_n8723_);
  not g_22719 (not_new_n4761_, new_n4761_);
  not g_22720 (not_new_n587__8235430, new_n587_);
  not g_22721 (not_new_n1601__1, new_n1601_);
  not g_22722 (not_new_n8911_, new_n8911_);
  not g_22723 (not_new_n2116_, new_n2116_);
  not g_22724 (new_n4236_, new_n705_);
  not g_22725 (not_new_n1320_, new_n1320_);
  or g_22726 (new_n6917_, not_new_n6511__0, not_new_n1071__24010);
  or g_22727 (new_n8281_, not_new_n8156_, not_new_n1053__57648010);
  not g_22728 (not_new_n1606__5, new_n1606_);
  not g_22729 (not_new_n4033_, new_n4033_);
  or g_22730 (new_n719_, not_new_n3264_, not_new_n3263_);
  not g_22731 (not_new_n7790_, new_n7790_);
  not g_22732 (not_new_n4741_, new_n4741_);
  not g_22733 (not_new_n1596__39098210485829880490, new_n1596_);
  not g_22734 (new_n5808_, new_n618_);
  not g_22735 (new_n8831_, new_n1031_);
  or g_22736 (new_n4462_, not_new_n4666_, not_new_n4665_);
  not g_22737 (new_n6084_, new_n5887_);
  not g_22738 (not_new_n9026_, new_n9026_);
  not g_22739 (new_n8613_, new_n1175_);
  not g_22740 (not_new_n9625__0, new_n9625_);
  or g_22741 (new_n6656_, not_new_n6472_, not_new_n1047__3430);
  and g_22742 (new_n9985_, new_n10086_, new_n10042_);
  not g_22743 (not_new_n1938__0, new_n1938_);
  or g_22744 (po165, not_new_n3557_, not_new_n3556_);
  not g_22745 (not_new_n8576_, new_n8576_);
  not g_22746 (not_new_n7439__1, new_n7439_);
  not g_22747 (not_new_n7640__0, new_n7640_);
  not g_22748 (not_new_n4839__1, new_n4839_);
  or g_22749 (new_n9734_, not_new_n9732_, not_new_n9733_);
  or g_22750 (new_n2101_, not_new_n6556_, not_new_n1580__8235430);
  or g_22751 (new_n6134_, not_new_n6084_, not_new_n6133_);
  or g_22752 (new_n2357_, not_new_n603__0, not_new_n632__1);
  not g_22753 (not_new_n2822_, new_n2822_);
  or g_22754 (new_n10210_, not_new_n1596__273687473400809163430, not_new_n618__4599865365447399609768010);
  not g_22755 (not_new_n4351__0, new_n4351_);
  not g_22756 (not_new_n1603__10, new_n1603_);
  not g_22757 (not_new_n8136_, new_n8136_);
  not g_22758 (not_new_n600__9, new_n600_);
  not g_22759 (not_new_n7307_, new_n7307_);
  or g_22760 (new_n7813_, not_new_n7773__0, not_new_n7619_);
  or g_22761 (new_n8396_, not_new_n8177_, not_new_n8282_);
  not g_22762 (not_new_n626__19773267430, new_n626_);
  or g_22763 (new_n9277_, not_new_n8972_, not_new_n8993_);
  not g_22764 (not_new_n4524_, new_n4524_);
  and g_22765 (new_n5038_, new_n5154_, new_n5083_);
  or g_22766 (new_n7666_, not_new_n7710_, not_new_n7931_);
  not g_22767 (new_n8250_, new_n1607_);
  or g_22768 (new_n5180_, not_new_n5179_, not_new_n4997_);
  or g_22769 (new_n8173_, not_new_n8372_, not_new_n8426_);
  not g_22770 (not_new_n4277_, new_n4277_);
  not g_22771 (not_new_n2968_, new_n2968_);
  or g_22772 (new_n3074_, not_new_n1055__2, not_new_n581__16284135979104490);
  not g_22773 (not_new_n3350_, new_n3350_);
  not g_22774 (not_new_n928__968890104070, new_n928_);
  not g_22775 (not_new_n5432__0, new_n5432_);
  not g_22776 (not_new_n6208_, new_n6208_);
  not g_22777 (not_new_n9512__1, new_n9512_);
  or g_22778 (po259, not_new_n3704_, not_new_n3705_);
  or g_22779 (new_n8979_, not_new_n9185_, not_new_n9184_);
  not g_22780 (not_new_n1037__8, new_n1037_);
  or g_22781 (new_n7804_, not_new_n7701_, not_new_n7803_);
  not g_22782 (new_n8555_, new_n8235_);
  or g_22783 (new_n8546_, not_new_n8292_, not_new_n8545_);
  not g_22784 (not_new_n4931_, new_n4931_);
  or g_22785 (new_n4714_, not_new_n4507_, not_new_n4508__0);
  or g_22786 (new_n7764_, not_new_n7752_, not_new_n7753__0);
  not g_22787 (not_pi032, pi032);
  or g_22788 (new_n8326_, not_new_n8286__0, not_new_n8126_);
  or g_22789 (new_n9654_, not_new_n9402__0, not_new_n9646_);
  not g_22790 (not_new_n1031__19773267430, new_n1031_);
  not g_22791 (not_new_n6074_, new_n6074_);
  not g_22792 (not_new_n928__8235430, new_n928_);
  or g_22793 (new_n8266_, not_new_n8455_, not_new_n8412_);
  not g_22794 (not_new_n1053__19773267430, new_n1053_);
  not g_22795 (not_new_n5630_, new_n5630_);
  not g_22796 (not_new_n8133__0, new_n8133_);
  or g_22797 (new_n5653_, not_pi147_3, not_new_n5473_);
  not g_22798 (not_new_n6622_, new_n6622_);
  and g_22799 (new_n9858_, new_n10095_, new_n10096_);
  or g_22800 (new_n3121_, not_new_n621__6, not_new_n581__541169560379521116689596608490);
  not g_22801 (not_new_n2856_, new_n2856_);
  and g_22802 (new_n8820_, new_n9020_, new_n9017_);
  not g_22803 (not_new_n8945_, new_n8945_);
  not g_22804 (not_new_n9326_, new_n9326_);
  not g_22805 (not_new_n4466__0, new_n4466_);
  not g_22806 (not_new_n621__70, new_n621_);
  or g_22807 (new_n1676_, not_new_n1631__3430, not_pi047);
  not g_22808 (not_new_n722_, new_n722_);
  or g_22809 (new_n8797_, not_new_n8711_, not_new_n8710_);
  or g_22810 (new_n6412_, not_new_n6245_, not_new_n1598__3430);
  not g_22811 (not_new_n1584__19773267430, new_n1584_);
  not g_22812 (not_po296_273687473400809163430, po296);
  not g_22813 (not_new_n5298_, new_n5298_);
  not g_22814 (new_n4733_, new_n1047_);
  not g_22815 (not_new_n7033__0, new_n7033_);
  or g_22816 (or_not_new_n5463__not_new_n5680__1, not_new_n5463_, not_new_n5680__1);
  or g_22817 (new_n2225_, not_pi154, not_new_n587__6782230728490);
  or g_22818 (new_n686_, not_new_n3026_, not_new_n1502_);
  or g_22819 (new_n4102_, not_pi252_0, not_new_n4169_);
  or g_22820 (new_n2537_, not_new_n2536_, not_new_n611__6);
  not g_22821 (not_new_n8947_, new_n8947_);
  not g_22822 (not_new_n5248_, new_n5248_);
  or g_22823 (new_n4576_, not_new_n1012__2, not_pi178_1);
  not g_22824 (not_new_n4171_, new_n4171_);
  not g_22825 (not_new_n581__93874803376477543056490, new_n581_);
  not g_22826 (not_new_n8135__0, new_n8135_);
  not g_22827 (new_n4276_, new_n654_);
  or g_22828 (new_n6952_, not_new_n6609_, not_new_n6642_);
  not g_22829 (not_new_n3467_, new_n3467_);
  and g_22830 (new_n6357_, and_new_n6417__new_n6418_, new_n6419_);
  not g_22831 (not_new_n3752_, new_n3752_);
  not g_22832 (not_new_n7934__0, new_n7934_);
  not g_22833 (not_new_n7863__0, new_n7863_);
  and g_22834 (new_n9467_, new_n9618_, new_n9338_);
  not g_22835 (not_new_n7750_, new_n7750_);
  not g_22836 (not_new_n1728__168070, new_n1728_);
  or g_22837 (new_n6744_, not_new_n6539_, not_new_n1597__24010);
  not g_22838 (new_n6812_, new_n6547_);
  not g_22839 (not_new_n6002_, new_n6002_);
  or g_22840 (or_not_new_n9361__not_new_n9358__0, not_new_n9358__0, not_new_n9361_);
  or g_22841 (new_n1919_, not_new_n1914_, not_new_n1256_);
  and g_22842 (new_n5022_, new_n5091_, new_n5023_);
  not g_22843 (new_n7628_, new_n625_);
  not g_22844 (not_new_n5891__0, new_n5891_);
  not g_22845 (not_new_n10104_, new_n10104_);
  not g_22846 (new_n6486_, new_n1039_);
  not g_22847 (not_new_n629__1, new_n629_);
  or g_22848 (or_not_new_n5291__not_new_n5290_, not_new_n5291_, not_new_n5290_);
  not g_22849 (not_new_n3147_, new_n3147_);
  or g_22850 (new_n6679_, not_new_n6473_, not_new_n6474__0);
  not g_22851 (not_new_n9646_, new_n9646_);
  not g_22852 (not_new_n1604__16284135979104490, new_n1604_);
  and g_22853 (and_new_n8723__new_n1174_, new_n1174_, new_n8723_);
  not g_22854 (not_new_n1631__4, key_gate_76);
  not g_22855 (not_new_n3184__332329305696010, new_n3184_);
  not g_22856 (not_new_n9503_, new_n9503_);
  and g_22857 (new_n1520_, and_new_n3061__new_n998_, new_n3059_);
  not g_22858 (not_new_n1353_, new_n1353_);
  not g_22859 (not_new_n10001_, new_n10001_);
  and g_22860 (new_n6364_, new_n6431_, and_new_n6433__new_n6432_);
  not g_22861 (not_new_n7313_, new_n7313_);
  not g_22862 (new_n8522_, new_n8226_);
  not g_22863 (not_new_n9809_, new_n9809_);
  not g_22864 (not_new_n5728_, new_n5728_);
  not g_22865 (not_new_n1576__1176490, new_n1576_);
  not g_22866 (not_new_n5028_, new_n5028_);
  not g_22867 (not_new_n4128__0, new_n4128_);
  or g_22868 (new_n6399_, not_new_n648__57648010, not_new_n6296_);
  not g_22869 (not_new_n8818_, new_n8818_);
  not g_22870 (not_new_n741__0, new_n741_);
  not g_22871 (not_pi149_0, pi149);
  or g_22872 (new_n7857_, not_new_n7854_, not_new_n7856_);
  and g_22873 (and_new_n2048__new_n2051_, new_n2051_, new_n2048_);
  not g_22874 (not_new_n944_, new_n944_);
  or g_22875 (new_n10057_, not_new_n10056_, not_new_n634__5585458640832840070);
  not g_22876 (not_new_n9523__0, new_n9523_);
  or g_22877 (new_n4193_, not_pi247_1, not_new_n4108_);
  not g_22878 (not_new_n1071__10, new_n1071_);
  and g_22879 (new_n6583_, new_n6725_, new_n6790_);
  not g_22880 (not_new_n7599__1, new_n7599_);
  not g_22881 (not_new_n6953_, new_n6953_);
  or g_22882 (new_n2542_, not_new_n2509__2, not_pi196);
  not g_22883 (not_new_n2209_, new_n2209_);
  and g_22884 (new_n6340_, new_n6373_, new_n6268_);
  not g_22885 (not_new_n5186_, new_n5186_);
  or g_22886 (new_n2302_, not_new_n587__16284135979104490, not_pi158);
  not g_22887 (not_new_n8443__0, new_n8443_);
  or g_22888 (new_n3815_, not_new_n6243_, not_new_n940__0);
  or g_22889 (new_n4331_, not_new_n708_, not_new_n4230_);
  or g_22890 (new_n5670_, not_new_n5668_, not_new_n5669_);
  not g_22891 (not_new_n7606__0, new_n7606_);
  or g_22892 (new_n4897_, not_new_n4809__0, not_new_n4824_);
  or g_22893 (po194, or_not_new_n1551__not_new_n1372_, not_new_n1371_);
  not g_22894 (not_new_n601__9, new_n601_);
  and g_22895 (and_new_n1451__new_n2679_, new_n2679_, new_n1451_);
  or g_22896 (new_n6935_, not_new_n6532__0, not_new_n1063__24010);
  not g_22897 (not_new_n8431_, new_n8431_);
  or g_22898 (new_n7816_, not_new_n7599__1, not_new_n631__332329305696010);
  or g_22899 (new_n5091_, new_n628_, new_n1039_);
  and g_22900 (new_n6328_, new_n6232_, new_n6261_);
  or g_22901 (new_n2033_, not_new_n2028_, not_new_n1280_);
  or g_22902 (new_n10078_, not_new_n631__32199057558131797268376070, not_new_n1043__2326305139872070);
  or g_22903 (new_n6044_, not_new_n5839_, not_new_n5882__1);
  not g_22904 (not_new_n6998_, new_n6998_);
  and g_22905 (new_n9980_, new_n10246_, and_new_n9879__new_n10247_);
  not g_22906 (not_new_n9628_, new_n9628_);
  not g_22907 (not_new_n5770_, new_n5770_);
  not g_22908 (not_new_n8949_, new_n8949_);
  not g_22909 (not_new_n10113_, new_n10113_);
  not g_22910 (not_new_n4080_, new_n4080_);
  not g_22911 (not_new_n4222_, new_n4222_);
  not g_22912 (not_new_n9613_, new_n9613_);
  not g_22913 (not_new_n9402_, new_n9402_);
  or g_22914 (new_n2502_, not_new_n4759__0, not_new_n597__113988951853731430);
  not g_22915 (not_new_n630__70, new_n630_);
  not g_22916 (new_n8103_, new_n634_);
  not g_22917 (not_new_n4194_, new_n4194_);
  or g_22918 (new_n7419_, not_new_n775__168070, not_new_n7121_);
  not g_22919 (not_new_n7643__1, new_n7643_);
  and g_22920 (new_n3923_, new_n4037_, new_n3949_);
  not g_22921 (not_new_n2836_, new_n2836_);
  not g_22922 (not_pi038_1, pi038);
  not g_22923 (new_n9002_, new_n8845_);
  not g_22924 (not_new_n602__6, new_n602_);
  not g_22925 (not_new_n635__1176490, new_n635_);
  not g_22926 (not_new_n635_, new_n635_);
  and g_22927 (and_and_and_not_pi056_1_not_pi055_1_not_pi054_1_not_pi053_1, not_pi053_1, and_and_not_pi056_1_not_pi055_1_not_pi054_1);
  not g_22928 (not_new_n1581__113988951853731430, new_n1581_);
  or g_22929 (new_n8377_, not_new_n8169_, not_new_n8170__0);
  not g_22930 (not_new_n2840_, new_n2840_);
  or g_22931 (new_n2622_, not_new_n2509__10, not_pi204);
  xor g_22932 (key_gate_108, new_n1678_, key_108);
  not g_22933 (not_new_n640__8235430, new_n640_);
  not g_22934 (not_new_n3998__0, key_gate_114);
  not g_22935 (new_n4026_, new_n3984_);
  not g_22936 (not_new_n4516_, new_n4516_);
  or g_22937 (new_n4666_, not_new_n4573_, not_new_n4664_);
  not g_22938 (not_new_n631__47475615099430, new_n631_);
  not g_22939 (new_n9942_, new_n621_);
  not g_22940 (not_new_n603__490, new_n603_);
  not g_22941 (not_new_n621__403536070, new_n621_);
  not g_22942 (not_new_n4185_, new_n4185_);
  xnor g_22943 (key_gate_27, not_new_n3979_, key_27);
  or g_22944 (new_n1703_, not_new_n1631__138412872010, not_pi056);
  or g_22945 (new_n9279_, not_new_n8872_, not_new_n645__47475615099430);
  not g_22946 (not_new_n3184__8235430, new_n3184_);
  not g_22947 (not_new_n1784_, new_n1784_);
  or g_22948 (new_n4636_, not_new_n1009__3, not_new_n4417_);
  not g_22949 (new_n9421_, new_n1596_);
  not g_22950 (not_new_n1055__5, new_n1055_);
  not g_22951 (not_new_n6137_, new_n6137_);
  or g_22952 (or_or_not_new_n1806__not_new_n1807__not_new_n1809_, not_new_n1809_, or_not_new_n1806__not_new_n1807_);
  not g_22953 (not_new_n8128_, new_n8128_);
  not g_22954 (not_pi187, pi187);
  not g_22955 (not_new_n618__168070, new_n618_);
  not g_22956 (new_n4972_, new_n1071_);
  not g_22957 (not_new_n1600__6, new_n1600_);
  not g_22958 (not_pi141_0, pi141);
  not g_22959 (not_new_n5996_, new_n5996_);
  not g_22960 (not_new_n1019__1, new_n1019_);
  and g_22961 (new_n1546_, new_n3604_, new_n3605_);
  and g_22962 (new_n1436_, new_n2609_, new_n2608_);
  or g_22963 (new_n8484_, not_new_n8117__0, not_new_n628__2326305139872070);
  not g_22964 (not_new_n6024_, new_n6024_);
  not g_22965 (not_pi064_16284135979104490, pi064);
  or g_22966 (new_n7672_, not_new_n7933_, not_new_n7652_);
  not g_22967 (not_new_n640__19773267430, new_n640_);
  or g_22968 (new_n5934_, not_new_n635__168070, not_new_n5743_);
  or g_22969 (new_n6081_, not_new_n5890__0, not_new_n5720_);
  not g_22970 (not_new_n8847_, new_n8847_);
  not g_22971 (not_new_n8678_, new_n8678_);
  and g_22972 (new_n6310_, new_n625_, new_n6300_);
  or g_22973 (new_n4126_, not_new_n4204_, not_new_n4203_);
  not g_22974 (not_new_n6308_, new_n6308_);
  not g_22975 (not_new_n6966_, new_n6966_);
  or g_22976 (new_n6024_, not_new_n638__8235430, not_new_n5786__0);
  not g_22977 (new_n3946_, pi059);
  not g_22978 (not_new_n9647__0, new_n9647_);
  or g_22979 (new_n7837_, not_new_n1061__8235430, not_new_n7657_);
  or g_22980 (new_n7015_, not_new_n7006_, not_new_n7276_);
  or g_22981 (new_n3846_, not_new_n1576__8, not_new_n619__7);
  not g_22982 (not_new_n1043__47475615099430, new_n1043_);
  not g_22983 (not_pi110, pi110);
  not g_22984 (not_new_n6974__47475615099430, new_n6974_);
  not g_22985 (not_new_n5617__0, new_n5617_);
  or g_22986 (new_n5221_, not_new_n5219__0, not_new_n5182__0);
  not g_22987 (not_new_n8779_, new_n8779_);
  not g_22988 (not_pi129, pi129);
  or g_22989 (new_n9157_, not_new_n9035_, not_new_n8828__1);
  not g_22990 (not_new_n626__2824752490, new_n626_);
  not g_22991 (not_new_n7666__1, new_n7666_);
  not g_22992 (not_new_n9756_, new_n9756_);
  or g_22993 (new_n6708_, not_new_n6524__0, not_new_n1055__8235430);
  not g_22994 (not_new_n2725_, new_n2725_);
  not g_22995 (not_new_n8581_, new_n8581_);
  not g_22996 (not_new_n1552_, new_n1552_);
  not g_22997 (not_new_n1051__57648010, new_n1051_);
  and g_22998 (new_n587_, new_n1030_, new_n3390_);
  or g_22999 (new_n929_, not_new_n1768__0, not_new_n1028_);
  not g_23000 (not_new_n5772__0, new_n5772_);
  or g_23001 (new_n6137_, not_new_n617__8235430, not_new_n5807__0);
  not g_23002 (not_pi266_1, pi266);
  not g_23003 (not_new_n7893_, new_n7893_);
  not g_23004 (not_new_n1059__490, new_n1059_);
  not g_23005 (not_new_n2675_, new_n2675_);
  not g_23006 (not_new_n1534__138412872010, key_gate_5);
  not g_23007 (not_new_n7173_, new_n7173_);
  or g_23008 (new_n9308_, not_new_n8976_, not_new_n8977_);
  not g_23009 (not_new_n617__8235430, new_n617_);
  not g_23010 (not_new_n5900__2, new_n5900_);
  not g_23011 (not_new_n2779_, new_n2779_);
  not g_23012 (not_new_n6757_, new_n6757_);
  not g_23013 (not_new_n3315__797922662976120010, new_n3315_);
  not g_23014 (not_new_n1067__5, new_n1067_);
  or g_23015 (po290, or_not_new_n2939__not_new_n1485_, not_new_n2938_);
  or g_23016 (or_or_not_new_n8696__not_new_n8690__not_new_n8689_, not_new_n8689_, or_not_new_n8696__not_new_n8690_);
  not g_23017 (not_new_n5697_, new_n5697_);
  or g_23018 (new_n9640_, not_new_n9473_, not_new_n9639_);
  not g_23019 (not_new_n7962_, new_n7962_);
  or g_23020 (new_n2952_, not_new_n602__6782230728490, not_new_n629__3);
  not g_23021 (not_new_n6531_, new_n6531_);
  or g_23022 (new_n2252_, not_new_n1581__6782230728490, not_new_n8181_);
  and g_23023 (new_n1294_, new_n2100_, new_n2101_);
  not g_23024 (not_new_n5888_, new_n5888_);
  not g_23025 (not_new_n4599_, new_n4599_);
  not g_23026 (not_new_n1613__8, new_n1613_);
  not g_23027 (new_n6503_, new_n630_);
  not g_23028 (not_new_n634__47475615099430, new_n634_);
  or g_23029 (new_n7056_, not_new_n7478_, not_new_n7479_);
  not g_23030 (not_new_n10231_, new_n10231_);
  or g_23031 (new_n6802_, not_new_n6635__0, not_new_n6458_);
  not g_23032 (not_new_n4979_, new_n4979_);
  or g_23033 (new_n9619_, not_new_n1602__47475615099430, not_new_n625__273687473400809163430);
  not g_23034 (not_new_n578_, new_n578_);
  not g_23035 (not_new_n647__4, new_n647_);
  not g_23036 (not_new_n3402_, new_n3402_);
  and g_23037 (new_n1451_, new_n1620_, new_n2677_);
  or g_23038 (new_n7835_, not_new_n7573_, not_new_n7775_);
  or g_23039 (new_n3174_, not_new_n1035__3, not_new_n928__113988951853731430);
  or g_23040 (new_n9182_, not_new_n8939_, not_new_n8899__2);
  not g_23041 (not_new_n1047_, new_n1047_);
  not g_23042 (not_new_n8810_, new_n8810_);
  not g_23043 (not_new_n608__3, new_n608_);
  not g_23044 (not_new_n8146__0, new_n8146_);
  not g_23045 (not_new_n928__4, new_n928_);
  not g_23046 (not_new_n1583__10, new_n1583_);
  not g_23047 (not_new_n1639_, key_gate_79);
  not g_23048 (new_n8655_, new_n1159_);
  not g_23049 (not_new_n629__8, new_n629_);
  not g_23050 (not_new_n7905_, new_n7905_);
  and g_23051 (new_n8695_, new_n8791_, new_n8694_);
  or g_23052 (new_n1968_, not_new_n1580__10, not_new_n6569_);
  not g_23053 (not_new_n1039__1176490, new_n1039_);
  and g_23054 (and_not_pi037_2_not_pi036_2, not_pi036_2, not_pi037_2);
  not g_23055 (not_new_n9348_, new_n9348_);
  not g_23056 (not_new_n2721_, new_n2721_);
  or g_23057 (new_n694_, not_new_n1518_, not_new_n3054_);
  not g_23058 (not_new_n643__2, new_n643_);
  or g_23059 (new_n1926_, not_new_n7594_, not_new_n1583__7);
  not g_23060 (not_new_n634__273687473400809163430, new_n634_);
  and g_23061 (new_n588_, new_n3393_, new_n3390_);
  not g_23062 (not_new_n3568_, new_n3568_);
  not g_23063 (not_new_n1536__16284135979104490, new_n1536_);
  not g_23064 (not_new_n6352_, new_n6352_);
  or g_23065 (new_n3744_, not_new_n3743_, not_new_n3742_);
  not g_23066 (not_new_n9479_, new_n9479_);
  not g_23067 (not_new_n633__9, new_n633_);
  not g_23068 (not_new_n9069_, new_n9069_);
  and g_23069 (new_n1303_, new_n2140_, and_new_n1302__new_n2141_);
  not g_23070 (not_new_n635__0, new_n635_);
  or g_23071 (new_n9225_, not_new_n8959__0, not_new_n619__2824752490);
  and g_23072 (new_n6362_, new_n6427_, new_n6428_);
  not g_23073 (not_new_n5049_, new_n5049_);
  not g_23074 (not_new_n8898__1, new_n8898_);
  not g_23075 (not_new_n994__70, new_n994_);
  or g_23076 (new_n4633_, not_new_n4632_, not_new_n4631_);
  not g_23077 (not_new_n631__113988951853731430, new_n631_);
  or g_23078 (new_n8730_, not_new_n1043__403536070, not_new_n8632_);
  or g_23079 (new_n3580_, not_pi156_0, not_new_n1538__332329305696010);
  and g_23080 (new_n1295_, new_n2102_, and_new_n1294__new_n2103_);
  or g_23081 (new_n6139_, not_new_n1597__3430, not_new_n5767__2);
  not g_23082 (not_po296_138412872010, po296);
  not g_23083 (not_pi101, pi101);
  or g_23084 (new_n8845_, not_new_n8927_, not_new_n8926_);
  or g_23085 (new_n9812_, not_new_n9404_, not_new_n646__2326305139872070);
  or g_23086 (new_n9428_, not_new_n9394_, not_new_n9667_);
  or g_23087 (new_n3779_, not_new_n1061__6, not_new_n643__10);
  or g_23088 (new_n2500_, not_new_n4761__0, not_new_n597__16284135979104490);
  not g_23089 (not_new_n630__968890104070, new_n630_);
  not g_23090 (not_new_n626__168070, new_n626_);
  not g_23091 (not_new_n9909_, new_n9909_);
  or g_23092 (new_n968_, not_new_n2191_, or_or_not_new_n1315__not_new_n1313__not_new_n2192_);
  not g_23093 (not_new_n7511_, new_n7511_);
  not g_23094 (not_new_n4645_, new_n4645_);
  not g_23095 (not_new_n6445_, new_n6445_);
  not g_23096 (not_new_n6982__1, new_n6982_);
  or g_23097 (new_n9670_, not_new_n9428_, not_new_n9669_);
  not g_23098 (not_new_n9357_, new_n9357_);
  not g_23099 (not_new_n9668__0, new_n9668_);
  not g_23100 (not_new_n617__4, new_n617_);
  not g_23101 (not_new_n8995__0, new_n8995_);
  not g_23102 (not_new_n644__403536070, new_n644_);
  not g_23103 (not_new_n632__168070, new_n632_);
  not g_23104 (not_new_n9506__1, new_n9506_);
  not g_23105 (not_new_n5732_, new_n5732_);
  not g_23106 (not_new_n7655__0, new_n7655_);
  or g_23107 (new_n2016_, not_new_n587__3430, not_pi143);
  or g_23108 (new_n4530_, new_n1005_, pi167);
  not g_23109 (not_new_n926__0, new_n926_);
  not g_23110 (not_new_n6481__0, new_n6481_);
  not g_23111 (new_n7887_, new_n7671_);
  not g_23112 (not_new_n2583_, new_n2583_);
  not g_23113 (not_new_n5822_, new_n5822_);
  or g_23114 (new_n6940_, not_new_n6520__0, not_new_n643__138412872010);
  not g_23115 (not_new_n7392_, new_n7392_);
  not g_23116 (not_new_n4937__1, new_n4937_);
  or g_23117 (new_n8330_, not_new_n8329_, not_new_n8286__1);
  not g_23118 (not_new_n9397__0, new_n9397_);
  not g_23119 (not_new_n1576__4, new_n1576_);
  not g_23120 (not_new_n9095_, new_n9095_);
  not g_23121 (not_new_n3292_, new_n3292_);
  not g_23122 (not_new_n6456_, new_n6456_);
  not g_23123 (not_new_n2754_, new_n2754_);
  not g_23124 (new_n5785_, new_n1065_);
  not g_23125 (not_new_n593_, new_n593_);
  not g_23126 (not_new_n9191_, new_n9191_);
  not g_23127 (not_new_n9423_, new_n9423_);
  not g_23128 (not_new_n4447_, new_n4447_);
  not g_23129 (not_new_n4711_, new_n4711_);
  not g_23130 (not_new_n585__168070, new_n585_);
  xnor g_23131 (key_gate_47, new_n1651_, key_47);
  not g_23132 (not_new_n1959_, new_n1959_);
  not g_23133 (not_new_n8610_, new_n8610_);
  or g_23134 (new_n4742_, or_not_new_n4831__not_new_n4789_, not_new_n4792_);
  not g_23135 (not_new_n1600__19773267430, new_n1600_);
  not g_23136 (new_n6444_, new_n620_);
  not g_23137 (new_n6302_, new_n1597_);
  not g_23138 (not_new_n5953_, new_n5953_);
  not g_23139 (not_new_n4337__0, new_n4337_);
  not g_23140 (not_new_n617__168070, new_n617_);
  not g_23141 (not_new_n8068_, new_n8068_);
  and g_23142 (new_n4801_, new_n4888_, new_n4889_);
  not g_23143 (not_new_n1534__16284135979104490, key_gate_5);
  not g_23144 (not_new_n1015__4, new_n1015_);
  not g_23145 (not_new_n5814_, new_n5814_);
  or g_23146 (new_n4008_, not_pi039_4, not_new_n3935_);
  or g_23147 (new_n6738_, not_new_n6503__0, not_new_n1601__8235430);
  not g_23148 (not_new_n7301_, new_n7301_);
  or g_23149 (new_n2849_, not_new_n2846_, not_new_n1616__70);
  not g_23150 (not_new_n2934_, new_n2934_);
  or g_23151 (new_n7368_, not_new_n7325_, not_new_n7339_);
  or g_23152 (new_n7546_, not_new_n7412__1, not_new_n732__1);
  or g_23153 (new_n10305_, not_new_n10018__0, not_new_n10017_);
  not g_23154 (not_new_n4145_, new_n4145_);
  or g_23155 (or_not_new_n5276__not_new_n5277_, not_new_n5277_, not_new_n5276_);
  not g_23156 (not_new_n1480_, new_n1480_);
  not g_23157 (not_new_n9719_, new_n9719_);
  not g_23158 (not_pi241, pi241);
  or g_23159 (new_n6028_, not_new_n5798__1, not_new_n1065__490);
  not g_23160 (not_new_n659_, new_n659_);
  or g_23161 (new_n2236_, not_new_n5012_, not_new_n1589__968890104070);
  not g_23162 (not_new_n7655_, new_n7655_);
  not g_23163 (not_new_n5778__0, new_n5778_);
  not g_23164 (not_new_n4254_, new_n4254_);
  buf g_23165 (po025, pi239);
  not g_23166 (not_new_n4147_, new_n4147_);
  not g_23167 (not_new_n9962_, new_n9962_);
  or g_23168 (new_n2750_, not_new_n4116__2, not_new_n3310__0);
  not g_23169 (not_new_n4514_, new_n4514_);
  or g_23170 (new_n2662_, not_pi208, not_new_n2509__24010);
  not g_23171 (not_pi146_2, pi146);
  not g_23172 (not_new_n2948_, new_n2948_);
  not g_23173 (not_new_n736__1, new_n736_);
  or g_23174 (new_n8767_, not_new_n8661_, not_new_n8720__0);
  not g_23175 (not_new_n9506__0, new_n9506_);
  or g_23176 (new_n4006_, not_new_n4005_, not_pi042_3);
  or g_23177 (new_n6881_, not_new_n6497__0, not_new_n621__2824752490);
  or g_23178 (new_n7496_, not_new_n7495_, not_new_n7494_);
  not g_23179 (not_new_n635__138412872010, new_n635_);
  not g_23180 (not_pi139, pi139);
  or g_23181 (new_n2578_, not_new_n4467__0, not_new_n610__6);
  or g_23182 (new_n5360_, not_new_n5359_, not_new_n5358_);
  not g_23183 (new_n3449_, new_n1051_);
  or g_23184 (new_n3158_, not_new_n3315__6782230728490, not_new_n643__5);
  or g_23185 (or_not_new_n2555__not_new_n2554_, not_new_n2555_, not_new_n2554_);
  or g_23186 (new_n3723_, not_new_n3721_, not_new_n3722_);
  not g_23187 (not_new_n1057__9, new_n1057_);
  not g_23188 (not_new_n631__168070, new_n631_);
  or g_23189 (new_n2425_, not_new_n1061__0, not_new_n598__3430);
  not g_23190 (not_new_n8121_, new_n8121_);
  not g_23191 (new_n8875_, new_n1604_);
  or g_23192 (new_n3126_, not_new_n928__3430, not_new_n1600__3);
  not g_23193 (not_pi178_1, pi178);
  not g_23194 (not_new_n1597__70, new_n1597_);
  not g_23195 (not_new_n5279_, new_n5279_);
  not g_23196 (not_new_n8827_, new_n8827_);
  or g_23197 (new_n2585_, not_new_n5491_, not_new_n605__7);
  not g_23198 (not_new_n1156_, new_n1156_);
  and g_23199 (new_n6342_, new_n6224_, new_n1065_);
  not g_23200 (not_new_n5674_, new_n5674_);
  not g_23201 (not_new_n5762_, new_n5762_);
  and g_23202 (new_n1198_, new_n1685_, new_n1683_);
  not g_23203 (not_new_n3284_, new_n3284_);
  not g_23204 (not_new_n3708_, new_n3708_);
  not g_23205 (not_new_n775_, new_n775_);
  not g_23206 (not_new_n643__168070, new_n643_);
  xor g_23207 (key_gate_125, new_n1632_, key_125);
  not g_23208 (not_new_n3484_, new_n3484_);
  or g_23209 (po192, or_not_new_n1549__not_new_n1368_, not_new_n1367_);
  not g_23210 (not_new_n1601__490, new_n1601_);
  or g_23211 (new_n10163_, new_n1599_, new_n622_);
  not g_23212 (not_new_n7744_, new_n7744_);
  or g_23213 (new_n2122_, not_new_n1589__8235430, not_new_n5016_);
  not g_23214 (not_new_n1583__16284135979104490, new_n1583_);
  or g_23215 (new_n10301_, not_new_n1601__13410686196639649008070, not_new_n9935_);
  or g_23216 (new_n6006_, not_new_n5769_, not_new_n629__168070);
  or g_23217 (new_n3146_, not_new_n3315__2824752490, not_new_n646__5);
  not g_23218 (new_n8826_, new_n624_);
  or g_23219 (new_n4588_, not_pi170_2, not_new_n4431_);
  or g_23220 (new_n3870_, not_new_n1576__2824752490, not_new_n646__490);
  not g_23221 (not_new_n1037__9, new_n1037_);
  not g_23222 (not_new_n8596__0, new_n8596_);
  or g_23223 (new_n2742_, not_new_n2735_, not_new_n1616__0);
  or g_23224 (new_n5592_, not_pi138_3, not_new_n5450__0);
  not g_23225 (not_new_n7460_, new_n7460_);
  not g_23226 (not_new_n1171_, new_n1171_);
  not g_23227 (not_new_n9501__0, new_n9501_);
  or g_23228 (new_n5684_, not_new_n5682_, not_new_n1015__6);
  and g_23229 (new_n7584_, new_n7581_, new_n7583_);
  not g_23230 (not_new_n1942_, new_n1942_);
  or g_23231 (new_n9202_, not_new_n634__2326305139872070, not_new_n8838__0);
  or g_23232 (new_n6131_, not_new_n5808__1, not_new_n1596__24010);
  and g_23233 (new_n1367_, and_new_n2404__new_n2403_, new_n2402_);
  not g_23234 (not_new_n682_, new_n682_);
  not g_23235 (not_new_n1581__57648010, new_n1581_);
  not g_23236 (new_n991_, new_n4227_);
  and g_23237 (new_n5844_, new_n5961_, new_n5713_);
  or g_23238 (new_n2987_, not_new_n943_, not_new_n1022_);
  or g_23239 (new_n3764_, not_new_n979_, not_new_n2285_);
  not g_23240 (not_new_n8260_, new_n8260_);
  not g_23241 (not_new_n4142_, new_n4142_);
  or g_23242 (new_n2120_, not_new_n6555_, not_new_n1580__57648010);
  not g_23243 (new_n5202_, new_n5065_);
  not g_23244 (not_new_n3703_, new_n3703_);
  not g_23245 (not_new_n4621_, new_n4621_);
  and g_23246 (new_n612_, pi275, new_n2737_);
  not g_23247 (not_new_n4141_, new_n4141_);
  not g_23248 (new_n7262_, new_n7137_);
  not g_23249 (not_new_n9767_, new_n9767_);
  or g_23250 (new_n6693_, not_new_n6691_, not_new_n6692_);
  not g_23251 (not_new_n7434_, new_n7434_);
  not g_23252 (not_new_n4494__0, new_n4494_);
  not g_23253 (not_new_n1538__19773267430, new_n1538_);
  not g_23254 (not_new_n1043__0, new_n1043_);
  and g_23255 (and_new_n5289__new_n5287_, new_n5287_, new_n5289_);
  not g_23256 (not_new_n6921_, new_n6921_);
  not g_23257 (not_new_n1067__138412872010, new_n1067_);
  not g_23258 (not_new_n4541_, new_n4541_);
  not g_23259 (not_new_n1597__8235430, new_n1597_);
  or g_23260 (new_n1155_, not_new_n3839_, not_new_n3840_);
  not g_23261 (not_new_n6562_, new_n6562_);
  or g_23262 (new_n8975_, not_new_n9173_, not_new_n8871_);
  not g_23263 (not_new_n3315__47475615099430, new_n3315_);
  or g_23264 (new_n7933_, not_new_n7735_, not_new_n7801__0);
  not g_23265 (not_new_n3175_, new_n3175_);
  or g_23266 (new_n9718_, not_new_n9512__1, not_new_n9379_);
  not g_23267 (new_n4997_, new_n640_);
  not g_23268 (not_new_n1301_, new_n1301_);
  not g_23269 (not_new_n1538__9, new_n1538_);
  not g_23270 (not_new_n1585_, new_n1585_);
  not g_23271 (new_n9630_, new_n9493_);
  and g_23272 (new_n1190_, new_n1661_, new_n1659_);
  not g_23273 (not_new_n639__2, new_n639_);
  not g_23274 (not_new_n738_, new_n738_);
  or g_23275 (new_n6557_, not_new_n6947_, not_new_n6946_);
  or g_23276 (new_n2766_, or_not_new_n2765__not_new_n2764_, not_new_n2763_);
  not g_23277 (not_new_n9228_, new_n9228_);
  not g_23278 (not_new_n4732_, new_n4732_);
  or g_23279 (new_n9510_, not_new_n1051__138412872010, not_new_n647__332329305696010);
  not g_23280 (not_new_n8212_, new_n8212_);
  not g_23281 (not_new_n5319_, new_n5319_);
  not g_23282 (not_new_n626_, new_n626_);
  and g_23283 (and_and_new_n1991__new_n1994__new_n1992_, new_n1992_, and_new_n1991__new_n1994_);
  not g_23284 (not_new_n5796_, new_n5796_);
  not g_23285 (not_new_n601__138412872010, new_n601_);
  not g_23286 (not_new_n1616__1, new_n1616_);
  or g_23287 (new_n9508_, not_new_n618__273687473400809163430, not_new_n9491_);
  not g_23288 (not_new_n984__968890104070, new_n984_);
  not g_23289 (new_n7924_, new_n7751_);
  not g_23290 (new_n6260_, new_n644_);
  or g_23291 (new_n1018_, not_new_n3357_, not_new_n3358_);
  not g_23292 (new_n1586_, new_n987_);
  not g_23293 (not_new_n9515__0, new_n9515_);
  not g_23294 (not_pi131_1, pi131);
  not g_23295 (not_new_n4940_, new_n4940_);
  not g_23296 (not_pi024_0, pi024);
  not g_23297 (not_new_n1594_, new_n1594_);
  not g_23298 (not_new_n6544__0, new_n6544_);
  and g_23299 (new_n6639_, new_n6939_, new_n6940_);
  not g_23300 (not_new_n2750_, new_n2750_);
  not g_23301 (not_new_n597__797922662976120010, new_n597_);
  or g_23302 (new_n8031_, not_new_n8030_, not_new_n7779_);
  or g_23303 (new_n6118_, not_new_n5753__1, not_new_n628__57648010);
  or g_23304 (new_n9162_, not_new_n8878__0, not_new_n9086__0);
  or g_23305 (new_n6883_, not_new_n6810_, not_new_n6624_);
  or g_23306 (new_n6783_, not_new_n6644__0, not_new_n6623_);
  and g_23307 (new_n1398_, new_n2481_, new_n2480_);
  or g_23308 (new_n7492_, not_new_n723__0, not_new_n7445__0);
  not g_23309 (not_new_n10077_, new_n10077_);
  or g_23310 (new_n1841_, not_new_n591__3, not_new_n4724_);
  or g_23311 (new_n2481_, not_new_n4771__0, not_new_n597__6782230728490);
  not g_23312 (not_new_n3995__0, new_n3995_);
  not g_23313 (not_new_n4811__0, new_n4811_);
  not g_23314 (not_new_n6204_, new_n6204_);
  not g_23315 (not_new_n4032__1, new_n4032_);
  not g_23316 (not_new_n4440_, new_n4440_);
  not g_23317 (not_new_n633_, new_n633_);
  not g_23318 (not_new_n7098_, new_n7098_);
  not g_23319 (not_pi012, pi012);
  not g_23320 (not_new_n10060_, new_n10060_);
  not g_23321 (not_new_n4999__2, new_n4999_);
  not g_23322 (not_new_n1055__7, new_n1055_);
  not g_23323 (not_new_n4945_, new_n4945_);
  not g_23324 (not_new_n3386_, new_n3386_);
  not g_23325 (not_new_n991_, new_n991_);
  not g_23326 (not_new_n591__16284135979104490, new_n591_);
  not g_23327 (not_new_n6914_, new_n6914_);
  not g_23328 (not_new_n7263_, new_n7263_);
  not g_23329 (not_new_n3473_, new_n3473_);
  not g_23330 (not_new_n599__3, new_n599_);
  not g_23331 (not_po298_3430, po298);
  not g_23332 (not_new_n6972_, new_n6972_);
  not g_23333 (not_new_n729__0, new_n729_);
  not g_23334 (not_new_n1003__5, new_n1003_);
  not g_23335 (not_new_n8880__0, new_n8880_);
  not g_23336 (not_new_n4970__0, new_n4970_);
  or g_23337 (new_n7283_, not_new_n7281_, not_new_n7092_);
  not g_23338 (not_new_n649_, new_n649_);
  or g_23339 (new_n3825_, not_new_n2988_, not_new_n1020__3);
  not g_23340 (not_pi201, pi201);
  not g_23341 (not_po296_2824752490, po296);
  or g_23342 (new_n4367_, not_new_n4260_, not_new_n694_);
  not g_23343 (new_n9895_, new_n1049_);
  not g_23344 (not_new_n7605__1, new_n7605_);
  not g_23345 (not_new_n1597__2326305139872070, new_n1597_);
  not g_23346 (not_new_n1589__24010, new_n1589_);
  or g_23347 (new_n9288_, not_new_n9074_, not_new_n9286_);
  or g_23348 (new_n3791_, not_new_n1065__6, not_new_n637__10);
  not g_23349 (not_new_n3128_, new_n3128_);
  not g_23350 (not_new_n8858__0, new_n8858_);
  not g_23351 (new_n1585_, new_n930_);
  not g_23352 (not_pi021_0, pi021);
  and g_23353 (and_new_n3001__new_n998_, new_n998_, new_n3001_);
  not g_23354 (not_new_n5516_, new_n5516_);
  not g_23355 (not_new_n4772_, new_n4772_);
  and g_23356 (new_n6309_, new_n631_, new_n6287_);
  not g_23357 (not_new_n602__9, new_n602_);
  not g_23358 (not_new_n2323_, new_n2323_);
  not g_23359 (not_new_n7761_, new_n7761_);
  or g_23360 (or_not_new_n2151__not_new_n2148_, not_new_n2148_, not_new_n2151_);
  not g_23361 (not_new_n618__2326305139872070, new_n618_);
  or g_23362 (new_n6703_, not_new_n6524_, not_new_n1055__1176490);
  not g_23363 (not_new_n10337_, new_n10337_);
  not g_23364 (not_new_n4118__1, new_n4118_);
  not g_23365 (not_new_n1983_, new_n1983_);
  not g_23366 (not_new_n4087_, new_n4087_);
  not g_23367 (not_new_n5265_, new_n5265_);
  or g_23368 (new_n9183_, not_new_n9090_, not_new_n8895_);
  not g_23369 (not_new_n4168__0, new_n4168_);
  or g_23370 (new_n6147_, not_new_n5805__0, not_new_n1599__70);
  not g_23371 (not_pi275, pi275);
  not g_23372 (not_new_n9233_, new_n9233_);
  xnor g_23373 (key_gate_103, new_n1687_, key_103);
  or g_23374 (new_n3732_, not_new_n3731_, not_new_n3730_);
  and g_23375 (new_n1276_, and_and_new_n2010__new_n2013__new_n2011_, new_n2012_);
  not g_23376 (not_new_n1019__6, new_n1019_);
  not g_23377 (not_new_n631__6782230728490, new_n631_);
  not g_23378 (not_new_n8926_, new_n8926_);
  or g_23379 (new_n6463_, not_new_n6773_, not_new_n6776_);
  or g_23380 (or_not_new_n4414__0_not_new_n1010__3, not_new_n1010__3, not_new_n4414__0);
  not g_23381 (not_new_n1061_, new_n1061_);
  not g_23382 (not_po298_8, po298);
  not g_23383 (not_new_n773_, new_n773_);
  not g_23384 (not_new_n3238_, new_n3238_);
  not g_23385 (not_new_n7531_, new_n7531_);
  or g_23386 (new_n3226_, not_new_n3185__403536070, not_new_n1065__4);
  not g_23387 (not_new_n9795_, new_n9795_);
  or g_23388 (new_n684_, not_new_n3020_, not_new_n1498_);
  not g_23389 (not_new_n6644_, new_n6644_);
  or g_23390 (new_n4334_, not_new_n4337_, or_or_not_new_n4234__not_new_n4336__not_new_n675_);
  or g_23391 (new_n6393_, not_new_n6272_, not_new_n636__57648010);
  not g_23392 (not_new_n1576__5, new_n1576_);
  or g_23393 (new_n5257_, not_new_n5135_, not_new_n4928__1);
  or g_23394 (new_n7065_, not_new_n7538_, not_new_n7537_);
  or g_23395 (new_n2701_, not_new_n606__57648010, not_new_n5475__0);
  or g_23396 (new_n5607_, not_new_n5497_, not_new_n5498__0);
  not g_23397 (not_new_n6501__0, new_n6501_);
  not g_23398 (not_new_n1061__168070, new_n1061_);
  or g_23399 (new_n9042_, not_new_n9040_, not_new_n8933_);
  or g_23400 (new_n579_, not_new_n641_, not_new_n9891_);
  or g_23401 (or_not_new_n6334__not_new_n6232__0, not_new_n6232__0, not_new_n6334_);
  or g_23402 (new_n8411_, not_new_n642__6782230728490, not_new_n8264__0);
  not g_23403 (not_new_n1576__6, new_n1576_);
  not g_23404 (not_new_n2509__70, new_n2509_);
  and g_23405 (new_n6445_, new_n6670_, new_n6669_);
  not g_23406 (not_new_n7409_, new_n7409_);
  not g_23407 (not_new_n8645_, new_n8645_);
  not g_23408 (not_new_n1039__19773267430, new_n1039_);
  not g_23409 (not_new_n618__39098210485829880490, new_n618_);
  or g_23410 (new_n3345_, not_pi050_0, not_new_n1534__24010);
  or g_23411 (new_n8969_, not_new_n9180_, not_new_n9178_);
  not g_23412 (new_n8353_, new_n8166_);
  or g_23413 (new_n2719_, not_new_n2716_, or_not_new_n2718__not_new_n2717_);
  or g_23414 (new_n2037_, not_new_n585__24010, not_new_n4132_);
  not g_23415 (not_new_n10030_, new_n10030_);
  not g_23416 (not_new_n587__113988951853731430, new_n587_);
  not g_23417 (new_n4437_, pi173);
  not g_23418 (not_new_n5784__0, new_n5784_);
  not g_23419 (not_new_n7752__1, new_n7752_);
  not g_23420 (not_new_n9872__0, new_n9872_);
  not g_23421 (not_new_n4753__0, new_n4753_);
  or g_23422 (new_n4464_, not_new_n4680_, not_new_n4679_);
  or g_23423 (new_n10208_, not_new_n10033__0, not_new_n10191_);
  not g_23424 (not_new_n2886_, new_n2886_);
  not g_23425 (new_n5441_, new_n1006_);
  not g_23426 (not_new_n1035__4, new_n1035_);
  not g_23427 (new_n9633_, new_n9491_);
  or g_23428 (new_n9447_, not_new_n9836_, not_new_n9837_);
  not g_23429 (new_n6794_, new_n6543_);
  or g_23430 (new_n4879_, not_new_n4787__1, not_new_n4833__1);
  or g_23431 (new_n7440_, not_new_n775__138412872010, not_new_n7128_);
  not g_23432 (not_new_n647__2824752490, new_n647_);
  or g_23433 (new_n8990_, new_n624_, new_n1041_);
  not g_23434 (not_new_n3184_, new_n3184_);
  not g_23435 (not_new_n9407_, new_n9407_);
  not g_23436 (not_new_n4159_, new_n4159_);
  and g_23437 (new_n5854_, new_n6015_, new_n6126_);
  not g_23438 (not_new_n605__2, new_n605_);
  not g_23439 (not_new_n625__1, new_n625_);
  not g_23440 (not_new_n10085_, new_n10085_);
  not g_23441 (not_new_n4998_, new_n4998_);
  not g_23442 (not_new_n5063_, new_n5063_);
  or g_23443 (new_n9557_, new_n624_, new_n1041_);
  not g_23444 (not_new_n3143_, new_n3143_);
  or g_23445 (new_n9851_, not_new_n1053__332329305696010, not_new_n9389_);
  not g_23446 (not_new_n6910_, new_n6910_);
  or g_23447 (new_n9725_, not_new_n9368_, not_new_n648__5585458640832840070);
  not g_23448 (not_new_n7360__1, new_n7360_);
  not g_23449 (not_new_n7541_, new_n7541_);
  not g_23450 (not_new_n923_, new_n923_);
  or g_23451 (or_not_new_n2854__not_new_n2853_, not_new_n2853_, not_new_n2854_);
  and g_23452 (new_n7095_, new_n7546_, and_new_n7159__new_n7547_);
  or g_23453 (new_n5572_, new_n1013_, pi145);
  and g_23454 (new_n8086_, new_n8079_, new_n8350_);
  not g_23455 (not_new_n9947__0, new_n9947_);
  not g_23456 (not_new_n7623_, new_n7623_);
  not g_23457 (not_new_n722__0, new_n722_);
  not g_23458 (not_new_n2002_, new_n2002_);
  not g_23459 (not_new_n6189_, new_n6189_);
  not g_23460 (not_new_n581__3, new_n581_);
  or g_23461 (new_n1825_, not_new_n586__3, not_pi165);
  not g_23462 (new_n1800_, new_n944_);
  not g_23463 (not_new_n2104_, new_n2104_);
  not g_23464 (not_new_n6618_, new_n6618_);
  and g_23465 (new_n5036_, new_n5149_, new_n5272_);
  and g_23466 (and_new_n6993__new_n7526_, new_n6993_, new_n7526_);
  not g_23467 (not_new_n7350_, new_n7350_);
  not g_23468 (not_new_n1603_, new_n1603_);
  not g_23469 (not_new_n7863_, new_n7863_);
  not g_23470 (not_new_n1031__490, new_n1031_);
  and g_23471 (and_new_n1746__new_n1747_, new_n1746_, new_n1747_);
  not g_23472 (new_n3937_, pi039);
  not g_23473 (not_po296_1915812313805664144010, po296);
  not g_23474 (not_new_n9378__0, new_n9378_);
  or g_23475 (new_n4204_, not_new_n4099_, not_new_n4168__0);
  or g_23476 (or_not_new_n1291__not_new_n1289_, not_new_n1289_, not_new_n1291_);
  not g_23477 (not_new_n586__19773267430, new_n586_);
  not g_23478 (not_new_n3184__1, new_n3184_);
  or g_23479 (new_n2798_, not_pi253_0, not_po296_367033682172941254412302110320336601888010);
  or g_23480 (new_n6560_, not_new_n6839_, not_new_n6840_);
  not g_23481 (not_new_n7605__0, new_n7605_);
  not g_23482 (not_new_n4375_, new_n4375_);
  not g_23483 (not_new_n4421__0, new_n4421_);
  not g_23484 (not_new_n6467_, new_n6467_);
  or g_23485 (new_n2158_, not_new_n6552_, not_new_n1580__2824752490);
  not g_23486 (not_new_n8412_, new_n8412_);
  or g_23487 (po057, key_gate_59, not_new_n1184_);
  not g_23488 (not_new_n698_, new_n698_);
  not g_23489 (not_new_n9293_, new_n9293_);
  not g_23490 (not_new_n1536__490, new_n1536_);
  not g_23491 (not_new_n9148_, new_n9148_);
  not g_23492 (not_new_n3111_, new_n3111_);
  not g_23493 (not_new_n624__113988951853731430, new_n624_);
  not g_23494 (not_new_n1961_, new_n1961_);
  not g_23495 (new_n7767_, new_n7597_);
  not g_23496 (new_n7325_, new_n7109_);
  not g_23497 (not_new_n5899__1, new_n5899_);
  or g_23498 (new_n4862_, not_new_n1598__7, not_new_n4768_);
  not g_23499 (not_new_n989__168070, new_n989_);
  not g_23500 (not_new_n5501_, new_n5501_);
  not g_23501 (not_new_n2867_, new_n2867_);
  not g_23502 (not_new_n3006_, new_n3006_);
  or g_23503 (or_or_not_new_n1561__not_new_n2464__not_new_n1391_, not_new_n1391_, or_not_new_n1561__not_new_n2464_);
  not g_23504 (not_pi145_1, pi145);
  or g_23505 (or_not_new_n1544__not_new_n1358_, not_new_n1358_, not_new_n1544_);
  or g_23506 (new_n1869_, not_new_n1583__4, not_new_n7686_);
  and g_23507 (new_n8660_, new_n8638_, new_n1055_);
  or g_23508 (new_n4564_, not_new_n1015__2, not_pi175_1);
  or g_23509 (new_n2911_, not_new_n4114__2, not_new_n3310__490);
  or g_23510 (new_n5595_, not_new_n5593_, not_new_n5547_);
  not g_23511 (not_new_n7482_, new_n7482_);
  not g_23512 (new_n8545_, new_n8233_);
  or g_23513 (new_n946_, not_new_n1830_, or_or_not_new_n1239__not_new_n1237__not_new_n1831_);
  not g_23514 (not_new_n2205_, new_n2205_);
  not g_23515 (not_new_n1069__1, new_n1069_);
  not g_23516 (not_new_n5834_, new_n5834_);
  not g_23517 (not_new_n601__6782230728490, new_n601_);
  and g_23518 (new_n4486_, new_n4636_, new_n4637_);
  or g_23519 (new_n3572_, not_new_n1538__138412872010, not_pi152_0);
  not g_23520 (not_new_n647__6782230728490, new_n647_);
  not g_23521 (new_n8066_, new_n7731_);
  not g_23522 (not_new_n1303_, new_n1303_);
  not g_23523 (not_new_n9250_, new_n9250_);
  or g_23524 (new_n6895_, not_new_n6506__0, not_new_n630__403536070);
  not g_23525 (not_new_n4020_, new_n4020_);
  not g_23526 (not_new_n7591_, new_n7591_);
  or g_23527 (new_n5385_, not_new_n1069__9, not_new_n4977_);
  or g_23528 (new_n2828_, not_new_n2825_, or_not_new_n2827__not_new_n2826_);
  or g_23529 (new_n10112_, new_n637_, new_n1065_);
  not g_23530 (not_new_n9499_, new_n9499_);
  not g_23531 (not_new_n7696_, new_n7696_);
  not g_23532 (not_new_n2952_, new_n2952_);
  not g_23533 (not_new_n6194_, new_n6194_);
  not g_23534 (not_new_n585__57648010, new_n585_);
  not g_23535 (not_new_n3384__4, new_n3384_);
  not g_23536 (not_new_n4665_, new_n4665_);
  and g_23537 (new_n6308_, new_n630_, new_n6257_);
  or g_23538 (new_n10319_, not_new_n640__113988951853731430, not_new_n9906__0);
  or g_23539 (po276, not_new_n2813_, or_not_new_n1479__not_new_n1480_);
  or g_23540 (new_n7953_, not_new_n648__968890104070, not_new_n7603__0);
  not g_23541 (not_pi077, pi077);
  not g_23542 (not_new_n1857_, new_n1857_);
  not g_23543 (not_new_n611__0, new_n611_);
  and g_23544 (new_n9860_, new_n10117_, new_n10118_);
  not g_23545 (not_new_n1065__113988951853731430, new_n1065_);
  or g_23546 (new_n2930_, not_new_n1616__2824752490, not_new_n2927_);
  or g_23547 (or_not_new_n3145__not_new_n3146_, not_new_n3146_, not_new_n3145_);
  or g_23548 (new_n1639_, key_gate_80, not_new_n596__1);
  not g_23549 (not_new_n9732_, new_n9732_);
  not g_23550 (not_new_n6503__1, new_n6503_);
  or g_23551 (new_n6370_, not_new_n6283_, not_new_n1605__5);
  not g_23552 (not_new_n6482__0, new_n6482_);
  not g_23553 (not_new_n599__70, new_n599_);
  not g_23554 (not_new_n989__2326305139872070, new_n989_);
  not g_23555 (not_new_n618__2, new_n618_);
  or g_23556 (new_n10324_, not_new_n1071__47475615099430, not_new_n9904_);
  not g_23557 (not_pi268_2, pi268);
  not g_23558 (not_pi167_3, pi167);
  not g_23559 (new_n8885_, new_n1067_);
  or g_23560 (new_n8999_, not_new_n8829_, not_new_n8828_);
  or g_23561 (new_n627_, or_or_not_new_n1958__not_new_n1959__not_new_n1961_, not_new_n1960_);
  not g_23562 (not_new_n3543_, new_n3543_);
  and g_23563 (new_n6341_, new_n6232_, new_n6388_);
  not g_23564 (new_n2057_, new_n637_);
  not g_23565 (not_new_n1047__3, new_n1047_);
  and g_23566 (and_new_n1033__new_n3404_, new_n3404_, new_n1033_);
  or g_23567 (new_n697_, not_new_n1521_, not_new_n3063_);
  not g_23568 (not_new_n1063__8235430, new_n1063_);
  not g_23569 (not_pi127, pi127);
  or g_23570 (po235, not_new_n3656_, not_new_n3657_);
  not g_23571 (not_new_n4280_, new_n4280_);
  not g_23572 (not_new_n8834_, new_n8834_);
  not g_23573 (not_new_n3110_, new_n3110_);
  not g_23574 (not_pi022_0, pi022);
  not g_23575 (new_n7351_, new_n7025_);
  not g_23576 (not_new_n1631__968890104070, key_gate_76);
  not g_23577 (not_new_n2152_, new_n2152_);
  or g_23578 (or_not_new_n1473__not_new_n2722_, not_new_n1473_, not_new_n2722_);
  or g_23579 (new_n963_, not_pi012, not_new_n1536_);
  not g_23580 (new_n7646_, new_n1059_);
  not g_23581 (not_new_n5578_, new_n5578_);
  or g_23582 (new_n4556_, not_new_n1017__2, not_pi173_1);
  or g_23583 (new_n1894_, not_new_n1589__5, not_new_n5005_);
  not g_23584 (new_n9390_, new_n1057_);
  or g_23585 (new_n3029_, not_new_n1027__1176490, not_new_n1162_);
  not g_23586 (not_new_n6534__0, new_n6534_);
  not g_23587 (not_new_n5977_, new_n5977_);
  not g_23588 (not_new_n5486__0, new_n5486_);
  or g_23589 (po160, not_new_n3547_, not_new_n3546_);
  and g_23590 (new_n9481_, new_n9330_, new_n9673_);
  not g_23591 (not_new_n1061__6, new_n1061_);
  not g_23592 (not_new_n4928__1, new_n4928_);
  not g_23593 (not_new_n6060_, new_n6060_);
  or g_23594 (new_n2756_, not_new_n994__4, not_new_n4129__1);
  not g_23595 (not_new_n7034__0, new_n7034_);
  not g_23596 (not_new_n2809_, new_n2809_);
  and g_23597 (new_n1275_, and_new_n1274__new_n2008_, new_n2007_);
  not g_23598 (not_new_n6288_, new_n6288_);
  or g_23599 (new_n4974_, not_new_n1071__8, not_new_n645__3430);
  not g_23600 (not_new_n6049_, new_n6049_);
  not g_23601 (not_pi156_0, pi156);
  not g_23602 (not_new_n1209_, new_n1209_);
  or g_23603 (new_n5011_, not_new_n5349_, not_new_n5350_);
  or g_23604 (new_n8485_, not_new_n8113__2, not_new_n1039__968890104070);
  not g_23605 (new_n10138_, new_n10016_);
  not g_23606 (not_new_n1288_, new_n1288_);
  not g_23607 (not_new_n7078_, new_n7078_);
  or g_23608 (new_n9665_, not_new_n9663_, not_new_n9479_);
  or g_23609 (or_not_new_n3375__2_not_new_n3387__1, not_new_n3387__1, not_new_n3375__2);
  not g_23610 (not_new_n755_, new_n755_);
  not g_23611 (not_new_n5984_, new_n5984_);
  or g_23612 (new_n654_, not_new_n3120_, or_not_new_n3122__not_new_n3121_);
  or g_23613 (new_n1709_, not_pi058, not_new_n1631__6782230728490);
  not g_23614 (not_new_n3307_, new_n3307_);
  or g_23615 (new_n8370_, not_new_n8367_, not_new_n8369_);
  not g_23616 (not_new_n9807_, new_n9807_);
  not g_23617 (not_new_n8676_, new_n8676_);
  or g_23618 (new_n7540_, not_new_n7001__0, not_new_n7034__0);
  not g_23619 (not_new_n9927_, new_n9927_);
  or g_23620 (new_n4819_, not_new_n4731_, not_new_n1047__7);
  not g_23621 (not_new_n9935__0, new_n9935_);
  and g_23622 (and_and_new_n1858__new_n1861__new_n1859_, and_new_n1858__new_n1861_, new_n1859_);
  or g_23623 (new_n9835_, not_new_n9834_, not_new_n9833_);
  not g_23624 (not_new_n626__273687473400809163430, new_n626_);
  not g_23625 (not_new_n6672_, new_n6672_);
  or g_23626 (new_n6916_, not_new_n6634__2, not_new_n6602_);
  or g_23627 (new_n2740_, not_new_n1598__1, not_new_n613_);
  or g_23628 (new_n8189_, not_new_n8582_, not_new_n8583_);
  and g_23629 (new_n9495_, new_n9784_, new_n9785_);
  not g_23630 (not_new_n1051__403536070, new_n1051_);
  not g_23631 (not_new_n1069__3, new_n1069_);
  xor g_23632 (key_gate_31, key_31, not_new_n3930_);
  or g_23633 (new_n10158_, not_new_n9947_, not_new_n10157_);
  not g_23634 (not_new_n645__5, new_n645_);
  not g_23635 (new_n7642_, new_n1065_);
  not g_23636 (not_new_n5333_, new_n5333_);
  or g_23637 (or_not_new_n5766__1_not_new_n6140_, not_new_n5766__1, not_new_n6140_);
  or g_23638 (new_n9852_, not_new_n641__19773267430, not_new_n9359_);
  not g_23639 (not_new_n5575_, new_n5575_);
  or g_23640 (new_n6851_, not_new_n6616_, not_new_n6820_);
  not g_23641 (not_new_n9402__1, new_n9402_);
  or g_23642 (new_n4542_, pi170, new_n1002_);
  not g_23643 (not_new_n6929_, new_n6929_);
  not g_23644 (new_n7117_, new_n763_);
  not g_23645 (not_new_n1189_, new_n1189_);
  and g_23646 (new_n4303_, new_n4358_, new_n4359_);
  not g_23647 (new_n9353_, new_n1041_);
  and g_23648 (and_and_new_n1217__new_n1218__new_n1220_, and_new_n1217__new_n1218_, new_n1220_);
  or g_23649 (new_n1879_, not_new_n4726_, not_new_n591__5);
  not g_23650 (new_n3366_, new_n1021_);
  not g_23651 (new_n9588_, new_n9505_);
  not g_23652 (not_new_n1536__2824752490, new_n1536_);
  or g_23653 (new_n6747_, not_new_n6498_, not_new_n6746_);
  not g_23654 (not_new_n7022_, new_n7022_);
  not g_23655 (not_new_n5592_, new_n5592_);
  or g_23656 (new_n6030_, not_new_n638__57648010, not_new_n5786__1);
  not g_23657 (not_new_n7545_, new_n7545_);
  not g_23658 (not_new_n1585__168070, new_n1585_);
  or g_23659 (new_n3091_, not_new_n634__5, not_new_n3315__3);
  not g_23660 (new_n6886_, new_n6594_);
  or g_23661 (new_n6214_, not_new_n6213_, not_new_n6070_);
  not g_23662 (not_new_n1065__19773267430, new_n1065_);
  not g_23663 (not_new_n4129__2, new_n4129_);
  not g_23664 (not_new_n8915_, new_n8915_);
  or g_23665 (new_n7746_, not_new_n7929_, not_new_n7921_);
  or g_23666 (new_n670_, or_not_new_n3173__not_new_n3172_, not_new_n3171_);
  not g_23667 (not_new_n3187_, new_n3187_);
  or g_23668 (new_n2597_, not_new_n2596_, not_new_n611__490);
  not g_23669 (not_new_n642__47475615099430, new_n642_);
  or g_23670 (new_n10147_, not_new_n10143_, not_new_n10145_);
  not g_23671 (not_new_n610__490, new_n610_);
  not g_23672 (not_pi237, pi237);
  or g_23673 (new_n2518_, not_new_n610__0, not_new_n4461__0);
  not g_23674 (not_new_n1843__0, new_n1843_);
  not g_23675 (not_new_n1434_, new_n1434_);
  not g_23676 (not_new_n8013_, new_n8013_);
  not g_23677 (not_new_n6455_, new_n6455_);
  not g_23678 (not_new_n9646__0, new_n9646_);
  or g_23679 (new_n2170_, not_new_n4125_, not_new_n585__19773267430);
  or g_23680 (new_n9517_, new_n631_, new_n1043_);
  not g_23681 (not_new_n602__8, new_n602_);
  or g_23682 (new_n3173_, not_new_n3315__113988951853731430, not_new_n647__6);
  or g_23683 (new_n5391_, not_new_n637__24010, not_new_n4981_);
  or g_23684 (new_n10303_, not_new_n1601__93874803376477543056490, not_new_n9935__0);
  not g_23685 (not_new_n9299_, new_n9299_);
  not g_23686 (not_new_n9951__2, new_n9951_);
  not g_23687 (not_new_n6776_, new_n6776_);
  or g_23688 (new_n2523_, not_new_n609__1, not_new_n4462_);
  or g_23689 (new_n3287_, not_new_n589__9095436801298611408202050198891430, not_new_n1063__5);
  not g_23690 (not_new_n5576_, new_n5576_);
  not g_23691 (not_new_n642_, new_n642_);
  or g_23692 (new_n7811_, not_new_n7810_, not_new_n7809_);
  not g_23693 (not_new_n8059_, new_n8059_);
  not g_23694 (new_n7921_, new_n7667_);
  not g_23695 (not_new_n596__19773267430, key_gate_88);
  not g_23696 (not_new_n9162_, new_n9162_);
  not g_23697 (not_new_n8349_, new_n8349_);
  and g_23698 (new_n1237_, new_n1832_, new_n1833_);
  not g_23699 (new_n9368_, new_n1049_);
  not g_23700 (not_pi147_3, pi147);
  not g_23701 (not_new_n614_, new_n614_);
  not g_23702 (not_new_n10305_, new_n10305_);
  not g_23703 (not_new_n6061_, new_n6061_);
  or g_23704 (new_n4341_, not_new_n4344_, or_or_not_new_n4240__not_new_n4343__not_new_n704_);
  not g_23705 (not_pi170_0, pi170);
  or g_23706 (or_not_new_n3914__not_new_n3969_, not_new_n3914_, not_new_n3969_);
  not g_23707 (not_new_n2596_, new_n2596_);
  not g_23708 (not_new_n3137_, new_n3137_);
  not g_23709 (not_new_n7660__0, new_n7660_);
  not g_23710 (not_new_n1004__0, new_n1004_);
  not g_23711 (not_new_n5541_, new_n5541_);
  not g_23712 (not_new_n1603__7, new_n1603_);
  and g_23713 (and_new_n1739__new_n1740_, new_n1739_, new_n1740_);
  or g_23714 (new_n7160_, not_new_n7039_, not_new_n725_);
  or g_23715 (new_n3708_, not_pi240, not_new_n989__332329305696010);
  not g_23716 (not_new_n9359_, new_n9359_);
  and g_23717 (new_n1370_, new_n2410_, new_n2411_);
  or g_23718 (new_n2419_, not_new_n9868__0, not_new_n599__490);
  not g_23719 (not_new_n600__24010, new_n600_);
  not g_23720 (not_new_n9236_, new_n9236_);
  not g_23721 (new_n5991_, new_n5901_);
  or g_23722 (new_n9773_, not_new_n1598__332329305696010, not_new_n9378__0);
  not g_23723 (not_new_n3412_, new_n3412_);
  and g_23724 (new_n5855_, new_n5729_, new_n6014_);
  or g_23725 (new_n1988_, not_new_n1591__10, not_new_n8921_);
  not g_23726 (not_new_n5121_, new_n5121_);
  not g_23727 (not_new_n3371_, new_n3371_);
  or g_23728 (new_n5333_, not_new_n4992__0, not_new_n1596__70);
  not g_23729 (not_new_n6003_, new_n6003_);
  not g_23730 (not_new_n9220_, new_n9220_);
  or g_23731 (new_n5630_, not_new_n5437_, not_new_n5526_);
  not g_23732 (not_new_n7766_, new_n7766_);
  not g_23733 (not_new_n3324__0, new_n3324_);
  or g_23734 (or_not_new_n2801__not_new_n2800_, not_new_n2801_, not_new_n2800_);
  not g_23735 (not_new_n8149__0, new_n8149_);
  not g_23736 (not_new_n1549_, new_n1549_);
  not g_23737 (new_n7128_, new_n755_);
  or g_23738 (new_n4147_, not_pi257_4, not_pi269_4);
  or g_23739 (po071, key_gate_123, not_new_n1198_);
  or g_23740 (new_n973_, not_new_n1536__4, not_pi007);
  not g_23741 (not_new_n1537__4, new_n1537_);
  and g_23742 (new_n775_, new_n3179_, new_n922_);
  not g_23743 (not_new_n8143__0, new_n8143_);
  not g_23744 (not_new_n647__2, new_n647_);
  or g_23745 (new_n8482_, not_new_n8451_, not_new_n8247_);
  or g_23746 (new_n5338_, not_new_n4949_, not_new_n1597__9);
  not g_23747 (not_new_n2557_, new_n2557_);
  or g_23748 (new_n5056_, not_new_n5109_, not_new_n5269_);
  or g_23749 (new_n6804_, not_new_n6459_, not_new_n6635__1);
  not g_23750 (not_new_n2525_, new_n2525_);
  or g_23751 (new_n7774_, not_new_n1047__168070, not_new_n7596_);
  or g_23752 (or_or_not_new_n1323__not_new_n1321__not_new_n2230_, or_not_new_n1323__not_new_n1321_, not_new_n2230_);
  not g_23753 (not_new_n2686_, new_n2686_);
  not g_23754 (not_new_n4225_, new_n4225_);
  not g_23755 (not_new_n4268_, new_n4268_);
  or g_23756 (new_n2846_, or_not_new_n2845__not_new_n2844_, not_new_n2843_);
  or g_23757 (new_n3392_, not_pi064_797922662976120010, not_new_n3928__0);
  not g_23758 (not_new_n1631__24010, key_gate_76);
  or g_23759 (new_n3426_, not_new_n1613__3, not_new_n1862_);
  not g_23760 (not_new_n4693_, new_n4693_);
  or g_23761 (new_n7981_, not_new_n1607__490, not_new_n7742_);
  not g_23762 (not_new_n1584__2, new_n1584_);
  not g_23763 (not_new_n3229_, new_n3229_);
  and g_23764 (new_n1273_, new_n2003_, new_n2004_);
  and g_23765 (new_n4293_, new_n674_, new_n4235_);
  not g_23766 (not_new_n621__2326305139872070, new_n621_);
  not g_23767 (not_new_n6653_, new_n6653_);
  not g_23768 (not_new_n606__2, new_n606_);
  and g_23769 (new_n9470_, and_new_n9717__new_n9715_, new_n9632_);
  or g_23770 (new_n3658_, not_new_n989__1, not_pi215);
  not g_23771 (not_new_n3311__24010, new_n3311_);
  or g_23772 (new_n3860_, not_new_n1576__168070, not_new_n625__490);
  or g_23773 (new_n4137_, not_new_n4225_, not_new_n4226_);
  not g_23774 (not_new_n10227_, new_n10227_);
  not g_23775 (not_new_n1061__8235430, new_n1061_);
  not g_23776 (not_new_n1964_, new_n1964_);
  not g_23777 (not_new_n632__6782230728490, new_n632_);
  and g_23778 (and_new_n1215__new_n1780_, new_n1780_, new_n1215_);
  and g_23779 (new_n9979_, new_n10051_, and_new_n10212__new_n10211_);
  and g_23780 (new_n6574_, new_n6573_, new_n6785_);
  xnor g_23781 (key_gate_26, key_26, not_new_n3915_);
  not g_23782 (not_new_n1045__797922662976120010, new_n1045_);
  or g_23783 (new_n7787_, not_new_n7600_, not_new_n635__2824752490);
  or g_23784 (new_n9422_, not_new_n9636_, not_new_n9382_);
  not g_23785 (not_new_n3873_, new_n3873_);
  not g_23786 (not_pi173, pi173);
  not g_23787 (not_new_n9384__0, new_n9384_);
  not g_23788 (not_new_n4320_, new_n4320_);
  not g_23789 (not_new_n1037__2326305139872070, new_n1037_);
  not g_23790 (not_new_n735__0, new_n735_);
  not g_23791 (new_n5739_, new_n634_);
  not g_23792 (not_new_n618__6, new_n618_);
  or g_23793 (new_n9226_, not_new_n1607__8235430, not_new_n8958__0);
  or g_23794 (or_or_not_new_n2537__not_new_n2541__not_new_n1423_, or_not_new_n2537__not_new_n2541_, not_new_n1423_);
  or g_23795 (new_n6949_, not_new_n636__2824752490, not_new_n6523__0);
  or g_23796 (new_n7309_, not_new_n7212__0, not_new_n6997__0);
  not g_23797 (not_new_n4136__1, new_n4136_);
  not g_23798 (not_new_n5579__0, new_n5579_);
  or g_23799 (new_n2891_, not_new_n2888_, or_not_new_n2890__not_new_n2889_);
  or g_23800 (new_n4007_, not_new_n4002_, not_pi040_4);
  not g_23801 (not_new_n9277_, new_n9277_);
  not g_23802 (not_new_n1924_, new_n1924_);
  or g_23803 (or_not_new_n1311__not_new_n1309_, not_new_n1309_, not_new_n1311_);
  or g_23804 (new_n2338_, not_new_n616__0, or_not_new_n1342__not_new_n1343_);
  not g_23805 (not_new_n606__3430, new_n606_);
  or g_23806 (new_n2077_, not_new_n638__0, not_new_n601__24010);
  not g_23807 (not_pi139_2, pi139);
  or g_23808 (new_n9803_, not_new_n9403__0, not_new_n640__2326305139872070);
  not g_23809 (new_n8988_, new_n8859_);
  or g_23810 (new_n9135_, not_new_n9066_, not_new_n8884__0);
  not g_23811 (not_new_n617__16284135979104490, new_n617_);
  not g_23812 (not_new_n1882_, new_n1882_);
  or g_23813 (new_n6930_, not_new_n6723_, not_new_n6929_);
  not g_23814 (not_new_n8892_, new_n8892_);
  not g_23815 (not_new_n603__138412872010, new_n603_);
  not g_23816 (not_new_n621__57648010, new_n621_);
  not g_23817 (not_new_n3387__5, new_n3387_);
  not g_23818 (not_new_n8714_, new_n8714_);
  not g_23819 (not_new_n8885__0, new_n8885_);
  or g_23820 (new_n6591_, not_new_n6868_, not_new_n6869_);
  or g_23821 (new_n2455_, not_new_n1604__0, not_new_n598__403536070);
  or g_23822 (new_n3898_, not_new_n10208_, not_new_n9952_);
  not g_23823 (not_new_n7606__2, new_n7606_);
  not g_23824 (not_new_n4036_, new_n4036_);
  not g_23825 (not_pi261_2, pi261);
  or g_23826 (new_n9951_, or_not_new_n10219__not_new_n10220_, not_new_n10109_);
  not g_23827 (not_new_n1594__9, new_n1594_);
  not g_23828 (new_n1579_, new_n986_);
  not g_23829 (not_new_n4976_, new_n4976_);
  not g_23830 (not_new_n3211_, new_n3211_);
  not g_23831 (not_new_n8264_, new_n8264_);
  and g_23832 (and_and_new_n3750__new_n3753__new_n3759_, and_new_n3750__new_n3753_, new_n3759_);
  not g_23833 (not_new_n2131_, new_n2131_);
  not g_23834 (not_new_n1583__332329305696010, new_n1583_);
  or g_23835 (new_n2182_, not_new_n593__2824752490, not_new_n625_);
  not g_23836 (new_n9378_, new_n621_);
  not g_23837 (new_n7840_, new_n7659_);
  or g_23838 (new_n6817_, not_new_n6613__2, not_new_n6581_);
  not g_23839 (not_new_n1623__0, new_n1623_);
  not g_23840 (not_new_n5138_, new_n5138_);
  not g_23841 (not_new_n1016__3, new_n1016_);
  not g_23842 (not_new_n5161_, new_n5161_);
  and g_23843 (and_new_n4937__new_n5303_, new_n5303_, new_n4937_);
  not g_23844 (not_new_n5296_, new_n5296_);
  not g_23845 (not_new_n4910_, new_n4910_);
  not g_23846 (not_new_n3315__113988951853731430, new_n3315_);
  and g_23847 (new_n3996_, new_n4068_, new_n4067_);
  or g_23848 (new_n4584_, new_n1011_, pi179);
  or g_23849 (new_n6868_, not_new_n6541__1, not_new_n1596__8235430);
  not g_23850 (not_new_n5472__0, new_n5472_);
  not g_23851 (not_pi175, pi175);
  not g_23852 (not_new_n9278_, new_n9278_);
  not g_23853 (not_new_n9890_, new_n9890_);
  not g_23854 (not_new_n7934_, new_n7934_);
  not g_23855 (not_new_n8245_, new_n8245_);
  or g_23856 (new_n7823_, not_new_n626__332329305696010, not_new_n7651_);
  not g_23857 (not_new_n2180_, new_n2180_);
  not g_23858 (not_new_n1536__1, new_n1536_);
  not g_23859 (not_new_n1002__3, new_n1002_);
  not g_23860 (not_new_n9806_, new_n9806_);
  not g_23861 (not_new_n5948_, new_n5948_);
  or g_23862 (new_n9560_, not_new_n9356__0, not_new_n9556_);
  not g_23863 (not_new_n617__24010, new_n617_);
  not g_23864 (not_new_n7989_, new_n7989_);
  or g_23865 (new_n2971_, not_new_n4120__1, not_new_n994__16284135979104490);
  and g_23866 (new_n8217_, new_n8284_, new_n8375_);
  and g_23867 (new_n6973_, new_n7191_, new_n7194_);
  not g_23868 (not_new_n8780_, new_n8780_);
  not g_23869 (not_new_n618__4, new_n618_);
  and g_23870 (new_n1306_, new_n2157_, new_n2158_);
  not g_23871 (not_new_n4480_, new_n4480_);
  not g_23872 (not_new_n2906_, new_n2906_);
  not g_23873 (not_new_n7672__0, new_n7672_);
  not g_23874 (not_new_n3852_, new_n3852_);
  not g_23875 (not_new_n7042__0, new_n7042_);
  not g_23876 (not_new_n3913__1, new_n3913_);
  not g_23877 (not_new_n644__5, new_n644_);
  not g_23878 (not_new_n624__16284135979104490, new_n624_);
  not g_23879 (not_new_n10316_, new_n10316_);
  not g_23880 (new_n5884_, new_n1607_);
  or g_23881 (new_n2539_, not_po296_1915812313805664144010, not_pi261);
  not g_23882 (not_new_n2537_, new_n2537_);
  and g_23883 (new_n1291_, new_n2083_, and_new_n1290__new_n2084_);
  not g_23884 (not_new_n8595__0, new_n8595_);
  or g_23885 (new_n979_, not_pi004, not_new_n1536__7);
  or g_23886 (new_n7944_, not_new_n7704_, not_new_n7943_);
  not g_23887 (not_new_n9586_, new_n9586_);
  or g_23888 (new_n1738_, not_pi082, not_new_n1728__6);
  not g_23889 (new_n1623_, new_n932_);
  not g_23890 (not_new_n3899_, new_n3899_);
  not g_23891 (not_new_n1069__403536070, new_n1069_);
  not g_23892 (new_n9635_, new_n9489_);
  not g_23893 (not_new_n1623_, new_n1623_);
  not g_23894 (new_n1591_, new_n936_);
  or g_23895 (new_n2324_, not_new_n1536__490, not_new_n2323_);
  not g_23896 (not_new_n3498_, new_n3498_);
  or g_23897 (new_n6806_, not_new_n6635__2, not_new_n6460_);
  or g_23898 (new_n2388_, not_new_n600__6, not_new_n4115__0);
  not g_23899 (not_new_n10057_, new_n10057_);
  not g_23900 (not_new_n611__10, new_n611_);
  or g_23901 (new_n9264_, not_new_n1602__968890104070, not_new_n8856_);
  and g_23902 (new_n8595_, new_n8668_, new_n8596_);
  not g_23903 (not_new_n3057_, new_n3057_);
  not g_23904 (not_new_n9126_, new_n9126_);
  not g_23905 (not_new_n8241_, new_n8241_);
  not g_23906 (not_new_n6149_, new_n6149_);
  or g_23907 (new_n4116_, not_new_n4183_, not_new_n4184_);
  not g_23908 (not_new_n6234__1, new_n6234_);
  not g_23909 (not_new_n6602_, new_n6602_);
  or g_23910 (new_n646_, or_or_not_new_n2091__not_new_n2092__not_new_n2094_, not_new_n2093_);
  not g_23911 (not_pi064_47475615099430, pi064);
  not g_23912 (not_new_n1597__6, new_n1597_);
  not g_23913 (not_pi062_1, pi062);
  not g_23914 (not_new_n1019__0, new_n1019_);
  and g_23915 (and_new_n1877__new_n1880_, new_n1880_, new_n1877_);
  not g_23916 (not_new_n3377_, new_n3377_);
  and g_23917 (new_n9862_, new_n10139_, new_n10140_);
  not g_23918 (not_new_n5263_, new_n5263_);
  not g_23919 (not_new_n1268_, new_n1268_);
  or g_23920 (new_n6096_, not_new_n648__1176490, not_new_n5746__0);
  not g_23921 (not_new_n9527_, new_n9527_);
  not g_23922 (not_new_n4841__0, new_n4841_);
  xnor g_23923 (key_gate_40, not_new_n1720_, key_40);
  or g_23924 (new_n4494_, not_new_n4571_, not_new_n4572_);
  not g_23925 (new_n8863_, new_n636_);
  or g_23926 (new_n5824_, not_new_n6209_, not_new_n6210_);
  not g_23927 (not_new_n1041__403536070, new_n1041_);
  not g_23928 (not_new_n1069__47475615099430, new_n1069_);
  or g_23929 (po227, not_new_n1443_, not_new_n1442_);
  buf g_23930 (po008, pi201);
  not g_23931 (not_new_n4498__0, new_n4498_);
  or g_23932 (new_n637_, not_new_n2055_, or_or_not_new_n2053__not_new_n2054__not_new_n2056_);
  or g_23933 (new_n3028_, not_new_n621__4, not_new_n3372__1176490);
  and g_23934 (new_n9977_, new_n1031_, new_n641_);
  not g_23935 (new_n5128_, new_n4946_);
  not g_23936 (not_new_n8984__1, new_n8984_);
  not g_23937 (not_new_n8820_, new_n8820_);
  not g_23938 (not_new_n5633_, new_n5633_);
  or g_23939 (new_n9138_, new_n637_, new_n1065_);
  or g_23940 (or_not_new_n1566__not_new_n2489_, not_new_n2489_, not_new_n1566_);
  not g_23941 (new_n4247_, new_n700_);
  not g_23942 (not_pi046_2, pi046);
  not g_23943 (not_new_n994__5, new_n994_);
  not g_23944 (not_new_n2338__0, new_n2338_);
  not g_23945 (not_new_n625__2824752490, new_n625_);
  or g_23946 (new_n1845_, not_pi134, not_new_n587__4);
  or g_23947 (po264, not_new_n3715_, not_new_n3714_);
  not g_23948 (not_new_n1600__10, new_n1600_);
  not g_23949 (not_new_n1598__5, new_n1598_);
  not g_23950 (not_new_n9465_, new_n9465_);
  not g_23951 (not_new_n5102__0, new_n5102_);
  not g_23952 (not_new_n591__490, new_n591_);
  not g_23953 (not_new_n629__7, new_n629_);
  not g_23954 (not_new_n631__32199057558131797268376070, new_n631_);
  or g_23955 (new_n6773_, not_new_n6611_, not_new_n6772_);
  not g_23956 (not_new_n5985_, new_n5985_);
  not g_23957 (not_new_n3905_, new_n3905_);
  not g_23958 (not_new_n1059__2, new_n1059_);
  or g_23959 (or_not_new_n3100__not_new_n3099_, not_new_n3100_, not_new_n3099_);
  not g_23960 (not_new_n6443__0, new_n6443_);
  not g_23961 (not_new_n10037_, new_n10037_);
  not g_23962 (not_new_n5798__1, new_n5798_);
  or g_23963 (or_not_new_n8696__not_new_n8690_, not_new_n8690_, not_new_n8696_);
  not g_23964 (new_n9878_, new_n634_);
  or g_23965 (new_n7565_, not_new_n6974__16284135979104490, not_new_n745__0);
  not g_23966 (not_new_n1053__332329305696010, new_n1053_);
  not g_23967 (not_new_n1631__10, key_gate_76);
  not g_23968 (not_new_n1607__57648010, new_n1607_);
  or g_23969 (or_not_new_n2756__not_new_n2755_, not_new_n2756_, not_new_n2755_);
  not g_23970 (new_n4414_, pi162);
  and g_23971 (new_n7572_, new_n7823_, new_n7822_);
  or g_23972 (new_n9207_, not_new_n8845__2, not_new_n9156_);
  not g_23973 (not_new_n4321_, new_n4321_);
  or g_23974 (new_n3069_, not_new_n1175_, not_new_n1027__113988951853731430);
  not g_23975 (not_new_n4019_, new_n4019_);
  or g_23976 (new_n10277_, not_new_n1596__13410686196639649008070, not_new_n9945__0);
  not g_23977 (not_pi141_2, pi141);
  or g_23978 (new_n4630_, not_pi164_2, not_new_n4420_);
  or g_23979 (new_n10197_, not_new_n10195_, not_new_n10005_);
  not g_23980 (not_new_n3496_, new_n3496_);
  not g_23981 (new_n7107_, new_n767_);
  not g_23982 (not_new_n5419_, new_n5419_);
  and g_23983 (new_n1567_, new_n3646_, new_n3647_);
  or g_23984 (new_n4182_, not_new_n4073_, not_new_n4154_);
  not g_23985 (not_new_n10013_, new_n10013_);
  or g_23986 (new_n7481_, not_new_n7042__0, not_new_n7011__0);
  not g_23987 (not_new_n9013_, new_n9013_);
  or g_23988 (new_n9211_, not_new_n8825_, not_new_n624__47475615099430);
  not g_23989 (not_new_n1588__2, new_n1588_);
  not g_23990 (new_n7120_, new_n764_);
  and g_23991 (new_n5880_, new_n6108_, new_n6107_);
  or g_23992 (new_n3142_, not_new_n632__6, not_new_n581__445676403263631959001900459745680070);
  not g_23993 (not_new_n2826_, new_n2826_);
  not g_23994 (not_new_n4129__0, new_n4129_);
  and g_23995 (new_n6329_, new_n6225_, new_n1063_);
  or g_23996 (new_n2075_, not_new_n4130_, not_new_n585__1176490);
  not g_23997 (not_new_n1728__5, new_n1728_);
  not g_23998 (not_new_n5018_, new_n5018_);
  not g_23999 (not_new_n5905_, new_n5905_);
  or g_24000 (new_n8542_, not_new_n8263_, not_new_n8232_);
  not g_24001 (not_new_n1588__332329305696010, new_n1588_);
  or g_24002 (new_n3778_, not_new_n3474_, not_new_n2019_);
  or g_24003 (new_n733_, not_new_n3294_, not_new_n3293_);
  or g_24004 (new_n5606_, not_new_n5605_, not_new_n5604_);
  not g_24005 (not_new_n598__16284135979104490, new_n598_);
  not g_24006 (not_new_n3146_, new_n3146_);
  not g_24007 (not_new_n1589__47475615099430, new_n1589_);
  or g_24008 (new_n4224_, not_new_n4081_, not_new_n4158_);
  or g_24009 (new_n2317_, not_new_n1596_, not_new_n1588__16284135979104490);
  or g_24010 (new_n1875_, not_new_n4919_, not_new_n1589__4);
  not g_24011 (new_n6070_, new_n5907_);
  not g_24012 (not_new_n8170_, new_n8170_);
  or g_24013 (new_n3824_, not_new_n1023__4, not_new_n998__0);
  not g_24014 (not_new_n8008_, new_n8008_);
  not g_24015 (not_new_n3090_, new_n3090_);
  not g_24016 (not_new_n585__1176490, new_n585_);
  not g_24017 (not_new_n7665__1, new_n7665_);
  not g_24018 (not_new_n3285_, new_n3285_);
  not g_24019 (not_new_n6974__6782230728490, new_n6974_);
  or g_24020 (po171, not_new_n3569_, not_new_n3568_);
  not g_24021 (not_new_n3989_, new_n3989_);
  not g_24022 (not_new_n5858_, new_n5858_);
  or g_24023 (new_n1837_, not_new_n5007_, not_new_n1589__2);
  not g_24024 (not_new_n9460_, new_n9460_);
  not g_24025 (not_new_n3930__0, key_gate_43);
  not g_24026 (not_new_n3202_, new_n3202_);
  or g_24027 (or_or_or_not_new_n2740__not_new_n2743__not_new_n2742__not_new_n2744_, or_or_not_new_n2740__not_new_n2743__not_new_n2742_, not_new_n2744_);
  and g_24028 (new_n6323_, new_n6373_, new_n6270_);
  not g_24029 (not_new_n643__19773267430, new_n643_);
  or g_24030 (new_n6631_, not_new_n6792_, not_new_n6802_);
  not g_24031 (not_new_n605__10, new_n605_);
  not g_24032 (new_n5518_, new_n5505_);
  not g_24033 (not_pi168_0, pi168);
  or g_24034 (new_n1923_, not_new_n4113_, not_new_n585__8);
  not g_24035 (not_new_n2347_, new_n2347_);
  not g_24036 (not_new_n6004_, new_n6004_);
  and g_24037 (new_n8224_, new_n8284_, new_n8256_);
  or g_24038 (new_n10264_, not_new_n10262_, not_new_n10082_);
  or g_24039 (new_n4361_, not_new_n696_, not_new_n4256_);
  not g_24040 (new_n6511_, new_n645_);
  not g_24041 (new_n6996_, new_n734_);
  not g_24042 (not_new_n8604_, new_n8604_);
  not g_24043 (new_n2123_, new_n961_);
  not g_24044 (new_n7366_, new_n7020_);
  and g_24045 (new_n6361_, new_n6423_, and_and_and_new_n6422__new_n6426__new_n6360__new_n6359_);
  or g_24046 (po260, not_new_n3707_, not_new_n3706_);
  not g_24047 (not_new_n1603__968890104070, new_n1603_);
  or g_24048 (new_n9017_, not_new_n9016_, not_new_n8928_);
  not g_24049 (not_new_n2262_, new_n2262_);
  or g_24050 (new_n2809_, not_new_n994__10, not_new_n2808_);
  not g_24051 (not_new_n6524__0, new_n6524_);
  not g_24052 (not_new_n581__24010, new_n581_);
  or g_24053 (new_n4815_, not_new_n4735__0, not_new_n4814__0);
  not g_24054 (not_new_n589__57648010, new_n589_);
  not g_24055 (new_n7653_, new_n636_);
  not g_24056 (not_new_n6443__10, new_n6443_);
  not g_24057 (not_new_n1867_, new_n1867_);
  xnor g_24058 (key_gate_99, not_new_n1693_, key_99);
  or g_24059 (new_n745_, not_new_n1533_, not_new_n3302_);
  and g_24060 (new_n7081_, new_n7227_, new_n7228_);
  not g_24061 (not_new_n9014_, new_n9014_);
  or g_24062 (new_n1743_, not_new_n1728__70, not_pi087);
  or g_24063 (new_n1994_, not_new_n1588__70, not_new_n1055_);
  not g_24064 (not_new_n7441_, new_n7441_);
  not g_24065 (not_new_n1580__2, new_n1580_);
  not g_24066 (not_new_n598__968890104070, new_n598_);
  not g_24067 (not_new_n1067__0, new_n1067_);
  not g_24068 (not_new_n644__6, new_n644_);
  not g_24069 (not_new_n8647_, new_n8647_);
  or g_24070 (new_n5220_, not_new_n5047_, not_new_n5219_);
  not g_24071 (not_pi164_0, pi164);
  and g_24072 (new_n8935_, new_n8800_, new_n8806_);
  not g_24073 (not_new_n10228_, new_n10228_);
  or g_24074 (new_n10309_, not_new_n9932__0, not_new_n625__4599865365447399609768010);
  not g_24075 (not_new_n1538__7, new_n1538_);
  not g_24076 (not_new_n9956_, new_n9956_);
  not g_24077 (not_new_n5118_, new_n5118_);
  or g_24078 (or_not_new_n3103__not_new_n3102_, not_new_n3103_, not_new_n3102_);
  not g_24079 (not_new_n5448_, new_n5448_);
  not g_24080 (new_n5275_, new_n4971_);
  not g_24081 (not_new_n10055_, new_n10055_);
  not g_24082 (not_new_n989__4, new_n989_);
  or g_24083 (new_n3204_, not_new_n3185__8, not_new_n1598__4);
  not g_24084 (not_new_n6280_, new_n6280_);
  xnor g_24085 (key_gate_80, not_new_n3929_, key_80);
  not g_24086 (not_new_n606__0, new_n606_);
  not g_24087 (not_new_n4777__0, new_n4777_);
  not g_24088 (not_new_n5910_, new_n5910_);
  not g_24089 (not_new_n3914__0, new_n3914_);
  not g_24090 (not_new_n5490__0, new_n5490_);
  not g_24091 (not_new_n8495_, new_n8495_);
  not g_24092 (new_n5744_, new_n1041_);
  not g_24093 (not_new_n6699_, new_n6699_);
  and g_24094 (new_n8704_, new_n8786_, and_new_n8789__new_n8784_);
  not g_24095 (not_new_n733__0, new_n733_);
  or g_24096 (new_n9848_, not_new_n9506__3, not_new_n9693_);
  not g_24097 (not_new_n631__1176490, new_n631_);
  not g_24098 (not_new_n6976__0, new_n6976_);
  or g_24099 (new_n5589_, not_new_n1002__6, not_new_n5451_);
  not g_24100 (not_new_n8256_, new_n8256_);
  and g_24101 (new_n4141_, pi272, pi246);
  not g_24102 (not_new_n1055__5585458640832840070, new_n1055_);
  not g_24103 (not_new_n1284_, new_n1284_);
  not g_24104 (not_new_n10009__0, new_n10009_);
  not g_24105 (not_new_n1027__70, new_n1027_);
  or g_24106 (new_n4954_, not_new_n629__3430, not_new_n1600__8);
  or g_24107 (new_n2889_, not_new_n602__8235430, not_new_n625__2);
  or g_24108 (new_n4863_, not_new_n4767__0, not_new_n4840_);
  not g_24109 (not_new_n994__8235430, new_n994_);
  or g_24110 (new_n4384_, not_new_n4311_, not_new_n4381_);
  not g_24111 (not_new_n2964_, new_n2964_);
  or g_24112 (new_n9545_, not_new_n9544_, not_new_n9456_);
  not g_24113 (not_new_n10042_, new_n10042_);
  not g_24114 (not_new_n627__5, new_n627_);
  or g_24115 (new_n2437_, not_new_n646__1, not_new_n603__1176490);
  not g_24116 (not_new_n1534__3430, key_gate_5);
  not g_24117 (new_n7451_, new_n7043_);
  not g_24118 (new_n7919_, new_n7668_);
  not g_24119 (not_new_n8354_, new_n8354_);
  or g_24120 (new_n3759_, not_new_n3757_, not_new_n3758_);
  or g_24121 (new_n1716_, not_po296_2326305139872070, not_pi004_0);
  or g_24122 (new_n1989_, not_new_n1589__10, not_new_n5021_);
  not g_24123 (not_new_n4122__0, new_n4122_);
  not g_24124 (not_new_n3915_, key_gate_66);
  not g_24125 (not_pi240, pi240);
  not g_24126 (not_new_n3972_, new_n3972_);
  not g_24127 (not_new_n7933_, new_n7933_);
  or g_24128 (new_n9789_, not_new_n9495_, not_new_n9416__0);
  not g_24129 (not_new_n3246_, new_n3246_);
  not g_24130 (not_new_n3920__0, new_n3920_);
  not g_24131 (not_new_n3372__5585458640832840070, new_n3372_);
  not g_24132 (not_new_n1023__3, new_n1023_);
  not g_24133 (not_new_n7345__0, new_n7345_);
  not g_24134 (not_new_n647__168070, new_n647_);
  not g_24135 (not_new_n5299_, new_n5299_);
  or g_24136 (new_n3752_, not_new_n2171_, not_new_n967_);
  not g_24137 (new_n8739_, new_n8616_);
  or g_24138 (new_n5313_, not_new_n5311_, not_new_n5312_);
  not g_24139 (not_new_n4016__0, new_n4016_);
  not g_24140 (new_n7644_, new_n1061_);
  not g_24141 (not_new_n1584__7, new_n1584_);
  not g_24142 (new_n2152_, new_n639_);
  not g_24143 (not_new_n1483_, new_n1483_);
  not g_24144 (not_new_n6118_, new_n6118_);
  not g_24145 (not_new_n646__3, new_n646_);
  not g_24146 (not_new_n8026_, new_n8026_);
  not g_24147 (not_new_n6025_, new_n6025_);
  or g_24148 (new_n2560_, not_new_n608__4, not_new_n1015__0);
  not g_24149 (not_new_n629__1176490, new_n629_);
  or g_24150 (new_n2125_, not_new_n593__8235430, not_new_n645_);
  not g_24151 (not_new_n3261_, new_n3261_);
  not g_24152 (not_new_n8690_, new_n8690_);
  or g_24153 (new_n9149_, not_new_n9148_, not_new_n8844_);
  or g_24154 (new_n5317_, not_new_n4924_, not_new_n1039__10);
  not g_24155 (not_pi097, pi097);
  not g_24156 (not_new_n1037__24010, new_n1037_);
  not g_24157 (not_new_n4130__2, new_n4130_);
  or g_24158 (new_n4127_, not_new_n4206_, not_new_n4205_);
  and g_24159 (new_n6239_, and_new_n6316__new_n6227_, new_n6229_);
  or g_24160 (new_n7374_, not_new_n7111_, not_new_n7110_);
  or g_24161 (new_n3868_, not_new_n1576__403536070, not_new_n645__490);
  not g_24162 (not_new_n7268_, new_n7268_);
  not g_24163 (not_new_n7575_, new_n7575_);
  and g_24164 (and_and_new_n6373__new_n6254__new_n6402_, new_n6402_, and_new_n6373__new_n6254_);
  or g_24165 (new_n2855_, or_not_new_n2854__not_new_n2853_, not_new_n2852_);
  or g_24166 (new_n3490_, not_pi114_0, not_new_n1537__1176490);
  not g_24167 (not_new_n1616_, new_n1616_);
  or g_24168 (new_n5115_, new_n1045_, new_n635_);
  not g_24169 (not_new_n4518_, new_n4518_);
  or g_24170 (new_n3881_, not_new_n636__70, not_new_n6443__332329305696010);
  or g_24171 (new_n5138_, not_new_n628__24010, not_new_n1039__9);
  or g_24172 (new_n4177_, not_new_n4144_, not_pi256_1);
  or g_24173 (new_n1057_, not_new_n3462_, not_new_n3463_);
  or g_24174 (po173, not_new_n3573_, not_new_n3572_);
  not g_24175 (not_new_n1015_, new_n1015_);
  not g_24176 (not_new_n626__32199057558131797268376070, new_n626_);
  not g_24177 (not_new_n4961_, new_n4961_);
  not g_24178 (not_new_n5613_, new_n5613_);
  not g_24179 (not_new_n9877_, new_n9877_);
  not g_24180 (not_new_n5088_, new_n5088_);
  not g_24181 (not_new_n6232__0, new_n6232_);
  or g_24182 (new_n7396_, not_new_n7177_, not_new_n7394_);
  and g_24183 (new_n1429_, new_n2570_, new_n2572_);
  not g_24184 (not_new_n635__3430, new_n635_);
  and g_24185 (and_not_pi034_2_not_pi033_4, not_pi034_2, not_pi033_4);
  not g_24186 (not_new_n5471_, new_n5471_);
  not g_24187 (not_new_n6627_, new_n6627_);
  xor g_24188 (key_gate_119, key_119, not_new_n3927_);
  not g_24189 (not_new_n8313_, new_n8313_);
  or g_24190 (new_n1177_, not_new_n3883_, not_new_n3884_);
  not g_24191 (new_n8823_, new_n1039_);
  not g_24192 (not_new_n7655__2, new_n7655_);
  not g_24193 (not_new_n593__2, new_n593_);
  not g_24194 (not_new_n9946_, new_n9946_);
  and g_24195 (new_n5839_, new_n5722_, new_n5721_);
  or g_24196 (new_n2081_, not_new_n1581__168070, not_new_n8095_);
  not g_24197 (not_new_n6443__113988951853731430, new_n6443_);
  not g_24198 (not_pi037, pi037);
  not g_24199 (not_new_n7739_, new_n7739_);
  not g_24200 (not_new_n5327_, new_n5327_);
  not g_24201 (not_new_n4157__1, new_n4157_);
  and g_24202 (new_n1386_, new_n2451_, new_n2450_);
  not g_24203 (not_new_n4208_, new_n4208_);
  or g_24204 (new_n3865_, not_new_n6443__57648010, not_new_n632__70);
  not g_24205 (not_new_n10287_, new_n10287_);
  or g_24206 (new_n5254_, not_new_n5114_, not_new_n5082__0);
  not g_24207 (not_new_n7055_, new_n7055_);
  not g_24208 (not_new_n1584__1176490, new_n1584_);
  not g_24209 (new_n8118_, new_n635_);
  not g_24210 (not_new_n976_, new_n976_);
  not g_24211 (not_new_n7700_, new_n7700_);
  not g_24212 (not_new_n1069__1176490, new_n1069_);
  not g_24213 (not_new_n3452_, new_n3452_);
  and g_24214 (new_n8249_, new_n8489_, new_n8488_);
  not g_24215 (not_new_n5827_, new_n5827_);
  not g_24216 (not_new_n1786_, new_n1786_);
  not g_24217 (not_new_n7354__1, new_n7354_);
  and g_24218 (new_n1345_, new_n590_, new_n1032_);
  not g_24219 (not_new_n1037__3430, new_n1037_);
  or g_24220 (new_n8429_, not_new_n8262__0, not_new_n8227_);
  not g_24221 (not_new_n3830_, new_n3830_);
  or g_24222 (new_n9831_, not_new_n9397_, not_new_n643__5585458640832840070);
  not g_24223 (not_new_n5288_, new_n5288_);
  not g_24224 (not_new_n597__5, new_n597_);
  and g_24225 (new_n7092_, new_n6964_, new_n7282_);
  not g_24226 (not_new_n2929_, new_n2929_);
  not g_24227 (not_new_n4410_, new_n4410_);
  or g_24228 (new_n1993_, not_new_n4808_, not_new_n591__70);
  not g_24229 (not_new_n10092_, new_n10092_);
  not g_24230 (not_new_n7018__2, new_n7018_);
  not g_24231 (not_new_n1611__2326305139872070, new_n1611_);
  not g_24232 (not_new_n1611__57648010, new_n1611_);
  and g_24233 (new_n4474_, new_n4594_, new_n4595_);
  not g_24234 (not_new_n4760__0, new_n4760_);
  not g_24235 (not_new_n8715__0, new_n8715_);
  or g_24236 (new_n641_, not_new_n1789_, or_or_not_new_n1787__not_new_n1788__not_new_n1790_);
  not g_24237 (not_new_n9393_, new_n9393_);
  not g_24238 (not_new_n9928_, new_n9928_);
  or g_24239 (new_n2155_, not_new_n1585__403536070, not_new_n5819_);
  not g_24240 (not_new_n7003_, new_n7003_);
  or g_24241 (new_n1865_, not_new_n588__5, not_pi103);
  not g_24242 (not_new_n639__8, new_n639_);
  not g_24243 (not_new_n4026_, new_n4026_);
  not g_24244 (not_new_n6495__0, new_n6495_);
  not g_24245 (not_new_n589__797922662976120010, new_n589_);
  or g_24246 (new_n2808_, not_new_n995_, not_new_n993_);
  and g_24247 (new_n1411_, new_n607_, new_n1028_);
  not g_24248 (new_n5270_, new_n4996_);
  not g_24249 (not_new_n1581__6, new_n1581_);
  or g_24250 (new_n9375_, not_new_n9550_, not_new_n9551_);
  or g_24251 (new_n1685_, not_pi050, not_new_n1631__1176490);
  not g_24252 (new_n1613_, new_n1537_);
  not g_24253 (not_new_n10325_, new_n10325_);
  or g_24254 (new_n6026_, not_new_n6025_, not_new_n5872_);
  or g_24255 (new_n8027_, not_new_n7723_, not_new_n7751_);
  or g_24256 (new_n9573_, not_new_n9516_, not_new_n9329_);
  not g_24257 (not_new_n1299_, new_n1299_);
  not g_24258 (not_new_n9853_, new_n9853_);
  not g_24259 (not_new_n4650_, new_n4650_);
  and g_24260 (new_n1239_, and_new_n1238__new_n1837_, new_n1836_);
  and g_24261 (new_n1278_, new_n2024_, new_n2025_);
  not g_24262 (not_new_n1041__2824752490, new_n1041_);
  not g_24263 (not_new_n632__9, new_n632_);
  not g_24264 (not_pi188, pi188);
  not g_24265 (new_n6480_, new_n632_);
  not g_24266 (not_po298_5585458640832840070, po298);
  or g_24267 (new_n9224_, not_new_n1607__1176490, not_new_n8958_);
  not g_24268 (not_new_n4111_, new_n4111_);
  not g_24269 (not_new_n10131_, new_n10131_);
  not g_24270 (not_new_n5605_, new_n5605_);
  not g_24271 (new_n6060_, new_n5896_);
  not g_24272 (not_new_n9397_, new_n9397_);
  or g_24273 (po229, not_new_n1447_, not_new_n1448_);
  not g_24274 (not_new_n629__968890104070, new_n629_);
  not g_24275 (not_new_n8993_, new_n8993_);
  or g_24276 (new_n3487_, not_pi015_0, not_new_n1536__797922662976120010);
  and g_24277 (new_n4811_, new_n4896_, new_n4897_);
  not g_24278 (not_new_n4053_, new_n4053_);
  not g_24279 (not_new_n9426__0, new_n9426_);
  not g_24280 (not_new_n4173__0, new_n4173_);
  or g_24281 (or_or_not_new_n1958__not_new_n1959__not_new_n1961_, not_new_n1961_, or_not_new_n1958__not_new_n1959_);
  or g_24282 (or_or_not_new_n1243__not_new_n1241__not_new_n1850_, or_not_new_n1243__not_new_n1241_, not_new_n1850_);
  and g_24283 (new_n1258_, new_n1930_, new_n1929_);
  and g_24284 (new_n7712_, new_n7866_, new_n7865_);
  not g_24285 (not_new_n600__138412872010, new_n600_);
  or g_24286 (new_n3207_, not_new_n622__7, not_new_n589__9);
  or g_24287 (new_n6101_, not_new_n5745__0, not_new_n634__8235430);
  not g_24288 (not_new_n1580__3430, new_n1580_);
  or g_24289 (new_n1881_, not_new_n1248_, not_new_n1876_);
  and g_24290 (new_n7704_, new_n7972_, and_new_n7605__new_n7973_);
  not g_24291 (not_new_n7740_, new_n7740_);
  or g_24292 (new_n5136_, not_new_n5095__0, not_new_n5092__0);
  or g_24293 (new_n8531_, not_new_n8138__1, not_new_n625__113988951853731430);
  not g_24294 (not_new_n5477_, new_n5477_);
  not g_24295 (not_new_n8437_, new_n8437_);
  or g_24296 (new_n5089_, new_n631_, new_n1043_);
  or g_24297 (new_n3698_, not_pi235, not_new_n989__19773267430);
  not g_24298 (not_new_n1607__3, new_n1607_);
  not g_24299 (new_n4442_, new_n1015_);
  not g_24300 (not_new_n1357_, new_n1357_);
  not g_24301 (not_new_n7009__0, new_n7009_);
  not g_24302 (not_new_n4491_, new_n4491_);
  or g_24303 (new_n6848_, not_new_n6489__0, not_new_n1041__24010);
  not g_24304 (not_new_n1607__70, new_n1607_);
  not g_24305 (not_pi136_1, pi136);
  not g_24306 (not_new_n2261_, new_n2261_);
  not g_24307 (not_new_n1373_, new_n1373_);
  or g_24308 (new_n10251_, not_new_n9900__2, not_new_n10200_);
  not g_24309 (not_new_n4077_, new_n4077_);
  not g_24310 (not_new_n7342__1, new_n7342_);
  not g_24311 (not_new_n1604__138412872010, new_n1604_);
  or g_24312 (new_n6211_, not_new_n1057__490, not_new_n5796__0);
  not g_24313 (not_new_n9764_, new_n9764_);
  and g_24314 (and_and_new_n1463__new_n1465__new_n1464_, and_new_n1463__new_n1465_, new_n1464_);
  and g_24315 (new_n6596_, new_n6461_, new_n6737_);
  or g_24316 (new_n653_, or_not_new_n3118__not_new_n3119_, not_new_n3117_);
  or g_24317 (new_n4848_, not_new_n4732_, not_new_n1051__7);
  and g_24318 (new_n9854_, new_n10040_, new_n10039_);
  or g_24319 (new_n4330_, not_new_n4233_, not_new_n676_);
  or g_24320 (new_n8498_, not_new_n8171__0, or_not_new_n618__2326305139872070_not_new_n8496_);
  or g_24321 (new_n6957_, not_new_n626__47475615099430, not_new_n6527__2);
  not g_24322 (not_new_n8141_, new_n8141_);
  not g_24323 (not_new_n7113_, new_n7113_);
  not g_24324 (not_new_n5967_, new_n5967_);
  not g_24325 (not_new_n3715_, new_n3715_);
  not g_24326 (not_new_n6289_, new_n6289_);
  or g_24327 (new_n3451_, not_new_n1957_, not_new_n1613__8);
  not g_24328 (not_new_n5814__0, new_n5814_);
  or g_24329 (new_n4468_, not_new_n4707_, not_new_n4708_);
  not g_24330 (not_new_n1612__968890104070, new_n1612_);
  or g_24331 (or_or_not_new_n1055__168070_not_new_n6325__not_new_n6373__1, not_new_n6373__1, or_not_new_n1055__168070_not_new_n6325_);
  or g_24332 (new_n7219_, not_new_n7424_, not_new_n7002_);
  or g_24333 (new_n9298_, not_new_n638__13410686196639649008070, not_new_n8857__0);
  not g_24334 (not_new_n621__6, new_n621_);
  not g_24335 (not_new_n4806__0, new_n4806_);
  or g_24336 (new_n5208_, not_new_n5066_, not_new_n5199_);
  and g_24337 (new_n5720_, new_n5918_, new_n6011_);
  not g_24338 (not_new_n7615_, new_n7615_);
  or g_24339 (new_n2191_, not_new_n639__0, not_new_n601__2824752490);
  not g_24340 (not_new_n634__3, new_n634_);
  or g_24341 (new_n4332_, not_new_n4237_, not_new_n707_);
  and g_24342 (new_n1236_, and_and_new_n1820__new_n1823__new_n1821_, new_n1822_);
  not g_24343 (not_new_n2790_, new_n2790_);
  not g_24344 (not_new_n9794_, new_n9794_);
  not g_24345 (not_new_n3886_, new_n3886_);
  not g_24346 (not_new_n989__5, new_n989_);
  not g_24347 (not_new_n7795__0, new_n7795_);
  not g_24348 (not_new_n6719_, new_n6719_);
  not g_24349 (not_pi058_2, pi058);
  or g_24350 (new_n6629_, not_new_n6754_, not_new_n6508_);
  or g_24351 (or_not_new_n2774__not_new_n2773_, not_new_n2773_, not_new_n2774_);
  not g_24352 (not_new_n10263_, new_n10263_);
  not g_24353 (not_new_n5757_, new_n5757_);
  not g_24354 (not_new_n6640__0, new_n6640_);
  not g_24355 (not_new_n1603__2326305139872070, new_n1603_);
  or g_24356 (new_n8327_, not_new_n1045__47475615099430, not_new_n8118__1);
  or g_24357 (new_n2950_, not_pi270_0, not_po296_85383234134508499009700170379408027452893070589186688070);
  not g_24358 (not_new_n2849_, new_n2849_);
  not g_24359 (new_n2704_, new_n992_);
  not g_24360 (not_pi265_0, pi265);
  not g_24361 (not_new_n942_, new_n942_);
  not g_24362 (not_new_n634__6, new_n634_);
  and g_24363 (new_n8937_, new_n9064_, new_n8809_);
  not g_24364 (not_new_n8193_, new_n8193_);
  not g_24365 (new_n4157_, new_n4080_);
  not g_24366 (not_new_n4958__0, new_n4958_);
  not g_24367 (not_new_n9906_, new_n9906_);
  or g_24368 (new_n2354_, not_new_n599_, not_new_n9954__0);
  or g_24369 (new_n8256_, not_new_n8216_, not_new_n8440_);
  not g_24370 (not_pi064_10, pi064);
  and g_24371 (new_n1469_, new_n3821_, and_and_new_n2707__new_n2708__new_n3822_);
  or g_24372 (or_not_new_n8713__not_new_n8715_, not_new_n8715_, not_new_n8713_);
  not g_24373 (not_new_n3264_, new_n3264_);
  or g_24374 (new_n9139_, not_new_n8978__0, not_new_n9056_);
  not g_24375 (not_pi013_0, pi013);
  not g_24376 (not_new_n1053__968890104070, new_n1053_);
  and g_24377 (new_n1455_, new_n2690_, and_new_n2692__new_n2691_);
  not g_24378 (not_pi064_968890104070, pi064);
  or g_24379 (new_n4704_, not_new_n1018__4, not_new_n4435__0);
  or g_24380 (new_n6095_, not_new_n5741__1, not_new_n1049__70);
  not g_24381 (not_new_n4783_, new_n4783_);
  not g_24382 (not_new_n8150__0, new_n8150_);
  not g_24383 (not_new_n6536__0, new_n6536_);
  not g_24384 (new_n5436_, new_n1008_);
  not g_24385 (new_n9898_, new_n1051_);
  not g_24386 (not_new_n642__6, new_n642_);
  not g_24387 (not_new_n597__968890104070, new_n597_);
  not g_24388 (not_new_n4762_, new_n4762_);
  not g_24389 (not_new_n7294_, new_n7294_);
  and g_24390 (new_n1217_, and_and_new_n1731__new_n1732__new_n1734_, new_n1733_);
  not g_24391 (not_new_n1952_, new_n1952_);
  not g_24392 (not_new_n4030_, new_n4030_);
  not g_24393 (not_new_n3236_, new_n3236_);
  not g_24394 (not_new_n3839_, new_n3839_);
  not g_24395 (not_new_n6486__1, new_n6486_);
  not g_24396 (not_new_n642__4, new_n642_);
  or g_24397 (new_n1816_, not_new_n6563_, not_new_n1580__2);
  not g_24398 (not_new_n9506_, new_n9506_);
  not g_24399 (not_new_n608__9, new_n608_);
  not g_24400 (not_new_n3226_, new_n3226_);
  or g_24401 (new_n2117_, not_new_n1585__8235430, not_new_n5822_);
  or g_24402 (new_n3773_, not_new_n1069__6, not_new_n646__10);
  not g_24403 (not_new_n648__70, new_n648_);
  not g_24404 (not_new_n8452_, new_n8452_);
  or g_24405 (new_n2307_, not_new_n1585__2326305139872070, not_new_n5816_);
  not g_24406 (not_new_n4094_, new_n4094_);
  not g_24407 (not_new_n4034_, new_n4034_);
  not g_24408 (not_new_n636__4, new_n636_);
  not g_24409 (not_new_n602__10, new_n602_);
  or g_24410 (new_n2590_, not_new_n608__7, not_new_n1018__0);
  not g_24411 (not_new_n644__1, new_n644_);
  not g_24412 (not_new_n7682_, new_n7682_);
  or g_24413 (new_n2100_, not_new_n1581__1176490, not_new_n8187_);
  not g_24414 (not_new_n7494_, new_n7494_);
  not g_24415 (not_new_n1572__0, new_n1572_);
  not g_24416 (not_new_n4088_, new_n4088_);
  not g_24417 (not_new_n4551_, new_n4551_);
  not g_24418 (not_new_n8859__0, new_n8859_);
  and g_24419 (and_not_pi056_1_not_pi055_1, not_pi056_1, not_pi055_1);
  or g_24420 (new_n4876_, not_new_n1035__7, not_new_n4786_);
  not g_24421 (not_new_n984__10, new_n984_);
  not g_24422 (not_new_n6594_, new_n6594_);
  or g_24423 (new_n4399_, not_new_n4396_, not_new_n4316_);
  not g_24424 (not_new_n8903_, new_n8903_);
  or g_24425 (new_n4568_, not_pi176_1, not_new_n1014__2);
  not g_24426 (not_new_n989__57648010, new_n989_);
  not g_24427 (not_new_n775__3, new_n775_);
  not g_24428 (not_new_n1047__138412872010, new_n1047_);
  not g_24429 (not_new_n3212_, new_n3212_);
  not g_24430 (not_new_n9697_, new_n9697_);
  not g_24431 (not_new_n1573_, new_n1573_);
  or g_24432 (new_n10077_, not_new_n10073_, not_new_n9888__0);
  or g_24433 (po076, key_gate_102, not_new_n1203_);
  not g_24434 (not_new_n603__1, new_n603_);
  not g_24435 (not_new_n7430__1, new_n7430_);
  not g_24436 (not_new_n8028_, new_n8028_);
  not g_24437 (not_new_n10168_, new_n10168_);
  or g_24438 (new_n965_, not_new_n1536__0, not_pi011);
  not g_24439 (new_n1588_, new_n920_);
  not g_24440 (not_new_n1611__16284135979104490, new_n1611_);
  not g_24441 (not_new_n7688_, new_n7688_);
  or g_24442 (new_n5649_, not_new_n1028__490, not_new_n5508__0);
  not g_24443 (not_new_n1536__1176490, new_n1536_);
  not g_24444 (not_new_n9789_, new_n9789_);
  not g_24445 (new_n8876_, new_n1069_);
  or g_24446 (new_n4131_, not_new_n4214_, not_new_n4213_);
  not g_24447 (not_new_n9246_, new_n9246_);
  not g_24448 (not_new_n5312_, new_n5312_);
  not g_24449 (new_n4287_, new_n713_);
  or g_24450 (or_not_new_n3167__not_new_n3166_, not_new_n3167_, not_new_n3166_);
  or g_24451 (new_n8422_, not_new_n8360_, not_new_n8361_);
  or g_24452 (new_n6538_, not_new_n621__403536070, not_new_n6497_);
  not g_24453 (not_new_n1010__3, new_n1010_);
  not g_24454 (not_new_n8514_, new_n8514_);
  not g_24455 (not_new_n1045__3, new_n1045_);
  not g_24456 (not_new_n725_, new_n725_);
  or g_24457 (new_n3719_, not_new_n981_, not_new_n2304_);
  not g_24458 (not_new_n9669_, new_n9669_);
  not g_24459 (not_new_n8884__0, new_n8884_);
  or g_24460 (new_n1665_, not_po296_10, not_pi021);
  not g_24461 (not_new_n2781_, new_n2781_);
  not g_24462 (not_new_n7660_, new_n7660_);
  not g_24463 (not_new_n6280__0, new_n6280_);
  not g_24464 (not_new_n2113_, new_n2113_);
  not g_24465 (not_new_n2997_, new_n2997_);
  not g_24466 (not_new_n640__16284135979104490, new_n640_);
  not g_24467 (not_po296_1070069044235980333563563003849377848070, po296);
  or g_24468 (new_n5736_, not_new_n5951_, not_new_n5953_);
  not g_24469 (new_n9916_, new_n1067_);
  not g_24470 (new_n4003_, new_n3936_);
  not g_24471 (not_new_n9960__0, new_n9960_);
  not g_24472 (not_new_n5145_, new_n5145_);
  or g_24473 (new_n3137_, not_new_n3315__8235430, not_new_n640__5);
  or g_24474 (or_not_new_n2989__not_new_n3826_, not_new_n3826_, not_new_n2989_);
  or g_24475 (new_n6063_, not_new_n5900__2, not_new_n5863_);
  not g_24476 (not_new_n5305_, new_n5305_);
  and g_24477 (new_n4903_, new_n5168_, new_n5167_);
  and g_24478 (and_new_n2219__new_n2222_, new_n2219_, new_n2222_);
  not g_24479 (not_pi015_0, pi015);
  not g_24480 (not_new_n3185__5, new_n3185_);
  not g_24481 (not_new_n3948_, new_n3948_);
  and g_24482 (new_n8925_, new_n1031_, new_n641_);
  not g_24483 (not_new_n1005__4, new_n1005_);
  and g_24484 (new_n5842_, new_n6095_, and_new_n5740__new_n6096_);
  not g_24485 (not_new_n5058_, new_n5058_);
  or g_24486 (new_n7373_, not_new_n7371_, not_new_n7372_);
  not g_24487 (new_n6283_, new_n620_);
  or g_24488 (new_n2505_, or_or_not_new_n1406__not_new_n1407__not_new_n1410_, not_new_n1409_);
  not g_24489 (not_new_n1599__4, new_n1599_);
  not g_24490 (not_new_n8881_, new_n8881_);
  or g_24491 (or_or_not_new_n6348__not_new_n6232__2_not_new_n6234__1, not_new_n6234__1, or_not_new_n6348__not_new_n6232__2);
  or g_24492 (new_n3737_, not_new_n624__10, not_new_n1041__6);
  not g_24493 (not_new_n8798_, new_n8798_);
  not g_24494 (not_new_n9932__0, new_n9932_);
  or g_24495 (new_n2601_, not_new_n5492__0, not_new_n606__8);
  not g_24496 (new_n4432_, pi170);
  not g_24497 (new_n7448_, new_n7041_);
  not g_24498 (not_new_n8161_, new_n8161_);
  not g_24499 (not_new_n623__1, new_n623_);
  not g_24500 (not_new_n5735_, new_n5735_);
  not g_24501 (not_new_n2095_, new_n2095_);
  or g_24502 (new_n2725_, not_new_n2724_, not_new_n994__0);
  and g_24503 (and_new_n2354__new_n2353_, new_n2354_, new_n2353_);
  or g_24504 (new_n922_, or_not_new_n1001__not_new_n1000_, not_new_n999_);
  or g_24505 (new_n2764_, not_new_n628__2, not_new_n602__3);
  not g_24506 (not_new_n8281__0, new_n8281_);
  not g_24507 (not_new_n9551_, new_n9551_);
  or g_24508 (or_or_not_new_n2910__not_new_n2913__not_new_n2912_, or_not_new_n2910__not_new_n2913_, not_new_n2912_);
  or g_24509 (new_n1705_, not_new_n596__968890104070, key_gate_124);
  not g_24510 (not_new_n8037_, new_n8037_);
  not g_24511 (not_new_n1589__5, new_n1589_);
  not g_24512 (not_new_n9739_, new_n9739_);
  not g_24513 (new_n6523_, new_n1057_);
  not g_24514 (not_new_n2561_, new_n2561_);
  or g_24515 (new_n2611_, not_new_n5476__0, not_new_n606__9);
  or g_24516 (new_n10121_, not_new_n10120_, not_new_n1604__2326305139872070);
  and g_24517 (new_n1183_, new_n1640_, new_n1638_);
  or g_24518 (new_n8454_, not_new_n8294_, not_new_n8112__1);
  or g_24519 (or_not_new_n2863__not_new_n2862_, not_new_n2863_, not_new_n2862_);
  or g_24520 (new_n5213_, not_new_n5209_, not_new_n5084_);
  or g_24521 (new_n7370_, not_new_n6975__0, not_new_n7019__0);
  not g_24522 (not_new_n5128_, new_n5128_);
  not g_24523 (not_new_n7844_, new_n7844_);
  not g_24524 (not_new_n1537__3, new_n1537_);
  or g_24525 (new_n6530_, not_new_n6786_, not_new_n6710_);
  not g_24526 (not_new_n1016__0, new_n1016_);
  not g_24527 (not_new_n619__1176490, new_n619_);
  not g_24528 (not_new_n1031__403536070, new_n1031_);
  or g_24529 (new_n9155_, not_new_n9011__0, not_new_n8859__0);
  and g_24530 (new_n9456_, new_n9730_, and_new_n9365__new_n9731_);
  or g_24531 (new_n8915_, not_new_n9283_, not_new_n9282_);
  not g_24532 (not_new_n3185__4, new_n3185_);
  or g_24533 (new_n5159_, not_new_n5155_, not_new_n5157_);
  or g_24534 (new_n3082_, not_new_n642__3, not_new_n3372__1915812313805664144010);
  not g_24535 (not_new_n9912_, new_n9912_);
  not g_24536 (not_new_n2114_, new_n2114_);
  not g_24537 (not_new_n5087__0, new_n5087_);
  not g_24538 (not_new_n4641_, new_n4641_);
  or g_24539 (new_n2113_, not_new_n585__57648010, not_new_n4128_);
  or g_24540 (new_n10151_, not_new_n617__13410686196639649008070, not_new_n1597__797922662976120010);
  not g_24541 (not_new_n640__8, new_n640_);
  not g_24542 (not_new_n587__2, new_n587_);
  or g_24543 (new_n5131_, not_new_n5130_, not_new_n5031_);
  not g_24544 (not_new_n606__9, new_n606_);
  or g_24545 (new_n8139_, not_new_n8140_, not_new_n639__968890104070);
  not g_24546 (not_new_n4796_, new_n4796_);
  and g_24547 (new_n7736_, new_n7957_, new_n7958_);
  not g_24548 (not_new_n8794__0, new_n8794_);
  not g_24549 (not_new_n7149_, new_n7149_);
  not g_24550 (not_new_n10243_, new_n10243_);
  or g_24551 (new_n3234_, not_new_n3185__968890104070, not_new_n1057__4);
  not g_24552 (not_pi179_3, pi179);
  not g_24553 (not_new_n9279_, new_n9279_);
  not g_24554 (new_n7357_, new_n7019_);
  not g_24555 (not_new_n4974__1, new_n4974_);
  or g_24556 (new_n3557_, not_new_n2071__0, not_new_n1612__24010);
  not g_24557 (not_new_n3934_, new_n3934_);
  or g_24558 (new_n6171_, not_new_n5779__0, not_new_n640__1176490);
  not g_24559 (new_n8628_, new_n1604_);
  not g_24560 (new_n10069_, new_n9902_);
  and g_24561 (new_n9461_, new_n9520_, new_n9569_);
  not g_24562 (not_new_n9486__0, new_n9486_);
  not g_24563 (not_new_n1597__138412872010, new_n1597_);
  not g_24564 (not_pi010, pi010);
  and g_24565 (new_n7114_, new_n7390_, new_n7391_);
  not g_24566 (not_new_n7746_, new_n7746_);
  not g_24567 (not_new_n3828_, new_n3828_);
  not g_24568 (not_new_n3932__0, key_gate_15);
  or g_24569 (po274, or_or_or_not_new_n2794__not_new_n2797__not_new_n2796__not_new_n2798_, not_new_n2795_);
  not g_24570 (not_new_n5452__1, new_n5452_);
  not g_24571 (not_new_n5398_, new_n5398_);
  not g_24572 (not_new_n605__6, new_n605_);
  not g_24573 (not_new_n10266_, new_n10266_);
  not g_24574 (not_new_n5887__0, new_n5887_);
  or g_24575 (new_n5297_, not_new_n4940_, not_new_n648__24010);
  or g_24576 (new_n9579_, new_n644_, new_n1059_);
  not g_24577 (not_new_n6742_, new_n6742_);
  or g_24578 (new_n3893_, not_new_n10209_, not_new_n10029_);
  not g_24579 (not_new_n3698_, new_n3698_);
  or g_24580 (or_or_not_new_n6354__not_new_n6373__8_not_new_n6355_, not_new_n6355_, or_not_new_n6354__not_new_n6373__8);
  not g_24581 (new_n5105_, new_n4937_);
  not g_24582 (new_n4030_, new_n3947_);
  not g_24583 (not_new_n963_, new_n963_);
  or g_24584 (new_n2507_, not_new_n1411_, not_new_n611__0);
  not g_24585 (not_new_n1259_, new_n1259_);
  or g_24586 (new_n8760_, not_new_n8639_, not_new_n1061__19773267430);
  not g_24587 (not_new_n1631__6, key_gate_76);
  not g_24588 (not_new_n4839__0, new_n4839_);
  not g_24589 (new_n7938_, new_n7760_);
  or g_24590 (new_n8050_, not_new_n8048_, not_new_n8049_);
  or g_24591 (new_n3373_, not_pi054_0, not_new_n1534__332329305696010);
  and g_24592 (new_n4309_, new_n4376_, new_n4377_);
  or g_24593 (new_n7918_, not_new_n7669_, not_new_n7581_);
  or g_24594 (new_n3432_, not_new_n1536__403536070, not_pi026_0);
  not g_24595 (not_pi257_4, pi257);
  not g_24596 (not_new_n9810_, new_n9810_);
  not g_24597 (new_n9355_, new_n631_);
  and g_24598 (po088, key_gate_101, pi067);
  not g_24599 (not_new_n4553_, new_n4553_);
  or g_24600 (new_n7821_, not_new_n7648_, not_new_n1055__2824752490);
  not g_24601 (not_new_n10201_, new_n10201_);
  not g_24602 (not_new_n6528__0, new_n6528_);
  not g_24603 (not_new_n4326_, new_n4326_);
  not g_24604 (not_new_n3315__7, new_n3315_);
  or g_24605 (po212, not_new_n2501_, or_not_new_n1570__not_new_n2502_);
  not g_24606 (new_n2028_, new_n956_);
  or g_24607 (new_n4543_, not_new_n4473_, not_new_n4542_);
  not g_24608 (not_new_n5163_, new_n5163_);
  not g_24609 (not_new_n1004__7, new_n1004_);
  or g_24610 (new_n5118_, not_new_n4937__0, not_new_n5102_);
  not g_24611 (not_new_n648__10, new_n648_);
  not g_24612 (not_new_n2986_, new_n2986_);
  not g_24613 (not_new_n3505_, new_n3505_);
  not g_24614 (not_new_n8815_, new_n8815_);
  or g_24615 (new_n8963_, not_new_n9188_, not_new_n8942_);
  not g_24616 (new_n5805_, new_n622_);
  or g_24617 (new_n2011_, not_new_n593__70, not_new_n644_);
  not g_24618 (not_pi177_3, pi177);
  not g_24619 (not_new_n6322_, new_n6322_);
  not g_24620 (not_new_n601__8, new_n601_);
  or g_24621 (or_or_or_not_new_n2982__not_new_n2985__not_new_n2984__not_new_n2986_, or_or_not_new_n2982__not_new_n2985__not_new_n2984_, not_new_n2986_);
  not g_24622 (not_new_n2910_, new_n2910_);
  not g_24623 (not_new_n1519_, new_n1519_);
  not g_24624 (not_new_n632__113988951853731430, new_n632_);
  or g_24625 (new_n621_, or_or_not_new_n2246__not_new_n2243__not_new_n2244_, not_new_n2245_);
  and g_24626 (new_n7717_, new_n7993_, and_new_n7662__new_n7994_);
  not g_24627 (not_new_n1207_, new_n1207_);
  not g_24628 (not_new_n636__16284135979104490, new_n636_);
  or g_24629 (new_n9775_, not_new_n9418_, not_new_n1599__968890104070);
  not g_24630 (not_new_n9930_, new_n9930_);
  or g_24631 (new_n6617_, not_new_n6819_, not_new_n6571_);
  not g_24632 (not_new_n9890__1, new_n9890_);
  or g_24633 (new_n7861_, not_new_n7624_, not_new_n622__2824752490);
  not g_24634 (new_n1600_, new_n971_);
  not g_24635 (not_new_n2866_, new_n2866_);
  not g_24636 (not_pi040_2, pi040);
  not g_24637 (not_new_n609__1176490, new_n609_);
  or g_24638 (new_n7179_, not_new_n6979_, not_new_n7360_);
  not g_24639 (not_new_n1536__47475615099430, new_n1536_);
  or g_24640 (new_n6601_, not_new_n6907_, not_new_n6908_);
  and g_24641 (and_new_n3375__new_n3387_, new_n3387_, new_n3375_);
  or g_24642 (new_n2279_, not_new_n1588__332329305696010, not_new_n1598_);
  not g_24643 (not_new_n5556_, new_n5556_);
  not g_24644 (not_new_n4450_, new_n4450_);
  or g_24645 (new_n5634_, not_new_n1008__6, not_new_n5632_);
  not g_24646 (not_pi064_57648010, pi064);
  and g_24647 (and_new_n3076__new_n998_, new_n998_, new_n3076_);
  and g_24648 (new_n8942_, and_new_n9189__new_n9187_, new_n9104_);
  not g_24649 (not_new_n1604__5, new_n1604_);
  or g_24650 (new_n10181_, not_new_n10001_, not_new_n10229_);
  not g_24651 (new_n1606_, new_n982_);
  not g_24652 (not_new_n9961_, new_n9961_);
  or g_24653 (new_n10196_, not_new_n626__1577753820348458066150427430, not_new_n1053__16284135979104490);
  or g_24654 (new_n10194_, not_new_n10004_, not_new_n10193_);
  not g_24655 (new_n5571_, new_n5513_);
  not g_24656 (not_new_n632__7, new_n632_);
  not g_24657 (new_n6749_, new_n6622_);
  not g_24658 (not_new_n1045__4, new_n1045_);
  not g_24659 (not_new_n4617_, new_n4617_);
  not g_24660 (not_new_n626__2326305139872070, new_n626_);
  not g_24661 (not_new_n9623__0, new_n9623_);
  not g_24662 (not_new_n928__138412872010, new_n928_);
  not g_24663 (not_new_n9432_, new_n9432_);
  or g_24664 (new_n3724_, not_new_n623__3, not_new_n1606__3);
  not g_24665 (not_new_n4337_, new_n4337_);
  or g_24666 (new_n7253_, not_new_n7451_, not_new_n7013_);
  or g_24667 (new_n4380_, not_new_n689_, not_new_n4271_);
  not g_24668 (not_new_n8262__0, new_n8262_);
  or g_24669 (new_n7208_, not_new_n6995_, not_new_n7415_);
  and g_24670 (new_n8229_, new_n625_, new_n8138_);
  not g_24671 (not_new_n1407_, new_n1407_);
  or g_24672 (or_not_new_n2665__not_new_n2664_, not_new_n2665_, not_new_n2664_);
  or g_24673 (new_n2777_, not_new_n3310__3, not_new_n4136__2);
  not g_24674 (not_new_n618__138412872010, new_n618_);
  or g_24675 (new_n704_, not_new_n1488_, not_new_n2994_);
  not g_24676 (not_new_n4306_, new_n4306_);
  or g_24677 (new_n7877_, not_new_n625__6782230728490, not_new_n7631__0);
  or g_24678 (new_n2139_, not_new_n6554_, not_new_n1580__403536070);
  not g_24679 (not_new_n1004__5, new_n1004_);
  not g_24680 (not_new_n8516_, new_n8516_);
  not g_24681 (not_new_n7652__0, new_n7652_);
  not g_24682 (not_pi196, pi196);
  not g_24683 (not_new_n5786_, new_n5786_);
  not g_24684 (not_new_n7195_, new_n7195_);
  not g_24685 (not_new_n591__3, new_n591_);
  not g_24686 (not_new_n7031__0, new_n7031_);
  not g_24687 (not_new_n1591__332329305696010, new_n1591_);
  or g_24688 (new_n4046_, not_pi044_3, not_new_n4012_);
  not g_24689 (not_new_n7759__2, new_n7759_);
  or g_24690 (or_not_new_n1547__not_new_n1364_, not_new_n1547_, not_new_n1364_);
  not g_24691 (not_new_n5987_, new_n5987_);
  or g_24692 (new_n3380_, not_pi066, not_new_n1535__0);
  or g_24693 (or_not_new_n1773__not_new_n1213_, not_new_n1213_, not_new_n1773_);
  not g_24694 (not_new_n1580__2824752490, new_n1580_);
  or g_24695 (new_n2621_, not_new_n5477__0, not_new_n606__10);
  or g_24696 (or_not_new_n1469__not_new_n3820_, not_new_n1469_, not_new_n3820_);
  not g_24697 (not_new_n3713_, new_n3713_);
  and g_24698 (new_n9488_, new_n9751_, new_n9752_);
  not g_24699 (not_new_n7248_, new_n7248_);
  not g_24700 (not_new_n2853_, new_n2853_);
  or g_24701 (new_n7515_, not_new_n7514_, not_new_n7513_);
  or g_24702 (new_n9374_, not_new_n9458_, not_new_n9554_);
  and g_24703 (new_n8219_, new_n8496_, new_n8381_);
  not g_24704 (not_new_n9494_, new_n9494_);
  or g_24705 (po265, not_new_n3717_, not_new_n3716_);
  and g_24706 (new_n1465_, new_n3747_, new_n3744_);
  not g_24707 (not_new_n5618_, new_n5618_);
  not g_24708 (not_new_n6569_, new_n6569_);
  not g_24709 (not_new_n6467__0, new_n6467_);
  not g_24710 (not_new_n4666_, new_n4666_);
  not g_24711 (not_new_n1612__797922662976120010, new_n1612_);
  not g_24712 (not_new_n600__6, new_n600_);
  not g_24713 (not_new_n2846_, new_n2846_);
  not g_24714 (new_n9486_, new_n619_);
  not g_24715 (not_new_n4966__0, new_n4966_);
  not g_24716 (not_new_n6891_, new_n6891_);
  not g_24717 (not_new_n1711_, key_gate_35);
  not g_24718 (not_new_n4760__1, new_n4760_);
  not g_24719 (not_new_n5865_, new_n5865_);
  not g_24720 (not_new_n4256_, new_n4256_);
  not g_24721 (new_n7781_, new_n7620_);
  or g_24722 (new_n2065_, not_new_n1589__24010, not_new_n5018_);
  or g_24723 (new_n7292_, not_new_n7153_, not_new_n7212_);
  not g_24724 (not_new_n3542_, new_n3542_);
  or g_24725 (new_n7782_, not_new_n7606_, not_new_n1039__57648010);
  not g_24726 (not_new_n8884__1, new_n8884_);
  not g_24727 (not_new_n9874__0, new_n9874_);
  not g_24728 (not_new_n5435__0, new_n5435_);
  not g_24729 (new_n4277_, new_n686_);
  or g_24730 (new_n5748_, not_new_n5750_, not_new_n632__1176490);
  not g_24731 (new_n4533_, new_n4477_);
  or g_24732 (new_n6441_, not_new_n6370__0, not_new_n6238_);
  not g_24733 (not_new_n9893_, new_n9893_);
  not g_24734 (not_new_n596__8235430, key_gate_88);
  not g_24735 (not_new_n9575_, new_n9575_);
  not g_24736 (not_new_n1047__7, new_n1047_);
  not g_24737 (not_new_n1049__19773267430, new_n1049_);
  not g_24738 (not_new_n4997__0, new_n4997_);
  or g_24739 (new_n9221_, not_new_n8821_, not_new_n632__2326305139872070);
  not g_24740 (not_new_n1275_, new_n1275_);
  and g_24741 (new_n5713_, new_n5935_, new_n5934_);
  not g_24742 (not_new_n9092__0, new_n9092_);
  or g_24743 (new_n2079_, not_new_n1585__168070, not_new_n5731_);
  not g_24744 (not_pi159_0, pi159);
  not g_24745 (not_new_n3267_, new_n3267_);
  not g_24746 (not_new_n638__93874803376477543056490, new_n638_);
  or g_24747 (new_n1882_, not_pi168, not_new_n586__6);
  not g_24748 (not_new_n3563_, new_n3563_);
  not g_24749 (not_new_n6992__0, new_n6992_);
  or g_24750 (or_or_or_not_new_n2892__not_new_n2895__not_new_n2894__not_new_n2896_, not_new_n2896_, or_or_not_new_n2892__not_new_n2895__not_new_n2894_);
  or g_24751 (new_n8516_, not_new_n622__968890104070, not_new_n8131__0);
  xnor g_24752 (key_gate_55, key_55, not_new_n3918_);
  not g_24753 (not_new_n632__490, new_n632_);
  or g_24754 (or_or_not_new_n6343__not_new_n6344__not_new_n6345_, or_not_new_n6343__not_new_n6344_, not_new_n6345_);
  or g_24755 (new_n3196_, not_new_n1041__4, not_new_n3185__4);
  not g_24756 (not_new_n8264__0, new_n8264_);
  or g_24757 (new_n5419_, not_new_n5418_, not_new_n5417_);
  or g_24758 (new_n7533_, not_new_n7002__0, not_new_n7035__0);
  not g_24759 (not_new_n8057_, new_n8057_);
  and g_24760 (po092, key_gate_101, pi071);
  not g_24761 (not_new_n1057__168070, new_n1057_);
  or g_24762 (new_n3678_, not_pi225, not_new_n989__70);
  or g_24763 (new_n8538_, not_new_n1604__403536070, not_new_n8141__0);
  not g_24764 (not_new_n5880_, new_n5880_);
  not g_24765 (not_pi135, pi135);
  not g_24766 (not_new_n1031__24010, new_n1031_);
  and g_24767 (new_n4808_, new_n4894_, new_n4895_);
  not g_24768 (not_new_n9103__0, new_n9103_);
  or g_24769 (new_n771_, not_new_n3198_, not_new_n3199_);
  not g_24770 (not_new_n775__24010, new_n775_);
  or g_24771 (new_n5243_, not_new_n5242_, not_new_n5052_);
  or g_24772 (new_n2319_, not_pi191, not_new_n586__113988951853731430);
  not g_24773 (not_new_n3581_, new_n3581_);
  not g_24774 (not_new_n1598__6782230728490, new_n1598_);
  and g_24775 (new_n5076_, new_n5404_, new_n5403_);
  or g_24776 (new_n5985_, not_new_n5798__0, not_new_n1065__70);
  not g_24777 (not_new_n7137__0, new_n7137_);
  or g_24778 (new_n982_, not_pi002, not_new_n1536__9);
  or g_24779 (new_n1918_, not_new_n1588__7, not_new_n1047_);
  not g_24780 (not_new_n7453_, new_n7453_);
  not g_24781 (not_new_n1681_, key_gate_72);
  not g_24782 (not_new_n4578_, new_n4578_);
  not g_24783 (not_new_n7459_, new_n7459_);
  or g_24784 (new_n4178_, not_new_n4079_, not_new_n4156_);
  not g_24785 (not_new_n9560_, new_n9560_);
  not g_24786 (not_new_n1071__6782230728490, new_n1071_);
  not g_24787 (not_po296_113988951853731430, po296);
  or g_24788 (new_n3362_, not_pi064_138412872010, not_pi033_2);
  not g_24789 (not_new_n4137__2, new_n4137_);
  not g_24790 (not_new_n1150__0, new_n1150_);
  or g_24791 (new_n2493_, not_new_n4119__0, not_new_n600__2326305139872070);
  or g_24792 (or_not_new_n5095__1_not_new_n4899__1, not_new_n5095__1, not_new_n4899__1);
  not g_24793 (not_new_n9097__0, new_n9097_);
  not g_24794 (not_new_n4900_, new_n4900_);
  or g_24795 (new_n9960_, not_new_n10272_, not_new_n10273_);
  and g_24796 (and_new_n6357__new_n6356_, new_n6357_, new_n6356_);
  or g_24797 (new_n3518_, not_pi125_0, not_new_n1537__2326305139872070);
  not g_24798 (not_new_n1584__16284135979104490, new_n1584_);
  not g_24799 (not_new_n3369_, new_n3369_);
  or g_24800 (new_n6644_, not_new_n6625_, not_new_n6592_);
  or g_24801 (new_n3150_, not_new_n928__19773267430, not_new_n1067__3);
  not g_24802 (not_new_n637__3, new_n637_);
  not g_24803 (not_new_n632__8, new_n632_);
  not g_24804 (not_new_n5950_, new_n5950_);
  not g_24805 (new_n6273_, new_n627_);
  or g_24806 (new_n6752_, not_new_n6644_, not_new_n6593_);
  not g_24807 (not_new_n8828__1, new_n8828_);
  or g_24808 (new_n3882_, not_new_n636__490, not_new_n1576__332329305696010);
  not g_24809 (not_new_n5580_, new_n5580_);
  or g_24810 (new_n1069_, not_new_n3492_, not_new_n3493_);
  or g_24811 (new_n3032_, not_new_n1027__8235430, not_new_n1163_);
  or g_24812 (new_n9676_, new_n1051_, new_n647_);
  not g_24813 (not_new_n7102_, new_n7102_);
  not g_24814 (not_new_n6329_, new_n6329_);
  not g_24815 (not_new_n633__2824752490, new_n633_);
  not g_24816 (not_new_n8941_, new_n8941_);
  not g_24817 (not_new_n8594_, new_n8594_);
  not g_24818 (not_new_n717_, new_n717_);
  not g_24819 (not_new_n3980_, new_n3980_);
  or g_24820 (po153, not_new_n3532_, not_new_n3533_);
  or g_24821 (new_n7982_, not_new_n7741_, not_new_n619__168070);
  not g_24822 (not_new_n4765__1, new_n4765_);
  not g_24823 (not_new_n1271_, new_n1271_);
  or g_24824 (new_n9700_, not_new_n9367_, not_new_n9334_);
  or g_24825 (new_n624_, or_or_not_new_n1825__not_new_n1826__not_new_n1828_, not_new_n1827_);
  or g_24826 (new_n2216_, not_new_n1591__138412872010, not_new_n8913_);
  or g_24827 (new_n10189_, not_new_n1059__113988951853731430, not_new_n644__273687473400809163430);
  not g_24828 (not_new_n7655__1, new_n7655_);
  or g_24829 (new_n9246_, not_new_n8889_, not_new_n622__47475615099430);
  not g_24830 (new_n6532_, new_n638_);
  not g_24831 (not_new_n5913_, new_n5913_);
  or g_24832 (new_n774_, not_new_n3242_, not_new_n1532_);
  and g_24833 (new_n7074_, new_n7376_, and_new_n6977__new_n7377_);
  not g_24834 (not_new_n3712_, new_n3712_);
  not g_24835 (not_new_n2953_, new_n2953_);
  not g_24836 (not_new_n1599__70, new_n1599_);
  not g_24837 (not_new_n5807_, new_n5807_);
  or g_24838 (new_n8980_, not_new_n618__113988951853731430, not_new_n8963_);
  xor g_24839 (key_gate_70, new_n3917_, key_70);
  not g_24840 (new_n1534_, pi064);
  not g_24841 (not_new_n8862_, new_n8862_);
  not g_24842 (not_new_n1348_, new_n1348_);
  not g_24843 (not_new_n8899__1, new_n8899_);
  or g_24844 (new_n10145_, new_n621_, new_n1598_);
  not g_24845 (not_new_n635__403536070, new_n635_);
  not g_24846 (not_new_n642__2824752490, new_n642_);
  not g_24847 (not_new_n6990_, new_n6990_);
  not g_24848 (not_new_n594__5, new_n594_);
  not g_24849 (not_new_n984__1176490, new_n984_);
  not g_24850 (not_new_n5048_, new_n5048_);
  not g_24851 (new_n4762_, new_n1596_);
  not g_24852 (not_new_n3456_, new_n3456_);
  not g_24853 (not_new_n8007_, new_n8007_);
  or g_24854 (new_n5298_, not_new_n1049__9, not_new_n4941_);
  or g_24855 (new_n3241_, not_new_n642__6, not_new_n589__332329305696010);
  not g_24856 (not_new_n1597__1176490, new_n1597_);
  not g_24857 (not_pi188_0, pi188);
  not g_24858 (not_new_n9358__1, new_n9358_);
  and g_24859 (new_n6963_, new_n7224_, new_n7223_);
  not g_24860 (not_new_n994__168070, new_n994_);
  or g_24861 (new_n8240_, not_new_n8579_, not_new_n8580_);
  not g_24862 (not_new_n7417_, new_n7417_);
  or g_24863 (new_n6423_, not_new_n1039__24010, or_or_not_new_n6334__not_new_n6232__0_not_new_n6235__0);
  not g_24864 (not_new_n4953_, new_n4953_);
  or g_24865 (new_n8199_, not_new_n8572_, not_new_n8573_);
  not g_24866 (new_n8639_, new_n1174_);
  not g_24867 (not_pi161_2, pi161);
  not g_24868 (not_pi039, pi039);
  or g_24869 (new_n7157_, not_new_n7018_, not_new_n7109_);
  not g_24870 (not_new_n5787__0, new_n5787_);
  or g_24871 (new_n6662_, not_new_n6634__1, not_new_n642__8235430);
  or g_24872 (new_n6025_, not_new_n6024_, not_new_n6023_);
  or g_24873 (new_n4580_, not_new_n1011__1, not_pi179_1);
  or g_24874 (new_n2220_, not_new_n629_, not_new_n593__138412872010);
  not g_24875 (not_pi100, pi100);
  not g_24876 (not_new_n5409_, new_n5409_);
  and g_24877 (and_and_new_n1222__new_n1223__new_n1225_, new_n1225_, and_new_n1222__new_n1223_);
  or g_24878 (new_n7016_, not_new_n7220_, not_new_n7221_);
  not g_24879 (not_new_n8563_, new_n8563_);
  not g_24880 (not_new_n8215_, new_n8215_);
  not g_24881 (not_new_n604__70, new_n604_);
  and g_24882 (and_new_n2325__new_n2332_, new_n2325_, new_n2332_);
  and g_24883 (new_n9459_, and_new_n9356__new_n9738_, new_n9737_);
  and g_24884 (new_n6325_, new_n6232_, new_n6273_);
  not g_24885 (not_new_n3845_, new_n3845_);
  or g_24886 (new_n717_, not_new_n3260_, not_new_n3259_);
  or g_24887 (new_n10044_, new_n642_, new_n1035_);
  or g_24888 (new_n8920_, not_new_n9316_, not_new_n9315_);
  and g_24889 (new_n586_, new_n1029_, new_n3393_);
  not g_24890 (not_new_n6066_, new_n6066_);
  and g_24891 (and_new_n2369__new_n2368_, new_n2369_, new_n2368_);
  and g_24892 (new_n1193_, new_n1668_, new_n1670_);
  or g_24893 (new_n4023_, not_new_n3913__1, not_new_n4017__0);
  not g_24894 (not_new_n6052_, new_n6052_);
  not g_24895 (not_new_n7308_, new_n7308_);
  or g_24896 (new_n3096_, not_new_n635__6, not_new_n581__13410686196639649008070);
  or g_24897 (new_n2555_, not_new_n605__4, not_new_n5488_);
  not g_24898 (not_new_n4776_, new_n4776_);
  or g_24899 (new_n8479_, not_new_n8120__0, not_new_n1041__57648010);
  not g_24900 (not_new_n7621__0, new_n7621_);
  not g_24901 (not_new_n8077_, new_n8077_);
  not g_24902 (not_new_n6506__0, new_n6506_);
  not g_24903 (not_new_n1598__403536070, new_n1598_);
  not g_24904 (not_new_n4706_, new_n4706_);
  or g_24905 (new_n3797_, not_new_n635__10, not_new_n1045__6);
  not g_24906 (not_new_n1411_, new_n1411_);
  not g_24907 (not_new_n1616__5, new_n1616_);
  not g_24908 (not_new_n9254_, new_n9254_);
  not g_24909 (not_new_n641__2824752490, new_n641_);
  or g_24910 (new_n7856_, not_new_n1601__19773267430, not_new_n7627__0);
  or g_24911 (new_n5487_, not_new_n5678_, not_new_n5677_);
  not g_24912 (not_new_n1576__0, new_n1576_);
  not g_24913 (not_pi248_3, pi248);
  not g_24914 (not_new_n633__0, new_n633_);
  not g_24915 (new_n2256_, new_n974_);
  not g_24916 (new_n4285_, new_n682_);
  or g_24917 (new_n8181_, not_new_n8518_, not_new_n8519_);
  not g_24918 (not_new_n9398_, new_n9398_);
  or g_24919 (po211, or_or_or_not_new_n2497__not_new_n1568__not_new_n2498__not_new_n2500_, not_new_n2499_);
endmodule

// Benchmark "b17" written by ABC on Sun Apr 23 00:34:15 2023

module b17 ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205,
    pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214,
    pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223,
    pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232,
    pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241,
    pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250,
    pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259,
    pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268,
    pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277,
    pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286,
    pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295,
    pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304,
    pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313,
    pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322,
    pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331,
    pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340,
    pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349,
    pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358,
    pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367,
    pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376,
    pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385,
    pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394,
    pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403,
    pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412,
    pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421,
    pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430,
    pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439,
    pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448,
    pi1449, pi1450, pi1451, pi1452,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232,
    po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241,
    po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250,
    po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259,
    po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268,
    po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277,
    po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286,
    po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295,
    po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304,
    po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313,
    po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322,
    po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331,
    po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340,
    po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349,
    po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358,
    po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367,
    po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376,
    po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385,
    po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394,
    po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403,
    po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412,
    po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421,
    po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430,
    po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439,
    po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448,
    po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457,
    po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466,
    po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475,
    po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484,
    po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493,
    po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502,
    po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204,
    pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213,
    pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222,
    pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231,
    pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240,
    pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249,
    pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258,
    pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267,
    pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276,
    pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285,
    pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294,
    pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303,
    pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312,
    pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321,
    pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330,
    pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339,
    pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348,
    pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357,
    pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366,
    pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375,
    pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384,
    pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393,
    pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402,
    pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411,
    pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420,
    pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429,
    pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438,
    pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447,
    pi1448, pi1449, pi1450, pi1451, pi1452;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231,
    po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240,
    po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249,
    po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258,
    po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267,
    po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276,
    po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285,
    po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294,
    po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303,
    po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312,
    po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321,
    po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330,
    po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339,
    po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348,
    po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357,
    po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366,
    po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375,
    po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384,
    po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393,
    po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402,
    po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411,
    po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420,
    po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429,
    po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438,
    po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447,
    po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456,
    po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465,
    po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474,
    po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483,
    po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492,
    po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501,
    po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510,
    po1511;
  wire new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n3010_, new_n3011_, new_n3012_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_,
    new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4434_, new_n4435_, new_n4439_, new_n4442_,
    new_n4443_, new_n4447_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_,
    new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_,
    new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_,
    new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_,
    new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_,
    new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_,
    new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_,
    new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_,
    new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_,
    new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_,
    new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_,
    new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_,
    new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_,
    new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_,
    new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_,
    new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_,
    new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_,
    new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_,
    new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_,
    new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_,
    new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_,
    new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_,
    new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_,
    new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_,
    new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_,
    new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_,
    new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_,
    new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_,
    new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_,
    new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_,
    new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_,
    new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_,
    new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_,
    new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_,
    new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_,
    new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_,
    new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_,
    new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_,
    new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_,
    new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_,
    new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_,
    new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_,
    new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_,
    new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_,
    new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_,
    new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_,
    new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_,
    new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_,
    new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_,
    new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_,
    new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_,
    new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_,
    new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8065_,
    new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_,
    new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_,
    new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_,
    new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_,
    new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_,
    new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_,
    new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_,
    new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_,
    new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_,
    new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_,
    new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_,
    new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_,
    new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_,
    new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_,
    new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_,
    new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_,
    new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_,
    new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_,
    new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_,
    new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_,
    new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_,
    new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_,
    new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_,
    new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_,
    new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_,
    new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_,
    new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_,
    new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_,
    new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_,
    new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_,
    new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_,
    new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_,
    new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_,
    new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_,
    new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_,
    new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_,
    new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_,
    new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_,
    new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_,
    new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_,
    new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_,
    new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_,
    new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_,
    new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_,
    new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_,
    new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_,
    new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_,
    new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_,
    new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_,
    new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_,
    new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_,
    new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_,
    new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8569_,
    new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_,
    new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_,
    new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_,
    new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_,
    new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_,
    new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_,
    new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_,
    new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_,
    new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_,
    new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_,
    new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_,
    new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_,
    new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_,
    new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_,
    new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_,
    new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_,
    new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_,
    new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_,
    new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_,
    new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_,
    new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_,
    new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_,
    new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_,
    new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_,
    new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_,
    new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_,
    new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_,
    new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_,
    new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_,
    new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_,
    new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_,
    new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_,
    new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_,
    new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_,
    new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_,
    new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_,
    new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_,
    new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_,
    new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_,
    new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_,
    new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_,
    new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_,
    new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_,
    new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n10283_, new_n10284_, new_n10285_, new_n10286_,
    new_n10287_, new_n10288_, new_n10289_, new_n10290_, new_n10291_,
    new_n10292_, new_n10293_, new_n10294_, new_n10295_, new_n10296_,
    new_n10297_, new_n10298_, new_n10299_, new_n10300_, new_n10301_,
    new_n10302_, new_n10303_, new_n10304_, new_n10305_, new_n10306_,
    new_n10307_, new_n10308_, new_n10309_, new_n10310_, new_n10311_,
    new_n10312_, new_n10313_, new_n10314_, new_n10315_, new_n10316_,
    new_n10317_, new_n10318_, new_n10319_, new_n10320_, new_n10321_,
    new_n10322_, new_n10323_, new_n10324_, new_n10325_, new_n10326_,
    new_n10327_, new_n10328_, new_n10329_, new_n10330_, new_n10331_,
    new_n10332_, new_n10333_, new_n10334_, new_n10335_, new_n10336_,
    new_n10337_, new_n10338_, new_n10339_, new_n10340_, new_n10341_,
    new_n10342_, new_n10343_, new_n10344_, new_n10345_, new_n10346_,
    new_n10347_, new_n10348_, new_n10349_, new_n10350_, new_n10351_,
    new_n10352_, new_n10353_, new_n10354_, new_n10355_, new_n10356_,
    new_n10357_, new_n10358_, new_n10359_, new_n10360_, new_n10361_,
    new_n10362_, new_n10363_, new_n10364_, new_n10365_, new_n10366_,
    new_n10367_, new_n10368_, new_n10369_, new_n10370_, new_n10371_,
    new_n10372_, new_n10373_, new_n10374_, new_n10375_, new_n10376_,
    new_n10377_, new_n10378_, new_n10379_, new_n10380_, new_n10381_,
    new_n10382_, new_n10383_, new_n10384_, new_n10385_, new_n10386_,
    new_n10387_, new_n10388_, new_n10389_, new_n10390_, new_n10391_,
    new_n10392_, new_n10393_, new_n10394_, new_n10395_, new_n10396_,
    new_n10397_, new_n10398_, new_n10399_, new_n10400_, new_n10401_,
    new_n10402_, new_n10403_, new_n10404_, new_n10405_, new_n10406_,
    new_n10407_, new_n10408_, new_n10409_, new_n10410_, new_n10411_,
    new_n10412_, new_n10413_, new_n10414_, new_n10415_, new_n10416_,
    new_n10417_, new_n10418_, new_n10419_, new_n10420_, new_n10421_,
    new_n10422_, new_n10423_, new_n10424_, new_n10425_, new_n10426_,
    new_n10427_, new_n10428_, new_n10429_, new_n10430_, new_n10431_,
    new_n10432_, new_n10433_, new_n10434_, new_n10435_, new_n10436_,
    new_n10437_, new_n10438_, new_n10439_, new_n10440_, new_n10441_,
    new_n10442_, new_n10443_, new_n10444_, new_n10445_, new_n10446_,
    new_n10447_, new_n10448_, new_n10449_, new_n10450_, new_n10451_,
    new_n10452_, new_n10453_, new_n10454_, new_n10455_, new_n10456_,
    new_n10457_, new_n10458_, new_n10459_, new_n10460_, new_n10461_,
    new_n10462_, new_n10463_, new_n10464_, new_n10465_, new_n10466_,
    new_n10467_, new_n10468_, new_n10469_, new_n10470_, new_n10471_,
    new_n10472_, new_n10473_, new_n10474_, new_n10475_, new_n10476_,
    new_n10477_, new_n10478_, new_n10479_, new_n10480_, new_n10481_,
    new_n10482_, new_n10483_, new_n10484_, new_n10485_, new_n10486_,
    new_n10487_, new_n10488_, new_n10489_, new_n10490_, new_n10491_,
    new_n10492_, new_n10493_, new_n10494_, new_n10495_, new_n10496_,
    new_n10497_, new_n10498_, new_n10499_, new_n10500_, new_n10501_,
    new_n10502_, new_n10503_, new_n10504_, new_n10505_, new_n10506_,
    new_n10507_, new_n10508_, new_n10509_, new_n10510_, new_n10511_,
    new_n10512_, new_n10513_, new_n10514_, new_n10515_, new_n10516_,
    new_n10517_, new_n10518_, new_n10519_, new_n10520_, new_n10521_,
    new_n10522_, new_n10523_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10530_, new_n10531_,
    new_n10532_, new_n10533_, new_n10534_, new_n10535_, new_n10536_,
    new_n10537_, new_n10538_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10590_, new_n10591_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10615_, new_n10616_,
    new_n10617_, new_n10618_, new_n10619_, new_n10620_, new_n10621_,
    new_n10622_, new_n10623_, new_n10624_, new_n10625_, new_n10630_,
    new_n10631_, new_n10635_, new_n10638_, new_n10639_, new_n10647_,
    new_n10648_, new_n10654_, new_n10655_, new_n10656_, new_n10657_,
    new_n10658_, new_n10659_, new_n10660_, new_n10661_, new_n10662_,
    new_n10663_, new_n10664_, new_n10665_, new_n10666_, new_n10667_,
    new_n10668_, new_n10669_, new_n10670_, new_n10671_, new_n10672_,
    new_n10673_, new_n10674_, new_n10675_, new_n10676_, new_n10677_,
    new_n10678_, new_n10679_, new_n10680_, new_n10681_, new_n10682_,
    new_n10683_, new_n10684_, new_n10685_, new_n10686_, new_n10687_,
    new_n10688_, new_n10689_, new_n10690_, new_n10691_, new_n10692_,
    new_n10693_, new_n10694_, new_n10695_, new_n10696_, new_n10697_,
    new_n10698_, new_n10699_, new_n10700_, new_n10701_, new_n10702_,
    new_n10703_, new_n10704_, new_n10705_, new_n10706_, new_n10707_,
    new_n10708_, new_n10709_, new_n10710_, new_n10711_, new_n10712_,
    new_n10713_, new_n10714_, new_n10715_, new_n10716_, new_n10717_,
    new_n10718_, new_n10719_, new_n10720_, new_n10721_, new_n10722_,
    new_n10723_, new_n10724_, new_n10725_, new_n10726_, new_n10727_,
    new_n10728_, new_n10729_, new_n10730_, new_n10731_, new_n10732_,
    new_n10733_, new_n10734_, new_n10735_, new_n10736_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10743_, new_n10744_, new_n10745_, new_n10746_, new_n10747_,
    new_n10748_, new_n10749_, new_n10750_, new_n10751_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10757_,
    new_n10758_, new_n10759_, new_n10760_, new_n10761_, new_n10762_,
    new_n10763_, new_n10764_, new_n10765_, new_n10766_, new_n10767_,
    new_n10768_, new_n10769_, new_n10770_, new_n10771_, new_n10772_,
    new_n10773_, new_n10774_, new_n10775_, new_n10776_, new_n10777_,
    new_n10778_, new_n10779_, new_n10780_, new_n10781_, new_n10782_,
    new_n10783_, new_n10784_, new_n10785_, new_n10786_, new_n10787_,
    new_n10788_, new_n10789_, new_n10790_, new_n10791_, new_n10792_,
    new_n10793_, new_n10794_, new_n10795_, new_n10796_, new_n10797_,
    new_n10798_, new_n10799_, new_n10800_, new_n10801_, new_n10802_,
    new_n10803_, new_n10804_, new_n10805_, new_n10806_, new_n10807_,
    new_n10808_, new_n10809_, new_n10810_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10863_, new_n10864_, new_n10865_, new_n10866_, new_n10867_,
    new_n10868_, new_n10869_, new_n10870_, new_n10871_, new_n10872_,
    new_n10873_, new_n10874_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10880_, new_n10881_, new_n10882_,
    new_n10883_, new_n10884_, new_n10885_, new_n10886_, new_n10887_,
    new_n10888_, new_n10889_, new_n10890_, new_n10891_, new_n10892_,
    new_n10893_, new_n10894_, new_n10895_, new_n10896_, new_n10897_,
    new_n10898_, new_n10899_, new_n10900_, new_n10901_, new_n10902_,
    new_n10903_, new_n10904_, new_n10905_, new_n10906_, new_n10907_,
    new_n10908_, new_n10909_, new_n10910_, new_n10911_, new_n10912_,
    new_n10913_, new_n10914_, new_n10915_, new_n10916_, new_n10917_,
    new_n10918_, new_n10919_, new_n10920_, new_n10921_, new_n10922_,
    new_n10923_, new_n10924_, new_n10925_, new_n10926_, new_n10927_,
    new_n10928_, new_n10929_, new_n10930_, new_n10931_, new_n10932_,
    new_n10933_, new_n10934_, new_n10935_, new_n10936_, new_n10937_,
    new_n10938_, new_n10939_, new_n10940_, new_n10941_, new_n10942_,
    new_n10943_, new_n10944_, new_n10945_, new_n10946_, new_n10947_,
    new_n10948_, new_n10949_, new_n10950_, new_n10951_, new_n10952_,
    new_n10953_, new_n10954_, new_n10955_, new_n10956_, new_n10957_,
    new_n10958_, new_n10959_, new_n10960_, new_n10961_, new_n10962_,
    new_n10963_, new_n10964_, new_n10965_, new_n10966_, new_n10967_,
    new_n10968_, new_n10969_, new_n10970_, new_n10971_, new_n10972_,
    new_n10973_, new_n10974_, new_n10975_, new_n10976_, new_n10977_,
    new_n10978_, new_n10979_, new_n10980_, new_n10981_, new_n10982_,
    new_n10983_, new_n10984_, new_n10985_, new_n10986_, new_n10987_,
    new_n10988_, new_n10989_, new_n10990_, new_n10991_, new_n10992_,
    new_n10993_, new_n10994_, new_n10995_, new_n10996_, new_n10997_,
    new_n10998_, new_n10999_, new_n11000_, new_n11001_, new_n11002_,
    new_n11003_, new_n11004_, new_n11005_, new_n11006_, new_n11007_,
    new_n11008_, new_n11009_, new_n11010_, new_n11011_, new_n11012_,
    new_n11013_, new_n11014_, new_n11015_, new_n11016_, new_n11017_,
    new_n11018_, new_n11019_, new_n11020_, new_n11021_, new_n11022_,
    new_n11023_, new_n11024_, new_n11025_, new_n11026_, new_n11027_,
    new_n11028_, new_n11029_, new_n11030_, new_n11031_, new_n11032_,
    new_n11033_, new_n11034_, new_n11035_, new_n11036_, new_n11037_,
    new_n11038_, new_n11039_, new_n11040_, new_n11041_, new_n11042_,
    new_n11043_, new_n11044_, new_n11045_, new_n11046_, new_n11047_,
    new_n11048_, new_n11049_, new_n11050_, new_n11051_, new_n11052_,
    new_n11053_, new_n11054_, new_n11055_, new_n11056_, new_n11057_,
    new_n11058_, new_n11059_, new_n11060_, new_n11061_, new_n11062_,
    new_n11063_, new_n11064_, new_n11065_, new_n11066_, new_n11067_,
    new_n11068_, new_n11069_, new_n11070_, new_n11071_, new_n11072_,
    new_n11073_, new_n11074_, new_n11075_, new_n11076_, new_n11077_,
    new_n11078_, new_n11079_, new_n11080_, new_n11081_, new_n11082_,
    new_n11083_, new_n11084_, new_n11085_, new_n11086_, new_n11087_,
    new_n11088_, new_n11089_, new_n11090_, new_n11091_, new_n11092_,
    new_n11093_, new_n11094_, new_n11095_, new_n11096_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11101_, new_n11102_,
    new_n11103_, new_n11104_, new_n11105_, new_n11106_, new_n11107_,
    new_n11108_, new_n11109_, new_n11110_, new_n11111_, new_n11112_,
    new_n11113_, new_n11114_, new_n11115_, new_n11116_, new_n11117_,
    new_n11118_, new_n11119_, new_n11120_, new_n11121_, new_n11122_,
    new_n11123_, new_n11124_, new_n11125_, new_n11126_, new_n11127_,
    new_n11128_, new_n11129_, new_n11130_, new_n11131_, new_n11132_,
    new_n11133_, new_n11134_, new_n11135_, new_n11136_, new_n11137_,
    new_n11138_, new_n11139_, new_n11140_, new_n11141_, new_n11142_,
    new_n11143_, new_n11144_, new_n11145_, new_n11146_, new_n11147_,
    new_n11148_, new_n11149_, new_n11150_, new_n11151_, new_n11152_,
    new_n11153_, new_n11154_, new_n11155_, new_n11156_, new_n11157_,
    new_n11158_, new_n11159_, new_n11160_, new_n11161_, new_n11162_,
    new_n11163_, new_n11164_, new_n11165_, new_n11166_, new_n11167_,
    new_n11168_, new_n11169_, new_n11170_, new_n11171_, new_n11172_,
    new_n11173_, new_n11174_, new_n11175_, new_n11176_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11205_, new_n11206_, new_n11207_,
    new_n11208_, new_n11209_, new_n11210_, new_n11211_, new_n11212_,
    new_n11213_, new_n11214_, new_n11215_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11236_, new_n11237_,
    new_n11238_, new_n11239_, new_n11240_, new_n11241_, new_n11242_,
    new_n11243_, new_n11244_, new_n11245_, new_n11246_, new_n11247_,
    new_n11248_, new_n11249_, new_n11250_, new_n11251_, new_n11252_,
    new_n11253_, new_n11254_, new_n11255_, new_n11256_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11262_,
    new_n11263_, new_n11264_, new_n11265_, new_n11266_, new_n11267_,
    new_n11268_, new_n11269_, new_n11270_, new_n11271_, new_n11272_,
    new_n11273_, new_n11274_, new_n11275_, new_n11276_, new_n11277_,
    new_n11278_, new_n11279_, new_n11280_, new_n11281_, new_n11282_,
    new_n11283_, new_n11284_, new_n11285_, new_n11286_, new_n11287_,
    new_n11288_, new_n11289_, new_n11290_, new_n11291_, new_n11292_,
    new_n11293_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11310_, new_n11311_, new_n11312_,
    new_n11313_, new_n11314_, new_n11315_, new_n11316_, new_n11317_,
    new_n11318_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11435_, new_n11436_, new_n11437_,
    new_n11438_, new_n11439_, new_n11440_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11451_, new_n11452_,
    new_n11453_, new_n11454_, new_n11455_, new_n11456_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11591_, new_n11592_,
    new_n11593_, new_n11594_, new_n11595_, new_n11596_, new_n11597_,
    new_n11598_, new_n11599_, new_n11600_, new_n11601_, new_n11602_,
    new_n11603_, new_n11604_, new_n11605_, new_n11606_, new_n11607_,
    new_n11608_, new_n11609_, new_n11610_, new_n11611_, new_n11612_,
    new_n11613_, new_n11614_, new_n11615_, new_n11616_, new_n11617_,
    new_n11618_, new_n11619_, new_n11620_, new_n11621_, new_n11622_,
    new_n11623_, new_n11624_, new_n11625_, new_n11626_, new_n11627_,
    new_n11628_, new_n11629_, new_n11630_, new_n11631_, new_n11632_,
    new_n11633_, new_n11634_, new_n11635_, new_n11636_, new_n11637_,
    new_n11638_, new_n11639_, new_n11640_, new_n11641_, new_n11642_,
    new_n11643_, new_n11644_, new_n11645_, new_n11646_, new_n11647_,
    new_n11648_, new_n11649_, new_n11650_, new_n11651_, new_n11652_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11663_, new_n11664_, new_n11665_, new_n11666_, new_n11667_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11878_, new_n11879_, new_n11880_, new_n11881_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11966_, new_n11967_,
    new_n11968_, new_n11969_, new_n11970_, new_n11971_, new_n11972_,
    new_n11973_, new_n11974_, new_n11975_, new_n11976_, new_n11977_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11988_, new_n11989_, new_n11990_, new_n11991_, new_n11992_,
    new_n11993_, new_n11994_, new_n11995_, new_n11996_, new_n11997_,
    new_n11998_, new_n11999_, new_n12000_, new_n12001_, new_n12002_,
    new_n12003_, new_n12004_, new_n12005_, new_n12006_, new_n12007_,
    new_n12008_, new_n12009_, new_n12010_, new_n12011_, new_n12012_,
    new_n12013_, new_n12014_, new_n12015_, new_n12016_, new_n12017_,
    new_n12018_, new_n12019_, new_n12020_, new_n12021_, new_n12022_,
    new_n12023_, new_n12024_, new_n12025_, new_n12026_, new_n12027_,
    new_n12028_, new_n12029_, new_n12030_, new_n12031_, new_n12032_,
    new_n12033_, new_n12034_, new_n12035_, new_n12036_, new_n12037_,
    new_n12038_, new_n12039_, new_n12040_, new_n12041_, new_n12042_,
    new_n12043_, new_n12044_, new_n12045_, new_n12046_, new_n12047_,
    new_n12048_, new_n12049_, new_n12050_, new_n12051_, new_n12052_,
    new_n12053_, new_n12054_, new_n12055_, new_n12056_, new_n12057_,
    new_n12058_, new_n12059_, new_n12060_, new_n12061_, new_n12062_,
    new_n12063_, new_n12064_, new_n12065_, new_n12066_, new_n12067_,
    new_n12068_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12073_, new_n12074_, new_n12075_, new_n12076_, new_n12077_,
    new_n12078_, new_n12079_, new_n12080_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12164_, new_n12165_, new_n12166_, new_n12167_,
    new_n12168_, new_n12169_, new_n12170_, new_n12171_, new_n12172_,
    new_n12173_, new_n12174_, new_n12175_, new_n12176_, new_n12177_,
    new_n12178_, new_n12179_, new_n12180_, new_n12181_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12226_, new_n12227_,
    new_n12228_, new_n12229_, new_n12230_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12238_, new_n12239_, new_n12240_, new_n12241_, new_n12242_,
    new_n12243_, new_n12244_, new_n12245_, new_n12246_, new_n12247_,
    new_n12248_, new_n12249_, new_n12250_, new_n12251_, new_n12252_,
    new_n12253_, new_n12254_, new_n12255_, new_n12256_, new_n12257_,
    new_n12258_, new_n12259_, new_n12260_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12290_, new_n12291_, new_n12292_,
    new_n12293_, new_n12294_, new_n12295_, new_n12296_, new_n12297_,
    new_n12298_, new_n12299_, new_n12300_, new_n12301_, new_n12302_,
    new_n12303_, new_n12304_, new_n12305_, new_n12306_, new_n12307_,
    new_n12308_, new_n12309_, new_n12310_, new_n12311_, new_n12312_,
    new_n12313_, new_n12314_, new_n12315_, new_n12316_, new_n12317_,
    new_n12318_, new_n12319_, new_n12320_, new_n12321_, new_n12322_,
    new_n12323_, new_n12324_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12417_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12428_, new_n12429_, new_n12430_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12438_, new_n12439_, new_n12440_, new_n12441_, new_n12442_,
    new_n12443_, new_n12444_, new_n12445_, new_n12446_, new_n12447_,
    new_n12448_, new_n12449_, new_n12450_, new_n12451_, new_n12452_,
    new_n12453_, new_n12454_, new_n12455_, new_n12456_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12463_, new_n12464_, new_n12465_, new_n12466_, new_n12467_,
    new_n12468_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12528_, new_n12529_, new_n12530_, new_n12531_, new_n12532_,
    new_n12533_, new_n12534_, new_n12535_, new_n12536_, new_n12537_,
    new_n12538_, new_n12539_, new_n12540_, new_n12541_, new_n12542_,
    new_n12543_, new_n12544_, new_n12545_, new_n12546_, new_n12547_,
    new_n12548_, new_n12549_, new_n12550_, new_n12551_, new_n12552_,
    new_n12553_, new_n12554_, new_n12555_, new_n12556_, new_n12557_,
    new_n12558_, new_n12559_, new_n12560_, new_n12561_, new_n12562_,
    new_n12563_, new_n12564_, new_n12565_, new_n12566_, new_n12567_,
    new_n12568_, new_n12569_, new_n12570_, new_n12571_, new_n12572_,
    new_n12573_, new_n12574_, new_n12575_, new_n12576_, new_n12577_,
    new_n12578_, new_n12579_, new_n12580_, new_n12581_, new_n12582_,
    new_n12583_, new_n12584_, new_n12585_, new_n12586_, new_n12587_,
    new_n12588_, new_n12589_, new_n12590_, new_n12591_, new_n12592_,
    new_n12593_, new_n12594_, new_n12595_, new_n12596_, new_n12597_,
    new_n12598_, new_n12599_, new_n12600_, new_n12601_, new_n12602_,
    new_n12603_, new_n12604_, new_n12605_, new_n12606_, new_n12607_,
    new_n12608_, new_n12609_, new_n12610_, new_n12611_, new_n12612_,
    new_n12613_, new_n12614_, new_n12615_, new_n12616_, new_n12617_,
    new_n12618_, new_n12619_, new_n12620_, new_n12621_, new_n12622_,
    new_n12623_, new_n12624_, new_n12625_, new_n12626_, new_n12627_,
    new_n12628_, new_n12629_, new_n12630_, new_n12631_, new_n12632_,
    new_n12633_, new_n12634_, new_n12635_, new_n12636_, new_n12637_,
    new_n12638_, new_n12639_, new_n12640_, new_n12641_, new_n12642_,
    new_n12643_, new_n12644_, new_n12645_, new_n12646_, new_n12647_,
    new_n12648_, new_n12649_, new_n12650_, new_n12651_, new_n12652_,
    new_n12653_, new_n12654_, new_n12655_, new_n12656_, new_n12657_,
    new_n12658_, new_n12659_, new_n12660_, new_n12661_, new_n12662_,
    new_n12663_, new_n12664_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12766_, new_n12767_,
    new_n12768_, new_n12769_, new_n12770_, new_n12771_, new_n12772_,
    new_n12773_, new_n12774_, new_n12775_, new_n12776_, new_n12777_,
    new_n12778_, new_n12779_, new_n12780_, new_n12781_, new_n12782_,
    new_n12783_, new_n12784_, new_n12785_, new_n12786_, new_n12787_,
    new_n12788_, new_n12789_, new_n12790_, new_n12791_, new_n12792_,
    new_n12793_, new_n12794_, new_n12795_, new_n12796_, new_n12797_,
    new_n12798_, new_n12799_, new_n12800_, new_n12801_, new_n12802_,
    new_n12803_, new_n12804_, new_n12805_, new_n12806_, new_n12807_,
    new_n12808_, new_n12809_, new_n12810_, new_n12811_, new_n12812_,
    new_n12813_, new_n12814_, new_n12815_, new_n12816_, new_n12817_,
    new_n12818_, new_n12819_, new_n12820_, new_n12821_, new_n12822_,
    new_n12823_, new_n12824_, new_n12825_, new_n12826_, new_n12827_,
    new_n12828_, new_n12829_, new_n12830_, new_n12831_, new_n12832_,
    new_n12833_, new_n12834_, new_n12835_, new_n12836_, new_n12837_,
    new_n12838_, new_n12839_, new_n12840_, new_n12841_, new_n12842_,
    new_n12843_, new_n12844_, new_n12845_, new_n12846_, new_n12847_,
    new_n12848_, new_n12849_, new_n12850_, new_n12851_, new_n12852_,
    new_n12853_, new_n12854_, new_n12855_, new_n12856_, new_n12857_,
    new_n12858_, new_n12859_, new_n12860_, new_n12861_, new_n12862_,
    new_n12863_, new_n12864_, new_n12865_, new_n12866_, new_n12867_,
    new_n12868_, new_n12869_, new_n12870_, new_n12871_, new_n12872_,
    new_n12873_, new_n12874_, new_n12875_, new_n12876_, new_n12877_,
    new_n12878_, new_n12879_, new_n12880_, new_n12881_, new_n12882_,
    new_n12883_, new_n12884_, new_n12885_, new_n12886_, new_n12887_,
    new_n12888_, new_n12889_, new_n12890_, new_n12891_, new_n12892_,
    new_n12893_, new_n12894_, new_n12895_, new_n12896_, new_n12897_,
    new_n12898_, new_n12899_, new_n12900_, new_n12901_, new_n12902_,
    new_n12903_, new_n12904_, new_n12905_, new_n12906_, new_n12907_,
    new_n12908_, new_n12909_, new_n12910_, new_n12911_, new_n12912_,
    new_n12913_, new_n12914_, new_n12915_, new_n12916_, new_n12917_,
    new_n12918_, new_n12919_, new_n12920_, new_n12921_, new_n12922_,
    new_n12923_, new_n12924_, new_n12925_, new_n12926_, new_n12927_,
    new_n12928_, new_n12929_, new_n12930_, new_n12931_, new_n12932_,
    new_n12933_, new_n12934_, new_n12935_, new_n12936_, new_n12937_,
    new_n12938_, new_n12939_, new_n12940_, new_n12941_, new_n12942_,
    new_n12943_, new_n12944_, new_n12945_, new_n12946_, new_n12947_,
    new_n12948_, new_n12949_, new_n12950_, new_n12951_, new_n12952_,
    new_n12953_, new_n12954_, new_n12955_, new_n12956_, new_n12957_,
    new_n12958_, new_n12959_, new_n12960_, new_n12961_, new_n12962_,
    new_n12963_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12993_, new_n12994_, new_n12995_, new_n12996_, new_n12997_,
    new_n12998_, new_n12999_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13009_, new_n13010_, new_n13011_, new_n13012_,
    new_n13013_, new_n13014_, new_n13015_, new_n13016_, new_n13017_,
    new_n13018_, new_n13019_, new_n13020_, new_n13021_, new_n13022_,
    new_n13023_, new_n13024_, new_n13025_, new_n13026_, new_n13027_,
    new_n13028_, new_n13029_, new_n13030_, new_n13031_, new_n13032_,
    new_n13033_, new_n13034_, new_n13035_, new_n13036_, new_n13037_,
    new_n13038_, new_n13039_, new_n13040_, new_n13041_, new_n13042_,
    new_n13043_, new_n13044_, new_n13045_, new_n13046_, new_n13047_,
    new_n13048_, new_n13049_, new_n13050_, new_n13051_, new_n13052_,
    new_n13053_, new_n13054_, new_n13055_, new_n13056_, new_n13057_,
    new_n13058_, new_n13059_, new_n13060_, new_n13061_, new_n13062_,
    new_n13063_, new_n13064_, new_n13065_, new_n13066_, new_n13067_,
    new_n13068_, new_n13069_, new_n13070_, new_n13071_, new_n13072_,
    new_n13073_, new_n13074_, new_n13075_, new_n13076_, new_n13077_,
    new_n13078_, new_n13079_, new_n13080_, new_n13081_, new_n13082_,
    new_n13083_, new_n13084_, new_n13085_, new_n13086_, new_n13087_,
    new_n13088_, new_n13089_, new_n13090_, new_n13091_, new_n13092_,
    new_n13093_, new_n13094_, new_n13095_, new_n13096_, new_n13097_,
    new_n13098_, new_n13099_, new_n13100_, new_n13101_, new_n13102_,
    new_n13103_, new_n13104_, new_n13105_, new_n13106_, new_n13107_,
    new_n13108_, new_n13109_, new_n13110_, new_n13111_, new_n13112_,
    new_n13113_, new_n13114_, new_n13115_, new_n13116_, new_n13117_,
    new_n13118_, new_n13119_, new_n13120_, new_n13121_, new_n13122_,
    new_n13123_, new_n13124_, new_n13125_, new_n13126_, new_n13127_,
    new_n13128_, new_n13129_, new_n13130_, new_n13131_, new_n13132_,
    new_n13133_, new_n13134_, new_n13135_, new_n13136_, new_n13137_,
    new_n13138_, new_n13139_, new_n13140_, new_n13141_, new_n13142_,
    new_n13143_, new_n13144_, new_n13145_, new_n13146_, new_n13147_,
    new_n13148_, new_n13149_, new_n13150_, new_n13151_, new_n13152_,
    new_n13153_, new_n13154_, new_n13155_, new_n13156_, new_n13157_,
    new_n13158_, new_n13159_, new_n13160_, new_n13161_, new_n13162_,
    new_n13163_, new_n13164_, new_n13165_, new_n13166_, new_n13167_,
    new_n13168_, new_n13169_, new_n13170_, new_n13171_, new_n13172_,
    new_n13173_, new_n13174_, new_n13175_, new_n13176_, new_n13177_,
    new_n13178_, new_n13179_, new_n13180_, new_n13181_, new_n13182_,
    new_n13183_, new_n13184_, new_n13185_, new_n13186_, new_n13187_,
    new_n13188_, new_n13189_, new_n13190_, new_n13191_, new_n13192_,
    new_n13193_, new_n13194_, new_n13195_, new_n13196_, new_n13197_,
    new_n13198_, new_n13199_, new_n13200_, new_n13201_, new_n13202_,
    new_n13203_, new_n13204_, new_n13205_, new_n13206_, new_n13207_,
    new_n13208_, new_n13209_, new_n13210_, new_n13211_, new_n13212_,
    new_n13213_, new_n13214_, new_n13215_, new_n13216_, new_n13217_,
    new_n13218_, new_n13219_, new_n13220_, new_n13221_, new_n13222_,
    new_n13223_, new_n13224_, new_n13225_, new_n13226_, new_n13227_,
    new_n13228_, new_n13229_, new_n13230_, new_n13231_, new_n13232_,
    new_n13233_, new_n13234_, new_n13235_, new_n13236_, new_n13237_,
    new_n13238_, new_n13239_, new_n13240_, new_n13241_, new_n13242_,
    new_n13243_, new_n13244_, new_n13245_, new_n13246_, new_n13247_,
    new_n13248_, new_n13249_, new_n13250_, new_n13251_, new_n13252_,
    new_n13253_, new_n13254_, new_n13255_, new_n13256_, new_n13257_,
    new_n13258_, new_n13259_, new_n13260_, new_n13261_, new_n13262_,
    new_n13263_, new_n13264_, new_n13265_, new_n13266_, new_n13267_,
    new_n13268_, new_n13269_, new_n13270_, new_n13271_, new_n13272_,
    new_n13273_, new_n13274_, new_n13275_, new_n13276_, new_n13277_,
    new_n13278_, new_n13279_, new_n13280_, new_n13281_, new_n13282_,
    new_n13283_, new_n13284_, new_n13285_, new_n13286_, new_n13287_,
    new_n13288_, new_n13289_, new_n13290_, new_n13291_, new_n13292_,
    new_n13293_, new_n13294_, new_n13295_, new_n13296_, new_n13297_,
    new_n13298_, new_n13299_, new_n13300_, new_n13301_, new_n13302_,
    new_n13303_, new_n13304_, new_n13305_, new_n13306_, new_n13307_,
    new_n13308_, new_n13309_, new_n13310_, new_n13311_, new_n13312_,
    new_n13313_, new_n13314_, new_n13315_, new_n13316_, new_n13317_,
    new_n13318_, new_n13319_, new_n13320_, new_n13321_, new_n13322_,
    new_n13323_, new_n13324_, new_n13325_, new_n13326_, new_n13327_,
    new_n13328_, new_n13329_, new_n13330_, new_n13331_, new_n13332_,
    new_n13333_, new_n13334_, new_n13335_, new_n13336_, new_n13337_,
    new_n13338_, new_n13339_, new_n13340_, new_n13341_, new_n13342_,
    new_n13343_, new_n13344_, new_n13345_, new_n13346_, new_n13347_,
    new_n13348_, new_n13349_, new_n13350_, new_n13351_, new_n13352_,
    new_n13353_, new_n13354_, new_n13355_, new_n13356_, new_n13357_,
    new_n13358_, new_n13359_, new_n13360_, new_n13361_, new_n13362_,
    new_n13363_, new_n13364_, new_n13365_, new_n13366_, new_n13367_,
    new_n13368_, new_n13369_, new_n13370_, new_n13371_, new_n13372_,
    new_n13373_, new_n13374_, new_n13375_, new_n13376_, new_n13377_,
    new_n13378_, new_n13379_, new_n13380_, new_n13381_, new_n13382_,
    new_n13383_, new_n13384_, new_n13385_, new_n13386_, new_n13387_,
    new_n13388_, new_n13389_, new_n13390_, new_n13391_, new_n13392_,
    new_n13393_, new_n13394_, new_n13395_, new_n13396_, new_n13397_,
    new_n13398_, new_n13399_, new_n13400_, new_n13401_, new_n13402_,
    new_n13403_, new_n13404_, new_n13405_, new_n13406_, new_n13407_,
    new_n13408_, new_n13409_, new_n13410_, new_n13411_, new_n13412_,
    new_n13413_, new_n13414_, new_n13415_, new_n13416_, new_n13417_,
    new_n13418_, new_n13419_, new_n13420_, new_n13421_, new_n13422_,
    new_n13423_, new_n13424_, new_n13425_, new_n13426_, new_n13427_,
    new_n13428_, new_n13429_, new_n13430_, new_n13431_, new_n13432_,
    new_n13433_, new_n13434_, new_n13435_, new_n13436_, new_n13437_,
    new_n13438_, new_n13439_, new_n13440_, new_n13441_, new_n13442_,
    new_n13443_, new_n13444_, new_n13445_, new_n13446_, new_n13447_,
    new_n13448_, new_n13449_, new_n13450_, new_n13451_, new_n13452_,
    new_n13453_, new_n13454_, new_n13455_, new_n13456_, new_n13457_,
    new_n13458_, new_n13459_, new_n13460_, new_n13461_, new_n13462_,
    new_n13463_, new_n13464_, new_n13465_, new_n13466_, new_n13467_,
    new_n13468_, new_n13469_, new_n13470_, new_n13471_, new_n13472_,
    new_n13473_, new_n13474_, new_n13475_, new_n13476_, new_n13477_,
    new_n13478_, new_n13479_, new_n13480_, new_n13481_, new_n13482_,
    new_n13483_, new_n13484_, new_n13485_, new_n13486_, new_n13487_,
    new_n13488_, new_n13489_, new_n13490_, new_n13491_, new_n13492_,
    new_n13493_, new_n13494_, new_n13495_, new_n13496_, new_n13497_,
    new_n13498_, new_n13499_, new_n13500_, new_n13501_, new_n13502_,
    new_n13503_, new_n13504_, new_n13505_, new_n13506_, new_n13507_,
    new_n13508_, new_n13509_, new_n13510_, new_n13511_, new_n13512_,
    new_n13513_, new_n13514_, new_n13515_, new_n13516_, new_n13517_,
    new_n13518_, new_n13519_, new_n13520_, new_n13521_, new_n13522_,
    new_n13523_, new_n13524_, new_n13525_, new_n13526_, new_n13527_,
    new_n13528_, new_n13529_, new_n13530_, new_n13531_, new_n13532_,
    new_n13533_, new_n13534_, new_n13535_, new_n13536_, new_n13537_,
    new_n13538_, new_n13539_, new_n13540_, new_n13541_, new_n13542_,
    new_n13543_, new_n13544_, new_n13545_, new_n13546_, new_n13547_,
    new_n13548_, new_n13549_, new_n13550_, new_n13551_, new_n13552_,
    new_n13553_, new_n13554_, new_n13555_, new_n13556_, new_n13557_,
    new_n13558_, new_n13559_, new_n13560_, new_n13561_, new_n13562_,
    new_n13563_, new_n13564_, new_n13565_, new_n13566_, new_n13567_,
    new_n13568_, new_n13569_, new_n13570_, new_n13571_, new_n13572_,
    new_n13573_, new_n13574_, new_n13575_, new_n13576_, new_n13577_,
    new_n13578_, new_n13579_, new_n13580_, new_n13581_, new_n13582_,
    new_n13583_, new_n13584_, new_n13585_, new_n13586_, new_n13587_,
    new_n13588_, new_n13589_, new_n13590_, new_n13591_, new_n13592_,
    new_n13593_, new_n13594_, new_n13595_, new_n13596_, new_n13597_,
    new_n13598_, new_n13599_, new_n13600_, new_n13601_, new_n13602_,
    new_n13603_, new_n13604_, new_n13605_, new_n13606_, new_n13607_,
    new_n13608_, new_n13609_, new_n13610_, new_n13611_, new_n13612_,
    new_n13613_, new_n13614_, new_n13615_, new_n13616_, new_n13617_,
    new_n13618_, new_n13619_, new_n13620_, new_n13621_, new_n13622_,
    new_n13623_, new_n13624_, new_n13625_, new_n13626_, new_n13627_,
    new_n13628_, new_n13629_, new_n13630_, new_n13631_, new_n13632_,
    new_n13633_, new_n13634_, new_n13635_, new_n13636_, new_n13637_,
    new_n13638_, new_n13639_, new_n13640_, new_n13641_, new_n13642_,
    new_n13643_, new_n13644_, new_n13645_, new_n13646_, new_n13647_,
    new_n13648_, new_n13649_, new_n13650_, new_n13651_, new_n13652_,
    new_n13653_, new_n13654_, new_n13655_, new_n13656_, new_n13657_,
    new_n13658_, new_n13659_, new_n13660_, new_n13661_, new_n13662_,
    new_n13663_, new_n13664_, new_n13665_, new_n13666_, new_n13667_,
    new_n13668_, new_n13669_, new_n13670_, new_n13671_, new_n13672_,
    new_n13673_, new_n13674_, new_n13675_, new_n13676_, new_n13677_,
    new_n13678_, new_n13679_, new_n13680_, new_n13681_, new_n13682_,
    new_n13683_, new_n13684_, new_n13685_, new_n13686_, new_n13687_,
    new_n13688_, new_n13689_, new_n13690_, new_n13691_, new_n13692_,
    new_n13693_, new_n13694_, new_n13695_, new_n13696_, new_n13697_,
    new_n13698_, new_n13699_, new_n13700_, new_n13701_, new_n13702_,
    new_n13703_, new_n13704_, new_n13705_, new_n13706_, new_n13707_,
    new_n13708_, new_n13709_, new_n13710_, new_n13711_, new_n13712_,
    new_n13713_, new_n13714_, new_n13715_, new_n13716_, new_n13717_,
    new_n13718_, new_n13719_, new_n13720_, new_n13721_, new_n13722_,
    new_n13723_, new_n13724_, new_n13725_, new_n13726_, new_n13727_,
    new_n13728_, new_n13729_, new_n13730_, new_n13731_, new_n13732_,
    new_n13733_, new_n13734_, new_n13735_, new_n13736_, new_n13737_,
    new_n13738_, new_n13739_, new_n13740_, new_n13741_, new_n13742_,
    new_n13743_, new_n13744_, new_n13745_, new_n13746_, new_n13747_,
    new_n13748_, new_n13749_, new_n13750_, new_n13751_, new_n13752_,
    new_n13753_, new_n13754_, new_n13755_, new_n13756_, new_n13757_,
    new_n13758_, new_n13759_, new_n13760_, new_n13761_, new_n13762_,
    new_n13763_, new_n13764_, new_n13765_, new_n13766_, new_n13767_,
    new_n13768_, new_n13769_, new_n13770_, new_n13771_, new_n13772_,
    new_n13773_, new_n13774_, new_n13775_, new_n13776_, new_n13777_,
    new_n13778_, new_n13779_, new_n13780_, new_n13781_, new_n13782_,
    new_n13783_, new_n13784_, new_n13785_, new_n13786_, new_n13787_,
    new_n13788_, new_n13789_, new_n13790_, new_n13791_, new_n13792_,
    new_n13793_, new_n13794_, new_n13795_, new_n13796_, new_n13797_,
    new_n13798_, new_n13799_, new_n13800_, new_n13801_, new_n13802_,
    new_n13803_, new_n13804_, new_n13805_, new_n13806_, new_n13807_,
    new_n13808_, new_n13809_, new_n13810_, new_n13811_, new_n13812_,
    new_n13813_, new_n13814_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13822_,
    new_n13823_, new_n13824_, new_n13825_, new_n13826_, new_n13827_,
    new_n13828_, new_n13829_, new_n13830_, new_n13831_, new_n13832_,
    new_n13833_, new_n13834_, new_n13835_, new_n13836_, new_n13837_,
    new_n13838_, new_n13839_, new_n13840_, new_n13841_, new_n13842_,
    new_n13843_, new_n13844_, new_n13845_, new_n13846_, new_n13847_,
    new_n13848_, new_n13849_, new_n13850_, new_n13851_, new_n13852_,
    new_n13853_, new_n13854_, new_n13855_, new_n13856_, new_n13857_,
    new_n13858_, new_n13859_, new_n13860_, new_n13861_, new_n13862_,
    new_n13863_, new_n13864_, new_n13865_, new_n13866_, new_n13867_,
    new_n13868_, new_n13869_, new_n13870_, new_n13871_, new_n13872_,
    new_n13873_, new_n13874_, new_n13875_, new_n13876_, new_n13877_,
    new_n13878_, new_n13879_, new_n13880_, new_n13881_, new_n13882_,
    new_n13883_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13889_, new_n13890_, new_n13891_, new_n13892_,
    new_n13893_, new_n13894_, new_n13895_, new_n13896_, new_n13897_,
    new_n13898_, new_n13899_, new_n13900_, new_n13901_, new_n13902_,
    new_n13903_, new_n13904_, new_n13905_, new_n13906_, new_n13907_,
    new_n13908_, new_n13909_, new_n13910_, new_n13911_, new_n13912_,
    new_n13913_, new_n13914_, new_n13915_, new_n13916_, new_n13917_,
    new_n13918_, new_n13919_, new_n13920_, new_n13921_, new_n13922_,
    new_n13923_, new_n13924_, new_n13925_, new_n13926_, new_n13927_,
    new_n13928_, new_n13929_, new_n13930_, new_n13931_, new_n13932_,
    new_n13933_, new_n13934_, new_n13935_, new_n13936_, new_n13937_,
    new_n13938_, new_n13939_, new_n13940_, new_n13941_, new_n13942_,
    new_n13943_, new_n13944_, new_n13945_, new_n13946_, new_n13947_,
    new_n13948_, new_n13949_, new_n13950_, new_n13951_, new_n13952_,
    new_n13953_, new_n13954_, new_n13955_, new_n13956_, new_n13957_,
    new_n13958_, new_n13959_, new_n13960_, new_n13961_, new_n13962_,
    new_n13963_, new_n13964_, new_n13965_, new_n13966_, new_n13967_,
    new_n13968_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14044_, new_n14045_, new_n14046_, new_n14047_,
    new_n14048_, new_n14049_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14055_, new_n14056_, new_n14057_,
    new_n14058_, new_n14059_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14066_, new_n14067_,
    new_n14068_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14206_, new_n14207_,
    new_n14208_, new_n14209_, new_n14210_, new_n14211_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14217_,
    new_n14218_, new_n14219_, new_n14220_, new_n14221_, new_n14222_,
    new_n14223_, new_n14224_, new_n14225_, new_n14226_, new_n14227_,
    new_n14228_, new_n14229_, new_n14230_, new_n14231_, new_n14232_,
    new_n14233_, new_n14234_, new_n14235_, new_n14236_, new_n14237_,
    new_n14238_, new_n14239_, new_n14240_, new_n14241_, new_n14242_,
    new_n14243_, new_n14244_, new_n14245_, new_n14246_, new_n14247_,
    new_n14248_, new_n14249_, new_n14250_, new_n14251_, new_n14252_,
    new_n14253_, new_n14254_, new_n14255_, new_n14256_, new_n14257_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14551_, new_n14552_,
    new_n14553_, new_n14554_, new_n14555_, new_n14556_, new_n14557_,
    new_n14558_, new_n14559_, new_n14560_, new_n14561_, new_n14562_,
    new_n14563_, new_n14564_, new_n14565_, new_n14566_, new_n14567_,
    new_n14568_, new_n14569_, new_n14570_, new_n14571_, new_n14572_,
    new_n14573_, new_n14574_, new_n14575_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14712_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14719_, new_n14720_, new_n14721_, new_n14722_,
    new_n14723_, new_n14724_, new_n14725_, new_n14726_, new_n14727_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14734_, new_n14735_, new_n14736_, new_n14737_,
    new_n14738_, new_n14739_, new_n14740_, new_n14741_, new_n14742_,
    new_n14743_, new_n14744_, new_n14745_, new_n14746_, new_n14747_,
    new_n14748_, new_n14749_, new_n14750_, new_n14751_, new_n14752_,
    new_n14753_, new_n14754_, new_n14755_, new_n14756_, new_n14757_,
    new_n14758_, new_n14759_, new_n14760_, new_n14761_, new_n14762_,
    new_n14763_, new_n14764_, new_n14765_, new_n14766_, new_n14767_,
    new_n14768_, new_n14769_, new_n14770_, new_n14771_, new_n14772_,
    new_n14773_, new_n14774_, new_n14775_, new_n14776_, new_n14777_,
    new_n14778_, new_n14779_, new_n14780_, new_n14781_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14818_, new_n14819_, new_n14820_, new_n14821_, new_n14822_,
    new_n14823_, new_n14824_, new_n14825_, new_n14826_, new_n14827_,
    new_n14828_, new_n14829_, new_n14830_, new_n14831_, new_n14832_,
    new_n14833_, new_n14834_, new_n14835_, new_n14836_, new_n14837_,
    new_n14838_, new_n14839_, new_n14840_, new_n14841_, new_n14842_,
    new_n14843_, new_n14844_, new_n14845_, new_n14846_, new_n14847_,
    new_n14848_, new_n14849_, new_n14850_, new_n14851_, new_n14852_,
    new_n14853_, new_n14854_, new_n14855_, new_n14856_, new_n14857_,
    new_n14858_, new_n14859_, new_n14860_, new_n14861_, new_n14862_,
    new_n14863_, new_n14864_, new_n14865_, new_n14866_, new_n14867_,
    new_n14868_, new_n14869_, new_n14870_, new_n14871_, new_n14872_,
    new_n14873_, new_n14874_, new_n14875_, new_n14876_, new_n14877_,
    new_n14878_, new_n14879_, new_n14880_, new_n14881_, new_n14882_,
    new_n14883_, new_n14884_, new_n14885_, new_n14886_, new_n14887_,
    new_n14888_, new_n14889_, new_n14890_, new_n14891_, new_n14892_,
    new_n14893_, new_n14894_, new_n14895_, new_n14896_, new_n14897_,
    new_n14898_, new_n14899_, new_n14900_, new_n14901_, new_n14902_,
    new_n14903_, new_n14904_, new_n14905_, new_n14906_, new_n14907_,
    new_n14908_, new_n14909_, new_n14910_, new_n14911_, new_n14912_,
    new_n14913_, new_n14914_, new_n14915_, new_n14916_, new_n14917_,
    new_n14918_, new_n14919_, new_n14920_, new_n14921_, new_n14922_,
    new_n14923_, new_n14924_, new_n14925_, new_n14926_, new_n14927_,
    new_n14928_, new_n14929_, new_n14930_, new_n14931_, new_n14932_,
    new_n14933_, new_n14934_, new_n14935_, new_n14936_, new_n14937_,
    new_n14938_, new_n14939_, new_n14940_, new_n14941_, new_n14942_,
    new_n14943_, new_n14944_, new_n14945_, new_n14946_, new_n14947_,
    new_n14948_, new_n14949_, new_n14950_, new_n14951_, new_n14952_,
    new_n14953_, new_n14954_, new_n14955_, new_n14956_, new_n14957_,
    new_n14958_, new_n14959_, new_n14960_, new_n14961_, new_n14962_,
    new_n14963_, new_n14964_, new_n14965_, new_n14966_, new_n14967_,
    new_n14968_, new_n14969_, new_n14970_, new_n14971_, new_n14972_,
    new_n14973_, new_n14974_, new_n14975_, new_n14976_, new_n14977_,
    new_n14978_, new_n14979_, new_n14980_, new_n14981_, new_n14982_,
    new_n14983_, new_n14984_, new_n14985_, new_n14986_, new_n14987_,
    new_n14988_, new_n14989_, new_n14990_, new_n14991_, new_n14992_,
    new_n14993_, new_n14994_, new_n14995_, new_n14996_, new_n14997_,
    new_n14998_, new_n14999_, new_n15000_, new_n15001_, new_n15002_,
    new_n15003_, new_n15004_, new_n15005_, new_n15006_, new_n15007_,
    new_n15008_, new_n15009_, new_n15010_, new_n15011_, new_n15012_,
    new_n15013_, new_n15014_, new_n15015_, new_n15016_, new_n15017_,
    new_n15018_, new_n15019_, new_n15020_, new_n15021_, new_n15022_,
    new_n15023_, new_n15024_, new_n15025_, new_n15026_, new_n15027_,
    new_n15028_, new_n15029_, new_n15030_, new_n15031_, new_n15032_,
    new_n15033_, new_n15034_, new_n15035_, new_n15036_, new_n15037_,
    new_n15038_, new_n15039_, new_n15040_, new_n15041_, new_n15042_,
    new_n15043_, new_n15044_, new_n15045_, new_n15046_, new_n15047_,
    new_n15048_, new_n15049_, new_n15050_, new_n15051_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15057_,
    new_n15058_, new_n15059_, new_n15060_, new_n15061_, new_n15062_,
    new_n15063_, new_n15064_, new_n15065_, new_n15066_, new_n15067_,
    new_n15068_, new_n15069_, new_n15070_, new_n15071_, new_n15072_,
    new_n15073_, new_n15074_, new_n15075_, new_n15076_, new_n15077_,
    new_n15078_, new_n15079_, new_n15080_, new_n15081_, new_n15082_,
    new_n15083_, new_n15084_, new_n15085_, new_n15086_, new_n15087_,
    new_n15088_, new_n15089_, new_n15090_, new_n15091_, new_n15092_,
    new_n15093_, new_n15094_, new_n15095_, new_n15096_, new_n15097_,
    new_n15098_, new_n15099_, new_n15100_, new_n15101_, new_n15102_,
    new_n15103_, new_n15104_, new_n15105_, new_n15106_, new_n15107_,
    new_n15108_, new_n15109_, new_n15110_, new_n15111_, new_n15112_,
    new_n15113_, new_n15114_, new_n15115_, new_n15116_, new_n15117_,
    new_n15118_, new_n15119_, new_n15120_, new_n15121_, new_n15122_,
    new_n15123_, new_n15124_, new_n15125_, new_n15126_, new_n15127_,
    new_n15128_, new_n15129_, new_n15130_, new_n15131_, new_n15132_,
    new_n15133_, new_n15134_, new_n15135_, new_n15136_, new_n15137_,
    new_n15138_, new_n15139_, new_n15140_, new_n15141_, new_n15142_,
    new_n15143_, new_n15144_, new_n15145_, new_n15146_, new_n15147_,
    new_n15148_, new_n15149_, new_n15150_, new_n15151_, new_n15152_,
    new_n15153_, new_n15154_, new_n15155_, new_n15156_, new_n15157_,
    new_n15158_, new_n15159_, new_n15160_, new_n15161_, new_n15162_,
    new_n15163_, new_n15164_, new_n15165_, new_n15166_, new_n15167_,
    new_n15168_, new_n15169_, new_n15170_, new_n15171_, new_n15172_,
    new_n15173_, new_n15174_, new_n15175_, new_n15176_, new_n15177_,
    new_n15178_, new_n15179_, new_n15180_, new_n15181_, new_n15182_,
    new_n15183_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15188_, new_n15189_, new_n15190_, new_n15191_, new_n15192_,
    new_n15193_, new_n15194_, new_n15195_, new_n15196_, new_n15197_,
    new_n15198_, new_n15199_, new_n15200_, new_n15201_, new_n15202_,
    new_n15203_, new_n15204_, new_n15205_, new_n15206_, new_n15207_,
    new_n15208_, new_n15209_, new_n15210_, new_n15211_, new_n15212_,
    new_n15213_, new_n15214_, new_n15215_, new_n15216_, new_n15217_,
    new_n15218_, new_n15219_, new_n15220_, new_n15221_, new_n15222_,
    new_n15223_, new_n15224_, new_n15225_, new_n15226_, new_n15227_,
    new_n15228_, new_n15229_, new_n15230_, new_n15231_, new_n15232_,
    new_n15233_, new_n15234_, new_n15235_, new_n15236_, new_n15237_,
    new_n15238_, new_n15239_, new_n15240_, new_n15241_, new_n15242_,
    new_n15243_, new_n15244_, new_n15245_, new_n15246_, new_n15247_,
    new_n15248_, new_n15249_, new_n15250_, new_n15251_, new_n15252_,
    new_n15253_, new_n15254_, new_n15255_, new_n15256_, new_n15257_,
    new_n15258_, new_n15259_, new_n15260_, new_n15261_, new_n15262_,
    new_n15263_, new_n15264_, new_n15265_, new_n15266_, new_n15267_,
    new_n15268_, new_n15269_, new_n15270_, new_n15271_, new_n15272_,
    new_n15273_, new_n15274_, new_n15275_, new_n15276_, new_n15277_,
    new_n15278_, new_n15279_, new_n15280_, new_n15281_, new_n15282_,
    new_n15283_, new_n15284_, new_n15285_, new_n15286_, new_n15287_,
    new_n15288_, new_n15289_, new_n15290_, new_n15291_, new_n15292_,
    new_n15293_, new_n15294_, new_n15295_, new_n15296_, new_n15297_,
    new_n15298_, new_n15299_, new_n15300_, new_n15301_, new_n15302_,
    new_n15303_, new_n15304_, new_n15305_, new_n15306_, new_n15307_,
    new_n15308_, new_n15309_, new_n15310_, new_n15311_, new_n15312_,
    new_n15313_, new_n15314_, new_n15315_, new_n15316_, new_n15317_,
    new_n15318_, new_n15319_, new_n15320_, new_n15321_, new_n15322_,
    new_n15323_, new_n15324_, new_n15325_, new_n15326_, new_n15327_,
    new_n15328_, new_n15329_, new_n15330_, new_n15331_, new_n15332_,
    new_n15333_, new_n15334_, new_n15335_, new_n15336_, new_n15337_,
    new_n15338_, new_n15339_, new_n15340_, new_n15341_, new_n15342_,
    new_n15343_, new_n15344_, new_n15345_, new_n15346_, new_n15347_,
    new_n15348_, new_n15349_, new_n15350_, new_n15351_, new_n15352_,
    new_n15353_, new_n15354_, new_n15355_, new_n15356_, new_n15357_,
    new_n15358_, new_n15359_, new_n15360_, new_n15361_, new_n15362_,
    new_n15363_, new_n15364_, new_n15365_, new_n15366_, new_n15367_,
    new_n15368_, new_n15369_, new_n15370_, new_n15371_, new_n15372_,
    new_n15373_, new_n15374_, new_n15375_, new_n15376_, new_n15377_,
    new_n15378_, new_n15379_, new_n15380_, new_n15381_, new_n15382_,
    new_n15383_, new_n15384_, new_n15385_, new_n15386_, new_n15387_,
    new_n15388_, new_n15389_, new_n15390_, new_n15391_, new_n15392_,
    new_n15393_, new_n15394_, new_n15395_, new_n15396_, new_n15397_,
    new_n15398_, new_n15399_, new_n15400_, new_n15401_, new_n15402_,
    new_n15403_, new_n15404_, new_n15405_, new_n15406_, new_n15407_,
    new_n15408_, new_n15409_, new_n15410_, new_n15411_, new_n15412_,
    new_n15413_, new_n15414_, new_n15415_, new_n15416_, new_n15417_,
    new_n15418_, new_n15419_, new_n15420_, new_n15421_, new_n15422_,
    new_n15423_, new_n15424_, new_n15425_, new_n15426_, new_n15427_,
    new_n15428_, new_n15429_, new_n15430_, new_n15431_, new_n15432_,
    new_n15433_, new_n15434_, new_n15435_, new_n15436_, new_n15437_,
    new_n15438_, new_n15439_, new_n15440_, new_n15441_, new_n15442_,
    new_n15443_, new_n15444_, new_n15445_, new_n15446_, new_n15447_,
    new_n15448_, new_n15449_, new_n15450_, new_n15451_, new_n15452_,
    new_n15453_, new_n15454_, new_n15455_, new_n15456_, new_n15457_,
    new_n15458_, new_n15459_, new_n15460_, new_n15461_, new_n15462_,
    new_n15463_, new_n15464_, new_n15465_, new_n15466_, new_n15467_,
    new_n15468_, new_n15469_, new_n15470_, new_n15471_, new_n15472_,
    new_n15473_, new_n15474_, new_n15475_, new_n15476_, new_n15477_,
    new_n15478_, new_n15479_, new_n15480_, new_n15481_, new_n15482_,
    new_n15483_, new_n15484_, new_n15485_, new_n15486_, new_n15487_,
    new_n15488_, new_n15489_, new_n15490_, new_n15491_, new_n15492_,
    new_n15493_, new_n15494_, new_n15495_, new_n15496_, new_n15497_,
    new_n15498_, new_n15499_, new_n15500_, new_n15501_, new_n15502_,
    new_n15503_, new_n15504_, new_n15505_, new_n15506_, new_n15507_,
    new_n15508_, new_n15509_, new_n15510_, new_n15511_, new_n15512_,
    new_n15513_, new_n15514_, new_n15515_, new_n15516_, new_n15517_,
    new_n15518_, new_n15519_, new_n15520_, new_n15521_, new_n15522_,
    new_n15523_, new_n15524_, new_n15525_, new_n15526_, new_n15527_,
    new_n15528_, new_n15529_, new_n15530_, new_n15531_, new_n15532_,
    new_n15533_, new_n15534_, new_n15535_, new_n15536_, new_n15537_,
    new_n15538_, new_n15539_, new_n15540_, new_n15541_, new_n15542_,
    new_n15543_, new_n15544_, new_n15545_, new_n15546_, new_n15547_,
    new_n15548_, new_n15549_, new_n15550_, new_n15551_, new_n15552_,
    new_n15553_, new_n15554_, new_n15555_, new_n15556_, new_n15557_,
    new_n15558_, new_n15559_, new_n15560_, new_n15561_, new_n15562_,
    new_n15563_, new_n15564_, new_n15565_, new_n15566_, new_n15567_,
    new_n15568_, new_n15569_, new_n15570_, new_n15571_, new_n15572_,
    new_n15573_, new_n15574_, new_n15575_, new_n15576_, new_n15577_,
    new_n15578_, new_n15579_, new_n15580_, new_n15581_, new_n15582_,
    new_n15583_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15590_, new_n15591_, new_n15592_,
    new_n15593_, new_n15594_, new_n15595_, new_n15596_, new_n15597_,
    new_n15598_, new_n15599_, new_n15600_, new_n15601_, new_n15602_,
    new_n15603_, new_n15604_, new_n15605_, new_n15606_, new_n15607_,
    new_n15608_, new_n15609_, new_n15610_, new_n15611_, new_n15612_,
    new_n15613_, new_n15614_, new_n15615_, new_n15616_, new_n15617_,
    new_n15618_, new_n15619_, new_n15620_, new_n15621_, new_n15622_,
    new_n15623_, new_n15624_, new_n15625_, new_n15626_, new_n15627_,
    new_n15628_, new_n15629_, new_n15630_, new_n15631_, new_n15632_,
    new_n15633_, new_n15634_, new_n15635_, new_n15636_, new_n15637_,
    new_n15638_, new_n15639_, new_n15640_, new_n15641_, new_n15642_,
    new_n15643_, new_n15644_, new_n15645_, new_n15646_, new_n15647_,
    new_n15648_, new_n15649_, new_n15650_, new_n15651_, new_n15652_,
    new_n15653_, new_n15654_, new_n15655_, new_n15656_, new_n15657_,
    new_n15658_, new_n15659_, new_n15660_, new_n15661_, new_n15662_,
    new_n15663_, new_n15664_, new_n15665_, new_n15666_, new_n15667_,
    new_n15668_, new_n15669_, new_n15670_, new_n15671_, new_n15672_,
    new_n15673_, new_n15674_, new_n15675_, new_n15676_, new_n15677_,
    new_n15678_, new_n15679_, new_n15680_, new_n15681_, new_n15682_,
    new_n15683_, new_n15684_, new_n15685_, new_n15686_, new_n15687_,
    new_n15688_, new_n15689_, new_n15690_, new_n15691_, new_n15692_,
    new_n15693_, new_n15694_, new_n15695_, new_n15696_, new_n15697_,
    new_n15698_, new_n15699_, new_n15700_, new_n15701_, new_n15702_,
    new_n15703_, new_n15704_, new_n15705_, new_n15706_, new_n15707_,
    new_n15708_, new_n15709_, new_n15710_, new_n15711_, new_n15712_,
    new_n15713_, new_n15714_, new_n15715_, new_n15716_, new_n15717_,
    new_n15718_, new_n15719_, new_n15720_, new_n15721_, new_n15722_,
    new_n15723_, new_n15724_, new_n15725_, new_n15726_, new_n15727_,
    new_n15728_, new_n15729_, new_n15730_, new_n15731_, new_n15732_,
    new_n15733_, new_n15734_, new_n15735_, new_n15736_, new_n15737_,
    new_n15738_, new_n15739_, new_n15740_, new_n15741_, new_n15742_,
    new_n15743_, new_n15744_, new_n15745_, new_n15746_, new_n15747_,
    new_n15748_, new_n15749_, new_n15750_, new_n15751_, new_n15752_,
    new_n15753_, new_n15754_, new_n15755_, new_n15756_, new_n15757_,
    new_n15758_, new_n15759_, new_n15760_, new_n15761_, new_n15762_,
    new_n15763_, new_n15764_, new_n15765_, new_n15766_, new_n15767_,
    new_n15768_, new_n15769_, new_n15770_, new_n15771_, new_n15772_,
    new_n15773_, new_n15774_, new_n15775_, new_n15776_, new_n15777_,
    new_n15778_, new_n15779_, new_n15780_, new_n15781_, new_n15782_,
    new_n15783_, new_n15784_, new_n15785_, new_n15786_, new_n15787_,
    new_n15788_, new_n15789_, new_n15790_, new_n15791_, new_n15792_,
    new_n15793_, new_n15794_, new_n15795_, new_n15796_, new_n15797_,
    new_n15798_, new_n15799_, new_n15800_, new_n15801_, new_n15802_,
    new_n15803_, new_n15804_, new_n15805_, new_n15806_, new_n15807_,
    new_n15808_, new_n15809_, new_n15810_, new_n15811_, new_n15812_,
    new_n15813_, new_n15814_, new_n15815_, new_n15816_, new_n15817_,
    new_n15818_, new_n15819_, new_n15820_, new_n15821_, new_n15822_,
    new_n15823_, new_n15824_, new_n15825_, new_n15826_, new_n15827_,
    new_n15828_, new_n15829_, new_n15830_, new_n15831_, new_n15832_,
    new_n15833_, new_n15834_, new_n15835_, new_n15836_, new_n15837_,
    new_n15838_, new_n15839_, new_n15840_, new_n15841_, new_n15842_,
    new_n15843_, new_n15844_, new_n15845_, new_n15846_, new_n15847_,
    new_n15848_, new_n15849_, new_n15850_, new_n15851_, new_n15852_,
    new_n15853_, new_n15854_, new_n15855_, new_n15856_, new_n15857_,
    new_n15858_, new_n15859_, new_n15860_, new_n15861_, new_n15862_,
    new_n15863_, new_n15864_, new_n15865_, new_n15866_, new_n15867_,
    new_n15868_, new_n15869_, new_n15870_, new_n15871_, new_n15872_,
    new_n15873_, new_n15874_, new_n15875_, new_n15876_, new_n15877_,
    new_n15878_, new_n15879_, new_n15880_, new_n15881_, new_n15882_,
    new_n15883_, new_n15884_, new_n15885_, new_n15886_, new_n15887_,
    new_n15888_, new_n15889_, new_n15890_, new_n15891_, new_n15892_,
    new_n15893_, new_n15894_, new_n15895_, new_n15896_, new_n15897_,
    new_n15898_, new_n15899_, new_n15900_, new_n15901_, new_n15902_,
    new_n15903_, new_n15904_, new_n15905_, new_n15906_, new_n15907_,
    new_n15908_, new_n15909_, new_n15910_, new_n15911_, new_n15912_,
    new_n15913_, new_n15914_, new_n15915_, new_n15916_, new_n15917_,
    new_n15918_, new_n15919_, new_n15920_, new_n15921_, new_n15922_,
    new_n15923_, new_n15924_, new_n15925_, new_n15926_, new_n15927_,
    new_n15928_, new_n15929_, new_n15930_, new_n15931_, new_n15932_,
    new_n15933_, new_n15934_, new_n15935_, new_n15936_, new_n15937_,
    new_n15938_, new_n15939_, new_n15940_, new_n15941_, new_n15942_,
    new_n15943_, new_n15944_, new_n15945_, new_n15946_, new_n15947_,
    new_n15948_, new_n15949_, new_n15950_, new_n15951_, new_n15952_,
    new_n15953_, new_n15954_, new_n15955_, new_n15956_, new_n15957_,
    new_n15958_, new_n15959_, new_n15960_, new_n15961_, new_n15962_,
    new_n15963_, new_n15964_, new_n15965_, new_n15966_, new_n15967_,
    new_n15968_, new_n15969_, new_n15970_, new_n15971_, new_n15972_,
    new_n15973_, new_n15974_, new_n15975_, new_n15976_, new_n15977_,
    new_n15978_, new_n15979_, new_n15980_, new_n15981_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16424_, new_n16425_, new_n16426_, new_n16427_, new_n16428_,
    new_n16429_, new_n16430_, new_n16431_, new_n16432_, new_n16433_,
    new_n16434_, new_n16435_, new_n16436_, new_n16437_, new_n16438_,
    new_n16439_, new_n16440_, new_n16441_, new_n16442_, new_n16443_,
    new_n16444_, new_n16445_, new_n16446_, new_n16447_, new_n16448_,
    new_n16449_, new_n16450_, new_n16451_, new_n16452_, new_n16453_,
    new_n16454_, new_n16455_, new_n16456_, new_n16457_, new_n16458_,
    new_n16459_, new_n16460_, new_n16461_, new_n16462_, new_n16463_,
    new_n16464_, new_n16465_, new_n16466_, new_n16467_, new_n16468_,
    new_n16469_, new_n16470_, new_n16471_, new_n16472_, new_n16473_,
    new_n16474_, new_n16475_, new_n16476_, new_n16477_, new_n16478_,
    new_n16479_, new_n16480_, new_n16481_, new_n16482_, new_n16483_,
    new_n16484_, new_n16485_, new_n16486_, new_n16487_, new_n16488_,
    new_n16489_, new_n16490_, new_n16491_, new_n16492_, new_n16493_,
    new_n16494_, new_n16495_, new_n16496_, new_n16497_, new_n16498_,
    new_n16499_, new_n16500_, new_n16501_, new_n16502_, new_n16503_,
    new_n16504_, new_n16505_, new_n16506_, new_n16507_, new_n16508_,
    new_n16509_, new_n16510_, new_n16511_, new_n16512_, new_n16513_,
    new_n16514_, new_n16515_, new_n16516_, new_n16517_, new_n16518_,
    new_n16519_, new_n16520_, new_n16521_, new_n16522_, new_n16523_,
    new_n16524_, new_n16525_, new_n16526_, new_n16527_, new_n16528_,
    new_n16529_, new_n16530_, new_n16531_, new_n16532_, new_n16533_,
    new_n16534_, new_n16535_, new_n16536_, new_n16537_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16571_, new_n16572_, new_n16573_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16584_, new_n16585_, new_n16586_, new_n16587_, new_n16588_,
    new_n16589_, new_n16590_, new_n16591_, new_n16592_, new_n16593_,
    new_n16594_, new_n16595_, new_n16596_, new_n16597_, new_n16598_,
    new_n16599_, new_n16600_, new_n16601_, new_n16602_, new_n16603_,
    new_n16604_, new_n16605_, new_n16606_, new_n16607_, new_n16608_,
    new_n16609_, new_n16610_, new_n16611_, new_n16612_, new_n16613_,
    new_n16614_, new_n16615_, new_n16616_, new_n16617_, new_n16618_,
    new_n16619_, new_n16620_, new_n16621_, new_n16622_, new_n16623_,
    new_n16624_, new_n16625_, new_n16626_, new_n16627_, new_n16628_,
    new_n16629_, new_n16630_, new_n16631_, new_n16632_, new_n16633_,
    new_n16634_, new_n16635_, new_n16636_, new_n16637_, new_n16638_,
    new_n16643_, new_n16644_, new_n16648_, new_n16651_, new_n16652_,
    new_n16660_, new_n16661_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16933_, new_n16934_, new_n16935_, new_n16936_,
    new_n16937_, new_n16938_, new_n16939_, new_n16940_, new_n16941_,
    new_n16942_, new_n16943_, new_n16944_, new_n16945_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16952_, new_n16953_, new_n16954_, new_n16955_, new_n16956_,
    new_n16957_, new_n16958_, new_n16959_, new_n16960_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16980_, new_n16981_,
    new_n16982_, new_n16983_, new_n16984_, new_n16985_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16992_, new_n16993_, new_n16994_, new_n16995_, new_n16996_,
    new_n16997_, new_n16998_, new_n16999_, new_n17000_, new_n17001_,
    new_n17002_, new_n17003_, new_n17004_, new_n17005_, new_n17006_,
    new_n17007_, new_n17008_, new_n17009_, new_n17010_, new_n17011_,
    new_n17012_, new_n17013_, new_n17014_, new_n17015_, new_n17016_,
    new_n17017_, new_n17018_, new_n17019_, new_n17020_, new_n17021_,
    new_n17022_, new_n17023_, new_n17024_, new_n17025_, new_n17026_,
    new_n17027_, new_n17028_, new_n17029_, new_n17030_, new_n17031_,
    new_n17032_, new_n17033_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17106_,
    new_n17107_, new_n17108_, new_n17109_, new_n17110_, new_n17111_,
    new_n17112_, new_n17113_, new_n17114_, new_n17115_, new_n17116_,
    new_n17117_, new_n17118_, new_n17119_, new_n17120_, new_n17121_,
    new_n17122_, new_n17123_, new_n17124_, new_n17125_, new_n17126_,
    new_n17127_, new_n17128_, new_n17129_, new_n17130_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17225_, new_n17226_,
    new_n17227_, new_n17228_, new_n17229_, new_n17230_, new_n17231_,
    new_n17232_, new_n17233_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17251_,
    new_n17252_, new_n17253_, new_n17254_, new_n17255_, new_n17256_,
    new_n17257_, new_n17258_, new_n17259_, new_n17260_, new_n17261_,
    new_n17262_, new_n17263_, new_n17264_, new_n17265_, new_n17266_,
    new_n17267_, new_n17268_, new_n17269_, new_n17270_, new_n17271_,
    new_n17272_, new_n17273_, new_n17274_, new_n17275_, new_n17276_,
    new_n17277_, new_n17278_, new_n17279_, new_n17280_, new_n17281_,
    new_n17282_, new_n17283_, new_n17284_, new_n17285_, new_n17286_,
    new_n17287_, new_n17288_, new_n17289_, new_n17290_, new_n17291_,
    new_n17292_, new_n17293_, new_n17294_, new_n17295_, new_n17296_,
    new_n17297_, new_n17298_, new_n17299_, new_n17300_, new_n17301_,
    new_n17302_, new_n17303_, new_n17304_, new_n17305_, new_n17306_,
    new_n17307_, new_n17308_, new_n17309_, new_n17310_, new_n17311_,
    new_n17312_, new_n17313_, new_n17314_, new_n17315_, new_n17316_,
    new_n17317_, new_n17318_, new_n17319_, new_n17320_, new_n17321_,
    new_n17322_, new_n17323_, new_n17324_, new_n17325_, new_n17326_,
    new_n17327_, new_n17328_, new_n17329_, new_n17330_, new_n17331_,
    new_n17332_, new_n17333_, new_n17334_, new_n17335_, new_n17336_,
    new_n17337_, new_n17338_, new_n17339_, new_n17340_, new_n17341_,
    new_n17342_, new_n17343_, new_n17344_, new_n17345_, new_n17346_,
    new_n17347_, new_n17348_, new_n17349_, new_n17350_, new_n17351_,
    new_n17352_, new_n17353_, new_n17354_, new_n17355_, new_n17356_,
    new_n17357_, new_n17358_, new_n17359_, new_n17360_, new_n17361_,
    new_n17362_, new_n17363_, new_n17364_, new_n17365_, new_n17366_,
    new_n17367_, new_n17368_, new_n17369_, new_n17370_, new_n17371_,
    new_n17372_, new_n17373_, new_n17374_, new_n17375_, new_n17376_,
    new_n17377_, new_n17378_, new_n17379_, new_n17380_, new_n17381_,
    new_n17382_, new_n17383_, new_n17384_, new_n17385_, new_n17386_,
    new_n17387_, new_n17388_, new_n17389_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17396_,
    new_n17397_, new_n17398_, new_n17399_, new_n17400_, new_n17401_,
    new_n17402_, new_n17403_, new_n17404_, new_n17405_, new_n17406_,
    new_n17407_, new_n17408_, new_n17409_, new_n17410_, new_n17411_,
    new_n17412_, new_n17413_, new_n17414_, new_n17415_, new_n17416_,
    new_n17417_, new_n17418_, new_n17419_, new_n17420_, new_n17421_,
    new_n17422_, new_n17423_, new_n17424_, new_n17425_, new_n17426_,
    new_n17427_, new_n17428_, new_n17429_, new_n17430_, new_n17431_,
    new_n17432_, new_n17433_, new_n17434_, new_n17435_, new_n17436_,
    new_n17437_, new_n17438_, new_n17439_, new_n17440_, new_n17441_,
    new_n17442_, new_n17443_, new_n17444_, new_n17445_, new_n17446_,
    new_n17447_, new_n17448_, new_n17449_, new_n17450_, new_n17451_,
    new_n17452_, new_n17453_, new_n17454_, new_n17455_, new_n17456_,
    new_n17457_, new_n17458_, new_n17459_, new_n17460_, new_n17461_,
    new_n17462_, new_n17463_, new_n17464_, new_n17465_, new_n17466_,
    new_n17467_, new_n17468_, new_n17469_, new_n17470_, new_n17471_,
    new_n17472_, new_n17473_, new_n17474_, new_n17475_, new_n17476_,
    new_n17477_, new_n17478_, new_n17479_, new_n17480_, new_n17481_,
    new_n17482_, new_n17483_, new_n17484_, new_n17485_, new_n17486_,
    new_n17487_, new_n17488_, new_n17489_, new_n17490_, new_n17491_,
    new_n17492_, new_n17493_, new_n17494_, new_n17495_, new_n17496_,
    new_n17497_, new_n17498_, new_n17499_, new_n17500_, new_n17501_,
    new_n17502_, new_n17503_, new_n17504_, new_n17505_, new_n17506_,
    new_n17507_, new_n17508_, new_n17509_, new_n17510_, new_n17511_,
    new_n17512_, new_n17513_, new_n17514_, new_n17515_, new_n17516_,
    new_n17517_, new_n17518_, new_n17519_, new_n17520_, new_n17521_,
    new_n17522_, new_n17523_, new_n17524_, new_n17525_, new_n17526_,
    new_n17527_, new_n17528_, new_n17529_, new_n17530_, new_n17531_,
    new_n17532_, new_n17533_, new_n17534_, new_n17535_, new_n17536_,
    new_n17537_, new_n17538_, new_n17539_, new_n17540_, new_n17541_,
    new_n17542_, new_n17543_, new_n17544_, new_n17545_, new_n17546_,
    new_n17547_, new_n17548_, new_n17549_, new_n17550_, new_n17551_,
    new_n17552_, new_n17553_, new_n17554_, new_n17555_, new_n17556_,
    new_n17557_, new_n17558_, new_n17559_, new_n17560_, new_n17561_,
    new_n17562_, new_n17563_, new_n17564_, new_n17565_, new_n17566_,
    new_n17567_, new_n17568_, new_n17569_, new_n17570_, new_n17571_,
    new_n17572_, new_n17573_, new_n17574_, new_n17575_, new_n17576_,
    new_n17577_, new_n17578_, new_n17579_, new_n17580_, new_n17581_,
    new_n17582_, new_n17583_, new_n17584_, new_n17585_, new_n17586_,
    new_n17587_, new_n17588_, new_n17589_, new_n17590_, new_n17591_,
    new_n17592_, new_n17593_, new_n17594_, new_n17595_, new_n17596_,
    new_n17597_, new_n17598_, new_n17599_, new_n17600_, new_n17601_,
    new_n17602_, new_n17603_, new_n17604_, new_n17605_, new_n17606_,
    new_n17607_, new_n17608_, new_n17609_, new_n17610_, new_n17611_,
    new_n17612_, new_n17613_, new_n17614_, new_n17615_, new_n17616_,
    new_n17617_, new_n17618_, new_n17619_, new_n17620_, new_n17621_,
    new_n17622_, new_n17623_, new_n17624_, new_n17625_, new_n17626_,
    new_n17627_, new_n17628_, new_n17629_, new_n17630_, new_n17631_,
    new_n17632_, new_n17633_, new_n17634_, new_n17635_, new_n17636_,
    new_n17637_, new_n17638_, new_n17639_, new_n17640_, new_n17641_,
    new_n17642_, new_n17643_, new_n17644_, new_n17645_, new_n17646_,
    new_n17647_, new_n17648_, new_n17649_, new_n17650_, new_n17651_,
    new_n17652_, new_n17653_, new_n17654_, new_n17655_, new_n17656_,
    new_n17657_, new_n17658_, new_n17659_, new_n17660_, new_n17661_,
    new_n17662_, new_n17663_, new_n17664_, new_n17665_, new_n17666_,
    new_n17667_, new_n17668_, new_n17669_, new_n17670_, new_n17671_,
    new_n17672_, new_n17673_, new_n17674_, new_n17675_, new_n17676_,
    new_n17677_, new_n17678_, new_n17679_, new_n17680_, new_n17681_,
    new_n17682_, new_n17683_, new_n17684_, new_n17685_, new_n17686_,
    new_n17687_, new_n17688_, new_n17689_, new_n17690_, new_n17691_,
    new_n17692_, new_n17693_, new_n17694_, new_n17695_, new_n17696_,
    new_n17697_, new_n17698_, new_n17699_, new_n17700_, new_n17701_,
    new_n17702_, new_n17703_, new_n17704_, new_n17705_, new_n17706_,
    new_n17707_, new_n17708_, new_n17709_, new_n17710_, new_n17711_,
    new_n17712_, new_n17713_, new_n17714_, new_n17715_, new_n17716_,
    new_n17717_, new_n17718_, new_n17719_, new_n17720_, new_n17721_,
    new_n17722_, new_n17723_, new_n17724_, new_n17725_, new_n17726_,
    new_n17727_, new_n17728_, new_n17729_, new_n17730_, new_n17731_,
    new_n17732_, new_n17733_, new_n17734_, new_n17735_, new_n17736_,
    new_n17737_, new_n17738_, new_n17739_, new_n17740_, new_n17741_,
    new_n17742_, new_n17743_, new_n17744_, new_n17745_, new_n17746_,
    new_n17747_, new_n17748_, new_n17749_, new_n17750_, new_n17751_,
    new_n17752_, new_n17753_, new_n17754_, new_n17755_, new_n17756_,
    new_n17757_, new_n17758_, new_n17759_, new_n17760_, new_n17761_,
    new_n17762_, new_n17763_, new_n17764_, new_n17765_, new_n17766_,
    new_n17767_, new_n17768_, new_n17769_, new_n17770_, new_n17771_,
    new_n17772_, new_n17773_, new_n17774_, new_n17775_, new_n17776_,
    new_n17777_, new_n17778_, new_n17779_, new_n17780_, new_n17781_,
    new_n17782_, new_n17783_, new_n17784_, new_n17785_, new_n17786_,
    new_n17787_, new_n17788_, new_n17789_, new_n17790_, new_n17791_,
    new_n17792_, new_n17793_, new_n17794_, new_n17795_, new_n17796_,
    new_n17797_, new_n17798_, new_n17799_, new_n17800_, new_n17801_,
    new_n17802_, new_n17803_, new_n17804_, new_n17805_, new_n17806_,
    new_n17807_, new_n17808_, new_n17809_, new_n17810_, new_n17811_,
    new_n17812_, new_n17813_, new_n17814_, new_n17815_, new_n17816_,
    new_n17817_, new_n17818_, new_n17819_, new_n17820_, new_n17821_,
    new_n17822_, new_n17823_, new_n17824_, new_n17825_, new_n17826_,
    new_n17827_, new_n17828_, new_n17829_, new_n17830_, new_n17831_,
    new_n17832_, new_n17833_, new_n17834_, new_n17835_, new_n17836_,
    new_n17837_, new_n17838_, new_n17839_, new_n17840_, new_n17841_,
    new_n17842_, new_n17843_, new_n17844_, new_n17845_, new_n17846_,
    new_n17847_, new_n17848_, new_n17849_, new_n17850_, new_n17851_,
    new_n17852_, new_n17853_, new_n17854_, new_n17855_, new_n17856_,
    new_n17857_, new_n17858_, new_n17859_, new_n17860_, new_n17861_,
    new_n17862_, new_n17863_, new_n17864_, new_n17865_, new_n17866_,
    new_n17867_, new_n17868_, new_n17869_, new_n17870_, new_n17871_,
    new_n17872_, new_n17873_, new_n17874_, new_n17875_, new_n17876_,
    new_n17877_, new_n17878_, new_n17879_, new_n17880_, new_n17881_,
    new_n17882_, new_n17883_, new_n17884_, new_n17885_, new_n17886_,
    new_n17887_, new_n17888_, new_n17889_, new_n17890_, new_n17891_,
    new_n17892_, new_n17893_, new_n17894_, new_n17895_, new_n17896_,
    new_n17897_, new_n17898_, new_n17899_, new_n17900_, new_n17901_,
    new_n17902_, new_n17903_, new_n17904_, new_n17905_, new_n17906_,
    new_n17907_, new_n17908_, new_n17909_, new_n17910_, new_n17911_,
    new_n17912_, new_n17913_, new_n17914_, new_n17915_, new_n17916_,
    new_n17917_, new_n17918_, new_n17919_, new_n17920_, new_n17921_,
    new_n17922_, new_n17923_, new_n17924_, new_n17925_, new_n17926_,
    new_n17927_, new_n17928_, new_n17929_, new_n17930_, new_n17931_,
    new_n17932_, new_n17933_, new_n17934_, new_n17935_, new_n17936_,
    new_n17937_, new_n17938_, new_n17939_, new_n17940_, new_n17941_,
    new_n17942_, new_n17943_, new_n17944_, new_n17945_, new_n17946_,
    new_n17947_, new_n17948_, new_n17949_, new_n17950_, new_n17951_,
    new_n17952_, new_n17953_, new_n17954_, new_n17955_, new_n17956_,
    new_n17957_, new_n17958_, new_n17959_, new_n17960_, new_n17961_,
    new_n17962_, new_n17963_, new_n17964_, new_n17965_, new_n17966_,
    new_n17967_, new_n17968_, new_n17969_, new_n17970_, new_n17971_,
    new_n17972_, new_n17973_, new_n17974_, new_n17975_, new_n17976_,
    new_n17977_, new_n17978_, new_n17979_, new_n17980_, new_n17981_,
    new_n17982_, new_n17983_, new_n17984_, new_n17985_, new_n17986_,
    new_n17987_, new_n17988_, new_n17989_, new_n17990_, new_n17991_,
    new_n17992_, new_n17993_, new_n17994_, new_n17995_, new_n17996_,
    new_n17997_, new_n17998_, new_n17999_, new_n18000_, new_n18001_,
    new_n18002_, new_n18003_, new_n18004_, new_n18005_, new_n18006_,
    new_n18007_, new_n18008_, new_n18009_, new_n18010_, new_n18011_,
    new_n18012_, new_n18013_, new_n18014_, new_n18015_, new_n18016_,
    new_n18017_, new_n18018_, new_n18019_, new_n18020_, new_n18021_,
    new_n18022_, new_n18023_, new_n18024_, new_n18025_, new_n18026_,
    new_n18027_, new_n18028_, new_n18029_, new_n18030_, new_n18031_,
    new_n18032_, new_n18033_, new_n18034_, new_n18035_, new_n18036_,
    new_n18037_, new_n18038_, new_n18039_, new_n18040_, new_n18041_,
    new_n18042_, new_n18043_, new_n18044_, new_n18045_, new_n18046_,
    new_n18047_, new_n18048_, new_n18049_, new_n18050_, new_n18051_,
    new_n18052_, new_n18053_, new_n18054_, new_n18055_, new_n18056_,
    new_n18057_, new_n18058_, new_n18059_, new_n18060_, new_n18061_,
    new_n18062_, new_n18063_, new_n18064_, new_n18065_, new_n18066_,
    new_n18067_, new_n18068_, new_n18069_, new_n18070_, new_n18071_,
    new_n18072_, new_n18073_, new_n18074_, new_n18075_, new_n18076_,
    new_n18077_, new_n18078_, new_n18079_, new_n18080_, new_n18081_,
    new_n18082_, new_n18083_, new_n18084_, new_n18085_, new_n18086_,
    new_n18087_, new_n18088_, new_n18089_, new_n18090_, new_n18091_,
    new_n18092_, new_n18093_, new_n18094_, new_n18095_, new_n18096_,
    new_n18097_, new_n18098_, new_n18099_, new_n18100_, new_n18101_,
    new_n18102_, new_n18103_, new_n18104_, new_n18105_, new_n18106_,
    new_n18107_, new_n18108_, new_n18109_, new_n18110_, new_n18111_,
    new_n18112_, new_n18113_, new_n18114_, new_n18115_, new_n18116_,
    new_n18117_, new_n18118_, new_n18119_, new_n18120_, new_n18121_,
    new_n18122_, new_n18123_, new_n18124_, new_n18125_, new_n18126_,
    new_n18127_, new_n18128_, new_n18129_, new_n18130_, new_n18131_,
    new_n18132_, new_n18133_, new_n18134_, new_n18135_, new_n18136_,
    new_n18137_, new_n18138_, new_n18139_, new_n18140_, new_n18141_,
    new_n18142_, new_n18143_, new_n18144_, new_n18145_, new_n18146_,
    new_n18147_, new_n18148_, new_n18149_, new_n18150_, new_n18151_,
    new_n18152_, new_n18153_, new_n18154_, new_n18155_, new_n18156_,
    new_n18157_, new_n18158_, new_n18159_, new_n18160_, new_n18161_,
    new_n18162_, new_n18163_, new_n18164_, new_n18165_, new_n18166_,
    new_n18167_, new_n18168_, new_n18169_, new_n18170_, new_n18171_,
    new_n18172_, new_n18173_, new_n18174_, new_n18175_, new_n18176_,
    new_n18177_, new_n18178_, new_n18179_, new_n18180_, new_n18181_,
    new_n18182_, new_n18183_, new_n18184_, new_n18185_, new_n18186_,
    new_n18187_, new_n18188_, new_n18189_, new_n18190_, new_n18191_,
    new_n18192_, new_n18193_, new_n18194_, new_n18195_, new_n18196_,
    new_n18197_, new_n18198_, new_n18199_, new_n18200_, new_n18201_,
    new_n18202_, new_n18203_, new_n18204_, new_n18205_, new_n18206_,
    new_n18207_, new_n18208_, new_n18209_, new_n18210_, new_n18211_,
    new_n18212_, new_n18213_, new_n18214_, new_n18215_, new_n18216_,
    new_n18217_, new_n18218_, new_n18219_, new_n18220_, new_n18221_,
    new_n18222_, new_n18223_, new_n18224_, new_n18225_, new_n18226_,
    new_n18227_, new_n18228_, new_n18229_, new_n18230_, new_n18231_,
    new_n18232_, new_n18233_, new_n18234_, new_n18235_, new_n18236_,
    new_n18237_, new_n18238_, new_n18239_, new_n18240_, new_n18241_,
    new_n18242_, new_n18243_, new_n18244_, new_n18245_, new_n18246_,
    new_n18247_, new_n18248_, new_n18249_, new_n18250_, new_n18251_,
    new_n18252_, new_n18253_, new_n18254_, new_n18255_, new_n18256_,
    new_n18257_, new_n18258_, new_n18259_, new_n18260_, new_n18261_,
    new_n18262_, new_n18263_, new_n18264_, new_n18265_, new_n18266_,
    new_n18267_, new_n18268_, new_n18269_, new_n18270_, new_n18271_,
    new_n18272_, new_n18273_, new_n18274_, new_n18275_, new_n18276_,
    new_n18277_, new_n18278_, new_n18279_, new_n18280_, new_n18281_,
    new_n18282_, new_n18283_, new_n18284_, new_n18285_, new_n18286_,
    new_n18287_, new_n18288_, new_n18289_, new_n18290_, new_n18291_,
    new_n18292_, new_n18293_, new_n18294_, new_n18295_, new_n18296_,
    new_n18297_, new_n18298_, new_n18299_, new_n18300_, new_n18301_,
    new_n18302_, new_n18303_, new_n18304_, new_n18305_, new_n18306_,
    new_n18307_, new_n18308_, new_n18309_, new_n18310_, new_n18311_,
    new_n18312_, new_n18313_, new_n18314_, new_n18315_, new_n18316_,
    new_n18317_, new_n18318_, new_n18319_, new_n18320_, new_n18321_,
    new_n18322_, new_n18323_, new_n18324_, new_n18325_, new_n18326_,
    new_n18327_, new_n18328_, new_n18329_, new_n18330_, new_n18331_,
    new_n18332_, new_n18333_, new_n18334_, new_n18335_, new_n18336_,
    new_n18337_, new_n18338_, new_n18339_, new_n18340_, new_n18341_,
    new_n18342_, new_n18343_, new_n18344_, new_n18345_, new_n18346_,
    new_n18347_, new_n18348_, new_n18349_, new_n18350_, new_n18351_,
    new_n18352_, new_n18353_, new_n18354_, new_n18355_, new_n18356_,
    new_n18357_, new_n18358_, new_n18359_, new_n18360_, new_n18361_,
    new_n18362_, new_n18363_, new_n18364_, new_n18365_, new_n18366_,
    new_n18367_, new_n18368_, new_n18369_, new_n18370_, new_n18371_,
    new_n18372_, new_n18373_, new_n18374_, new_n18375_, new_n18376_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18393_, new_n18394_, new_n18395_, new_n18396_,
    new_n18397_, new_n18398_, new_n18399_, new_n18400_, new_n18401_,
    new_n18402_, new_n18403_, new_n18404_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18409_, new_n18410_, new_n18411_,
    new_n18412_, new_n18413_, new_n18414_, new_n18415_, new_n18416_,
    new_n18417_, new_n18418_, new_n18419_, new_n18420_, new_n18421_,
    new_n18422_, new_n18423_, new_n18424_, new_n18425_, new_n18426_,
    new_n18427_, new_n18428_, new_n18429_, new_n18430_, new_n18431_,
    new_n18432_, new_n18433_, new_n18434_, new_n18435_, new_n18436_,
    new_n18437_, new_n18438_, new_n18439_, new_n18440_, new_n18441_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18511_,
    new_n18512_, new_n18513_, new_n18514_, new_n18515_, new_n18516_,
    new_n18517_, new_n18518_, new_n18519_, new_n18520_, new_n18521_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18528_, new_n18529_, new_n18530_, new_n18531_,
    new_n18532_, new_n18533_, new_n18534_, new_n18535_, new_n18536_,
    new_n18537_, new_n18538_, new_n18539_, new_n18540_, new_n18541_,
    new_n18542_, new_n18543_, new_n18544_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18549_, new_n18550_, new_n18551_,
    new_n18552_, new_n18553_, new_n18554_, new_n18555_, new_n18556_,
    new_n18557_, new_n18558_, new_n18559_, new_n18560_, new_n18561_,
    new_n18562_, new_n18563_, new_n18564_, new_n18565_, new_n18566_,
    new_n18567_, new_n18568_, new_n18569_, new_n18570_, new_n18571_,
    new_n18572_, new_n18573_, new_n18574_, new_n18575_, new_n18576_,
    new_n18577_, new_n18578_, new_n18579_, new_n18580_, new_n18581_,
    new_n18582_, new_n18583_, new_n18584_, new_n18585_, new_n18586_,
    new_n18587_, new_n18588_, new_n18589_, new_n18590_, new_n18591_,
    new_n18592_, new_n18593_, new_n18594_, new_n18595_, new_n18596_,
    new_n18597_, new_n18598_, new_n18599_, new_n18600_, new_n18601_,
    new_n18602_, new_n18603_, new_n18604_, new_n18605_, new_n18606_,
    new_n18607_, new_n18608_, new_n18609_, new_n18610_, new_n18611_,
    new_n18612_, new_n18613_, new_n18614_, new_n18615_, new_n18616_,
    new_n18617_, new_n18618_, new_n18619_, new_n18620_, new_n18621_,
    new_n18622_, new_n18623_, new_n18624_, new_n18625_, new_n18626_,
    new_n18627_, new_n18628_, new_n18629_, new_n18630_, new_n18631_,
    new_n18632_, new_n18633_, new_n18634_, new_n18635_, new_n18636_,
    new_n18637_, new_n18638_, new_n18639_, new_n18640_, new_n18641_,
    new_n18642_, new_n18643_, new_n18644_, new_n18645_, new_n18646_,
    new_n18647_, new_n18648_, new_n18649_, new_n18650_, new_n18651_,
    new_n18652_, new_n18653_, new_n18654_, new_n18655_, new_n18656_,
    new_n18657_, new_n18658_, new_n18659_, new_n18660_, new_n18661_,
    new_n18662_, new_n18663_, new_n18664_, new_n18665_, new_n18666_,
    new_n18667_, new_n18668_, new_n18669_, new_n18670_, new_n18671_,
    new_n18672_, new_n18673_, new_n18674_, new_n18675_, new_n18676_,
    new_n18677_, new_n18678_, new_n18679_, new_n18680_, new_n18681_,
    new_n18682_, new_n18683_, new_n18684_, new_n18685_, new_n18686_,
    new_n18687_, new_n18688_, new_n18689_, new_n18690_, new_n18691_,
    new_n18692_, new_n18693_, new_n18694_, new_n18695_, new_n18696_,
    new_n18697_, new_n18698_, new_n18699_, new_n18700_, new_n18701_,
    new_n18702_, new_n18703_, new_n18704_, new_n18705_, new_n18706_,
    new_n18707_, new_n18708_, new_n18709_, new_n18710_, new_n18711_,
    new_n18712_, new_n18713_, new_n18714_, new_n18715_, new_n18716_,
    new_n18717_, new_n18718_, new_n18719_, new_n18720_, new_n18721_,
    new_n18722_, new_n18723_, new_n18724_, new_n18725_, new_n18726_,
    new_n18727_, new_n18728_, new_n18729_, new_n18730_, new_n18731_,
    new_n18732_, new_n18733_, new_n18734_, new_n18735_, new_n18736_,
    new_n18737_, new_n18738_, new_n18739_, new_n18740_, new_n18741_,
    new_n18742_, new_n18743_, new_n18744_, new_n18745_, new_n18746_,
    new_n18747_, new_n18748_, new_n18749_, new_n18750_, new_n18751_,
    new_n18752_, new_n18753_, new_n18754_, new_n18755_, new_n18756_,
    new_n18757_, new_n18758_, new_n18759_, new_n18760_, new_n18761_,
    new_n18762_, new_n18763_, new_n18764_, new_n18765_, new_n18766_,
    new_n18767_, new_n18768_, new_n18769_, new_n18770_, new_n18771_,
    new_n18772_, new_n18773_, new_n18774_, new_n18775_, new_n18776_,
    new_n18777_, new_n18778_, new_n18779_, new_n18780_, new_n18781_,
    new_n18782_, new_n18783_, new_n18784_, new_n18785_, new_n18786_,
    new_n18787_, new_n18788_, new_n18789_, new_n18790_, new_n18791_,
    new_n18792_, new_n18793_, new_n18794_, new_n18795_, new_n18796_,
    new_n18797_, new_n18798_, new_n18799_, new_n18800_, new_n18801_,
    new_n18802_, new_n18803_, new_n18804_, new_n18805_, new_n18806_,
    new_n18807_, new_n18808_, new_n18809_, new_n18810_, new_n18811_,
    new_n18812_, new_n18813_, new_n18814_, new_n18815_, new_n18816_,
    new_n18817_, new_n18818_, new_n18819_, new_n18820_, new_n18821_,
    new_n18822_, new_n18823_, new_n18824_, new_n18825_, new_n18826_,
    new_n18827_, new_n18828_, new_n18829_, new_n18830_, new_n18831_,
    new_n18832_, new_n18833_, new_n18834_, new_n18835_, new_n18836_,
    new_n18837_, new_n18838_, new_n18839_, new_n18840_, new_n18841_,
    new_n18842_, new_n18843_, new_n18844_, new_n18845_, new_n18846_,
    new_n18847_, new_n18848_, new_n18849_, new_n18850_, new_n18851_,
    new_n18852_, new_n18853_, new_n18854_, new_n18855_, new_n18856_,
    new_n18857_, new_n18858_, new_n18859_, new_n18860_, new_n18861_,
    new_n18862_, new_n18863_, new_n18864_, new_n18865_, new_n18866_,
    new_n18867_, new_n18868_, new_n18869_, new_n18870_, new_n18871_,
    new_n18872_, new_n18873_, new_n18874_, new_n18875_, new_n18876_,
    new_n18877_, new_n18878_, new_n18879_, new_n18880_, new_n18881_,
    new_n18882_, new_n18883_, new_n18884_, new_n18885_, new_n18886_,
    new_n18887_, new_n18888_, new_n18889_, new_n18890_, new_n18891_,
    new_n18892_, new_n18893_, new_n18894_, new_n18895_, new_n18896_,
    new_n18897_, new_n18898_, new_n18899_, new_n18900_, new_n18901_,
    new_n18902_, new_n18903_, new_n18904_, new_n18905_, new_n18906_,
    new_n18907_, new_n18908_, new_n18909_, new_n18910_, new_n18911_,
    new_n18912_, new_n18913_, new_n18914_, new_n18915_, new_n18916_,
    new_n18917_, new_n18918_, new_n18919_, new_n18920_, new_n18921_,
    new_n18922_, new_n18923_, new_n18924_, new_n18925_, new_n18926_,
    new_n18927_, new_n18928_, new_n18929_, new_n18930_, new_n18931_,
    new_n18932_, new_n18933_, new_n18934_, new_n18935_, new_n18936_,
    new_n18937_, new_n18938_, new_n18939_, new_n18940_, new_n18941_,
    new_n18942_, new_n18943_, new_n18944_, new_n18945_, new_n18946_,
    new_n18947_, new_n18948_, new_n18949_, new_n18950_, new_n18951_,
    new_n18952_, new_n18953_, new_n18954_, new_n18955_, new_n18956_,
    new_n18957_, new_n18958_, new_n18959_, new_n18960_, new_n18961_,
    new_n18962_, new_n18963_, new_n18964_, new_n18965_, new_n18966_,
    new_n18967_, new_n18968_, new_n18969_, new_n18970_, new_n18971_,
    new_n18972_, new_n18973_, new_n18974_, new_n18975_, new_n18976_,
    new_n18977_, new_n18978_, new_n18979_, new_n18980_, new_n18981_,
    new_n18982_, new_n18983_, new_n18984_, new_n18985_, new_n18986_,
    new_n18987_, new_n18988_, new_n18989_, new_n18990_, new_n18991_,
    new_n18992_, new_n18993_, new_n18994_, new_n18995_, new_n18996_,
    new_n18997_, new_n18998_, new_n18999_, new_n19000_, new_n19001_,
    new_n19002_, new_n19003_, new_n19004_, new_n19005_, new_n19006_,
    new_n19007_, new_n19008_, new_n19009_, new_n19010_, new_n19011_,
    new_n19012_, new_n19013_, new_n19014_, new_n19015_, new_n19016_,
    new_n19017_, new_n19018_, new_n19019_, new_n19020_, new_n19021_,
    new_n19022_, new_n19023_, new_n19024_, new_n19025_, new_n19026_,
    new_n19027_, new_n19028_, new_n19029_, new_n19030_, new_n19031_,
    new_n19032_, new_n19033_, new_n19034_, new_n19035_, new_n19036_,
    new_n19037_, new_n19038_, new_n19039_, new_n19040_, new_n19041_,
    new_n19042_, new_n19043_, new_n19044_, new_n19045_, new_n19046_,
    new_n19047_, new_n19048_, new_n19049_, new_n19050_, new_n19051_,
    new_n19052_, new_n19053_, new_n19054_, new_n19055_, new_n19056_,
    new_n19057_, new_n19058_, new_n19059_, new_n19060_, new_n19061_,
    new_n19062_, new_n19063_, new_n19064_, new_n19065_, new_n19066_,
    new_n19067_, new_n19068_, new_n19069_, new_n19070_, new_n19071_,
    new_n19072_, new_n19073_, new_n19074_, new_n19075_, new_n19076_,
    new_n19077_, new_n19078_, new_n19079_, new_n19080_, new_n19081_,
    new_n19082_, new_n19083_, new_n19084_, new_n19085_, new_n19086_,
    new_n19087_, new_n19088_, new_n19089_, new_n19090_, new_n19091_,
    new_n19092_, new_n19093_, new_n19094_, new_n19095_, new_n19096_,
    new_n19097_, new_n19098_, new_n19099_, new_n19100_, new_n19101_,
    new_n19102_, new_n19103_, new_n19104_, new_n19105_, new_n19106_,
    new_n19107_, new_n19108_, new_n19109_, new_n19110_, new_n19111_,
    new_n19112_, new_n19113_, new_n19114_, new_n19115_, new_n19116_,
    new_n19117_, new_n19118_, new_n19119_, new_n19120_, new_n19121_,
    new_n19122_, new_n19123_, new_n19124_, new_n19125_, new_n19126_,
    new_n19127_, new_n19128_, new_n19129_, new_n19130_, new_n19131_,
    new_n19132_, new_n19133_, new_n19134_, new_n19135_, new_n19136_,
    new_n19137_, new_n19138_, new_n19139_, new_n19140_, new_n19141_,
    new_n19142_, new_n19143_, new_n19144_, new_n19145_, new_n19146_,
    new_n19147_, new_n19148_, new_n19149_, new_n19150_, new_n19151_,
    new_n19152_, new_n19153_, new_n19154_, new_n19155_, new_n19156_,
    new_n19157_, new_n19158_, new_n19159_, new_n19160_, new_n19161_,
    new_n19162_, new_n19163_, new_n19164_, new_n19165_, new_n19166_,
    new_n19167_, new_n19168_, new_n19169_, new_n19170_, new_n19171_,
    new_n19172_, new_n19173_, new_n19174_, new_n19175_, new_n19176_,
    new_n19177_, new_n19178_, new_n19179_, new_n19180_, new_n19181_,
    new_n19182_, new_n19183_, new_n19184_, new_n19185_, new_n19186_,
    new_n19187_, new_n19188_, new_n19189_, new_n19190_, new_n19191_,
    new_n19192_, new_n19193_, new_n19194_, new_n19195_, new_n19196_,
    new_n19197_, new_n19198_, new_n19199_, new_n19200_, new_n19201_,
    new_n19202_, new_n19203_, new_n19204_, new_n19205_, new_n19206_,
    new_n19207_, new_n19208_, new_n19209_, new_n19210_, new_n19211_,
    new_n19212_, new_n19213_, new_n19214_, new_n19215_, new_n19216_,
    new_n19217_, new_n19218_, new_n19219_, new_n19220_, new_n19221_,
    new_n19222_, new_n19223_, new_n19224_, new_n19225_, new_n19226_,
    new_n19227_, new_n19228_, new_n19229_, new_n19230_, new_n19231_,
    new_n19232_, new_n19233_, new_n19234_, new_n19235_, new_n19236_,
    new_n19237_, new_n19238_, new_n19239_, new_n19240_, new_n19241_,
    new_n19242_, new_n19243_, new_n19244_, new_n19245_, new_n19246_,
    new_n19247_, new_n19248_, new_n19249_, new_n19250_, new_n19251_,
    new_n19252_, new_n19253_, new_n19254_, new_n19255_, new_n19256_,
    new_n19257_, new_n19258_, new_n19259_, new_n19260_, new_n19261_,
    new_n19262_, new_n19263_, new_n19264_, new_n19265_, new_n19266_,
    new_n19267_, new_n19268_, new_n19269_, new_n19270_, new_n19271_,
    new_n19272_, new_n19273_, new_n19274_, new_n19275_, new_n19276_,
    new_n19277_, new_n19278_, new_n19279_, new_n19280_, new_n19281_,
    new_n19282_, new_n19283_, new_n19284_, new_n19285_, new_n19286_,
    new_n19287_, new_n19288_, new_n19289_, new_n19290_, new_n19291_,
    new_n19292_, new_n19293_, new_n19294_, new_n19295_, new_n19296_,
    new_n19297_, new_n19298_, new_n19299_, new_n19300_, new_n19301_,
    new_n19302_, new_n19303_, new_n19304_, new_n19305_, new_n19306_,
    new_n19307_, new_n19308_, new_n19309_, new_n19310_, new_n19311_,
    new_n19312_, new_n19313_, new_n19314_, new_n19315_, new_n19316_,
    new_n19317_, new_n19318_, new_n19319_, new_n19320_, new_n19321_,
    new_n19322_, new_n19323_, new_n19324_, new_n19325_, new_n19326_,
    new_n19327_, new_n19328_, new_n19329_, new_n19330_, new_n19331_,
    new_n19332_, new_n19333_, new_n19334_, new_n19335_, new_n19336_,
    new_n19337_, new_n19338_, new_n19339_, new_n19340_, new_n19341_,
    new_n19342_, new_n19343_, new_n19344_, new_n19345_, new_n19346_,
    new_n19347_, new_n19348_, new_n19349_, new_n19350_, new_n19351_,
    new_n19352_, new_n19353_, new_n19354_, new_n19355_, new_n19356_,
    new_n19357_, new_n19358_, new_n19359_, new_n19360_, new_n19361_,
    new_n19362_, new_n19363_, new_n19364_, new_n19365_, new_n19366_,
    new_n19367_, new_n19368_, new_n19369_, new_n19370_, new_n19371_,
    new_n19372_, new_n19373_, new_n19374_, new_n19375_, new_n19376_,
    new_n19377_, new_n19378_, new_n19379_, new_n19380_, new_n19381_,
    new_n19382_, new_n19383_, new_n19384_, new_n19385_, new_n19386_,
    new_n19387_, new_n19388_, new_n19389_, new_n19390_, new_n19391_,
    new_n19392_, new_n19393_, new_n19394_, new_n19395_, new_n19396_,
    new_n19397_, new_n19398_, new_n19399_, new_n19400_, new_n19401_,
    new_n19402_, new_n19403_, new_n19404_, new_n19405_, new_n19406_,
    new_n19407_, new_n19408_, new_n19409_, new_n19410_, new_n19411_,
    new_n19412_, new_n19413_, new_n19414_, new_n19415_, new_n19416_,
    new_n19417_, new_n19418_, new_n19419_, new_n19420_, new_n19421_,
    new_n19422_, new_n19423_, new_n19424_, new_n19425_, new_n19426_,
    new_n19427_, new_n19428_, new_n19429_, new_n19430_, new_n19431_,
    new_n19432_, new_n19433_, new_n19434_, new_n19435_, new_n19436_,
    new_n19437_, new_n19438_, new_n19439_, new_n19440_, new_n19441_,
    new_n19442_, new_n19443_, new_n19444_, new_n19445_, new_n19446_,
    new_n19447_, new_n19448_, new_n19449_, new_n19450_, new_n19451_,
    new_n19452_, new_n19453_, new_n19454_, new_n19455_, new_n19456_,
    new_n19457_, new_n19458_, new_n19459_, new_n19460_, new_n19461_,
    new_n19462_, new_n19463_, new_n19464_, new_n19465_, new_n19466_,
    new_n19467_, new_n19468_, new_n19469_, new_n19470_, new_n19471_,
    new_n19472_, new_n19473_, new_n19474_, new_n19475_, new_n19476_,
    new_n19477_, new_n19478_, new_n19479_, new_n19480_, new_n19481_,
    new_n19482_, new_n19483_, new_n19484_, new_n19485_, new_n19486_,
    new_n19487_, new_n19488_, new_n19489_, new_n19490_, new_n19491_,
    new_n19492_, new_n19493_, new_n19494_, new_n19495_, new_n19496_,
    new_n19497_, new_n19498_, new_n19499_, new_n19500_, new_n19501_,
    new_n19502_, new_n19503_, new_n19504_, new_n19505_, new_n19506_,
    new_n19507_, new_n19508_, new_n19509_, new_n19510_, new_n19511_,
    new_n19512_, new_n19513_, new_n19514_, new_n19515_, new_n19516_,
    new_n19517_, new_n19518_, new_n19519_, new_n19520_, new_n19521_,
    new_n19522_, new_n19523_, new_n19524_, new_n19525_, new_n19526_,
    new_n19527_, new_n19528_, new_n19529_, new_n19530_, new_n19531_,
    new_n19532_, new_n19533_, new_n19534_, new_n19535_, new_n19536_,
    new_n19537_, new_n19538_, new_n19539_, new_n19540_, new_n19541_,
    new_n19542_, new_n19543_, new_n19544_, new_n19545_, new_n19546_,
    new_n19547_, new_n19548_, new_n19549_, new_n19550_, new_n19551_,
    new_n19552_, new_n19553_, new_n19554_, new_n19555_, new_n19556_,
    new_n19557_, new_n19558_, new_n19559_, new_n19560_, new_n19561_,
    new_n19562_, new_n19563_, new_n19564_, new_n19565_, new_n19566_,
    new_n19567_, new_n19568_, new_n19569_, new_n19570_, new_n19571_,
    new_n19572_, new_n19573_, new_n19574_, new_n19575_, new_n19576_,
    new_n19577_, new_n19578_, new_n19579_, new_n19580_, new_n19581_,
    new_n19582_, new_n19583_, new_n19584_, new_n19585_, new_n19586_,
    new_n19587_, new_n19588_, new_n19589_, new_n19590_, new_n19591_,
    new_n19592_, new_n19593_, new_n19594_, new_n19595_, new_n19596_,
    new_n19597_, new_n19598_, new_n19599_, new_n19600_, new_n19601_,
    new_n19602_, new_n19603_, new_n19604_, new_n19605_, new_n19606_,
    new_n19607_, new_n19608_, new_n19609_, new_n19610_, new_n19611_,
    new_n19612_, new_n19613_, new_n19614_, new_n19615_, new_n19616_,
    new_n19617_, new_n19618_, new_n19619_, new_n19620_, new_n19621_,
    new_n19622_, new_n19623_, new_n19624_, new_n19625_, new_n19626_,
    new_n19627_, new_n19628_, new_n19629_, new_n19630_, new_n19631_,
    new_n19632_, new_n19633_, new_n19634_, new_n19635_, new_n19636_,
    new_n19637_, new_n19638_, new_n19639_, new_n19640_, new_n19641_,
    new_n19642_, new_n19643_, new_n19644_, new_n19645_, new_n19646_,
    new_n19647_, new_n19648_, new_n19649_, new_n19650_, new_n19651_,
    new_n19652_, new_n19653_, new_n19654_, new_n19655_, new_n19656_,
    new_n19657_, new_n19658_, new_n19659_, new_n19660_, new_n19661_,
    new_n19662_, new_n19663_, new_n19664_, new_n19665_, new_n19666_,
    new_n19667_, new_n19668_, new_n19669_, new_n19670_, new_n19671_,
    new_n19672_, new_n19673_, new_n19674_, new_n19675_, new_n19676_,
    new_n19677_, new_n19678_, new_n19679_, new_n19680_, new_n19681_,
    new_n19682_, new_n19683_, new_n19684_, new_n19685_, new_n19686_,
    new_n19687_, new_n19688_, new_n19689_, new_n19690_, new_n19691_,
    new_n19692_, new_n19693_, new_n19694_, new_n19695_, new_n19696_,
    new_n19697_, new_n19698_, new_n19699_, new_n19700_, new_n19701_,
    new_n19702_, new_n19703_, new_n19704_, new_n19705_, new_n19706_,
    new_n19707_, new_n19708_, new_n19709_, new_n19710_, new_n19711_,
    new_n19712_, new_n19713_, new_n19714_, new_n19715_, new_n19716_,
    new_n19717_, new_n19718_, new_n19719_, new_n19720_, new_n19721_,
    new_n19722_, new_n19723_, new_n19724_, new_n19725_, new_n19726_,
    new_n19727_, new_n19728_, new_n19729_, new_n19730_, new_n19731_,
    new_n19732_, new_n19733_, new_n19734_, new_n19735_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19842_, new_n19843_, new_n19844_, new_n19845_, new_n19846_,
    new_n19847_, new_n19848_, new_n19849_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20153_, new_n20154_, new_n20155_, new_n20156_,
    new_n20157_, new_n20158_, new_n20159_, new_n20160_, new_n20161_,
    new_n20162_, new_n20163_, new_n20164_, new_n20165_, new_n20166_,
    new_n20167_, new_n20168_, new_n20169_, new_n20170_, new_n20171_,
    new_n20172_, new_n20173_, new_n20174_, new_n20175_, new_n20176_,
    new_n20177_, new_n20178_, new_n20179_, new_n20180_, new_n20181_,
    new_n20182_, new_n20183_, new_n20184_, new_n20185_, new_n20186_,
    new_n20187_, new_n20188_, new_n20189_, new_n20190_, new_n20191_,
    new_n20192_, new_n20193_, new_n20194_, new_n20195_, new_n20196_,
    new_n20197_, new_n20198_, new_n20199_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20296_,
    new_n20297_, new_n20298_, new_n20299_, new_n20300_, new_n20301_,
    new_n20302_, new_n20303_, new_n20304_, new_n20305_, new_n20306_,
    new_n20307_, new_n20308_, new_n20309_, new_n20310_, new_n20311_,
    new_n20312_, new_n20313_, new_n20314_, new_n20315_, new_n20316_,
    new_n20317_, new_n20318_, new_n20319_, new_n20320_, new_n20321_,
    new_n20322_, new_n20323_, new_n20324_, new_n20325_, new_n20326_,
    new_n20327_, new_n20328_, new_n20329_, new_n20330_, new_n20331_,
    new_n20332_, new_n20333_, new_n20334_, new_n20335_, new_n20336_,
    new_n20337_, new_n20338_, new_n20339_, new_n20340_, new_n20341_,
    new_n20342_, new_n20343_, new_n20344_, new_n20345_, new_n20346_,
    new_n20347_, new_n20348_, new_n20349_, new_n20350_, new_n20351_,
    new_n20352_, new_n20353_, new_n20354_, new_n20355_, new_n20356_,
    new_n20357_, new_n20358_, new_n20359_, new_n20360_, new_n20361_,
    new_n20362_, new_n20363_, new_n20364_, new_n20365_, new_n20366_,
    new_n20367_, new_n20368_, new_n20369_, new_n20370_, new_n20371_,
    new_n20372_, new_n20373_, new_n20374_, new_n20375_, new_n20376_,
    new_n20377_, new_n20378_, new_n20379_, new_n20380_, new_n20381_,
    new_n20382_, new_n20383_, new_n20384_, new_n20385_, new_n20386_,
    new_n20387_, new_n20388_, new_n20389_, new_n20390_, new_n20391_,
    new_n20392_, new_n20393_, new_n20394_, new_n20395_, new_n20396_,
    new_n20397_, new_n20398_, new_n20399_, new_n20400_, new_n20401_,
    new_n20402_, new_n20403_, new_n20404_, new_n20405_, new_n20406_,
    new_n20407_, new_n20408_, new_n20409_, new_n20410_, new_n20411_,
    new_n20412_, new_n20413_, new_n20414_, new_n20415_, new_n20416_,
    new_n20417_, new_n20418_, new_n20419_, new_n20420_, new_n20421_,
    new_n20422_, new_n20423_, new_n20424_, new_n20425_, new_n20426_,
    new_n20427_, new_n20428_, new_n20429_, new_n20430_, new_n20431_,
    new_n20432_, new_n20433_, new_n20434_, new_n20435_, new_n20436_,
    new_n20437_, new_n20438_, new_n20439_, new_n20440_, new_n20441_,
    new_n20442_, new_n20443_, new_n20444_, new_n20445_, new_n20446_,
    new_n20447_, new_n20448_, new_n20449_, new_n20450_, new_n20451_,
    new_n20452_, new_n20453_, new_n20454_, new_n20455_, new_n20456_,
    new_n20457_, new_n20458_, new_n20459_, new_n20460_, new_n20461_,
    new_n20462_, new_n20463_, new_n20464_, new_n20465_, new_n20466_,
    new_n20467_, new_n20468_, new_n20469_, new_n20470_, new_n20471_,
    new_n20472_, new_n20473_, new_n20474_, new_n20475_, new_n20476_,
    new_n20477_, new_n20478_, new_n20479_, new_n20480_, new_n20481_,
    new_n20482_, new_n20483_, new_n20484_, new_n20485_, new_n20486_,
    new_n20487_, new_n20488_, new_n20489_, new_n20490_, new_n20491_,
    new_n20492_, new_n20493_, new_n20494_, new_n20495_, new_n20496_,
    new_n20497_, new_n20498_, new_n20499_, new_n20500_, new_n20501_,
    new_n20502_, new_n20503_, new_n20504_, new_n20505_, new_n20506_,
    new_n20507_, new_n20508_, new_n20509_, new_n20510_, new_n20511_,
    new_n20512_, new_n20513_, new_n20514_, new_n20515_, new_n20516_,
    new_n20517_, new_n20518_, new_n20519_, new_n20520_, new_n20521_,
    new_n20522_, new_n20523_, new_n20524_, new_n20525_, new_n20526_,
    new_n20527_, new_n20528_, new_n20529_, new_n20530_, new_n20531_,
    new_n20532_, new_n20533_, new_n20534_, new_n20535_, new_n20536_,
    new_n20537_, new_n20538_, new_n20539_, new_n20540_, new_n20541_,
    new_n20542_, new_n20543_, new_n20544_, new_n20545_, new_n20546_,
    new_n20547_, new_n20548_, new_n20549_, new_n20550_, new_n20551_,
    new_n20552_, new_n20553_, new_n20554_, new_n20555_, new_n20556_,
    new_n20557_, new_n20558_, new_n20559_, new_n20560_, new_n20561_,
    new_n20562_, new_n20563_, new_n20564_, new_n20565_, new_n20566_,
    new_n20567_, new_n20568_, new_n20569_, new_n20570_, new_n20571_,
    new_n20572_, new_n20573_, new_n20574_, new_n20575_, new_n20576_,
    new_n20577_, new_n20578_, new_n20579_, new_n20580_, new_n20581_,
    new_n20582_, new_n20583_, new_n20584_, new_n20585_, new_n20586_,
    new_n20587_, new_n20588_, new_n20589_, new_n20590_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20677_, new_n20678_, new_n20679_, new_n20680_, new_n20681_,
    new_n20682_, new_n20683_, new_n20684_, new_n20685_, new_n20686_,
    new_n20687_, new_n20688_, new_n20689_, new_n20690_, new_n20691_,
    new_n20692_, new_n20693_, new_n20694_, new_n20695_, new_n20696_,
    new_n20697_, new_n20698_, new_n20699_, new_n20700_, new_n20701_,
    new_n20702_, new_n20703_, new_n20704_, new_n20705_, new_n20706_,
    new_n20707_, new_n20708_, new_n20709_, new_n20710_, new_n20711_,
    new_n20712_, new_n20713_, new_n20714_, new_n20715_, new_n20716_,
    new_n20717_, new_n20718_, new_n20719_, new_n20720_, new_n20721_,
    new_n20722_, new_n20723_, new_n20724_, new_n20725_, new_n20726_,
    new_n20727_, new_n20728_, new_n20729_, new_n20730_, new_n20731_,
    new_n20732_, new_n20733_, new_n20734_, new_n20735_, new_n20736_,
    new_n20737_, new_n20738_, new_n20739_, new_n20740_, new_n20741_,
    new_n20742_, new_n20743_, new_n20744_, new_n20745_, new_n20746_,
    new_n20747_, new_n20748_, new_n20749_, new_n20750_, new_n20751_,
    new_n20752_, new_n20753_, new_n20754_, new_n20755_, new_n20756_,
    new_n20757_, new_n20758_, new_n20759_, new_n20760_, new_n20761_,
    new_n20762_, new_n20763_, new_n20764_, new_n20765_, new_n20766_,
    new_n20767_, new_n20768_, new_n20769_, new_n20770_, new_n20771_,
    new_n20772_, new_n20773_, new_n20774_, new_n20775_, new_n20776_,
    new_n20777_, new_n20778_, new_n20779_, new_n20780_, new_n20781_,
    new_n20782_, new_n20783_, new_n20784_, new_n20785_, new_n20786_,
    new_n20787_, new_n20788_, new_n20789_, new_n20790_, new_n20791_,
    new_n20792_, new_n20793_, new_n20794_, new_n20795_, new_n20796_,
    new_n20797_, new_n20798_, new_n20799_, new_n20800_, new_n20801_,
    new_n20802_, new_n20803_, new_n20804_, new_n20805_, new_n20806_,
    new_n20807_, new_n20808_, new_n20809_, new_n20810_, new_n20811_,
    new_n20812_, new_n20813_, new_n20814_, new_n20815_, new_n20816_,
    new_n20817_, new_n20818_, new_n20819_, new_n20820_, new_n20821_,
    new_n20822_, new_n20823_, new_n20824_, new_n20825_, new_n20826_,
    new_n20827_, new_n20828_, new_n20829_, new_n20830_, new_n20831_,
    new_n20832_, new_n20833_, new_n20834_, new_n20835_, new_n20836_,
    new_n20837_, new_n20838_, new_n20839_, new_n20840_, new_n20841_,
    new_n20842_, new_n20843_, new_n20844_, new_n20845_, new_n20846_,
    new_n20847_, new_n20848_, new_n20849_, new_n20850_, new_n20851_,
    new_n20852_, new_n20853_, new_n20854_, new_n20855_, new_n20856_,
    new_n20857_, new_n20858_, new_n20859_, new_n20860_, new_n20861_,
    new_n20862_, new_n20863_, new_n20864_, new_n20865_, new_n20866_,
    new_n20867_, new_n20868_, new_n20869_, new_n20870_, new_n20871_,
    new_n20872_, new_n20873_, new_n20874_, new_n20875_, new_n20876_,
    new_n20877_, new_n20878_, new_n20879_, new_n20880_, new_n20881_,
    new_n20882_, new_n20883_, new_n20884_, new_n20885_, new_n20886_,
    new_n20887_, new_n20888_, new_n20889_, new_n20890_, new_n20891_,
    new_n20892_, new_n20893_, new_n20894_, new_n20895_, new_n20896_,
    new_n20897_, new_n20898_, new_n20899_, new_n20900_, new_n20901_,
    new_n20902_, new_n20903_, new_n20904_, new_n20905_, new_n20906_,
    new_n20907_, new_n20908_, new_n20909_, new_n20910_, new_n20911_,
    new_n20912_, new_n20913_, new_n20914_, new_n20915_, new_n20916_,
    new_n20917_, new_n20918_, new_n20919_, new_n20920_, new_n20921_,
    new_n20922_, new_n20923_, new_n20924_, new_n20925_, new_n20926_,
    new_n20927_, new_n20928_, new_n20929_, new_n20930_, new_n20931_,
    new_n20932_, new_n20933_, new_n20934_, new_n20935_, new_n20936_,
    new_n20937_, new_n20938_, new_n20939_, new_n20940_, new_n20941_,
    new_n20942_, new_n20943_, new_n20944_, new_n20945_, new_n20946_,
    new_n20947_, new_n20948_, new_n20949_, new_n20950_, new_n20951_,
    new_n20952_, new_n20953_, new_n20954_, new_n20955_, new_n20956_,
    new_n20957_, new_n20958_, new_n20959_, new_n20960_, new_n20961_,
    new_n20962_, new_n20963_, new_n20964_, new_n20965_, new_n20966_,
    new_n20967_, new_n20968_, new_n20969_, new_n20970_, new_n20971_,
    new_n20972_, new_n20973_, new_n20974_, new_n20975_, new_n20976_,
    new_n20977_, new_n20978_, new_n20979_, new_n20980_, new_n20981_,
    new_n20982_, new_n20983_, new_n20984_, new_n20985_, new_n20986_,
    new_n20987_, new_n20988_, new_n20989_, new_n20990_, new_n20991_,
    new_n20992_, new_n20993_, new_n20994_, new_n20995_, new_n20996_,
    new_n20997_, new_n20998_, new_n20999_, new_n21000_, new_n21001_,
    new_n21002_, new_n21003_, new_n21004_, new_n21005_, new_n21006_,
    new_n21007_, new_n21008_, new_n21009_, new_n21010_, new_n21011_,
    new_n21012_, new_n21013_, new_n21014_, new_n21015_, new_n21016_,
    new_n21017_, new_n21018_, new_n21019_, new_n21020_, new_n21021_,
    new_n21022_, new_n21023_, new_n21024_, new_n21025_, new_n21026_,
    new_n21027_, new_n21028_, new_n21029_, new_n21030_, new_n21031_,
    new_n21032_, new_n21033_, new_n21034_, new_n21035_, new_n21036_,
    new_n21037_, new_n21038_, new_n21039_, new_n21040_, new_n21041_,
    new_n21042_, new_n21043_, new_n21044_, new_n21045_, new_n21046_,
    new_n21047_, new_n21048_, new_n21049_, new_n21050_, new_n21051_,
    new_n21052_, new_n21053_, new_n21054_, new_n21055_, new_n21056_,
    new_n21057_, new_n21058_, new_n21059_, new_n21060_, new_n21061_,
    new_n21062_, new_n21063_, new_n21064_, new_n21065_, new_n21066_,
    new_n21067_, new_n21068_, new_n21069_, new_n21070_, new_n21071_,
    new_n21072_, new_n21073_, new_n21074_, new_n21075_, new_n21076_,
    new_n21077_, new_n21078_, new_n21079_, new_n21080_, new_n21081_,
    new_n21082_, new_n21083_, new_n21084_, new_n21085_, new_n21086_,
    new_n21087_, new_n21088_, new_n21089_, new_n21090_, new_n21091_,
    new_n21092_, new_n21093_, new_n21094_, new_n21095_, new_n21096_,
    new_n21097_, new_n21098_, new_n21099_, new_n21100_, new_n21101_,
    new_n21102_, new_n21103_, new_n21104_, new_n21105_, new_n21106_,
    new_n21107_, new_n21108_, new_n21109_, new_n21110_, new_n21111_,
    new_n21112_, new_n21113_, new_n21114_, new_n21115_, new_n21116_,
    new_n21117_, new_n21118_, new_n21119_, new_n21120_, new_n21121_,
    new_n21122_, new_n21123_, new_n21124_, new_n21125_, new_n21126_,
    new_n21127_, new_n21128_, new_n21129_, new_n21130_, new_n21131_,
    new_n21132_, new_n21133_, new_n21134_, new_n21135_, new_n21136_,
    new_n21137_, new_n21138_, new_n21139_, new_n21140_, new_n21141_,
    new_n21142_, new_n21143_, new_n21144_, new_n21145_, new_n21146_,
    new_n21147_, new_n21148_, new_n21149_, new_n21150_, new_n21151_,
    new_n21152_, new_n21153_, new_n21154_, new_n21155_, new_n21156_,
    new_n21157_, new_n21158_, new_n21159_, new_n21160_, new_n21161_,
    new_n21162_, new_n21163_, new_n21164_, new_n21165_, new_n21166_,
    new_n21167_, new_n21168_, new_n21169_, new_n21170_, new_n21171_,
    new_n21172_, new_n21173_, new_n21174_, new_n21175_, new_n21176_,
    new_n21177_, new_n21178_, new_n21179_, new_n21180_, new_n21181_,
    new_n21182_, new_n21183_, new_n21184_, new_n21185_, new_n21186_,
    new_n21187_, new_n21188_, new_n21189_, new_n21190_, new_n21191_,
    new_n21192_, new_n21193_, new_n21194_, new_n21195_, new_n21196_,
    new_n21197_, new_n21198_, new_n21199_, new_n21200_, new_n21201_,
    new_n21202_, new_n21203_, new_n21204_, new_n21205_, new_n21206_,
    new_n21207_, new_n21208_, new_n21209_, new_n21210_, new_n21211_,
    new_n21212_, new_n21213_, new_n21214_, new_n21215_, new_n21216_,
    new_n21217_, new_n21218_, new_n21219_, new_n21220_, new_n21221_,
    new_n21222_, new_n21223_, new_n21224_, new_n21225_, new_n21226_,
    new_n21227_, new_n21228_, new_n21229_, new_n21230_, new_n21231_,
    new_n21232_, new_n21233_, new_n21234_, new_n21235_, new_n21236_,
    new_n21237_, new_n21238_, new_n21239_, new_n21240_, new_n21241_,
    new_n21242_, new_n21243_, new_n21244_, new_n21245_, new_n21246_,
    new_n21247_, new_n21248_, new_n21249_, new_n21250_, new_n21251_,
    new_n21252_, new_n21253_, new_n21254_, new_n21255_, new_n21256_,
    new_n21257_, new_n21258_, new_n21259_, new_n21260_, new_n21261_,
    new_n21262_, new_n21263_, new_n21264_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21270_, new_n21271_,
    new_n21272_, new_n21273_, new_n21274_, new_n21275_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21377_, new_n21378_, new_n21379_, new_n21380_, new_n21381_,
    new_n21382_, new_n21383_, new_n21384_, new_n21385_, new_n21386_,
    new_n21387_, new_n21388_, new_n21389_, new_n21390_, new_n21391_,
    new_n21392_, new_n21393_, new_n21394_, new_n21395_, new_n21396_,
    new_n21397_, new_n21398_, new_n21399_, new_n21400_, new_n21401_,
    new_n21402_, new_n21403_, new_n21404_, new_n21405_, new_n21406_,
    new_n21407_, new_n21408_, new_n21409_, new_n21410_, new_n21411_,
    new_n21412_, new_n21413_, new_n21414_, new_n21415_, new_n21416_,
    new_n21417_, new_n21418_, new_n21419_, new_n21420_, new_n21421_,
    new_n21422_, new_n21423_, new_n21424_, new_n21425_, new_n21426_,
    new_n21427_, new_n21428_, new_n21429_, new_n21430_, new_n21431_,
    new_n21432_, new_n21433_, new_n21434_, new_n21435_, new_n21436_,
    new_n21437_, new_n21438_, new_n21439_, new_n21440_, new_n21441_,
    new_n21442_, new_n21443_, new_n21444_, new_n21445_, new_n21446_,
    new_n21447_, new_n21448_, new_n21449_, new_n21450_, new_n21451_,
    new_n21452_, new_n21453_, new_n21454_, new_n21455_, new_n21456_,
    new_n21457_, new_n21458_, new_n21459_, new_n21460_, new_n21461_,
    new_n21462_, new_n21463_, new_n21464_, new_n21465_, new_n21466_,
    new_n21467_, new_n21468_, new_n21469_, new_n21470_, new_n21471_,
    new_n21472_, new_n21473_, new_n21474_, new_n21475_, new_n21476_,
    new_n21477_, new_n21478_, new_n21479_, new_n21480_, new_n21481_,
    new_n21482_, new_n21483_, new_n21484_, new_n21485_, new_n21486_,
    new_n21487_, new_n21488_, new_n21489_, new_n21490_, new_n21491_,
    new_n21492_, new_n21493_, new_n21494_, new_n21495_, new_n21496_,
    new_n21497_, new_n21498_, new_n21499_, new_n21500_, new_n21501_,
    new_n21502_, new_n21503_, new_n21504_, new_n21505_, new_n21506_,
    new_n21507_, new_n21508_, new_n21509_, new_n21510_, new_n21511_,
    new_n21512_, new_n21513_, new_n21514_, new_n21515_, new_n21516_,
    new_n21517_, new_n21518_, new_n21519_, new_n21520_, new_n21521_,
    new_n21522_, new_n21523_, new_n21524_, new_n21525_, new_n21526_,
    new_n21527_, new_n21528_, new_n21529_, new_n21530_, new_n21531_,
    new_n21532_, new_n21533_, new_n21534_, new_n21535_, new_n21536_,
    new_n21537_, new_n21538_, new_n21539_, new_n21540_, new_n21541_,
    new_n21542_, new_n21543_, new_n21544_, new_n21545_, new_n21546_,
    new_n21547_, new_n21548_, new_n21549_, new_n21550_, new_n21551_,
    new_n21552_, new_n21553_, new_n21554_, new_n21555_, new_n21556_,
    new_n21557_, new_n21558_, new_n21559_, new_n21560_, new_n21561_,
    new_n21562_, new_n21563_, new_n21564_, new_n21565_, new_n21566_,
    new_n21567_, new_n21568_, new_n21569_, new_n21570_, new_n21571_,
    new_n21572_, new_n21573_, new_n21574_, new_n21575_, new_n21576_,
    new_n21577_, new_n21578_, new_n21579_, new_n21580_, new_n21581_,
    new_n21582_, new_n21583_, new_n21584_, new_n21585_, new_n21586_,
    new_n21587_, new_n21588_, new_n21589_, new_n21590_, new_n21591_,
    new_n21592_, new_n21593_, new_n21594_, new_n21595_, new_n21596_,
    new_n21597_, new_n21598_, new_n21599_, new_n21600_, new_n21601_,
    new_n21602_, new_n21603_, new_n21604_, new_n21605_, new_n21606_,
    new_n21607_, new_n21608_, new_n21609_, new_n21610_, new_n21611_,
    new_n21612_, new_n21613_, new_n21614_, new_n21615_, new_n21616_,
    new_n21617_, new_n21618_, new_n21619_, new_n21620_, new_n21621_,
    new_n21622_, new_n21623_, new_n21624_, new_n21625_, new_n21626_,
    new_n21627_, new_n21628_, new_n21629_, new_n21630_, new_n21631_,
    new_n21632_, new_n21633_, new_n21634_, new_n21635_, new_n21636_,
    new_n21637_, new_n21638_, new_n21639_, new_n21640_, new_n21641_,
    new_n21642_, new_n21643_, new_n21644_, new_n21645_, new_n21646_,
    new_n21647_, new_n21648_, new_n21649_, new_n21650_, new_n21651_,
    new_n21652_, new_n21653_, new_n21654_, new_n21655_, new_n21656_,
    new_n21657_, new_n21658_, new_n21659_, new_n21660_, new_n21661_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21670_, new_n21671_,
    new_n21672_, new_n21673_, new_n21674_, new_n21675_, new_n21676_,
    new_n21677_, new_n21678_, new_n21679_, new_n21680_, new_n21681_,
    new_n21682_, new_n21683_, new_n21684_, new_n21685_, new_n21686_,
    new_n21687_, new_n21688_, new_n21689_, new_n21690_, new_n21691_,
    new_n21692_, new_n21693_, new_n21694_, new_n21695_, new_n21696_,
    new_n21697_, new_n21698_, new_n21699_, new_n21700_, new_n21701_,
    new_n21702_, new_n21703_, new_n21704_, new_n21705_, new_n21706_,
    new_n21707_, new_n21708_, new_n21709_, new_n21710_, new_n21711_,
    new_n21712_, new_n21713_, new_n21714_, new_n21715_, new_n21716_,
    new_n21717_, new_n21718_, new_n21719_, new_n21720_, new_n21721_,
    new_n21722_, new_n21723_, new_n21724_, new_n21725_, new_n21726_,
    new_n21727_, new_n21728_, new_n21729_, new_n21730_, new_n21731_,
    new_n21732_, new_n21733_, new_n21734_, new_n21735_, new_n21736_,
    new_n21737_, new_n21738_, new_n21739_, new_n21740_, new_n21741_,
    new_n21742_, new_n21743_, new_n21744_, new_n21745_, new_n21746_,
    new_n21747_, new_n21748_, new_n21749_, new_n21750_, new_n21751_,
    new_n21752_, new_n21753_, new_n21754_, new_n21755_, new_n21756_,
    new_n21757_, new_n21758_, new_n21759_, new_n21760_, new_n21761_,
    new_n21762_, new_n21763_, new_n21764_, new_n21765_, new_n21766_,
    new_n21767_, new_n21768_, new_n21769_, new_n21770_, new_n21771_,
    new_n21772_, new_n21773_, new_n21774_, new_n21775_, new_n21776_,
    new_n21777_, new_n21778_, new_n21779_, new_n21780_, new_n21781_,
    new_n21782_, new_n21783_, new_n21784_, new_n21785_, new_n21786_,
    new_n21787_, new_n21788_, new_n21789_, new_n21790_, new_n21791_,
    new_n21792_, new_n21793_, new_n21794_, new_n21795_, new_n21796_,
    new_n21797_, new_n21798_, new_n21799_, new_n21800_, new_n21801_,
    new_n21802_, new_n21803_, new_n21804_, new_n21805_, new_n21806_,
    new_n21807_, new_n21808_, new_n21809_, new_n21810_, new_n21811_,
    new_n21812_, new_n21813_, new_n21814_, new_n21815_, new_n21816_,
    new_n21817_, new_n21818_, new_n21819_, new_n21820_, new_n21821_,
    new_n21822_, new_n21823_, new_n21824_, new_n21825_, new_n21826_,
    new_n21827_, new_n21828_, new_n21829_, new_n21830_, new_n21831_,
    new_n21832_, new_n21833_, new_n21834_, new_n21835_, new_n21836_,
    new_n21837_, new_n21838_, new_n21839_, new_n21840_, new_n21841_,
    new_n21842_, new_n21843_, new_n21844_, new_n21845_, new_n21846_,
    new_n21847_, new_n21848_, new_n21849_, new_n21850_, new_n21851_,
    new_n21852_, new_n21853_, new_n21854_, new_n21855_, new_n21856_,
    new_n21857_, new_n21858_, new_n21859_, new_n21860_, new_n21861_,
    new_n21862_, new_n21863_, new_n21864_, new_n21865_, new_n21866_,
    new_n21867_, new_n21868_, new_n21869_, new_n21870_, new_n21871_,
    new_n21872_, new_n21873_, new_n21874_, new_n21875_, new_n21876_,
    new_n21877_, new_n21878_, new_n21879_, new_n21880_, new_n21881_,
    new_n21882_, new_n21883_, new_n21884_, new_n21885_, new_n21886_,
    new_n21887_, new_n21888_, new_n21889_, new_n21890_, new_n21891_,
    new_n21892_, new_n21893_, new_n21894_, new_n21895_, new_n21896_,
    new_n21897_, new_n21898_, new_n21899_, new_n21900_, new_n21901_,
    new_n21902_, new_n21903_, new_n21904_, new_n21905_, new_n21906_,
    new_n21907_, new_n21908_, new_n21909_, new_n21910_, new_n21911_,
    new_n21912_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22014_, new_n22015_, new_n22016_,
    new_n22017_, new_n22018_, new_n22019_, new_n22020_, new_n22021_,
    new_n22022_, new_n22023_, new_n22024_, new_n22025_, new_n22026_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22035_, new_n22036_,
    new_n22037_, new_n22038_, new_n22039_, new_n22040_, new_n22041_,
    new_n22042_, new_n22043_, new_n22044_, new_n22045_, new_n22046_,
    new_n22047_, new_n22048_, new_n22049_, new_n22050_, new_n22051_,
    new_n22052_, new_n22053_, new_n22054_, new_n22055_, new_n22056_,
    new_n22057_, new_n22058_, new_n22059_, new_n22060_, new_n22061_,
    new_n22062_, new_n22063_, new_n22064_, new_n22065_, new_n22066_,
    new_n22067_, new_n22068_, new_n22069_, new_n22070_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22143_, new_n22144_, new_n22145_, new_n22146_,
    new_n22147_, new_n22148_, new_n22149_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22156_,
    new_n22157_, new_n22158_, new_n22159_, new_n22160_, new_n22161_,
    new_n22162_, new_n22163_, new_n22164_, new_n22165_, new_n22166_,
    new_n22167_, new_n22168_, new_n22169_, new_n22170_, new_n22171_,
    new_n22172_, new_n22173_, new_n22174_, new_n22175_, new_n22176_,
    new_n22177_, new_n22178_, new_n22179_, new_n22180_, new_n22181_,
    new_n22182_, new_n22183_, new_n22184_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22303_, new_n22304_, new_n22305_, new_n22306_,
    new_n22307_, new_n22308_, new_n22309_, new_n22310_, new_n22311_,
    new_n22312_, new_n22313_, new_n22314_, new_n22315_, new_n22316_,
    new_n22317_, new_n22318_, new_n22319_, new_n22320_, new_n22321_,
    new_n22322_, new_n22323_, new_n22324_, new_n22325_, new_n22326_,
    new_n22327_, new_n22328_, new_n22329_, new_n22330_, new_n22331_,
    new_n22332_, new_n22333_, new_n22334_, new_n22335_, new_n22336_,
    new_n22337_, new_n22338_, new_n22339_, new_n22340_, new_n22341_,
    new_n22342_, new_n22343_, new_n22344_, new_n22345_, new_n22346_,
    new_n22347_, new_n22348_, new_n22349_, new_n22350_, new_n22351_,
    new_n22352_, new_n22353_, new_n22354_, new_n22355_, new_n22356_,
    new_n22357_, new_n22358_, new_n22359_, new_n22360_, new_n22361_,
    new_n22362_, new_n22363_, new_n22364_, new_n22365_, new_n22366_,
    new_n22367_, new_n22368_, new_n22369_, new_n22370_, new_n22371_,
    new_n22372_, new_n22373_, new_n22374_, new_n22375_, new_n22376_,
    new_n22377_, new_n22378_, new_n22379_, new_n22380_, new_n22381_,
    new_n22382_, new_n22383_, new_n22384_, new_n22385_, new_n22386_,
    new_n22387_, new_n22388_, new_n22389_, new_n22390_, new_n22391_,
    new_n22392_, new_n22393_, new_n22394_, new_n22395_, new_n22396_,
    new_n22397_, new_n22398_, new_n22399_, new_n22400_, new_n22401_,
    new_n22402_, new_n22403_, new_n22404_, new_n22405_, new_n22406_,
    new_n22407_, new_n22408_, new_n22409_, new_n22410_, new_n22411_,
    new_n22412_, new_n22413_, new_n22414_, new_n22415_, new_n22416_,
    new_n22417_, new_n22418_, new_n22419_, new_n22420_, new_n22421_,
    new_n22422_, new_n22423_, new_n22424_, new_n22425_, new_n22426_,
    new_n22427_, new_n22428_, new_n22429_, new_n22430_, new_n22431_,
    new_n22432_, new_n22433_, new_n22434_, new_n22435_, new_n22436_,
    new_n22437_, new_n22438_, new_n22439_, new_n22440_, new_n22441_,
    new_n22442_, new_n22443_, new_n22444_, new_n22445_, new_n22446_,
    new_n22447_, new_n22448_, new_n22449_, new_n22450_, new_n22451_,
    new_n22452_, new_n22453_, new_n22454_, new_n22455_, new_n22456_,
    new_n22457_, new_n22458_, new_n22459_, new_n22460_, new_n22461_,
    new_n22462_, new_n22463_, new_n22464_, new_n22465_, new_n22466_,
    new_n22467_, new_n22468_, new_n22469_, new_n22470_, new_n22471_,
    new_n22472_, new_n22473_, new_n22474_, new_n22475_, new_n22476_,
    new_n22477_, new_n22478_, new_n22479_, new_n22480_, new_n22481_,
    new_n22482_, new_n22483_, new_n22484_, new_n22485_, new_n22486_,
    new_n22487_, new_n22488_, new_n22489_, new_n22490_, new_n22491_,
    new_n22492_, new_n22493_, new_n22494_, new_n22495_, new_n22496_,
    new_n22497_, new_n22498_, new_n22499_, new_n22500_, new_n22501_,
    new_n22502_, new_n22503_, new_n22504_, new_n22505_, new_n22506_,
    new_n22507_, new_n22508_, new_n22509_, new_n22510_, new_n22511_,
    new_n22512_, new_n22513_, new_n22514_, new_n22515_, new_n22516_,
    new_n22517_, new_n22518_, new_n22519_, new_n22520_, new_n22521_,
    new_n22522_, new_n22523_, new_n22524_, new_n22525_, new_n22526_,
    new_n22527_, new_n22528_, new_n22529_, new_n22530_, new_n22531_,
    new_n22532_, new_n22533_, new_n22534_, new_n22535_, new_n22536_,
    new_n22537_, new_n22538_, new_n22539_, new_n22540_, new_n22541_,
    new_n22542_, new_n22543_, new_n22544_, new_n22545_, new_n22546_,
    new_n22547_, new_n22548_, new_n22549_, new_n22550_, new_n22551_,
    new_n22552_, new_n22553_, new_n22554_, new_n22555_, new_n22556_,
    new_n22557_, new_n22558_, new_n22559_, new_n22560_, new_n22561_,
    new_n22562_, new_n22563_, new_n22564_, new_n22565_, new_n22566_,
    new_n22567_, new_n22568_, new_n22569_, new_n22570_, new_n22571_,
    new_n22572_, new_n22573_, new_n22574_, new_n22575_, new_n22576_,
    new_n22577_, new_n22578_, new_n22579_, new_n22580_, new_n22581_,
    new_n22582_, new_n22583_, new_n22584_, new_n22585_, new_n22586_,
    new_n22587_, new_n22588_, new_n22589_, new_n22590_, new_n22591_,
    new_n22592_, new_n22593_, new_n22594_, new_n22595_, new_n22596_,
    new_n22597_, new_n22598_, new_n22599_, new_n22600_, new_n22601_,
    new_n22602_, new_n22603_, new_n22604_, new_n22605_, new_n22606_,
    new_n22607_, new_n22608_, new_n22609_, new_n22610_, new_n22611_,
    new_n22612_, new_n22613_, new_n22614_, new_n22615_, new_n22616_,
    new_n22617_, new_n22618_, new_n22619_, new_n22620_, new_n22621_,
    new_n22622_, new_n22623_, new_n22624_, new_n22625_, new_n22626_,
    new_n22627_, new_n22628_, new_n22629_, new_n22630_, new_n22631_,
    new_n22632_, new_n22633_, new_n22634_, new_n22635_, new_n22636_,
    new_n22637_, new_n22638_, new_n22639_, new_n22640_, new_n22641_,
    new_n22642_, new_n22643_, new_n22644_, new_n22645_, new_n22646_,
    new_n22647_, new_n22648_, new_n22649_, new_n22650_, new_n22651_,
    new_n22652_, new_n22653_, new_n22654_, new_n22655_, new_n22656_,
    new_n22657_, new_n22658_, new_n22659_, new_n22660_, new_n22661_,
    new_n22662_, new_n22663_, new_n22664_, new_n22665_, new_n22666_,
    new_n22667_, new_n22668_, new_n22669_, new_n22670_, new_n22671_,
    new_n22672_, new_n22673_, new_n22674_, new_n22675_, new_n22676_,
    new_n22677_, new_n22678_, new_n22679_, new_n22680_, new_n22681_,
    new_n22682_, new_n22683_, new_n22684_, new_n22685_, new_n22686_,
    new_n22687_, new_n22688_, new_n22689_, new_n22690_, new_n22691_,
    new_n22692_, new_n22693_, new_n22694_, new_n22695_, new_n22696_,
    new_n22697_, new_n22698_, new_n22699_, new_n22700_, new_n22701_,
    new_n22702_, new_n22703_, new_n22704_, new_n22705_, new_n22706_,
    new_n22707_, new_n22708_, new_n22709_, new_n22710_, new_n22711_,
    new_n22712_, new_n22713_, new_n22714_, new_n22715_, new_n22716_,
    new_n22717_, new_n22718_, new_n22719_, new_n22720_, new_n22721_,
    new_n22722_, new_n22723_, new_n22724_, new_n22725_, new_n22726_,
    new_n22727_, new_n22728_, new_n22729_, new_n22730_, new_n22731_,
    new_n22732_, new_n22733_, new_n22734_, new_n22735_, new_n22736_,
    new_n22737_, new_n22738_, new_n22739_, new_n22740_, new_n22741_,
    new_n22742_, new_n22743_, new_n22744_, new_n22745_, new_n22746_,
    new_n22747_, new_n22748_, new_n22749_, new_n22750_, new_n22751_,
    new_n22752_, new_n22753_, new_n22754_, new_n22755_, new_n22756_,
    new_n22757_, new_n22758_, new_n22759_, new_n22760_, new_n22761_,
    new_n22762_, new_n22763_, new_n22764_, new_n22765_, new_n22766_,
    new_n22767_, new_n22768_, new_n22769_, new_n22770_, new_n22771_,
    new_n22772_, new_n22773_, new_n22774_, new_n22775_, new_n22776_,
    new_n22777_, new_n22778_, new_n22779_, new_n22780_, new_n22781_,
    new_n22782_, new_n22783_, new_n22784_, new_n22785_, new_n22786_,
    new_n22787_, new_n22788_, new_n22789_, new_n22790_, new_n22791_,
    new_n22792_, new_n22793_, new_n22794_, new_n22795_, new_n22796_,
    new_n22797_, new_n22798_, new_n22799_, new_n22800_, new_n22801_,
    new_n22802_, new_n22803_, new_n22804_, new_n22805_, new_n22806_,
    new_n22807_, new_n22808_, new_n22809_, new_n22810_, new_n22811_,
    new_n22812_, new_n22813_, new_n22814_, new_n22815_, new_n22816_,
    new_n22817_, new_n22818_, new_n22819_, new_n22820_, new_n22821_,
    new_n22822_, new_n22823_, new_n22824_, new_n22825_, new_n22826_,
    new_n22827_, new_n22828_, new_n22829_, new_n22830_, new_n22831_,
    new_n22832_, new_n22833_, new_n22834_, new_n22835_, new_n22836_,
    new_n22837_, new_n22838_, new_n22839_, new_n22840_, new_n22841_,
    new_n22842_, new_n22843_, new_n22844_, new_n22845_, new_n22846_,
    new_n22847_, new_n22848_, new_n22849_, new_n22850_, new_n22851_,
    new_n22852_, new_n22853_, new_n22854_, new_n22855_, new_n22856_,
    new_n22857_, new_n22858_, new_n22859_, new_n22860_, new_n22861_,
    new_n22862_, new_n22863_, new_n22864_, new_n22865_, new_n22866_,
    new_n22867_, new_n22868_, new_n22869_, new_n22870_, new_n22871_,
    new_n22872_, new_n22873_, new_n22874_, new_n22875_, new_n22876_,
    new_n22877_, new_n22878_, new_n22879_, new_n22880_, new_n22881_,
    new_n22882_, new_n22883_, new_n22884_, new_n22885_, new_n22886_,
    new_n22887_, new_n22888_, new_n22889_, new_n22890_, new_n22891_,
    new_n22892_, new_n22893_, new_n22894_, new_n22895_, new_n22896_,
    new_n22897_, new_n22898_, new_n22899_, new_n22900_, new_n22901_,
    new_n22902_, new_n22903_, new_n22904_, new_n22905_, new_n22906_,
    new_n22907_, new_n22908_, new_n22909_, new_n22910_, new_n22911_,
    new_n22912_, new_n22913_, new_n22914_, new_n22915_, new_n22916_,
    new_n22917_, new_n22918_, new_n22919_, new_n22920_, new_n22921_,
    new_n22922_, new_n22923_, new_n22924_, new_n22925_, new_n22926_,
    new_n22927_, new_n22928_, new_n22929_, new_n22930_, new_n22931_,
    new_n22932_, new_n22933_, new_n22934_, new_n22935_, new_n22936_,
    new_n22937_, new_n22938_, new_n22939_, new_n22940_, new_n22941_,
    new_n22942_, new_n22943_, new_n22944_, new_n22945_, new_n22946_,
    new_n22947_, new_n22948_, new_n22949_, new_n22950_, new_n22951_,
    new_n22952_, new_n22953_, new_n22954_, new_n22955_, new_n22956_,
    new_n22957_, new_n22958_, new_n22959_, new_n22960_, new_n22961_,
    new_n22962_, new_n22963_, new_n22964_, new_n22965_, new_n22966_,
    new_n22967_, new_n22968_, new_n22969_, new_n22970_, new_n22971_,
    new_n22972_, new_n22973_, new_n22974_, new_n22975_, new_n22976_,
    new_n22977_, new_n22978_, new_n22979_, new_n22980_, new_n22981_,
    new_n22982_, new_n22983_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23001_,
    new_n23002_, new_n23003_, new_n23004_, new_n23005_, new_n23006_,
    new_n23007_, new_n23008_, new_n23009_, new_n23010_, new_n23011_,
    new_n23012_, new_n23013_, new_n23014_, new_n23015_, new_n23016_,
    new_n23017_, new_n23018_, new_n23019_, new_n23020_, new_n23021_,
    new_n23022_, new_n23023_, new_n23024_, new_n23025_, new_n23026_,
    new_n23027_, new_n23028_, new_n23029_, new_n23030_, new_n23031_,
    new_n23032_, new_n23033_, new_n23034_, new_n23035_, new_n23036_,
    new_n23037_, new_n23038_, new_n23039_, new_n23040_, new_n23041_,
    new_n23042_, new_n23043_, new_n23044_, new_n23045_, new_n23046_,
    new_n23047_, new_n23048_, new_n23049_, new_n23050_, new_n23051_,
    new_n23052_, new_n23053_, new_n23054_, new_n23055_, new_n23056_,
    new_n23057_, new_n23058_, new_n23059_, new_n23060_, new_n23061_,
    new_n23062_, new_n23063_, new_n23064_, new_n23065_, new_n23066_,
    new_n23067_, new_n23068_, new_n23069_, new_n23070_, new_n23071_,
    new_n23072_, new_n23073_, new_n23074_, new_n23075_, new_n23076_,
    new_n23077_, new_n23078_, new_n23079_, new_n23080_, new_n23081_,
    new_n23082_, new_n23083_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23089_, new_n23090_, new_n23091_,
    new_n23092_, new_n23093_, new_n23094_, new_n23095_, new_n23096_,
    new_n23097_, new_n23098_, new_n23099_, new_n23100_, new_n23101_,
    new_n23102_, new_n23103_, new_n23104_, new_n23105_, new_n23106_,
    new_n23107_, new_n23108_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23116_,
    new_n23117_, new_n23118_, new_n23119_, new_n23120_, new_n23121_,
    new_n23122_, new_n23123_, new_n23124_, new_n23125_, new_n23126_,
    new_n23127_, new_n23128_, new_n23129_, new_n23130_, new_n23131_,
    new_n23132_, new_n23133_, new_n23134_, new_n23135_, new_n23136_,
    new_n23137_, new_n23138_, new_n23139_, new_n23140_, new_n23141_,
    new_n23142_, new_n23143_, new_n23144_, new_n23145_, new_n23146_,
    new_n23147_, new_n23148_, new_n23149_, new_n23150_, new_n23151_,
    new_n23152_, new_n23153_, new_n23154_, new_n23155_, new_n23156_,
    new_n23157_, new_n23158_, new_n23159_, new_n23160_, new_n23161_,
    new_n23162_, new_n23163_, new_n23164_, new_n23165_, new_n23166_,
    new_n23167_, new_n23168_, new_n23169_, new_n23170_, new_n23171_,
    new_n23172_, new_n23173_, new_n23174_, new_n23175_, new_n23176_,
    new_n23177_, new_n23178_, new_n23179_, new_n23180_, new_n23181_,
    new_n23182_, new_n23183_, new_n23184_, new_n23185_, new_n23186_,
    new_n23187_, new_n23188_, new_n23189_, new_n23190_, new_n23191_,
    new_n23192_, new_n23193_, new_n23194_, new_n23195_, new_n23196_,
    new_n23197_, new_n23198_, new_n23199_, new_n23200_, new_n23201_,
    new_n23202_, new_n23203_, new_n23204_, new_n23205_, new_n23206_,
    new_n23207_, new_n23208_, new_n23209_, new_n23210_, new_n23211_,
    new_n23212_, new_n23213_, new_n23214_, new_n23215_, new_n23216_,
    new_n23217_, new_n23218_, new_n23219_, new_n23220_, new_n23221_,
    new_n23222_, new_n23223_, new_n23224_, new_n23225_, new_n23226_,
    new_n23227_, new_n23228_, new_n23229_, new_n23230_, new_n23231_,
    new_n23232_, new_n23233_, new_n23234_, new_n23235_, new_n23236_,
    new_n23237_, new_n23238_, new_n23239_, new_n23240_, new_n23241_,
    new_n23242_, new_n23243_, new_n23244_, new_n23245_, new_n23246_,
    new_n23247_, new_n23248_, new_n23249_, new_n23250_, new_n23251_,
    new_n23252_, new_n23253_, new_n23254_, new_n23255_, new_n23256_,
    new_n23257_, new_n23258_, new_n23259_, new_n23260_, new_n23261_,
    new_n23262_, new_n23263_, new_n23264_, new_n23265_, new_n23266_,
    new_n23267_, new_n23268_, new_n23269_, new_n23270_, new_n23271_,
    new_n23272_, new_n23273_, new_n23274_, new_n23275_, new_n23276_,
    new_n23277_, new_n23278_, new_n23279_, new_n23280_, new_n23281_,
    new_n23282_, new_n23283_, new_n23284_, new_n23285_, new_n23286_,
    new_n23287_, new_n23288_, new_n23289_, new_n23290_, new_n23291_,
    new_n23292_, new_n23293_, new_n23294_, new_n23295_, new_n23296_,
    new_n23297_, new_n23298_, new_n23299_, new_n23300_, new_n23301_,
    new_n23302_, new_n23303_, new_n23304_, new_n23305_, new_n23306_,
    new_n23307_, new_n23308_, new_n23309_, new_n23310_, new_n23311_,
    new_n23312_, new_n23313_, new_n23314_, new_n23315_, new_n23316_,
    new_n23317_, new_n23318_, new_n23319_, new_n23320_, new_n23321_,
    new_n23322_, new_n23323_, new_n23324_, new_n23325_, new_n23326_,
    new_n23327_, new_n23328_, new_n23329_, new_n23330_, new_n23331_,
    new_n23332_, new_n23333_, new_n23334_, new_n23335_, new_n23336_,
    new_n23337_, new_n23338_, new_n23339_, new_n23340_, new_n23341_,
    new_n23342_, new_n23343_, new_n23344_, new_n23345_, new_n23346_,
    new_n23347_, new_n23348_, new_n23349_, new_n23350_, new_n23351_,
    new_n23352_, new_n23353_, new_n23354_, new_n23355_, new_n23356_,
    new_n23357_, new_n23358_, new_n23359_, new_n23360_, new_n23361_,
    new_n23362_, new_n23363_, new_n23364_, new_n23365_, new_n23366_,
    new_n23367_, new_n23368_, new_n23369_, new_n23370_, new_n23371_,
    new_n23372_, new_n23373_, new_n23374_, new_n23375_, new_n23376_,
    new_n23377_, new_n23378_, new_n23379_, new_n23380_, new_n23381_,
    new_n23382_, new_n23383_, new_n23384_, new_n23385_, new_n23386_,
    new_n23387_, new_n23388_, new_n23389_, new_n23390_, new_n23391_,
    new_n23392_, new_n23393_, new_n23394_, new_n23395_, new_n23396_,
    new_n23397_, new_n23398_, new_n23399_, new_n23400_, new_n23401_,
    new_n23402_, new_n23403_, new_n23404_, new_n23405_, new_n23406_,
    new_n23407_, new_n23408_, new_n23409_, new_n23410_, new_n23411_,
    new_n23412_, new_n23413_, new_n23414_, new_n23415_, new_n23416_,
    new_n23417_, new_n23418_, new_n23419_, new_n23420_, new_n23421_,
    new_n23422_, new_n23423_, new_n23424_, new_n23425_, new_n23426_,
    new_n23427_, new_n23428_, new_n23429_, new_n23430_, new_n23431_,
    new_n23432_, new_n23433_, new_n23434_, new_n23435_, new_n23436_,
    new_n23437_, new_n23438_, new_n23439_, new_n23440_, new_n23441_,
    new_n23442_, new_n23443_, new_n23444_, new_n23445_, new_n23446_,
    new_n23447_, new_n23448_, new_n23449_, new_n23450_, new_n23451_,
    new_n23452_, new_n23453_, new_n23454_, new_n23455_, new_n23456_,
    new_n23457_, new_n23458_, new_n23459_, new_n23460_, new_n23461_,
    new_n23462_, new_n23463_, new_n23464_, new_n23465_, new_n23466_,
    new_n23467_, new_n23468_, new_n23469_, new_n23470_, new_n23471_,
    new_n23472_, new_n23473_, new_n23474_, new_n23475_, new_n23476_,
    new_n23477_, new_n23478_, new_n23479_, new_n23480_, new_n23481_,
    new_n23482_, new_n23483_, new_n23484_, new_n23485_, new_n23486_,
    new_n23487_, new_n23488_, new_n23489_, new_n23490_, new_n23491_,
    new_n23492_, new_n23493_, new_n23494_, new_n23495_, new_n23496_,
    new_n23497_, new_n23498_, new_n23499_, new_n23500_, new_n23501_,
    new_n23502_, new_n23503_, new_n23504_, new_n23505_, new_n23506_,
    new_n23507_, new_n23508_, new_n23509_, new_n23510_, new_n23511_,
    new_n23512_, new_n23513_, new_n23514_, new_n23515_, new_n23516_,
    new_n23517_, new_n23518_, new_n23519_, new_n23520_, new_n23521_,
    new_n23522_, new_n23523_, new_n23524_, new_n23525_, new_n23526_,
    new_n23527_, new_n23528_, new_n23529_, new_n23530_, new_n23531_,
    new_n23532_, new_n23533_, new_n23534_, new_n23535_, new_n23536_,
    new_n23537_, new_n23538_, new_n23539_, new_n23540_, new_n23541_,
    new_n23542_, new_n23543_, new_n23544_, new_n23545_, new_n23546_,
    new_n23547_, new_n23548_, new_n23549_, new_n23550_, new_n23551_,
    new_n23552_, new_n23553_, new_n23554_, new_n23555_, new_n23556_,
    new_n23557_, new_n23558_, new_n23559_, new_n23560_, new_n23561_,
    new_n23562_, new_n23563_, new_n23564_, new_n23565_, new_n23566_,
    new_n23567_, new_n23568_, new_n23569_, new_n23570_, new_n23571_,
    new_n23572_, new_n23573_, new_n23574_, new_n23575_, new_n23576_,
    new_n23577_, new_n23578_, new_n23579_, new_n23580_, new_n23581_,
    new_n23582_, new_n23583_, new_n23584_, new_n23585_, new_n23586_,
    new_n23587_, new_n23588_, new_n23589_, new_n23590_, new_n23591_,
    new_n23592_, new_n23593_, new_n23594_, new_n23595_, new_n23596_,
    new_n23597_, new_n23598_, new_n23599_, new_n23600_, new_n23601_,
    new_n23602_, new_n23603_, new_n23604_, new_n23605_, new_n23606_,
    new_n23607_, new_n23608_, new_n23609_, new_n23610_, new_n23611_,
    new_n23612_, new_n23613_, new_n23614_, new_n23615_, new_n23616_,
    new_n23617_, new_n23618_, new_n23619_, new_n23620_, new_n23621_,
    new_n23622_, new_n23623_, new_n23624_, new_n23625_, new_n23626_,
    new_n23627_, new_n23628_, new_n23629_, new_n23630_, new_n23631_,
    new_n23632_, new_n23633_, new_n23634_, new_n23635_, new_n23636_,
    new_n23637_, new_n23638_, new_n23639_, new_n23640_, new_n23641_,
    new_n23642_, new_n23643_, new_n23644_, new_n23645_, new_n23646_,
    new_n23647_, new_n23648_, new_n23649_, new_n23650_, new_n23651_,
    new_n23652_, new_n23653_, new_n23654_, new_n23655_, new_n23656_,
    new_n23657_, new_n23658_, new_n23659_, new_n23660_, new_n23661_,
    new_n23662_, new_n23663_, new_n23664_, new_n23665_, new_n23666_,
    new_n23667_, new_n23668_, new_n23669_, new_n23670_, new_n23671_,
    new_n23672_, new_n23673_, new_n23674_, new_n23675_, new_n23676_,
    new_n23677_, new_n23678_, new_n23679_, new_n23680_, new_n23681_,
    new_n23682_, new_n23683_, new_n23684_, new_n23685_, new_n23686_,
    new_n23687_, new_n23688_, new_n23689_, new_n23690_, new_n23691_,
    new_n23692_, new_n23693_, new_n23694_, new_n23695_, new_n23696_,
    new_n23697_, new_n23698_, new_n23699_, new_n23700_, new_n23701_,
    new_n23702_, new_n23703_, new_n23704_, new_n23705_, new_n23706_,
    new_n23707_, new_n23708_, new_n23709_, new_n23710_, new_n23711_,
    new_n23712_, new_n23713_, new_n23714_, new_n23715_, new_n23716_,
    new_n23717_, new_n23718_, new_n23719_, new_n23720_, new_n23721_,
    new_n23722_, new_n23723_, new_n23724_, new_n23725_, new_n23726_,
    new_n23727_, new_n23728_, new_n23729_, new_n23730_, new_n23731_,
    new_n23732_, new_n23733_, new_n23734_, new_n23735_, new_n23736_,
    new_n23737_, new_n23738_, new_n23739_, new_n23740_, new_n23741_,
    new_n23742_, new_n23743_, new_n23744_, new_n23745_, new_n23746_,
    new_n23747_, new_n23748_, new_n23749_, new_n23750_, new_n23751_,
    new_n23752_, new_n23753_, new_n23754_, new_n23755_, new_n23756_,
    new_n23757_, new_n23758_, new_n23759_, new_n23760_, new_n23761_,
    new_n23762_, new_n23763_, new_n23764_, new_n23765_, new_n23766_,
    new_n23767_, new_n23768_, new_n23769_, new_n23770_, new_n23771_,
    new_n23772_, new_n23773_, new_n23774_, new_n23775_, new_n23776_,
    new_n23777_, new_n23778_, new_n23779_, new_n23780_, new_n23781_,
    new_n23782_, new_n23783_, new_n23784_, new_n23785_, new_n23786_,
    new_n23787_, new_n23788_, new_n23789_, new_n23790_, new_n23791_,
    new_n23792_, new_n23793_, new_n23794_, new_n23795_, new_n23796_,
    new_n23797_, new_n23798_, new_n23799_, new_n23800_, new_n23801_,
    new_n23802_, new_n23803_, new_n23804_, new_n23805_, new_n23806_,
    new_n23807_, new_n23808_, new_n23809_, new_n23810_, new_n23811_,
    new_n23812_, new_n23813_, new_n23814_, new_n23815_, new_n23816_,
    new_n23817_, new_n23818_, new_n23819_, new_n23820_, new_n23821_,
    new_n23822_, new_n23823_, new_n23824_, new_n23825_, new_n23826_,
    new_n23827_, new_n23828_, new_n23829_, new_n23830_, new_n23831_,
    new_n23832_, new_n23833_, new_n23834_, new_n23835_, new_n23836_,
    new_n23837_, new_n23838_, new_n23839_, new_n23840_, new_n23841_,
    new_n23842_, new_n23843_, new_n23844_, new_n23845_, new_n23846_,
    new_n23847_, new_n23848_, new_n23849_, new_n23850_, new_n23851_,
    new_n23852_, new_n23853_, new_n23854_, new_n23855_, new_n23856_,
    new_n23857_, new_n23858_, new_n23859_, new_n23860_, new_n23861_,
    new_n23862_, new_n23863_, new_n23864_, new_n23865_, new_n23866_,
    new_n23867_, new_n23868_, new_n23869_, new_n23870_, new_n23871_,
    new_n23872_, new_n23873_, new_n23874_, new_n23875_, new_n23876_,
    new_n23877_, new_n23878_, new_n23879_, new_n23880_, new_n23881_,
    new_n23882_, new_n23883_, new_n23884_, new_n23885_, new_n23886_,
    new_n23887_, new_n23888_, new_n23889_, new_n23890_, new_n23891_,
    new_n23892_, new_n23893_, new_n23894_, new_n23895_, new_n23896_,
    new_n23897_, new_n23898_, new_n23899_, new_n23900_, new_n23901_,
    new_n23902_, new_n23903_, new_n23904_, new_n23905_, new_n23906_,
    new_n23907_, new_n23908_, new_n23909_, new_n23910_, new_n23911_,
    new_n23912_, new_n23913_, new_n23914_, new_n23915_, new_n23916_,
    new_n23917_, new_n23918_, new_n23919_, new_n23920_, new_n23921_,
    new_n23922_, new_n23923_, new_n23924_, new_n23925_, new_n23926_,
    new_n23927_, new_n23928_, new_n23929_, new_n23930_, new_n23931_,
    new_n23932_, new_n23933_, new_n23934_, new_n23935_, new_n23936_,
    new_n23937_, new_n23938_, new_n23939_, new_n23940_, new_n23941_,
    new_n23942_, new_n23943_, new_n23944_, new_n23945_, new_n23946_,
    new_n23947_, new_n23948_, new_n23949_, new_n23950_, new_n23951_,
    new_n23952_, new_n23953_, new_n23954_, new_n23955_, new_n23956_,
    new_n23957_, new_n23958_, new_n23959_, new_n23960_, new_n23961_,
    new_n23962_, new_n23963_, new_n23964_, new_n23965_, new_n23966_,
    new_n23967_, new_n23968_, new_n23969_, new_n23970_, new_n23971_,
    new_n23972_, new_n23973_, new_n23974_, new_n23975_, new_n23976_,
    new_n23977_, new_n23978_, new_n23979_, new_n23980_, new_n23981_,
    new_n23982_, new_n23983_, new_n23984_, new_n23985_, new_n23986_,
    new_n23987_, new_n23988_, new_n23989_, new_n23990_, new_n23991_,
    new_n23992_, new_n23993_, new_n23994_, new_n23995_, new_n23996_,
    new_n23997_, new_n23998_, new_n23999_, new_n24000_, new_n24001_,
    new_n24002_, new_n24003_, new_n24004_, new_n24005_, new_n24006_,
    new_n24007_, new_n24008_, new_n24009_, new_n24010_, new_n24011_,
    new_n24012_, new_n24013_, new_n24014_, new_n24015_, new_n24016_,
    new_n24017_, new_n24018_, new_n24019_, new_n24020_, new_n24021_,
    new_n24022_, new_n24023_, new_n24024_, new_n24025_, new_n24026_,
    new_n24027_, new_n24028_, new_n24029_, new_n24030_, new_n24031_,
    new_n24032_, new_n24033_, new_n24034_, new_n24035_, new_n24036_,
    new_n24037_, new_n24038_, new_n24039_, new_n24040_, new_n24041_,
    new_n24042_, new_n24043_, new_n24044_, new_n24045_, new_n24046_,
    new_n24047_, new_n24048_, new_n24049_, new_n24050_, new_n24051_,
    new_n24052_, new_n24053_, new_n24054_, new_n24055_, new_n24056_,
    new_n24057_, new_n24058_, new_n24059_, new_n24060_, new_n24061_,
    new_n24062_, new_n24063_, new_n24064_, new_n24065_, new_n24066_,
    new_n24067_, new_n24068_, new_n24069_, new_n24070_, new_n24071_,
    new_n24072_, new_n24073_, new_n24074_, new_n24075_, new_n24076_,
    new_n24077_, new_n24078_, new_n24079_, new_n24080_, new_n24081_,
    new_n24082_, new_n24083_, new_n24084_, new_n24085_, new_n24086_,
    new_n24087_, new_n24088_, new_n24089_, new_n24090_, new_n24091_,
    new_n24092_, new_n24093_, new_n24094_, new_n24095_, new_n24096_,
    new_n24097_, new_n24098_, new_n24099_, new_n24100_, new_n24101_,
    new_n24102_, new_n24103_, new_n24104_, new_n24105_, new_n24106_,
    new_n24107_, new_n24108_, new_n24109_, new_n24110_, new_n24111_,
    new_n24112_, new_n24113_, new_n24114_, new_n24115_, new_n24116_,
    new_n24117_, new_n24118_, new_n24119_, new_n24120_, new_n24121_,
    new_n24122_, new_n24123_, new_n24124_, new_n24125_, new_n24126_,
    new_n24127_, new_n24128_, new_n24129_, new_n24130_, new_n24131_,
    new_n24132_, new_n24133_, new_n24134_, new_n24135_, new_n24136_,
    new_n24137_, new_n24138_, new_n24139_, new_n24140_, new_n24141_,
    new_n24142_, new_n24143_, new_n24144_, new_n24145_, new_n24146_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24164_, new_n24165_, new_n24166_,
    new_n24167_, new_n24168_, new_n24169_, new_n24170_, new_n24171_,
    new_n24172_, new_n24173_, new_n24174_, new_n24175_, new_n24176_,
    new_n24177_, new_n24178_, new_n24179_, new_n24180_, new_n24181_,
    new_n24182_, new_n24183_, new_n24184_, new_n24185_, new_n24186_,
    new_n24187_, new_n24188_, new_n24189_, new_n24190_, new_n24191_,
    new_n24192_, new_n24193_, new_n24194_, new_n24195_, new_n24196_,
    new_n24197_, new_n24198_, new_n24199_, new_n24200_, new_n24201_,
    new_n24202_, new_n24203_, new_n24204_, new_n24205_, new_n24206_,
    new_n24207_, new_n24208_, new_n24209_, new_n24210_, new_n24211_,
    new_n24212_, new_n24213_, new_n24214_, new_n24215_, new_n24216_,
    new_n24217_, new_n24218_, new_n24219_, new_n24220_, new_n24221_,
    new_n24222_, new_n24223_, new_n24224_, new_n24225_, new_n24226_,
    new_n24227_, new_n24228_, new_n24229_, new_n24230_, new_n24231_,
    new_n24232_, new_n24233_, new_n24234_, new_n24235_, new_n24236_,
    new_n24237_, new_n24238_, new_n24239_, new_n24240_, new_n24241_,
    new_n24242_, new_n24243_, new_n24244_, new_n24245_, new_n24246_,
    new_n24247_, new_n24248_, new_n24249_, new_n24250_, new_n24251_,
    new_n24252_, new_n24253_, new_n24254_, new_n24255_, new_n24256_,
    new_n24257_, new_n24258_, new_n24259_, new_n24260_, new_n24261_,
    new_n24262_, new_n24263_, new_n24264_, new_n24265_, new_n24266_,
    new_n24267_, new_n24268_, new_n24269_, new_n24270_, new_n24271_,
    new_n24272_, new_n24273_, new_n24274_, new_n24275_, new_n24276_,
    new_n24277_, new_n24278_, new_n24279_, new_n24280_, new_n24281_,
    new_n24282_, new_n24283_, new_n24284_, new_n24285_, new_n24286_,
    new_n24287_, new_n24288_, new_n24289_, new_n24290_, new_n24291_,
    new_n24292_, new_n24293_, new_n24294_, new_n24295_, new_n24296_,
    new_n24297_, new_n24298_, new_n24299_, new_n24300_, new_n24301_,
    new_n24302_, new_n24303_, new_n24304_, new_n24305_, new_n24306_,
    new_n24307_, new_n24308_, new_n24309_, new_n24310_, new_n24311_,
    new_n24312_, new_n24313_, new_n24314_, new_n24315_, new_n24316_,
    new_n24317_, new_n24318_, new_n24319_, new_n24320_, new_n24321_,
    new_n24322_, new_n24323_, new_n24324_, new_n24325_, new_n24326_,
    new_n24327_, new_n24328_, new_n24329_, new_n24330_, new_n24331_,
    new_n24332_, new_n24333_, new_n24334_, new_n24335_, new_n24336_,
    new_n24337_, new_n24338_, new_n24339_, new_n24340_, new_n24341_,
    new_n24342_, new_n24343_, new_n24344_, new_n24345_, new_n24346_,
    new_n24347_, new_n24348_, new_n24349_, new_n24350_, new_n24351_,
    new_n24352_, new_n24353_, new_n24354_, new_n24355_, new_n24356_,
    new_n24357_, new_n24358_, new_n24359_, new_n24360_, new_n24361_,
    new_n24362_, new_n24363_, new_n24364_, new_n24365_, new_n24366_,
    new_n24367_, new_n24368_, new_n24369_, new_n24370_, new_n24371_,
    new_n24372_, new_n24373_, new_n24374_, new_n24375_, new_n24376_,
    new_n24377_, new_n24378_, new_n24379_, new_n24380_, new_n24381_,
    new_n24382_, new_n24383_, new_n24384_, new_n24385_, new_n24386_,
    new_n24387_, new_n24388_, new_n24389_, new_n24390_, new_n24391_,
    new_n24392_, new_n24393_, new_n24394_, new_n24395_, new_n24396_,
    new_n24397_, new_n24398_, new_n24399_, new_n24400_, new_n24401_,
    new_n24402_, new_n24403_, new_n24404_, new_n24405_, new_n24406_,
    new_n24407_, new_n24408_, new_n24409_, new_n24410_, new_n24411_,
    new_n24412_, new_n24413_, new_n24414_, new_n24415_, new_n24416_,
    new_n24417_, new_n24418_, new_n24419_, new_n24420_, new_n24421_,
    new_n24422_, new_n24423_, new_n24424_, new_n24425_, new_n24426_,
    new_n24427_, new_n24428_, new_n24429_, new_n24430_, new_n24431_,
    new_n24432_, new_n24433_, new_n24434_, new_n24435_, new_n24436_,
    new_n24437_, new_n24438_, new_n24439_, new_n24440_, new_n24441_,
    new_n24442_, new_n24443_, new_n24444_, new_n24445_, new_n24446_,
    new_n24447_, new_n24448_, new_n24449_, new_n24450_, new_n24451_,
    new_n24452_, new_n24453_, new_n24454_, new_n24455_, new_n24456_,
    new_n24457_, new_n24458_, new_n24459_, new_n24460_, new_n24461_,
    new_n24462_, new_n24463_, new_n24464_, new_n24465_, new_n24466_,
    new_n24467_, new_n24468_, new_n24469_, new_n24470_, new_n24471_,
    new_n24472_, new_n24473_, new_n24474_, new_n24475_, new_n24476_,
    new_n24477_, new_n24478_, new_n24479_, new_n24480_, new_n24481_,
    new_n24482_, new_n24483_, new_n24484_, new_n24485_, new_n24486_,
    new_n24487_, new_n24488_, new_n24489_, new_n24490_, new_n24491_,
    new_n24492_, new_n24493_, new_n24494_, new_n24495_, new_n24496_,
    new_n24497_, new_n24498_, new_n24499_, new_n24500_, new_n24501_,
    new_n24502_, new_n24503_, new_n24504_, new_n24505_, new_n24506_,
    new_n24507_, new_n24508_, new_n24509_, new_n24510_, new_n24511_,
    new_n24512_, new_n24513_, new_n24514_, new_n24515_, new_n24516_,
    new_n24517_, new_n24518_, new_n24519_, new_n24520_, new_n24521_,
    new_n24522_, new_n24523_, new_n24524_, new_n24525_, new_n24526_,
    new_n24527_, new_n24528_, new_n24529_, new_n24530_, new_n24531_,
    new_n24532_, new_n24533_, new_n24534_, new_n24535_, new_n24536_,
    new_n24537_, new_n24538_, new_n24539_, new_n24540_, new_n24541_,
    new_n24542_, new_n24543_, new_n24544_, new_n24545_, new_n24546_,
    new_n24547_, new_n24548_, new_n24549_, new_n24550_, new_n24551_,
    new_n24552_, new_n24553_, new_n24554_, new_n24555_, new_n24556_,
    new_n24557_, new_n24558_, new_n24559_, new_n24560_, new_n24561_,
    new_n24562_, new_n24563_, new_n24564_, new_n24565_, new_n24566_,
    new_n24567_, new_n24568_, new_n24569_, new_n24570_, new_n24571_,
    new_n24572_, new_n24573_, new_n24574_, new_n24575_, new_n24576_,
    new_n24577_, new_n24578_, new_n24579_, new_n24580_, new_n24581_,
    new_n24582_, new_n24583_, new_n24584_, new_n24585_, new_n24586_,
    new_n24587_, new_n24588_, new_n24589_, new_n24590_, new_n24591_,
    new_n24592_, new_n24593_, new_n24594_, new_n24595_, new_n24596_,
    new_n24597_, new_n24598_, new_n24599_, new_n24600_, new_n24601_,
    new_n24602_, new_n24603_, new_n24604_, new_n24605_, new_n24606_,
    new_n24607_, new_n24608_, new_n24609_, new_n24610_, new_n24611_,
    new_n24612_, new_n24613_, new_n24614_, new_n24615_, new_n24616_,
    new_n24617_, new_n24618_, new_n24619_, new_n24620_, new_n24621_,
    new_n24622_, new_n24623_, new_n24624_, new_n24625_, new_n24626_,
    new_n24627_, new_n24628_, new_n24629_, new_n24630_, new_n24631_,
    new_n24632_, new_n24633_, new_n24634_, new_n24635_, new_n24636_,
    new_n24637_, new_n24638_, new_n24639_, new_n24640_, new_n24641_,
    new_n24642_, new_n24643_, new_n24644_, new_n24645_, new_n24646_,
    new_n24647_, new_n24648_, new_n24649_, new_n24650_, new_n24651_,
    new_n24652_, new_n24653_, new_n24654_, new_n24655_, new_n24656_,
    new_n24657_, new_n24658_, new_n24659_, new_n24660_, new_n24661_,
    new_n24662_, new_n24663_, new_n24664_, new_n24665_, new_n24666_,
    new_n24667_, new_n24668_, new_n24669_, new_n24670_, new_n24671_,
    new_n24672_, new_n24673_, new_n24674_, new_n24675_, new_n24676_,
    new_n24677_, new_n24678_, new_n24679_, new_n24680_, new_n24681_,
    new_n24682_, new_n24683_, new_n24684_, new_n24685_, new_n24686_,
    new_n24687_, new_n24688_, new_n24689_, new_n24690_, new_n24691_,
    new_n24692_, new_n24693_, new_n24694_, new_n24695_, new_n24696_,
    new_n24697_, new_n24698_, new_n24699_, new_n24700_, new_n24701_,
    new_n24702_, new_n24703_, new_n24704_, new_n24705_, new_n24706_,
    new_n24707_, new_n24708_, new_n24709_, new_n24710_, new_n24711_,
    new_n24712_, new_n24713_, new_n24714_, new_n24715_, new_n24716_,
    new_n24717_, new_n24718_, new_n24719_, new_n24720_, new_n24721_,
    new_n24722_, new_n24723_, new_n24724_, new_n24725_, new_n24726_,
    new_n24727_, new_n24728_, new_n24729_, new_n24730_, new_n24731_,
    new_n24732_, new_n24733_, new_n24734_, new_n24735_, new_n24736_,
    new_n24737_, new_n24738_, new_n24739_, new_n24740_, new_n24741_,
    new_n24742_, new_n24743_, new_n24744_, new_n24745_, new_n24746_,
    new_n24747_, new_n24748_, new_n24749_, new_n24750_, new_n24751_,
    new_n24752_, new_n24753_, new_n24754_, new_n24755_, new_n24756_,
    new_n24757_, new_n24758_, new_n24759_, new_n24760_, new_n24761_,
    new_n24762_, new_n24763_, new_n24764_, new_n24765_, new_n24766_,
    new_n24767_, new_n24768_, new_n24769_, new_n24770_, new_n24771_,
    new_n24772_, new_n24773_, new_n24774_, new_n24775_, new_n24776_,
    new_n24777_, new_n24778_, new_n24779_, new_n24780_, new_n24781_,
    new_n24782_, new_n24783_, new_n24784_, new_n24785_, new_n24786_,
    new_n24787_, new_n24788_, new_n24789_, new_n24790_, new_n24791_,
    new_n24792_, new_n24793_, new_n24794_, new_n24795_, new_n24796_,
    new_n24797_, new_n24798_, new_n24799_, new_n24800_, new_n24801_,
    new_n24802_, new_n24803_, new_n24804_, new_n24805_, new_n24806_,
    new_n24807_, new_n24808_, new_n24809_, new_n24810_, new_n24811_,
    new_n24812_, new_n24813_, new_n24814_, new_n24815_, new_n24816_,
    new_n24817_, new_n24818_, new_n24819_, new_n24820_, new_n24821_,
    new_n24822_, new_n24823_, new_n24824_, new_n24825_, new_n24826_,
    new_n24827_, new_n24828_, new_n24829_, new_n24830_, new_n24831_,
    new_n24832_, new_n24833_, new_n24834_, new_n24835_, new_n24836_,
    new_n24837_, new_n24838_, new_n24839_, new_n24840_, new_n24841_,
    new_n24842_, new_n24843_, new_n24844_, new_n24845_, new_n24846_,
    new_n24847_, new_n24848_, new_n24849_, new_n24850_, new_n24851_,
    new_n24852_, new_n24853_, new_n24854_, new_n24855_, new_n24856_,
    new_n24857_, new_n24858_, new_n24859_, new_n24860_, new_n24861_,
    new_n24862_, new_n24863_, new_n24864_, new_n24865_, new_n24866_,
    new_n24867_, new_n24868_, new_n24869_, new_n24870_, new_n24871_,
    new_n24872_, new_n24873_, new_n24874_, new_n24875_, new_n24876_,
    new_n24877_, new_n24878_, new_n24879_, new_n24880_, new_n24881_,
    new_n24882_, new_n24883_, new_n24884_, new_n24885_, new_n24886_,
    new_n24887_, new_n24888_, new_n24889_, new_n24890_, new_n24891_,
    new_n24892_, new_n24893_, new_n24894_, new_n24895_, new_n24896_,
    new_n24897_, new_n24898_, new_n24899_, new_n24900_, new_n24901_,
    new_n24902_, new_n24903_, new_n24904_, new_n24905_, new_n24906_,
    new_n24907_, new_n24908_, new_n24909_, new_n24910_, new_n24911_,
    new_n24912_, new_n24913_, new_n24914_, new_n24915_, new_n24916_,
    new_n24917_, new_n24918_, new_n24919_, new_n24920_, new_n24921_,
    new_n24922_, new_n24923_, new_n24924_, new_n24925_, new_n24926_,
    new_n24927_, new_n24928_, new_n24929_, new_n24930_, new_n24931_,
    new_n24932_, new_n24933_, new_n24934_, new_n24935_, new_n24936_,
    new_n24937_, new_n24938_, new_n24939_, new_n24940_, new_n24941_,
    new_n24942_, new_n24943_, new_n24944_, new_n24945_, new_n24946_,
    new_n24947_, new_n24948_, new_n24949_, new_n24950_, new_n24951_,
    new_n24952_, new_n24953_, new_n24954_, new_n24955_, new_n24956_,
    new_n24957_, new_n24958_, new_n24959_, new_n24960_, new_n24961_,
    new_n24962_, new_n24963_, new_n24964_, new_n24965_, new_n24966_,
    new_n24967_, new_n24968_, new_n24969_, new_n24970_, new_n24971_,
    new_n24972_, new_n24973_, new_n24974_, new_n24975_, new_n24976_,
    new_n24977_, new_n24978_, new_n24979_, new_n24980_, new_n24981_,
    new_n24982_, new_n24983_, new_n24984_, new_n24985_, new_n24986_,
    new_n24987_, new_n24988_, new_n24989_, new_n24990_, new_n24991_,
    new_n24992_, new_n24993_, new_n24994_, new_n24995_, new_n24996_,
    new_n24997_, new_n24998_, new_n24999_, new_n25000_, new_n25001_,
    new_n25002_, new_n25003_, new_n25004_, new_n25005_, new_n25006_,
    new_n25007_, new_n25008_, new_n25009_, new_n25010_, new_n25011_,
    new_n25012_, new_n25013_, new_n25014_, new_n25015_, new_n25016_,
    new_n25017_, new_n25018_, new_n25019_, new_n25020_, new_n25021_,
    new_n25022_, new_n25023_, new_n25024_, new_n25025_, new_n25026_,
    new_n25027_, new_n25028_, new_n25029_, new_n25030_, new_n25031_,
    new_n25032_, new_n25033_, new_n25034_, new_n25035_, new_n25036_,
    new_n25037_, new_n25038_, new_n25039_, new_n25040_, new_n25041_,
    new_n25042_, new_n25043_, new_n25044_, new_n25045_, new_n25046_,
    new_n25047_, new_n25048_, new_n25049_, new_n25050_, new_n25051_,
    new_n25052_, new_n25053_, new_n25054_, new_n25055_, new_n25056_,
    new_n25057_, new_n25058_, new_n25059_, new_n25060_, new_n25061_,
    new_n25062_, new_n25063_, new_n25064_, new_n25065_, new_n25066_,
    new_n25067_, new_n25068_, new_n25069_, new_n25070_, new_n25071_,
    new_n25072_, new_n25073_, new_n25074_, new_n25075_, new_n25076_,
    new_n25077_, new_n25078_, new_n25079_, new_n25080_, new_n25081_,
    new_n25082_, new_n25083_, new_n25084_, new_n25085_, new_n25086_,
    new_n25087_, new_n25088_, new_n25089_, new_n25090_, new_n25091_,
    new_n25092_, new_n25093_, new_n25094_, new_n25095_, new_n25096_,
    new_n25097_, new_n25098_, new_n25099_, new_n25100_, new_n25101_,
    new_n25102_, new_n25103_, new_n25104_, new_n25105_, new_n25106_,
    new_n25107_, new_n25108_, new_n25109_, new_n25110_, new_n25111_,
    new_n25112_, new_n25113_, new_n25114_, new_n25115_, new_n25116_,
    new_n25117_, new_n25118_, new_n25119_, new_n25120_, new_n25121_,
    new_n25122_, new_n25123_, new_n25124_, new_n25125_, new_n25126_,
    new_n25127_, new_n25128_, new_n25129_, new_n25130_, new_n25131_,
    new_n25132_, new_n25133_, new_n25134_, new_n25135_, new_n25136_,
    new_n25137_, new_n25138_, new_n25139_, new_n25140_, new_n25141_,
    new_n25142_, new_n25143_, new_n25144_, new_n25145_, new_n25146_,
    new_n25147_, new_n25148_, new_n25149_, new_n25150_, new_n25151_,
    new_n25152_, new_n25153_, new_n25154_, new_n25155_, new_n25156_,
    new_n25157_, new_n25158_, new_n25159_, new_n25160_, new_n25161_,
    new_n25162_, new_n25163_, new_n25164_, new_n25165_, new_n25166_,
    new_n25167_, new_n25168_, new_n25169_, new_n25170_, new_n25171_,
    new_n25172_, new_n25173_, new_n25174_, new_n25175_, new_n25176_,
    new_n25177_, new_n25178_, new_n25179_, new_n25180_, new_n25181_,
    new_n25182_, new_n25183_, new_n25184_, new_n25185_, new_n25186_,
    new_n25187_, new_n25188_, new_n25189_, new_n25190_, new_n25191_,
    new_n25192_, new_n25193_, new_n25194_, new_n25195_, new_n25196_,
    new_n25197_, new_n25198_, new_n25199_, new_n25200_, new_n25201_,
    new_n25202_, new_n25203_, new_n25204_, new_n25205_, new_n25206_,
    new_n25207_, new_n25208_, new_n25209_, new_n25210_, new_n25211_,
    new_n25212_, new_n25213_, new_n25214_, new_n25215_, new_n25216_,
    new_n25217_, new_n25218_, new_n25219_, new_n25220_, new_n25221_,
    new_n25222_, new_n25223_, new_n25224_, new_n25225_, new_n25226_,
    new_n25227_, new_n25228_, new_n25229_, new_n25230_, new_n25231_,
    new_n25232_, new_n25233_, new_n25234_, new_n25235_, new_n25236_,
    new_n25237_, new_n25238_, new_n25239_, new_n25240_, new_n25241_,
    new_n25242_, new_n25243_, new_n25244_, new_n25245_, new_n25246_,
    new_n25247_, new_n25248_, new_n25249_, new_n25250_, new_n25251_,
    new_n25252_, new_n25253_, new_n25254_, new_n25255_, new_n25256_,
    new_n25257_, new_n25258_, new_n25259_, new_n25260_, new_n25261_,
    new_n25262_, new_n25263_, new_n25264_, new_n25265_, new_n25266_,
    new_n25267_, new_n25268_, new_n25269_, new_n25270_, new_n25271_,
    new_n25272_, new_n25273_, new_n25274_, new_n25275_, new_n25276_,
    new_n25277_, new_n25278_, new_n25279_, new_n25280_, new_n25281_,
    new_n25282_, new_n25283_, new_n25284_, new_n25285_, new_n25286_,
    new_n25287_, new_n25288_, new_n25289_, new_n25290_, new_n25291_,
    new_n25292_, new_n25293_, new_n25294_, new_n25295_, new_n25296_,
    new_n25297_, new_n25298_, new_n25299_, new_n25300_, new_n25301_,
    new_n25302_, new_n25303_, new_n25304_, new_n25305_, new_n25306_,
    new_n25307_, new_n25308_, new_n25309_, new_n25310_, new_n25311_,
    new_n25312_, new_n25313_, new_n25314_, new_n25315_, new_n25316_,
    new_n25317_, new_n25318_, new_n25319_, new_n25320_, new_n25321_,
    new_n25322_, new_n25323_, new_n25324_, new_n25325_, new_n25326_,
    new_n25327_, new_n25328_, new_n25329_, new_n25330_, new_n25331_,
    new_n25332_, new_n25333_, new_n25334_, new_n25335_, new_n25336_,
    new_n25337_, new_n25338_, new_n25339_, new_n25340_, new_n25341_,
    new_n25342_, new_n25343_, new_n25344_, new_n25345_, new_n25346_,
    new_n25347_, new_n25348_, new_n25349_, new_n25350_, new_n25351_,
    new_n25352_, new_n25353_, new_n25354_, new_n25355_, new_n25356_,
    new_n25357_, new_n25358_, new_n25359_, new_n25360_, new_n25361_,
    new_n25362_, new_n25363_, new_n25364_, new_n25365_, new_n25366_,
    new_n25367_, new_n25368_, new_n25369_, new_n25370_, new_n25371_,
    new_n25372_, new_n25373_, new_n25374_, new_n25375_, new_n25376_,
    new_n25377_, new_n25378_, new_n25379_, new_n25380_, new_n25381_,
    new_n25382_, new_n25383_, new_n25384_, new_n25385_, new_n25386_,
    new_n25387_, new_n25388_, new_n25389_, new_n25390_, new_n25391_,
    new_n25392_, new_n25393_, new_n25394_, new_n25395_, new_n25396_,
    new_n25397_, new_n25398_, new_n25399_, new_n25400_, new_n25401_,
    new_n25402_, new_n25403_, new_n25404_, new_n25405_, new_n25406_,
    new_n25407_, new_n25408_, new_n25409_, new_n25410_, new_n25411_,
    new_n25412_, new_n25413_, new_n25414_, new_n25415_, new_n25416_,
    new_n25417_, new_n25418_, new_n25419_, new_n25420_, new_n25421_,
    new_n25422_, new_n25423_, new_n25424_, new_n25425_, new_n25426_,
    new_n25427_, new_n25428_, new_n25429_, new_n25430_, new_n25431_,
    new_n25432_, new_n25433_, new_n25434_, new_n25435_, new_n25436_,
    new_n25437_, new_n25438_, new_n25439_, new_n25440_, new_n25441_,
    new_n25442_, new_n25443_, new_n25444_, new_n25445_, new_n25446_,
    new_n25447_, new_n25448_, new_n25449_, new_n25450_, new_n25451_,
    new_n25452_, new_n25453_, new_n25454_, new_n25455_, new_n25456_,
    new_n25457_, new_n25458_, new_n25459_, new_n25460_, new_n25461_,
    new_n25462_, new_n25463_, new_n25464_, new_n25465_, new_n25466_,
    new_n25467_, new_n25468_, new_n25469_, new_n25470_, new_n25471_,
    new_n25472_, new_n25473_, new_n25474_, new_n25475_, new_n25476_,
    new_n25477_, new_n25478_, new_n25479_, new_n25480_, new_n25481_,
    new_n25482_, new_n25483_, new_n25484_, new_n25485_, new_n25486_,
    new_n25487_, new_n25488_, new_n25489_, new_n25490_, new_n25491_,
    new_n25492_, new_n25493_, new_n25494_, new_n25495_, new_n25496_,
    new_n25497_, new_n25498_, new_n25499_, new_n25500_, new_n25501_,
    new_n25502_, new_n25503_, new_n25504_, new_n25505_, new_n25506_,
    new_n25507_, new_n25508_, new_n25509_, new_n25510_, new_n25511_,
    new_n25512_, new_n25513_, new_n25514_, new_n25515_, new_n25516_,
    new_n25517_, new_n25518_, new_n25519_, new_n25520_, new_n25521_,
    new_n25522_, new_n25523_, new_n25524_, new_n25525_, new_n25526_,
    new_n25527_, new_n25528_, new_n25529_, new_n25530_, new_n25531_,
    new_n25532_, new_n25533_, new_n25534_, new_n25535_, new_n25536_,
    new_n25537_, new_n25538_, new_n25539_, new_n25540_, new_n25541_,
    new_n25542_, new_n25543_, new_n25544_, new_n25545_, new_n25546_,
    new_n25547_, new_n25548_, new_n25549_, new_n25550_, new_n25551_,
    new_n25552_, new_n25553_, new_n25554_, new_n25555_, new_n25556_,
    new_n25557_, new_n25558_, new_n25559_, new_n25560_, new_n25561_,
    new_n25562_, new_n25563_, new_n25564_, new_n25565_, new_n25566_,
    new_n25567_, new_n25568_, new_n25569_, new_n25570_, new_n25571_,
    new_n25572_, new_n25573_, new_n25574_, new_n25575_, new_n25576_,
    new_n25577_, new_n25578_, new_n25579_, new_n25580_, new_n25581_,
    new_n25582_, new_n25583_, new_n25584_, new_n25585_, new_n25586_,
    new_n25587_, new_n25588_, new_n25589_, new_n25590_, new_n25591_,
    new_n25592_, new_n25593_, new_n25594_, new_n25595_, new_n25596_,
    new_n25597_, new_n25598_, new_n25599_, new_n25600_, new_n25601_,
    new_n25602_, new_n25603_, new_n25604_, new_n25605_, new_n25606_,
    new_n25607_, new_n25608_, new_n25609_, new_n25610_, new_n25611_,
    new_n25612_, new_n25613_, new_n25614_, new_n25615_, new_n25616_,
    new_n25617_, new_n25618_, new_n25619_, new_n25620_, new_n25621_,
    new_n25622_, new_n25623_, new_n25624_, new_n25625_, new_n25626_,
    new_n25627_, new_n25628_, new_n25629_, new_n25630_, new_n25631_,
    new_n25632_, new_n25633_, new_n25634_, new_n25635_, new_n25636_,
    new_n25637_, new_n25638_, new_n25639_, new_n25640_, new_n25641_,
    new_n25642_, new_n25643_, new_n25644_, new_n25645_, new_n25646_,
    new_n25647_, new_n25648_, new_n25649_, new_n25650_, new_n25651_,
    new_n25652_, new_n25653_, new_n25654_, new_n25655_, new_n25656_,
    new_n25657_, new_n25658_, new_n25659_, new_n25660_, new_n25661_,
    new_n25662_, new_n25663_, new_n25664_, new_n25665_, new_n25666_,
    new_n25667_, new_n25668_, new_n25669_, new_n25670_, new_n25671_,
    new_n25672_, new_n25673_, new_n25674_, new_n25675_, new_n25676_,
    new_n25677_, new_n25678_, new_n25679_, new_n25680_, new_n25681_,
    new_n25682_, new_n25683_, new_n25684_, new_n25685_, new_n25686_,
    new_n25687_, new_n25688_, new_n25689_, new_n25690_, new_n25691_,
    new_n25692_, new_n25693_, new_n25694_, new_n25695_, new_n25696_,
    new_n25697_, new_n25698_, new_n25699_, new_n25700_, new_n25701_,
    new_n25702_, new_n25703_, new_n25704_, new_n25705_, new_n25706_,
    new_n25707_, new_n25708_, new_n25709_, new_n25710_, new_n25711_,
    new_n25712_, new_n25713_, new_n25714_, new_n25715_, new_n25716_,
    new_n25717_, new_n25718_, new_n25719_, new_n25720_, new_n25721_,
    new_n25722_, new_n25723_, new_n25724_, new_n25725_, new_n25726_,
    new_n25727_, new_n25728_, new_n25729_, new_n25730_, new_n25731_,
    new_n25732_, new_n25733_, new_n25734_, new_n25735_, new_n25736_,
    new_n25737_, new_n25738_, new_n25739_, new_n25740_, new_n25741_,
    new_n25742_, new_n25743_, new_n25744_, new_n25745_, new_n25746_,
    new_n25747_, new_n25748_, new_n25749_, new_n25750_, new_n25751_,
    new_n25752_, new_n25753_, new_n25754_, new_n25755_, new_n25756_,
    new_n25757_, new_n25758_, new_n25759_, new_n25760_, new_n25761_,
    new_n25762_, new_n25763_, new_n25764_, new_n25765_, new_n25766_,
    new_n25767_, new_n25768_, new_n25769_, new_n25770_, new_n25771_,
    new_n25772_, new_n25773_, new_n25774_, new_n25775_, new_n25776_,
    new_n25777_, new_n25778_, new_n25779_, new_n25780_, new_n25781_,
    new_n25782_, new_n25783_, new_n25784_, new_n25785_, new_n25786_,
    new_n25787_, new_n25788_, new_n25789_, new_n25790_, new_n25791_,
    new_n25792_, new_n25793_, new_n25794_, new_n25795_, new_n25796_,
    new_n25797_, new_n25798_, new_n25799_, new_n25800_, new_n25801_,
    new_n25802_, new_n25803_, new_n25804_, new_n25805_, new_n25806_,
    new_n25807_, new_n25808_, new_n25809_, new_n25810_, new_n25811_,
    new_n25812_, new_n25813_, new_n25814_, new_n25815_, new_n25816_,
    new_n25817_, new_n25818_, new_n25819_, new_n25820_, new_n25821_,
    new_n25822_, new_n25823_, new_n25824_, new_n25825_, new_n25826_,
    new_n25827_, new_n25828_, new_n25829_, new_n25830_, new_n25831_,
    new_n25832_, new_n25833_, new_n25834_, new_n25835_, new_n25836_,
    new_n25837_, new_n25838_, new_n25839_, new_n25840_, new_n25841_,
    new_n25842_, new_n25843_, new_n25844_, new_n25845_, new_n25846_,
    new_n25847_, new_n25848_, new_n25849_, new_n25850_, new_n25851_,
    new_n25852_, new_n25853_, new_n25854_, new_n25855_, new_n25856_,
    new_n25857_, new_n25858_, new_n25859_, new_n25860_, new_n25861_,
    new_n25862_, new_n25863_, new_n25864_, new_n25865_, new_n25866_,
    new_n25867_, new_n25868_, new_n25869_, new_n25870_, new_n25871_,
    new_n25872_, new_n25873_, new_n25874_, new_n25875_, new_n25876_,
    new_n25877_, new_n25878_, new_n25879_, new_n25880_, new_n25881_,
    new_n25882_, new_n25883_, new_n25884_, new_n25885_, new_n25886_,
    new_n25887_, new_n25888_, new_n25889_, new_n25890_, new_n25891_,
    new_n25892_, new_n25893_, new_n25894_, new_n25895_, new_n25896_,
    new_n25897_, new_n25898_, new_n25899_, new_n25900_, new_n25901_,
    new_n25902_, new_n25903_, new_n25904_, new_n25905_, new_n25906_,
    new_n25907_, new_n25908_, new_n25909_, new_n25910_, new_n25911_,
    new_n25912_, new_n25913_, new_n25914_, new_n25915_, new_n25916_,
    new_n25917_, new_n25918_, new_n25919_, new_n25920_, new_n25921_,
    new_n25922_, new_n25923_, new_n25924_, new_n25925_, new_n25926_,
    new_n25927_, new_n25928_, new_n25929_, new_n25930_, new_n25931_,
    new_n25932_, new_n25933_, new_n25934_, new_n25935_, new_n25936_,
    new_n25937_, new_n25938_, new_n25939_, new_n25940_, new_n25941_,
    new_n25942_, new_n25943_, new_n25944_, new_n25945_, new_n25946_,
    new_n25947_, new_n25948_, new_n25949_, new_n25950_, new_n25951_,
    new_n25952_, new_n25953_, new_n25954_, new_n25955_, new_n25956_,
    new_n25957_, new_n25958_, new_n25959_, new_n25960_, new_n25961_,
    new_n25962_, new_n25963_, new_n25964_, new_n25965_, new_n25966_,
    new_n25967_, new_n25968_, new_n25969_, new_n25970_, new_n25971_,
    new_n25972_, new_n25973_, new_n25974_, new_n25975_, new_n25976_,
    new_n25977_, new_n25978_, new_n25979_, new_n25980_, new_n25981_,
    new_n25982_, new_n25983_, new_n25984_, new_n25985_, new_n25986_,
    new_n25987_, new_n25988_, new_n25989_, new_n25990_, new_n25991_,
    new_n25992_, new_n25993_, new_n25994_, new_n25995_, new_n25996_,
    new_n25997_, new_n25998_, new_n25999_, new_n26000_, new_n26001_,
    new_n26002_, new_n26003_, new_n26004_, new_n26005_, new_n26006_,
    new_n26007_, new_n26008_, new_n26009_, new_n26010_, new_n26011_,
    new_n26012_, new_n26013_, new_n26014_, new_n26015_, new_n26016_,
    new_n26017_, new_n26018_, new_n26019_, new_n26020_, new_n26021_,
    new_n26022_, new_n26023_, new_n26024_, new_n26025_, new_n26026_,
    new_n26027_, new_n26028_, new_n26029_, new_n26030_, new_n26031_,
    new_n26032_, new_n26033_, new_n26034_, new_n26035_, new_n26036_,
    new_n26037_, new_n26038_, new_n26039_, new_n26040_, new_n26041_,
    new_n26042_, new_n26043_, new_n26044_, new_n26045_, new_n26046_,
    new_n26047_, new_n26048_, new_n26049_, new_n26050_, new_n26051_,
    new_n26052_, new_n26053_, new_n26054_, new_n26055_, new_n26056_,
    new_n26057_, new_n26058_, new_n26059_, new_n26060_, new_n26061_,
    new_n26062_, new_n26063_, new_n26064_, new_n26065_, new_n26066_,
    new_n26067_, new_n26068_, new_n26069_, new_n26070_, new_n26071_,
    new_n26072_, new_n26073_, new_n26074_, new_n26075_, new_n26076_,
    new_n26077_, new_n26078_, new_n26079_, new_n26080_, new_n26081_,
    new_n26082_, new_n26083_, new_n26084_, new_n26085_, new_n26086_,
    new_n26087_, new_n26088_, new_n26089_, new_n26090_, new_n26091_,
    new_n26092_, new_n26093_, new_n26094_, new_n26095_, new_n26096_,
    new_n26097_, new_n26098_, new_n26099_, new_n26100_, new_n26101_,
    new_n26102_, new_n26103_, new_n26104_, new_n26105_, new_n26106_,
    new_n26107_, new_n26108_, new_n26109_, new_n26110_, new_n26111_,
    new_n26112_, new_n26113_, new_n26114_, new_n26115_, new_n26116_,
    new_n26117_, new_n26118_, new_n26119_, new_n26120_, new_n26121_,
    new_n26122_, new_n26123_, new_n26124_, new_n26125_, new_n26126_,
    new_n26127_, new_n26128_, new_n26129_, new_n26130_, new_n26131_,
    new_n26132_, new_n26133_, new_n26134_, new_n26135_, new_n26136_,
    new_n26137_, new_n26138_, new_n26139_, new_n26140_, new_n26141_,
    new_n26142_, new_n26143_, new_n26144_, new_n26145_, new_n26146_,
    new_n26147_, new_n26148_, new_n26149_, new_n26150_, new_n26151_,
    new_n26152_, new_n26153_, new_n26154_, new_n26155_, new_n26156_,
    new_n26157_, new_n26158_, new_n26159_, new_n26160_, new_n26161_,
    new_n26162_, new_n26163_, new_n26164_, new_n26165_, new_n26166_,
    new_n26167_, new_n26168_, new_n26169_, new_n26170_, new_n26171_,
    new_n26172_, new_n26173_, new_n26174_, new_n26175_, new_n26176_,
    new_n26177_, new_n26178_, new_n26179_, new_n26180_, new_n26181_,
    new_n26182_, new_n26183_, new_n26184_, new_n26185_, new_n26186_,
    new_n26187_, new_n26188_, new_n26189_, new_n26190_, new_n26191_,
    new_n26192_, new_n26193_, new_n26194_, new_n26195_, new_n26196_,
    new_n26197_, new_n26198_, new_n26199_, new_n26200_, new_n26201_,
    new_n26202_, new_n26203_, new_n26204_, new_n26205_, new_n26206_,
    new_n26207_, new_n26208_, new_n26209_, new_n26210_, new_n26211_,
    new_n26212_, new_n26213_, new_n26214_, new_n26215_, new_n26216_,
    new_n26217_, new_n26218_, new_n26219_, new_n26220_, new_n26221_,
    new_n26222_, new_n26223_, new_n26224_, new_n26225_, new_n26226_,
    new_n26227_, new_n26228_, new_n26229_, new_n26230_, new_n26231_,
    new_n26232_, new_n26233_, new_n26234_, new_n26235_, new_n26236_,
    new_n26237_, new_n26238_, new_n26239_, new_n26240_, new_n26241_,
    new_n26242_, new_n26243_, new_n26244_, new_n26245_, new_n26246_,
    new_n26247_, new_n26248_, new_n26249_, new_n26250_, new_n26251_,
    new_n26252_, new_n26253_, new_n26254_, new_n26255_, new_n26256_,
    new_n26257_, new_n26258_, new_n26259_, new_n26260_, new_n26261_,
    new_n26262_, new_n26263_, new_n26264_, new_n26265_, new_n26266_,
    new_n26267_, new_n26268_, new_n26269_, new_n26270_, new_n26271_,
    new_n26272_, new_n26273_, new_n26274_, new_n26275_, new_n26276_,
    new_n26277_, new_n26278_, new_n26279_, new_n26280_, new_n26281_,
    new_n26282_, new_n26283_, new_n26284_, new_n26285_, new_n26286_,
    new_n26287_, new_n26288_, new_n26289_, new_n26290_, new_n26291_,
    new_n26292_, new_n26293_, new_n26294_, new_n26295_, new_n26296_,
    new_n26297_, new_n26298_, new_n26299_, new_n26300_, new_n26301_,
    new_n26302_, new_n26303_, new_n26304_, new_n26305_, new_n26306_,
    new_n26307_, new_n26308_, new_n26309_, new_n26310_, new_n26311_,
    new_n26312_, new_n26313_, new_n26314_, new_n26315_, new_n26316_,
    new_n26317_, new_n26318_, new_n26319_, new_n26320_, new_n26321_,
    new_n26322_, new_n26323_, new_n26324_, new_n26325_, new_n26326_,
    new_n26327_, new_n26328_, new_n26329_, new_n26330_, new_n26331_,
    new_n26332_, new_n26333_, new_n26334_, new_n26335_, new_n26336_,
    new_n26337_, new_n26338_, new_n26339_, new_n26340_, new_n26341_,
    new_n26342_, new_n26343_, new_n26344_, new_n26345_, new_n26346_,
    new_n26347_, new_n26348_, new_n26349_, new_n26350_, new_n26351_,
    new_n26352_, new_n26353_, new_n26354_, new_n26355_, new_n26356_,
    new_n26357_, new_n26358_, new_n26359_, new_n26360_, new_n26361_,
    new_n26362_, new_n26363_, new_n26364_, new_n26365_, new_n26366_,
    new_n26367_, new_n26368_, new_n26369_, new_n26370_, new_n26371_,
    new_n26372_, new_n26373_, new_n26374_, new_n26375_, new_n26376_,
    new_n26377_, new_n26378_, new_n26379_, new_n26380_, new_n26381_,
    new_n26382_, new_n26383_, new_n26384_, new_n26385_, new_n26386_,
    new_n26387_, new_n26388_, new_n26389_, new_n26390_, new_n26391_,
    new_n26392_, new_n26393_, new_n26394_, new_n26395_, new_n26396_,
    new_n26397_, new_n26398_, new_n26399_, new_n26400_, new_n26401_,
    new_n26402_, new_n26403_, new_n26404_, new_n26405_, new_n26406_,
    new_n26407_, new_n26408_, new_n26409_, new_n26410_, new_n26411_,
    new_n26412_, new_n26413_, new_n26414_, new_n26415_, new_n26416_,
    new_n26417_, new_n26418_, new_n26419_, new_n26420_, new_n26421_,
    new_n26422_, new_n26423_, new_n26424_, new_n26425_, new_n26426_,
    new_n26427_, new_n26428_, new_n26429_, new_n26430_, new_n26431_,
    new_n26432_, new_n26433_, new_n26434_, new_n26435_, new_n26436_,
    new_n26437_, new_n26438_, new_n26439_, new_n26440_, new_n26441_,
    new_n26442_, new_n26443_, new_n26444_, new_n26445_, new_n26446_,
    new_n26447_, new_n26448_, new_n26449_, new_n26450_, new_n26451_,
    new_n26452_, new_n26453_, new_n26454_, new_n26455_, new_n26456_,
    new_n26457_, new_n26458_, new_n26459_, new_n26460_, new_n26461_,
    new_n26462_, new_n26463_, new_n26464_, new_n26465_, new_n26466_,
    new_n26467_, new_n26468_, new_n26469_, new_n26470_, new_n26471_,
    new_n26472_, new_n26473_, new_n26474_, new_n26475_, new_n26476_,
    new_n26477_, new_n26478_, new_n26479_, new_n26480_, new_n26481_,
    new_n26482_, new_n26483_, new_n26484_, new_n26485_, new_n26486_,
    new_n26487_, new_n26488_, new_n26489_, new_n26490_, new_n26491_,
    new_n26492_, new_n26493_, new_n26494_, new_n26495_, new_n26496_,
    new_n26497_, new_n26498_, new_n26499_, new_n26500_, new_n26501_,
    new_n26502_, new_n26503_, new_n26504_, new_n26505_, new_n26506_,
    new_n26507_, new_n26508_, new_n26509_, new_n26510_, new_n26511_,
    new_n26512_, new_n26513_, new_n26514_, new_n26515_, new_n26516_,
    new_n26517_, new_n26518_, new_n26519_, new_n26520_, new_n26521_,
    new_n26522_, new_n26523_, new_n26524_, new_n26525_, new_n26526_,
    new_n26527_, new_n26528_, new_n26529_, new_n26530_, new_n26531_,
    new_n26532_, new_n26533_, new_n26534_, new_n26535_, new_n26536_,
    new_n26537_, new_n26538_, new_n26539_, new_n26540_, new_n26541_,
    new_n26542_, new_n26543_, new_n26544_, new_n26545_, new_n26546_,
    new_n26547_, new_n26548_, new_n26549_, new_n26550_, new_n26551_,
    new_n26552_, new_n26553_, new_n26554_, new_n26555_, new_n26556_,
    new_n26557_, new_n26558_, new_n26559_, new_n26560_, new_n26561_,
    new_n26562_, new_n26563_, new_n26564_, new_n26565_, new_n26566_,
    new_n26567_, new_n26568_, new_n26569_, new_n26570_, new_n26571_,
    new_n26572_, new_n26573_, new_n26574_, new_n26575_, new_n26576_,
    new_n26577_, new_n26578_, new_n26579_, new_n26580_, new_n26581_,
    new_n26582_, new_n26583_, new_n26584_, new_n26585_, new_n26586_,
    new_n26587_, new_n26588_, new_n26589_, new_n26590_, new_n26591_,
    new_n26592_, new_n26593_, new_n26594_, new_n26595_, new_n26596_,
    new_n26597_, new_n26598_, new_n26599_, new_n26600_, new_n26601_,
    new_n26602_, new_n26603_, new_n26604_, new_n26605_, new_n26606_,
    new_n26607_, new_n26608_, new_n26609_, new_n26610_, new_n26611_,
    new_n26612_, new_n26613_, new_n26614_, new_n26615_, new_n26616_,
    new_n26617_, new_n26618_, new_n26619_, new_n26620_, new_n26621_,
    new_n26622_, new_n26623_, new_n26624_, new_n26625_, new_n26626_,
    new_n26627_, new_n26628_, new_n26629_, new_n26630_, new_n26631_,
    new_n26632_, new_n26633_, new_n26634_, new_n26635_, new_n26636_,
    new_n26637_, new_n26638_, new_n26639_, new_n26640_, new_n26641_,
    new_n26642_, new_n26643_, new_n26644_, new_n26645_, new_n26646_,
    new_n26647_, new_n26648_, new_n26649_, new_n26650_, new_n26651_,
    new_n26652_, new_n26653_, new_n26654_, new_n26655_, new_n26656_,
    new_n26657_, new_n26658_, new_n26659_, new_n26660_, new_n26661_,
    new_n26662_, new_n26663_, new_n26664_, new_n26665_, new_n26666_,
    new_n26667_, new_n26668_, new_n26669_, new_n26670_, new_n26671_,
    new_n26672_, new_n26673_, new_n26674_, new_n26675_, new_n26676_,
    new_n26677_, new_n26678_, new_n26679_, new_n26680_, new_n26681_,
    new_n26682_, new_n26683_, new_n26684_, new_n26685_, new_n26686_,
    new_n26687_, new_n26688_, new_n26689_, new_n26690_, new_n26691_,
    new_n26692_, new_n26693_, new_n26694_, new_n26695_, new_n26696_,
    new_n26697_, new_n26698_, new_n26699_, new_n26700_, new_n26701_,
    new_n26702_, new_n26703_, new_n26704_, new_n26705_, new_n26706_,
    new_n26707_, new_n26708_, new_n26709_, new_n26710_, new_n26711_,
    new_n26712_, new_n26713_, new_n26714_, new_n26715_, new_n26716_,
    new_n26717_, new_n26718_, new_n26719_, new_n26720_, new_n26721_,
    new_n26722_, new_n26723_, new_n26724_, new_n26725_, new_n26726_,
    new_n26727_, new_n26728_, new_n26729_, new_n26730_, new_n26731_,
    new_n26732_, new_n26733_, new_n26734_, new_n26735_, new_n26736_,
    new_n26737_, new_n26738_, new_n26739_, new_n26740_, new_n26741_,
    new_n26742_, new_n26743_, new_n26744_, new_n26745_, new_n26746_,
    new_n26747_, new_n26748_, new_n26749_, new_n26750_, new_n26751_,
    new_n26752_, new_n26753_, new_n26754_, new_n26755_, new_n26756_,
    new_n26757_, new_n26758_, new_n26759_, new_n26760_, new_n26761_,
    new_n26762_, new_n26763_, new_n26764_, new_n26765_, new_n26766_,
    new_n26767_, new_n26768_, new_n26769_, new_n26770_, new_n26771_,
    new_n26772_, new_n26773_, new_n26774_, new_n26775_, new_n26776_,
    new_n26777_, new_n26778_, new_n26779_, new_n26780_, new_n26781_,
    new_n26782_, new_n26783_, new_n26784_, new_n26785_, new_n26786_,
    new_n26787_, new_n26788_, new_n26789_, new_n26790_, new_n26791_,
    new_n26792_, new_n26793_, new_n26794_, new_n26795_, new_n26796_,
    new_n26797_, new_n26798_, new_n26799_, new_n26800_, new_n26801_,
    new_n26802_, new_n26803_, new_n26804_, new_n26805_, new_n26806_,
    new_n26807_, new_n26808_, new_n26809_, new_n26810_, new_n26811_,
    new_n26812_, new_n26813_, new_n26814_, new_n26815_, new_n26816_,
    new_n26817_, new_n26818_, new_n26819_, new_n26820_, new_n26821_,
    new_n26822_, new_n26823_, new_n26824_, new_n26825_, new_n26826_,
    new_n26827_, new_n26828_, new_n26829_, new_n26830_, new_n26831_,
    new_n26832_, new_n26833_, new_n26834_, new_n26835_, new_n26836_,
    new_n26837_, new_n26838_, new_n26839_, new_n26840_, new_n26841_,
    new_n26842_, new_n26843_, new_n26844_, new_n26845_, new_n26846_,
    new_n26847_, new_n26848_, new_n26849_, new_n26850_, new_n26851_,
    new_n26852_, new_n26853_, new_n26854_, new_n26855_, new_n26856_,
    new_n26857_, new_n26858_, new_n26859_, new_n26860_, new_n26861_,
    new_n26862_, new_n26863_, new_n26864_, new_n26865_, new_n26866_,
    new_n26867_, new_n26868_, new_n26869_, new_n26870_, new_n26871_,
    new_n26872_, new_n26873_, new_n26874_, new_n26875_, new_n26876_,
    new_n26877_, new_n26878_, new_n26879_, new_n26880_, new_n26881_,
    new_n26882_, new_n26883_, new_n26884_, new_n26885_, new_n26886_,
    new_n26887_, new_n26888_, new_n26889_, new_n26890_, new_n26891_,
    new_n26892_, new_n26893_, new_n26894_, new_n26895_, new_n26896_,
    new_n26897_, new_n26898_, new_n26899_, new_n26900_, new_n26901_,
    new_n26902_, new_n26903_, new_n26904_, new_n26905_, new_n26906_,
    new_n26907_, new_n26908_, new_n26909_, new_n26910_, new_n26911_,
    new_n26912_, new_n26913_, new_n26914_, new_n26915_, new_n26916_,
    new_n26917_, new_n26918_, new_n26919_, new_n26920_, new_n26921_,
    new_n26922_, new_n26923_, new_n26924_, new_n26925_, new_n26926_,
    new_n26927_, new_n26928_, new_n26929_, new_n26930_, new_n26931_,
    new_n26932_, new_n26933_, new_n26934_, new_n26935_, new_n26936_,
    new_n26937_, new_n26938_, new_n26939_, new_n26940_, new_n26941_,
    new_n26942_, new_n26943_, new_n26944_, new_n26945_, new_n26946_,
    new_n26947_, new_n26948_, new_n26949_, new_n26950_, new_n26951_,
    new_n26952_, new_n26953_, new_n26954_, new_n26955_, new_n26956_,
    new_n26957_, new_n26958_, new_n26959_, new_n26960_, new_n26961_,
    new_n26962_, new_n26963_, new_n26964_, new_n26965_, new_n26966_,
    new_n26967_, new_n26968_, new_n26969_, new_n26970_, new_n26971_,
    new_n26972_, new_n26973_, new_n26974_, new_n26975_, new_n26976_,
    new_n26977_, new_n26978_, new_n26979_, new_n26980_, new_n26981_,
    new_n26982_, new_n26983_, new_n26984_, new_n26985_, new_n26986_,
    new_n26987_, new_n26988_, new_n26989_, new_n26990_, new_n26991_,
    new_n26992_, new_n26993_, new_n26994_, new_n26995_, new_n26996_,
    new_n26997_, new_n26998_, new_n26999_, new_n27000_, new_n27001_,
    new_n27002_, new_n27003_, new_n27004_, new_n27005_, new_n27006_,
    new_n27007_, new_n27008_, new_n27009_, new_n27010_, new_n27011_,
    new_n27012_, new_n27013_, new_n27014_, new_n27015_, new_n27016_,
    new_n27017_, new_n27018_, new_n27019_, new_n27020_, new_n27021_,
    new_n27022_, new_n27023_, new_n27024_, new_n27025_, new_n27026_,
    new_n27027_, new_n27028_, new_n27029_, new_n27030_, new_n27031_,
    new_n27032_, new_n27033_, new_n27034_, new_n27035_, new_n27036_,
    new_n27037_, new_n27038_, new_n27039_, new_n27040_, new_n27041_,
    new_n27042_, new_n27043_, new_n27044_, new_n27045_, new_n27046_,
    new_n27047_, new_n27048_, new_n27049_, new_n27050_, new_n27051_,
    new_n27052_, new_n27053_, new_n27054_, new_n27055_, new_n27056_,
    new_n27057_, new_n27058_, new_n27059_, new_n27060_, new_n27061_,
    new_n27062_, new_n27063_, new_n27064_, new_n27065_, new_n27066_,
    new_n27067_, new_n27068_, new_n27069_, new_n27070_, new_n27071_,
    new_n27072_, new_n27073_, new_n27074_, new_n27075_, new_n27076_,
    new_n27077_, new_n27078_, new_n27079_, new_n27080_, new_n27081_,
    new_n27082_, new_n27083_, new_n27084_, new_n27085_, new_n27086_,
    new_n27087_, new_n27088_, new_n27089_, new_n27090_, new_n27091_,
    new_n27092_, new_n27093_, new_n27094_, new_n27095_, new_n27096_,
    new_n27097_, new_n27098_, new_n27099_, new_n27100_, new_n27101_,
    new_n27102_, new_n27103_, new_n27104_, new_n27105_, new_n27106_,
    new_n27107_, new_n27108_, new_n27109_, new_n27110_, new_n27111_,
    new_n27112_, new_n27113_, new_n27114_, new_n27115_, new_n27116_,
    new_n27117_, new_n27118_, new_n27119_, new_n27120_, new_n27121_,
    new_n27122_, new_n27123_, new_n27124_, new_n27125_, new_n27126_,
    new_n27127_, new_n27128_, new_n27129_, new_n27130_, new_n27131_,
    new_n27132_, new_n27133_, new_n27134_, new_n27135_, new_n27136_,
    new_n27137_, new_n27138_, new_n27139_, new_n27140_, new_n27141_,
    new_n27142_, new_n27143_, new_n27144_, new_n27145_, new_n27146_,
    new_n27147_, new_n27148_, new_n27149_, new_n27150_, new_n27151_,
    new_n27152_, new_n27153_, new_n27154_, new_n27155_, new_n27156_,
    new_n27157_, new_n27158_, new_n27159_, new_n27160_, new_n27161_,
    new_n27162_, new_n27163_, new_n27164_, new_n27165_, new_n27166_,
    new_n27167_, new_n27168_, new_n27169_, new_n27170_, new_n27171_,
    new_n27172_, new_n27173_, new_n27174_, new_n27175_, new_n27176_,
    new_n27177_, new_n27178_, new_n27179_, new_n27180_, new_n27181_,
    new_n27182_, new_n27183_, new_n27184_, new_n27185_, new_n27186_,
    new_n27187_, new_n27188_, new_n27189_, new_n27190_, new_n27191_,
    new_n27192_, new_n27193_, new_n27194_, new_n27195_, new_n27196_,
    new_n27197_, new_n27198_, new_n27199_, new_n27200_, new_n27201_,
    new_n27202_, new_n27203_, new_n27204_, new_n27205_, new_n27206_,
    new_n27207_, new_n27208_, new_n27209_, new_n27210_, new_n27211_,
    new_n27212_, new_n27213_, new_n27214_, new_n27215_, new_n27216_,
    new_n27217_, new_n27218_, new_n27219_, new_n27220_, new_n27221_,
    new_n27222_, new_n27223_, new_n27224_, new_n27225_, new_n27226_,
    new_n27227_, new_n27228_, new_n27229_, new_n27230_, new_n27231_,
    new_n27232_, new_n27233_, new_n27234_, new_n27235_, new_n27236_,
    new_n27237_, new_n27238_, new_n27239_, new_n27240_, new_n27241_,
    new_n27242_, new_n27243_, new_n27244_, new_n27245_, new_n27246_,
    new_n27247_, new_n27248_, new_n27249_, new_n27250_, new_n27251_,
    new_n27252_, new_n27253_, new_n27254_, new_n27255_, new_n27256_,
    new_n27257_, new_n27258_, new_n27259_, new_n27260_, new_n27261_,
    new_n27262_, new_n27263_, new_n27264_, new_n27265_, new_n27266_,
    new_n27267_, new_n27268_, new_n27269_, new_n27270_, new_n27271_,
    new_n27272_, new_n27273_, new_n27274_, new_n27275_, new_n27276_,
    new_n27277_, new_n27278_, new_n27279_, new_n27280_, new_n27281_,
    new_n27282_, new_n27283_, new_n27284_, new_n27285_, new_n27286_,
    new_n27287_, new_n27288_, new_n27289_, new_n27290_, new_n27291_,
    new_n27292_, new_n27293_, new_n27294_, new_n27295_, new_n27296_,
    new_n27297_, new_n27298_, new_n27299_, new_n27300_, new_n27301_,
    new_n27302_, new_n27303_, new_n27304_, new_n27305_, new_n27306_,
    new_n27307_, new_n27308_, new_n27309_, new_n27310_, new_n27311_,
    new_n27312_, new_n27313_, new_n27314_, new_n27315_, new_n27316_,
    new_n27317_, new_n27318_, new_n27319_, new_n27320_, new_n27321_,
    new_n27322_, new_n27323_, new_n27324_, new_n27325_, new_n27326_,
    new_n27327_, new_n27328_, new_n27329_, new_n27330_, new_n27331_,
    new_n27332_, new_n27333_, new_n27334_, new_n27335_, new_n27336_,
    new_n27337_, new_n27338_, new_n27339_, new_n27340_, new_n27341_,
    new_n27342_, new_n27343_, new_n27344_, new_n27345_, new_n27346_,
    new_n27347_, new_n27348_, new_n27349_, new_n27350_, new_n27351_,
    new_n27352_, new_n27353_, new_n27354_, new_n27355_, new_n27356_,
    new_n27357_, new_n27358_, new_n27359_, new_n27360_, new_n27361_,
    new_n27362_, new_n27363_, new_n27364_, new_n27365_, new_n27366_,
    new_n27367_, new_n27368_, new_n27369_, new_n27370_, new_n27371_,
    new_n27372_, new_n27373_, new_n27374_, new_n27375_, new_n27376_,
    new_n27377_, new_n27378_, new_n27379_, new_n27380_, new_n27381_,
    new_n27382_, new_n27383_, new_n27384_, new_n27385_, new_n27386_,
    new_n27387_, new_n27388_, new_n27389_, new_n27390_, new_n27391_,
    new_n27392_, new_n27393_, new_n27394_, new_n27395_, new_n27396_,
    new_n27397_, new_n27398_, new_n27399_, new_n27400_, new_n27401_,
    new_n27402_, new_n27403_, new_n27404_, new_n27405_, new_n27406_,
    new_n27407_, new_n27408_, new_n27409_, new_n27410_, new_n27411_,
    new_n27412_, new_n27413_, new_n27414_, new_n27415_, new_n27416_,
    new_n27417_, new_n27418_, new_n27419_, new_n27420_, new_n27421_,
    new_n27422_, new_n27423_, new_n27424_, new_n27425_, new_n27426_,
    new_n27427_, new_n27428_, new_n27429_, new_n27430_, new_n27431_,
    new_n27432_, new_n27433_, new_n27434_, new_n27435_, new_n27436_,
    new_n27437_, new_n27438_, new_n27439_, new_n27440_, new_n27441_,
    new_n27442_, new_n27443_, new_n27444_, new_n27445_, new_n27446_,
    new_n27447_, new_n27448_, new_n27449_, new_n27450_, new_n27451_,
    new_n27452_, new_n27453_, new_n27454_, new_n27455_, new_n27456_,
    new_n27457_, new_n27458_, new_n27459_, new_n27460_, new_n27461_,
    new_n27462_, new_n27463_, new_n27464_, new_n27465_, new_n27466_,
    new_n27467_, new_n27468_, new_n27469_, new_n27470_, new_n27471_,
    new_n27472_, new_n27473_, new_n27474_, new_n27475_, new_n27476_,
    new_n27477_, new_n27478_, new_n27479_, new_n27480_, new_n27481_,
    new_n27482_, new_n27483_, new_n27484_, new_n27485_, new_n27486_,
    new_n27487_, new_n27488_, new_n27489_, new_n27490_, new_n27491_,
    new_n27492_, new_n27493_, new_n27494_, new_n27495_, new_n27496_,
    new_n27497_, new_n27498_, new_n27499_, new_n27500_, new_n27501_,
    new_n27502_, new_n27503_, new_n27504_, new_n27505_, new_n27506_,
    new_n27507_, new_n27508_, new_n27509_, new_n27510_, new_n27511_,
    new_n27512_, new_n27513_, new_n27514_, new_n27515_, new_n27516_,
    new_n27517_, new_n27518_, new_n27519_, new_n27520_, new_n27521_,
    new_n27522_, new_n27523_, new_n27524_, new_n27525_, new_n27526_,
    new_n27527_, new_n27528_, new_n27529_, new_n27530_, new_n27531_,
    new_n27532_, new_n27533_, new_n27534_, new_n27535_, new_n27536_,
    new_n27537_, new_n27538_, new_n27539_, new_n27540_, new_n27541_,
    new_n27542_, new_n27543_, new_n27544_, new_n27545_, new_n27546_,
    new_n27547_, new_n27548_, new_n27549_, new_n27550_, new_n27551_,
    new_n27552_, new_n27553_, new_n27554_, new_n27555_, new_n27556_,
    new_n27557_, new_n27558_, new_n27559_, new_n27560_, new_n27561_,
    new_n27562_, new_n27563_, new_n27564_, new_n27565_, new_n27566_,
    new_n27567_, new_n27568_, new_n27569_, new_n27570_, new_n27571_,
    new_n27572_, new_n27573_, new_n27574_, new_n27575_, new_n27576_,
    new_n27577_, new_n27578_, new_n27579_, new_n27580_, new_n27581_,
    new_n27582_, new_n27583_, new_n27584_, new_n27585_, new_n27586_,
    new_n27587_, new_n27588_, new_n27589_, new_n27590_, new_n27591_,
    new_n27592_, new_n27593_, new_n27594_, new_n27595_, new_n27596_,
    new_n27597_, new_n27598_, new_n27599_, new_n27600_, new_n27601_,
    new_n27602_, new_n27603_, new_n27604_, new_n27605_, new_n27606_,
    new_n27607_, new_n27608_, new_n27609_, new_n27610_, new_n27611_,
    new_n27612_, new_n27613_, new_n27614_, new_n27615_, new_n27616_,
    new_n27617_, new_n27618_, new_n27619_, new_n27620_, new_n27621_,
    new_n27622_, new_n27623_, new_n27624_, new_n27625_, new_n27626_,
    new_n27627_, new_n27628_, new_n27629_, new_n27630_, new_n27631_,
    new_n27632_, new_n27633_, new_n27634_, new_n27635_, new_n27636_,
    new_n27637_, new_n27638_, new_n27639_, new_n27640_, new_n27641_,
    new_n27642_, new_n27643_, new_n27644_, new_n27645_, new_n27646_,
    new_n27647_, new_n27648_, new_n27649_, new_n27650_, new_n27651_,
    new_n27652_, new_n27653_, new_n27654_, new_n27655_, new_n27656_,
    new_n27657_, new_n27658_, new_n27659_, new_n27660_, new_n27661_,
    new_n27662_, new_n27663_, new_n27664_, new_n27665_, new_n27666_,
    new_n27667_, new_n27668_, new_n27669_, new_n27670_, new_n27671_,
    new_n27672_, new_n27673_, new_n27674_, new_n27675_, new_n27676_,
    new_n27677_, new_n27678_, new_n27679_, new_n27680_, new_n27681_,
    new_n27682_, new_n27683_, new_n27684_, new_n27685_, new_n27686_,
    new_n27687_, new_n27688_, new_n27689_, new_n27690_, new_n27691_,
    new_n27692_, new_n27693_, new_n27694_, new_n27695_, new_n27696_,
    new_n27697_, new_n27698_, new_n27699_, new_n27700_, new_n27701_,
    new_n27702_, new_n27703_, new_n27704_, new_n27705_, new_n27706_,
    new_n27707_, new_n27708_, new_n27709_, new_n27710_, new_n27711_,
    new_n27712_, new_n27713_, new_n27714_, new_n27715_, new_n27716_,
    new_n27717_, new_n27718_, new_n27719_, new_n27720_, new_n27721_,
    new_n27722_, new_n27723_, new_n27724_, new_n27725_, new_n27726_,
    new_n27727_, new_n27728_, new_n27729_, new_n27730_, new_n27731_,
    new_n27732_, new_n27733_, new_n27734_, new_n27735_, new_n27736_,
    new_n27737_, new_n27738_, new_n27739_, new_n27740_, new_n27741_,
    new_n27742_, new_n27743_, new_n27744_, new_n27745_, new_n27746_,
    new_n27747_, new_n27748_, new_n27749_, new_n27750_, new_n27751_,
    new_n27752_, new_n27753_, new_n27754_, new_n27755_, new_n27756_,
    new_n27757_, new_n27758_, new_n27759_, new_n27760_, new_n27761_,
    new_n27762_, new_n27763_, new_n27764_, new_n27765_, new_n27766_,
    new_n27767_, new_n27768_, new_n27769_, new_n27770_, new_n27771_,
    new_n27772_, new_n27773_, new_n27774_, new_n27775_, new_n27776_,
    new_n27777_, new_n27778_, new_n27779_, new_n27780_, new_n27781_,
    new_n27782_, new_n27783_, new_n27784_, new_n27785_, new_n27786_,
    new_n27787_, new_n27788_, new_n27789_, new_n27790_, new_n27791_,
    new_n27792_, new_n27793_, new_n27794_, new_n27795_, new_n27796_,
    new_n27797_, new_n27798_, new_n27799_, new_n27800_, new_n27801_,
    new_n27802_, new_n27803_, new_n27804_, new_n27805_, new_n27806_,
    new_n27807_, new_n27808_, new_n27809_, new_n27810_, new_n27811_,
    new_n27812_, new_n27813_, new_n27814_, new_n27815_, new_n27816_,
    new_n27817_, new_n27818_, new_n27819_, new_n27820_, new_n27821_,
    new_n27822_, new_n27823_, new_n27824_, new_n27825_, new_n27826_,
    new_n27827_, new_n27828_, new_n27829_, new_n27830_, new_n27831_,
    new_n27832_, new_n27833_, new_n27834_, new_n27835_, new_n27836_,
    new_n27837_, new_n27838_, new_n27839_, new_n27840_, new_n27841_,
    new_n27842_, new_n27843_, new_n27844_, new_n27845_, new_n27846_,
    new_n27847_, new_n27848_, new_n27849_, new_n27850_, new_n27851_,
    new_n27852_, new_n27853_, new_n27854_, new_n27855_, new_n27856_,
    new_n27857_, new_n27858_, new_n27859_, new_n27860_, new_n27861_,
    new_n27862_, new_n27863_, new_n27864_, new_n27865_, new_n27866_,
    new_n27867_, new_n27868_, new_n27869_, new_n27870_, new_n27871_,
    new_n27872_, new_n27873_, new_n27874_, new_n27875_, new_n27876_,
    new_n27877_, new_n27878_, new_n27879_, new_n27880_, new_n27881_,
    new_n27882_, new_n27883_, new_n27884_, new_n27885_, new_n27886_,
    new_n27887_, new_n27888_, new_n27889_, new_n27890_, new_n27891_,
    new_n27892_, new_n27893_, new_n27894_, new_n27895_, new_n27896_,
    new_n27897_, new_n27898_, new_n27899_, new_n27900_, new_n27901_,
    new_n27902_, new_n27903_, new_n27904_, new_n27905_, new_n27906_,
    new_n27907_, new_n27908_, new_n27909_, new_n27910_, new_n27911_,
    new_n27912_, new_n27913_, new_n27914_, new_n27915_, new_n27916_,
    new_n27917_, new_n27918_, new_n27919_, new_n27920_, new_n27921_,
    new_n27922_, new_n27923_, new_n27924_, new_n27925_, new_n27926_,
    new_n27927_, new_n27928_, new_n27929_, new_n27930_, new_n27931_,
    new_n27932_, new_n27933_, new_n27934_, new_n27935_, new_n27936_,
    new_n27937_, new_n27938_, new_n27939_, new_n27940_, new_n27941_,
    new_n27942_, new_n27943_, new_n27944_, new_n27945_, new_n27946_,
    new_n27947_, new_n27948_, new_n27949_, new_n27950_, new_n27951_,
    new_n27952_, new_n27953_, new_n27954_, new_n27955_, new_n27956_,
    new_n27957_, new_n27958_, new_n27959_, new_n27960_, new_n27961_,
    new_n27962_, new_n27963_, new_n27964_, new_n27965_, new_n27966_,
    new_n27967_, new_n27968_, new_n27969_, new_n27970_, new_n27971_,
    new_n27972_, new_n27973_, new_n27974_, new_n27975_, new_n27976_,
    new_n27977_, new_n27978_, new_n27979_, new_n27980_, new_n27981_,
    new_n27982_, new_n27983_, new_n27984_, new_n27985_, new_n27986_,
    new_n27987_, new_n27988_, new_n27989_, new_n27990_, new_n27991_,
    new_n27992_, new_n27993_, new_n27994_, new_n27995_, new_n27996_,
    new_n27997_, new_n27998_, new_n27999_, new_n28000_, new_n28001_,
    new_n28002_, new_n28003_, new_n28004_, new_n28005_, new_n28006_,
    new_n28007_, new_n28008_, new_n28009_, new_n28010_, new_n28011_,
    new_n28012_, new_n28013_, new_n28014_, new_n28015_, new_n28016_,
    new_n28017_, new_n28018_, new_n28019_, new_n28020_, new_n28021_,
    new_n28022_, new_n28023_, new_n28024_, new_n28025_, new_n28026_,
    new_n28027_, new_n28028_, new_n28029_, new_n28030_, new_n28031_,
    new_n28032_, new_n28033_, new_n28034_, new_n28035_, new_n28036_,
    new_n28037_, new_n28038_, new_n28039_, new_n28040_, new_n28041_,
    new_n28042_, new_n28043_, new_n28044_, new_n28045_, new_n28046_,
    new_n28047_, new_n28048_, new_n28049_, new_n28050_, new_n28051_,
    new_n28052_, new_n28053_, new_n28054_, new_n28055_, new_n28056_,
    new_n28057_, new_n28058_, new_n28059_, new_n28060_, new_n28061_,
    new_n28062_, new_n28063_, new_n28064_, new_n28065_, new_n28066_,
    new_n28067_, new_n28068_, new_n28069_, new_n28070_, new_n28071_,
    new_n28072_, new_n28073_, new_n28074_, new_n28075_, new_n28076_,
    new_n28077_, new_n28078_, new_n28079_, new_n28080_, new_n28081_,
    new_n28082_, new_n28083_, new_n28084_, new_n28085_, new_n28086_,
    new_n28087_, new_n28088_, new_n28089_, new_n28090_, new_n28091_,
    new_n28092_, new_n28093_, new_n28094_, new_n28095_, new_n28096_,
    new_n28097_, new_n28098_, new_n28099_, new_n28100_, new_n28101_,
    new_n28102_, new_n28103_, new_n28104_, new_n28105_, new_n28106_,
    new_n28107_, new_n28108_, new_n28109_, new_n28110_, new_n28111_,
    new_n28112_, new_n28113_, new_n28114_, new_n28115_, new_n28116_,
    new_n28117_, new_n28118_, new_n28119_, new_n28120_, new_n28121_,
    new_n28122_, new_n28123_, new_n28124_, new_n28125_, new_n28126_,
    new_n28127_, new_n28128_, new_n28129_, new_n28130_, new_n28131_,
    new_n28132_, new_n28133_, new_n28134_, new_n28135_, new_n28136_,
    new_n28137_, new_n28138_, new_n28139_, new_n28140_, new_n28141_,
    new_n28142_, new_n28143_, new_n28144_, new_n28145_, new_n28146_,
    new_n28147_, new_n28148_, new_n28149_, new_n28150_, new_n28151_,
    new_n28152_, new_n28153_, new_n28154_, new_n28155_, new_n28156_,
    new_n28157_, new_n28158_, new_n28159_, new_n28160_, new_n28161_,
    new_n28162_, new_n28163_, new_n28164_, new_n28165_, new_n28166_,
    new_n28167_, new_n28168_, new_n28169_, new_n28170_, new_n28171_,
    new_n28172_, new_n28173_, new_n28174_, new_n28175_, new_n28176_,
    new_n28177_, new_n28178_, new_n28179_, new_n28180_, new_n28181_,
    new_n28182_, new_n28183_, new_n28184_, new_n28185_, new_n28186_,
    new_n28187_, new_n28188_, new_n28189_, new_n28190_, new_n28191_,
    new_n28192_, new_n28193_, new_n28194_, new_n28195_, new_n28196_,
    new_n28197_, new_n28198_, new_n28199_, new_n28200_, new_n28201_,
    new_n28202_, new_n28203_, new_n28204_, new_n28205_, new_n28206_,
    new_n28207_, new_n28208_, new_n28209_, new_n28210_, new_n28211_,
    new_n28212_, new_n28213_, new_n28214_, new_n28215_, new_n28216_,
    new_n28217_, new_n28218_, new_n28219_, new_n28220_, new_n28221_,
    new_n28222_, new_n28223_, new_n28224_, new_n28225_, new_n28226_,
    new_n28227_, new_n28228_, new_n28229_, new_n28230_, new_n28231_,
    new_n28232_, new_n28233_, new_n28234_, new_n28235_, new_n28236_,
    new_n28237_, new_n28238_, new_n28239_, new_n28240_, new_n28241_,
    new_n28242_, new_n28243_, new_n28244_, new_n28245_, new_n28246_,
    new_n28247_, new_n28248_, new_n28249_, new_n28250_, new_n28251_,
    new_n28252_, new_n28253_, new_n28254_, new_n28255_, new_n28256_,
    new_n28257_, new_n28258_, new_n28259_, new_n28260_, new_n28261_,
    new_n28262_, new_n28263_, new_n28264_, new_n28265_, new_n28266_,
    new_n28267_, new_n28268_, new_n28269_, new_n28270_, new_n28271_,
    new_n28272_, new_n28273_, new_n28274_, new_n28275_, new_n28276_,
    new_n28277_, new_n28278_, new_n28279_, new_n28280_, new_n28281_,
    new_n28282_, new_n28283_, new_n28284_, new_n28285_, new_n28286_,
    new_n28287_, new_n28288_, new_n28289_, new_n28290_, new_n28291_,
    new_n28292_, new_n28293_, new_n28294_, new_n28295_, new_n28296_,
    new_n28297_, new_n28298_, new_n28299_, new_n28300_, new_n28301_,
    new_n28302_, new_n28303_, new_n28304_, new_n28305_, new_n28306_,
    new_n28307_, new_n28308_, new_n28309_, new_n28310_, new_n28311_,
    new_n28312_, new_n28313_, new_n28314_, new_n28315_, new_n28316_,
    new_n28317_, new_n28318_, new_n28319_, new_n28320_, new_n28321_,
    new_n28322_, new_n28323_, new_n28324_, new_n28325_, new_n28326_,
    new_n28327_, new_n28328_, new_n28329_, new_n28330_, new_n28331_,
    new_n28332_, new_n28333_, new_n28334_, new_n28335_, new_n28336_,
    new_n28337_, new_n28338_, new_n28339_, new_n28340_, new_n28341_,
    new_n28342_, new_n28343_, new_n28344_, new_n28345_, new_n28346_,
    new_n28347_, new_n28348_, new_n28349_, new_n28350_, new_n28351_,
    new_n28352_, new_n28353_, new_n28354_, new_n28355_, new_n28356_,
    new_n28357_, new_n28358_, new_n28359_, new_n28360_, new_n28361_,
    new_n28362_, new_n28363_, new_n28364_, new_n28365_, new_n28366_,
    new_n28367_, new_n28368_, new_n28369_, new_n28370_, new_n28371_,
    new_n28372_, new_n28373_, new_n28374_, new_n28375_, new_n28376_,
    new_n28377_, new_n28378_, new_n28379_, new_n28380_, new_n28381_,
    new_n28382_, new_n28383_, new_n28384_, new_n28385_, new_n28386_,
    new_n28387_, new_n28388_, new_n28389_, new_n28390_, new_n28391_,
    new_n28392_, new_n28393_, new_n28394_, new_n28395_, new_n28396_,
    new_n28397_, new_n28398_, new_n28399_, new_n28400_, new_n28401_,
    new_n28402_, new_n28403_, new_n28404_, new_n28405_, new_n28406_,
    new_n28407_, new_n28408_, new_n28409_, new_n28410_, new_n28411_,
    new_n28412_, new_n28413_, new_n28414_, new_n28415_, new_n28416_,
    new_n28417_, new_n28418_, new_n28419_, new_n28420_, new_n28421_,
    new_n28422_, new_n28423_, new_n28424_, new_n28425_, new_n28426_,
    new_n28427_, new_n28428_, new_n28429_, new_n28430_, new_n28431_,
    new_n28432_, new_n28433_, new_n28434_, new_n28435_, new_n28436_,
    new_n28437_, new_n28438_, new_n28439_, new_n28440_, new_n28441_,
    new_n28442_, new_n28443_, new_n28444_, new_n28445_, new_n28446_,
    new_n28447_, new_n28448_, new_n28449_, new_n28450_, new_n28451_,
    new_n28452_, new_n28453_, new_n28454_, new_n28455_, new_n28456_,
    new_n28457_, new_n28458_, new_n28459_, new_n28460_, new_n28461_,
    new_n28462_, new_n28463_, new_n28464_, new_n28465_, new_n28466_,
    new_n28467_, new_n28468_, new_n28469_, new_n28470_, new_n28471_,
    new_n28472_, new_n28473_, new_n28474_, new_n28475_, new_n28476_,
    new_n28477_, new_n28478_, new_n28479_, new_n28480_, new_n28481_,
    new_n28482_, new_n28483_, new_n28484_, new_n28485_, new_n28486_,
    new_n28487_, new_n28488_, new_n28489_, new_n28490_, new_n28491_,
    new_n28492_, new_n28493_, new_n28494_, new_n28495_, new_n28496_,
    new_n28497_, new_n28498_, new_n28499_, new_n28500_, new_n28501_,
    new_n28502_, new_n28503_, new_n28504_, new_n28505_, new_n28506_,
    new_n28507_, new_n28508_, new_n28509_, new_n28510_, new_n28511_,
    new_n28512_, new_n28513_, new_n28514_, new_n28515_, new_n28516_,
    new_n28517_, new_n28518_, new_n28519_, new_n28520_, new_n28521_,
    new_n28522_, new_n28523_, new_n28524_, new_n28525_, new_n28526_,
    new_n28527_, new_n28528_, new_n28529_, new_n28530_, new_n28531_,
    new_n28532_, new_n28533_, new_n28534_, new_n28535_, new_n28536_,
    new_n28537_, new_n28538_, new_n28539_, new_n28540_, new_n28541_,
    new_n28542_, new_n28543_, new_n28544_, new_n28545_, new_n28546_,
    new_n28547_, new_n28548_, new_n28549_, new_n28550_, new_n28551_,
    new_n28552_, new_n28553_, new_n28554_, new_n28555_, new_n28556_,
    new_n28557_, new_n28558_, new_n28559_, new_n28560_, new_n28561_,
    new_n28562_, new_n28563_, new_n28564_, new_n28565_, new_n28566_,
    new_n28567_, new_n28568_, new_n28569_, new_n28570_, new_n28571_,
    new_n28572_, new_n28573_, new_n28574_, new_n28575_, new_n28576_,
    new_n28577_, new_n28578_, new_n28579_, new_n28580_, new_n28581_,
    new_n28582_, new_n28583_, new_n28584_, new_n28585_, new_n28586_,
    new_n28587_, new_n28588_, new_n28589_, new_n28590_, new_n28591_,
    new_n28592_, new_n28593_, new_n28594_, new_n28595_, new_n28596_,
    new_n28597_, new_n28598_, new_n28599_, new_n28600_, new_n28601_,
    new_n28602_, new_n28603_, new_n28604_, new_n28605_, new_n28606_,
    new_n28607_, new_n28608_, new_n28609_, new_n28610_, new_n28611_,
    new_n28612_, new_n28613_, new_n28614_, new_n28615_, new_n28616_,
    new_n28617_, new_n28618_, new_n28619_, new_n28620_, new_n28621_,
    new_n28622_, new_n28623_, new_n28624_, new_n28625_, new_n28626_,
    new_n28627_, new_n28628_, new_n28629_, new_n28630_, new_n28631_,
    new_n28632_, new_n28633_, new_n28634_, new_n28635_, new_n28636_,
    new_n28637_, new_n28638_, new_n28639_, new_n28640_, new_n28641_,
    new_n28642_, new_n28643_, new_n28644_, new_n28645_, new_n28646_,
    new_n28647_, new_n28648_, new_n28649_, new_n28650_, new_n28651_,
    new_n28652_, new_n28653_, new_n28654_, new_n28655_, new_n28656_,
    new_n28657_, new_n28658_, new_n28659_, new_n28660_, new_n28661_,
    new_n28662_, new_n28663_, new_n28664_, new_n28665_, new_n28666_,
    new_n28667_, new_n28668_, new_n28669_, new_n28670_, new_n28671_,
    new_n28672_, new_n28673_, new_n28674_, new_n28675_, new_n28676_,
    new_n28677_, new_n28678_, new_n28679_, new_n28680_, new_n28681_,
    new_n28682_, new_n28683_, new_n28684_, new_n28685_, new_n28686_,
    new_n28687_, new_n28688_, new_n28689_, new_n28690_, new_n28691_,
    new_n28692_, new_n28693_, new_n28694_, new_n28695_, new_n28696_,
    new_n28697_, new_n28698_, new_n28699_, new_n28700_, new_n28701_,
    new_n28702_, new_n28703_, new_n28704_, new_n28705_, new_n28706_,
    new_n28707_, new_n28708_, new_n28709_, new_n28710_, new_n28711_,
    new_n28712_, new_n28713_, new_n28714_, new_n28715_, new_n28716_,
    new_n28717_, new_n28718_, new_n28719_, new_n28720_, new_n28721_,
    new_n28722_, new_n28723_, new_n28724_, new_n28725_, new_n28726_,
    new_n28727_, new_n28728_, new_n28729_, new_n28730_, new_n28731_,
    new_n28732_, new_n28733_, new_n28734_, new_n28735_, new_n28736_,
    new_n28737_, new_n28738_, new_n28739_, new_n28740_, new_n28741_,
    new_n28742_, new_n28743_, new_n28744_, new_n28745_, new_n28746_,
    new_n28747_, new_n28748_, new_n28749_, new_n28750_, new_n28751_,
    new_n28752_, new_n28753_, new_n28754_, new_n28755_, new_n28756_,
    new_n28757_, new_n28758_, new_n28759_, new_n28760_, new_n28761_,
    new_n28762_, new_n28763_, new_n28764_, new_n28765_, new_n28766_,
    new_n28767_, new_n28768_, new_n28769_, new_n28770_, new_n28771_,
    new_n28772_, new_n28773_, new_n28774_, new_n28775_, new_n28776_,
    new_n28777_, new_n28778_, new_n28779_, new_n28780_, new_n28781_,
    new_n28782_, new_n28783_, new_n28784_, new_n28785_, new_n28786_,
    new_n28787_, new_n28788_, new_n28789_, new_n28790_, new_n28791_,
    new_n28792_, new_n28793_, new_n28794_, new_n28795_, new_n28796_,
    new_n28797_, new_n28798_, new_n28799_, new_n28800_, new_n28801_,
    new_n28802_, new_n28803_, new_n28804_, new_n28805_, new_n28806_,
    new_n28807_, new_n28808_, new_n28809_, new_n28810_, new_n28811_,
    new_n28812_, new_n28813_, new_n28814_, new_n28815_, new_n28816_,
    new_n28817_, new_n28818_, new_n28819_, new_n28820_, new_n28821_,
    new_n28822_, new_n28823_, new_n28824_, new_n28825_, new_n28826_,
    new_n28827_, new_n28828_, new_n28829_, new_n28830_, new_n28831_,
    new_n28832_, new_n28833_, new_n28834_, new_n28835_, new_n28836_,
    new_n28837_, new_n28838_, new_n28839_, new_n28840_, new_n28841_,
    new_n28842_, new_n28843_, new_n28844_, new_n28845_, new_n28846_,
    new_n28847_, new_n28848_, new_n28849_, new_n28850_, new_n28851_,
    new_n28852_, new_n28853_, new_n28854_, new_n28855_, new_n28856_,
    new_n28857_, new_n28858_, new_n28859_, new_n28860_, new_n28861_,
    new_n28862_, new_n28863_, new_n28864_, new_n28865_, new_n28866_,
    new_n28867_, new_n28868_, new_n28869_, new_n28870_, new_n28871_,
    new_n28872_, new_n28873_, new_n28874_, new_n28875_, new_n28876_,
    new_n28877_, new_n28878_, new_n28879_, new_n28880_, new_n28881_,
    new_n28882_, new_n28883_, new_n28884_, new_n28885_, new_n28886_,
    new_n28887_, new_n28888_, new_n28889_, new_n28890_, new_n28891_,
    new_n28892_, new_n28893_, new_n28894_, new_n28895_, new_n28896_,
    new_n28897_, new_n28898_, new_n28899_, new_n28900_, new_n28901_,
    new_n28902_, new_n28903_, new_n28904_, new_n28905_, new_n28906_,
    new_n28907_, new_n28908_, new_n28909_, new_n28910_, new_n28911_,
    new_n28912_, new_n28913_, new_n28914_, new_n28915_, new_n28916_,
    new_n28917_, new_n28918_, new_n28919_, new_n28920_, new_n28921_,
    new_n28922_, new_n28923_, new_n28924_, new_n28925_, new_n28926_,
    new_n28927_, new_n28928_, new_n28929_, new_n28930_, new_n28931_,
    new_n28932_, new_n28933_, new_n28934_, new_n28935_, new_n28936_,
    new_n28937_, new_n28938_, new_n28939_, new_n28940_, new_n28941_,
    new_n28942_, new_n28943_, new_n28944_, new_n28945_, new_n28946_,
    new_n28947_, new_n28948_, new_n28949_, new_n28950_, new_n28951_,
    new_n28952_, new_n28953_, new_n28954_, new_n28955_, new_n28956_,
    new_n28957_, new_n28958_, new_n28959_, new_n28960_, new_n28961_,
    new_n28962_, new_n28963_, new_n28964_, new_n28965_, new_n28966_,
    new_n28967_, new_n28968_, new_n28969_, new_n28970_, new_n28971_,
    new_n28972_, new_n28973_, new_n28974_, new_n28975_, new_n28976_,
    new_n28977_, new_n28978_, new_n28979_, new_n28980_, new_n28981_,
    new_n28982_, new_n28983_, new_n28984_, new_n28985_, new_n28986_,
    new_n28987_, new_n28988_, new_n28989_, new_n28990_, new_n28991_,
    new_n28992_, new_n28993_, new_n28994_, new_n28995_, new_n28996_,
    new_n28997_, new_n28998_, new_n28999_, new_n29000_, new_n29001_,
    new_n29002_, new_n29003_, new_n29004_, new_n29005_, new_n29006_,
    new_n29007_, new_n29008_, new_n29009_, new_n29010_, new_n29011_,
    new_n29012_, new_n29013_, new_n29014_, new_n29015_, new_n29016_,
    new_n29017_, new_n29018_, new_n29019_, new_n29020_, new_n29021_,
    new_n29022_, new_n29023_, new_n29024_, new_n29025_, new_n29026_,
    new_n29027_, new_n29028_, new_n29029_, new_n29030_, new_n29031_,
    new_n29032_, new_n29033_, new_n29034_, new_n29035_, new_n29036_,
    new_n29037_, new_n29038_, new_n29039_, new_n29040_, new_n29041_,
    new_n29042_, new_n29043_, new_n29044_, new_n29045_, new_n29046_,
    new_n29047_, new_n29048_, new_n29049_, new_n29050_, new_n29051_,
    new_n29052_, new_n29053_, new_n29054_, new_n29055_, new_n29056_,
    new_n29057_, new_n29058_, new_n29059_, new_n29060_, new_n29061_,
    new_n29062_, new_n29063_, new_n29064_, new_n29065_, new_n29066_,
    new_n29067_, new_n29068_, new_n29069_, new_n29070_, new_n29071_,
    new_n29072_, new_n29073_, new_n29074_, new_n29075_, new_n29076_,
    new_n29077_, new_n29078_, new_n29079_, new_n29080_, new_n29081_,
    new_n29082_, new_n29083_, new_n29084_, new_n29085_, new_n29086_,
    new_n29087_, new_n29088_, new_n29089_, new_n29090_, new_n29091_,
    new_n29092_, new_n29093_, new_n29094_, new_n29095_, new_n29096_,
    new_n29097_, new_n29098_, new_n29099_, new_n29100_, new_n29101_,
    new_n29102_, new_n29103_, new_n29104_, new_n29105_, new_n29106_,
    new_n29107_, new_n29108_, new_n29109_, new_n29110_, new_n29111_,
    new_n29112_, new_n29113_, new_n29114_, new_n29115_, new_n29116_,
    new_n29117_, new_n29118_, new_n29119_, new_n29120_, new_n29121_,
    new_n29122_, new_n29123_, new_n29124_, new_n29125_, new_n29126_,
    new_n29127_, new_n29128_, new_n29129_, new_n29130_, new_n29131_,
    new_n29132_, new_n29133_, new_n29134_, new_n29135_, new_n29136_,
    new_n29137_, new_n29138_, new_n29139_, new_n29140_, new_n29141_,
    new_n29142_, new_n29143_, new_n29144_, new_n29145_, new_n29146_,
    new_n29147_, new_n29148_, new_n29149_, new_n29150_, new_n29151_,
    new_n29152_, new_n29153_, new_n29154_, new_n29155_, new_n29156_,
    new_n29157_, new_n29158_, new_n29159_, new_n29160_, new_n29161_,
    new_n29162_, new_n29163_, new_n29164_, new_n29165_, new_n29166_,
    new_n29167_, new_n29168_, new_n29169_, new_n29170_, new_n29171_,
    new_n29172_, new_n29173_, new_n29174_, new_n29175_, new_n29176_,
    new_n29177_, new_n29178_, new_n29179_, new_n29180_, new_n29181_,
    new_n29182_, new_n29183_, new_n29184_, new_n29185_, new_n29186_,
    new_n29187_, new_n29188_, new_n29189_, new_n29190_, new_n29191_,
    new_n29192_, new_n29193_, new_n29194_, new_n29195_, new_n29196_,
    new_n29197_, new_n29198_, new_n29199_, new_n29200_, new_n29201_,
    new_n29202_, new_n29203_, new_n29204_, new_n29205_, new_n29206_,
    new_n29207_, new_n29208_, new_n29209_, new_n29210_, new_n29211_,
    new_n29212_, new_n29213_, new_n29214_, new_n29215_, new_n29216_,
    new_n29217_, new_n29218_, new_n29219_, new_n29220_, new_n29221_,
    new_n29222_, new_n29223_, new_n29224_, new_n29225_, new_n29226_,
    new_n29227_, new_n29228_, new_n29229_, new_n29230_, new_n29231_,
    new_n29232_, new_n29233_, new_n29234_, new_n29235_, new_n29236_,
    new_n29237_, new_n29238_, new_n29239_, new_n29240_, new_n29241_,
    new_n29242_, new_n29243_, new_n29244_, new_n29245_, new_n29246_,
    new_n29247_, new_n29248_, new_n29249_, new_n29250_, new_n29251_,
    new_n29252_, new_n29253_, new_n29254_, new_n29255_, new_n29256_,
    new_n29257_, new_n29258_, new_n29259_, new_n29260_, new_n29261_,
    new_n29262_, new_n29263_, new_n29264_, new_n29265_, new_n29266_,
    new_n29267_, new_n29268_, new_n29269_, new_n29270_, new_n29271_,
    new_n29272_, new_n29273_, new_n29274_, new_n29275_, new_n29276_,
    new_n29277_, new_n29278_, new_n29279_, new_n29280_, new_n29281_,
    new_n29282_, new_n29283_, new_n29284_, new_n29285_, new_n29286_,
    new_n29287_, new_n29288_, new_n29289_, new_n29290_, new_n29291_,
    new_n29292_, new_n29293_, new_n29294_, new_n29295_, new_n29296_,
    new_n29297_, new_n29298_, new_n29299_, new_n29300_, new_n29301_,
    new_n29302_, new_n29303_, new_n29304_, new_n29305_, new_n29306_,
    new_n29307_, new_n29308_, new_n29309_, new_n29310_, new_n29311_,
    new_n29312_, new_n29313_, new_n29314_, new_n29315_, new_n29316_,
    new_n29317_, new_n29318_, new_n29319_, new_n29320_, new_n29321_,
    new_n29322_, new_n29323_, new_n29324_, new_n29325_, new_n29326_,
    new_n29327_, new_n29328_, new_n29329_, new_n29330_, new_n29331_,
    new_n29332_, new_n29333_, new_n29334_, new_n29335_, new_n29336_,
    new_n29337_, new_n29338_, new_n29339_, new_n29340_, new_n29341_,
    new_n29342_, new_n29343_, new_n29344_, new_n29345_, new_n29346_,
    new_n29347_, new_n29348_, new_n29349_, new_n29350_, new_n29351_,
    new_n29352_, new_n29353_, new_n29354_, new_n29355_, new_n29356_,
    new_n29357_, new_n29358_, new_n29359_, new_n29360_, new_n29361_,
    new_n29362_, new_n29363_, new_n29364_, new_n29365_, new_n29366_,
    new_n29367_, new_n29368_, new_n29369_, new_n29370_, new_n29371_,
    new_n29372_, new_n29373_, new_n29374_, new_n29375_, new_n29376_,
    new_n29377_, new_n29378_, new_n29379_, new_n29380_, new_n29381_,
    new_n29382_, new_n29383_, new_n29384_, new_n29385_, new_n29386_,
    new_n29387_, new_n29388_, new_n29389_, new_n29390_, new_n29391_,
    new_n29392_, new_n29393_, new_n29394_, new_n29395_, new_n29396_,
    new_n29397_, new_n29398_, new_n29399_, new_n29400_, new_n29401_,
    new_n29402_, new_n29403_, new_n29404_, new_n29405_, new_n29406_,
    new_n29407_, new_n29408_, new_n29409_, new_n29410_, new_n29411_,
    new_n29412_, new_n29413_, new_n29414_, new_n29415_, new_n29416_,
    new_n29417_, new_n29418_, new_n29419_, new_n29420_, new_n29421_,
    new_n29422_, new_n29423_, new_n29424_, new_n29425_, new_n29426_,
    new_n29427_, new_n29428_, new_n29429_, new_n29430_, new_n29431_,
    new_n29432_, new_n29433_, new_n29434_, new_n29435_, new_n29436_,
    new_n29437_, new_n29438_, new_n29439_, new_n29440_, new_n29441_,
    new_n29442_, new_n29443_, new_n29444_, new_n29445_, new_n29446_,
    new_n29447_, new_n29448_, new_n29449_, new_n29450_, new_n29451_,
    new_n29452_, new_n29453_, new_n29454_, new_n29455_, new_n29456_,
    new_n29457_, new_n29458_, new_n29459_, new_n29460_, new_n29461_,
    new_n29462_, new_n29463_, new_n29464_, new_n29465_, new_n29466_,
    new_n29467_, new_n29468_, new_n29469_, new_n29470_, new_n29471_,
    new_n29472_, new_n29473_, new_n29474_, new_n29475_, new_n29476_,
    new_n29477_, new_n29478_, new_n29479_, new_n29480_, new_n29481_,
    new_n29482_, new_n29483_, new_n29484_, new_n29485_, new_n29486_,
    new_n29487_, new_n29488_, new_n29489_, new_n29490_, new_n29491_,
    new_n29492_, new_n29493_, new_n29494_, new_n29495_, new_n29496_,
    new_n29497_, new_n29498_, new_n29499_, new_n29500_, new_n29501_,
    new_n29502_, new_n29503_, new_n29504_, new_n29505_, new_n29506_,
    new_n29507_, new_n29508_, new_n29509_, new_n29510_, new_n29511_,
    new_n29512_, new_n29513_, new_n29514_, new_n29515_, new_n29516_,
    new_n29517_, new_n29518_, new_n29519_, new_n29520_, new_n29521_,
    new_n29522_, new_n29523_, new_n29524_, new_n29525_, new_n29526_,
    new_n29527_, new_n29528_, new_n29529_, new_n29530_, new_n29531_,
    new_n29532_, new_n29533_, new_n29534_, new_n29535_, new_n29536_,
    new_n29537_, new_n29538_, new_n29539_, new_n29540_, new_n29541_,
    new_n29542_, new_n29543_, new_n29544_, new_n29545_, new_n29546_,
    new_n29547_, new_n29548_, new_n29549_, new_n29550_, new_n29551_,
    new_n29552_, new_n29553_, new_n29554_, new_n29555_, new_n29556_,
    new_n29557_, new_n29558_, new_n29559_, new_n29560_, new_n29561_,
    new_n29562_, new_n29563_, new_n29564_, new_n29565_, new_n29566_,
    new_n29567_, new_n29568_, new_n29569_, new_n29570_, new_n29571_,
    new_n29572_, new_n29573_, new_n29574_, new_n29575_, new_n29576_,
    new_n29577_, new_n29578_, new_n29579_, new_n29580_, new_n29581_,
    new_n29582_, new_n29583_, new_n29584_, new_n29585_, new_n29586_,
    new_n29587_, new_n29588_, new_n29589_, new_n29590_, new_n29591_,
    new_n29592_, new_n29593_, new_n29594_, new_n29595_, new_n29596_,
    new_n29597_, new_n29598_, new_n29599_, new_n29600_, new_n29601_,
    new_n29602_, new_n29603_, new_n29604_, new_n29605_, new_n29606_,
    new_n29607_, new_n29608_, new_n29609_, new_n29610_, new_n29611_,
    new_n29612_, new_n29613_, new_n29614_, new_n29615_, new_n29616_,
    new_n29617_, new_n29618_, new_n29619_, new_n29620_, new_n29621_,
    new_n29622_, new_n29623_, new_n29624_, new_n29625_, new_n29626_,
    new_n29627_, new_n29628_, new_n29629_, new_n29630_, new_n29631_,
    new_n29632_, new_n29633_, new_n29634_, new_n29635_, new_n29636_,
    new_n29637_, new_n29638_, new_n29639_, new_n29640_, new_n29641_,
    new_n29642_, new_n29643_, new_n29644_, new_n29645_, new_n29646_,
    new_n29647_, new_n29648_, new_n29649_, new_n29650_, new_n29651_,
    new_n29652_, new_n29653_, new_n29654_, new_n29655_, new_n29656_,
    new_n29657_, new_n29658_, new_n29659_, new_n29660_, new_n29661_,
    new_n29662_, new_n29663_, new_n29664_, new_n29665_, new_n29666_,
    new_n29667_, new_n29668_, new_n29669_, new_n29670_, new_n29671_,
    new_n29672_, new_n29673_, new_n29674_, new_n29675_, new_n29676_,
    new_n29677_, new_n29678_, new_n29679_, new_n29680_, new_n29681_,
    new_n29682_, new_n29683_, new_n29684_, new_n29685_, new_n29686_,
    new_n29687_, new_n29688_, new_n29689_, new_n29690_, new_n29691_,
    new_n29692_, new_n29693_, new_n29694_, new_n29695_, new_n29696_,
    new_n29697_, new_n29698_, new_n29699_, new_n29700_, new_n29701_,
    new_n29702_, new_n29703_, new_n29704_, new_n29705_, new_n29706_,
    new_n29707_, new_n29708_, new_n29709_, new_n29710_, new_n29711_,
    new_n29712_, new_n29713_, new_n29714_, new_n29715_, new_n29716_,
    new_n29717_, new_n29718_, new_n29719_, new_n29720_, new_n29721_,
    new_n29722_, new_n29723_, new_n29724_, new_n29725_, new_n29726_,
    new_n29727_, new_n29728_, new_n29729_, new_n29730_, new_n29731_,
    new_n29732_, new_n29733_, new_n29734_, new_n29735_, new_n29736_,
    new_n29737_, new_n29738_, new_n29739_, new_n29740_, new_n29741_,
    new_n29742_, new_n29743_, new_n29744_, new_n29745_, new_n29746_,
    new_n29747_, new_n29748_, new_n29749_, new_n29750_, new_n29751_,
    new_n29752_, new_n29753_, new_n29754_, new_n29755_, new_n29756_,
    new_n29757_, new_n29758_, new_n29759_, new_n29760_, new_n29761_,
    new_n29762_, new_n29763_, new_n29764_, new_n29765_, new_n29766_,
    new_n29767_, new_n29768_, new_n29769_, new_n29770_, new_n29771_,
    new_n29772_, new_n29773_, new_n29774_, new_n29775_, new_n29776_,
    new_n29777_, new_n29778_, new_n29779_, new_n29780_, new_n29781_,
    new_n29782_, new_n29783_, new_n29784_, new_n29785_, new_n29786_,
    new_n29787_, new_n29788_, new_n29789_, new_n29790_, new_n29791_,
    new_n29792_, new_n29793_, new_n29794_, new_n29795_, new_n29796_,
    new_n29797_, new_n29798_, new_n29799_, new_n29800_, new_n29801_,
    new_n29802_, new_n29803_, new_n29804_, new_n29805_, new_n29806_,
    new_n29807_, new_n29808_, new_n29809_, new_n29810_, new_n29811_,
    new_n29812_, new_n29813_, new_n29814_, new_n29815_, new_n29816_,
    new_n29817_, new_n29818_, new_n29819_, new_n29820_, new_n29821_,
    new_n29822_, new_n29823_, new_n29824_, new_n29825_, new_n29826_,
    new_n29827_, new_n29828_, new_n29829_, new_n29830_, new_n29831_,
    new_n29832_, new_n29833_, new_n29834_, new_n29835_, new_n29836_,
    new_n29837_, new_n29838_, new_n29839_, new_n29840_, new_n29841_,
    new_n29842_, new_n29843_, new_n29844_, new_n29845_, new_n29846_,
    new_n29847_, new_n29848_, new_n29849_, new_n29850_, new_n29851_,
    new_n29852_, new_n29853_, new_n29854_, new_n29855_, new_n29856_,
    new_n29857_, new_n29858_, new_n29859_, new_n29860_, new_n29861_,
    new_n29862_, new_n29863_, new_n29864_, new_n29865_, new_n29866_,
    new_n29867_, new_n29868_, new_n29869_, new_n29870_, new_n29871_,
    new_n29872_, new_n29873_, new_n29874_, new_n29875_, new_n29876_,
    new_n29877_, new_n29878_, new_n29879_, new_n29880_, new_n29881_,
    new_n29882_, new_n29883_, new_n29884_, new_n29885_, new_n29886_,
    new_n29887_, new_n29888_, new_n29889_, new_n29890_, new_n29891_,
    new_n29892_, new_n29893_, new_n29894_, new_n29895_, new_n29896_,
    new_n29897_, new_n29898_, new_n29899_, new_n29900_, new_n29901_,
    new_n29902_, new_n29903_, new_n29904_, new_n29905_, new_n29906_,
    new_n29907_, new_n29908_, new_n29909_, new_n29910_, new_n29911_,
    new_n29912_, new_n29913_, new_n29914_, new_n29915_, new_n29916_,
    new_n29917_, new_n29918_, new_n29919_, new_n29920_, new_n29921_,
    new_n29922_, new_n29923_, new_n29924_, new_n29925_, new_n29926_,
    new_n29927_, new_n29928_, new_n29929_, new_n29930_, new_n29931_,
    new_n29932_, new_n29933_, new_n29934_, new_n29935_, new_n29936_,
    new_n29937_, new_n29938_, new_n29939_, new_n29940_, new_n29941_,
    new_n29942_, new_n29943_, new_n29944_, new_n29945_, new_n29946_,
    new_n29947_, new_n29948_, new_n29949_, new_n29950_, new_n29951_,
    new_n29952_, new_n29953_, new_n29954_, new_n29955_, new_n29956_,
    new_n29957_, new_n29958_, new_n29959_, new_n29960_, new_n29961_,
    new_n29962_, new_n29963_, new_n29964_, new_n29965_, new_n29966_,
    new_n29967_, new_n29968_, new_n29969_, new_n29970_, new_n29971_,
    new_n29972_, new_n29973_, new_n29974_, new_n29975_, new_n29976_,
    new_n29977_, new_n29978_, new_n29979_, new_n29980_, new_n29981_,
    new_n29982_, new_n29983_, new_n29984_, new_n29985_, new_n29986_,
    new_n29987_, new_n29988_, new_n29989_, new_n29990_, new_n29991_,
    new_n29992_, new_n29993_, new_n29994_, new_n29995_, new_n29996_,
    new_n29997_, new_n29998_, new_n29999_, new_n30000_, new_n30001_,
    new_n30002_, new_n30003_, new_n30004_, new_n30005_, new_n30006_,
    new_n30007_, new_n30008_, new_n30009_, new_n30010_, new_n30011_,
    new_n30012_, new_n30013_, new_n30014_, new_n30015_, new_n30016_,
    new_n30017_, new_n30018_, new_n30019_, new_n30020_, new_n30021_,
    new_n30022_, new_n30023_, new_n30024_, new_n30025_, new_n30026_,
    new_n30027_, new_n30028_, new_n30029_, new_n30030_, new_n30031_,
    new_n30032_, new_n30033_, new_n30034_, new_n30035_, new_n30036_,
    new_n30037_, new_n30038_, new_n30039_, new_n30040_, new_n30041_,
    new_n30042_, new_n30043_, new_n30044_, new_n30045_, new_n30046_,
    new_n30047_, new_n30048_, new_n30049_, new_n30050_, new_n30051_,
    new_n30052_, new_n30053_, new_n30054_, new_n30055_, new_n30056_,
    new_n30057_, new_n30058_, new_n30059_, new_n30060_, new_n30061_,
    new_n30062_, new_n30063_, new_n30064_, new_n30065_, new_n30066_,
    new_n30067_, new_n30068_, new_n30069_, new_n30070_, new_n30071_,
    new_n30072_, new_n30073_, new_n30074_, new_n30075_, new_n30076_,
    new_n30077_, new_n30078_, new_n30079_, new_n30080_, new_n30081_,
    new_n30082_, new_n30083_, new_n30084_, new_n30085_, new_n30086_,
    new_n30087_, new_n30088_, new_n30089_, new_n30090_, new_n30091_,
    new_n30092_, new_n30093_, new_n30094_, new_n30095_, new_n30096_,
    new_n30097_, new_n30098_, new_n30099_, new_n30100_, new_n30101_,
    new_n30102_, new_n30103_, new_n30104_, new_n30105_, new_n30106_,
    new_n30107_, new_n30108_, new_n30109_, new_n30110_, new_n30111_,
    new_n30112_, new_n30113_, new_n30114_, new_n30115_, new_n30116_,
    new_n30117_, new_n30118_, new_n30119_, new_n30120_, new_n30121_,
    new_n30122_, new_n30123_, new_n30124_, new_n30125_, new_n30126_,
    new_n30127_, new_n30128_, new_n30129_, new_n30130_, new_n30131_,
    new_n30132_, new_n30133_, new_n30134_, new_n30135_, new_n30136_,
    new_n30137_, new_n30138_, new_n30139_, new_n30140_, new_n30141_,
    new_n30142_, new_n30143_, new_n30144_, new_n30145_, new_n30146_,
    new_n30147_, new_n30148_, new_n30149_, new_n30150_, new_n30151_,
    new_n30152_, new_n30153_, new_n30154_, new_n30155_, new_n30156_,
    new_n30157_, new_n30158_, new_n30159_, new_n30160_, new_n30161_,
    new_n30162_, new_n30163_, new_n30164_, new_n30165_, new_n30166_,
    new_n30167_, new_n30168_, new_n30169_, new_n30170_, new_n30171_,
    new_n30172_, new_n30173_, new_n30174_, new_n30175_, new_n30176_,
    new_n30177_, new_n30178_, new_n30179_, new_n30180_, new_n30181_,
    new_n30182_, new_n30183_, new_n30184_, new_n30185_, new_n30186_,
    new_n30187_, new_n30188_, new_n30189_, new_n30190_, new_n30191_,
    new_n30192_, new_n30193_, new_n30194_, new_n30195_, new_n30196_,
    new_n30197_, new_n30198_, new_n30199_, new_n30200_, new_n30201_,
    new_n30202_, new_n30203_, new_n30204_, new_n30205_, new_n30206_,
    new_n30207_, new_n30208_, new_n30209_, new_n30210_, new_n30211_,
    new_n30212_, new_n30213_, new_n30214_, new_n30215_, new_n30216_,
    new_n30217_, new_n30218_, new_n30219_, new_n30220_, new_n30221_,
    new_n30222_, new_n30223_, new_n30224_, new_n30225_, new_n30226_,
    new_n30227_, new_n30228_, new_n30229_, new_n30230_, new_n30231_,
    new_n30232_, new_n30233_, new_n30234_, new_n30235_, new_n30236_,
    new_n30237_, new_n30238_, new_n30239_, new_n30240_, new_n30241_,
    new_n30242_, new_n30243_, new_n30244_, new_n30245_, new_n30246_,
    new_n30247_, new_n30248_, new_n30249_, new_n30250_, new_n30251_,
    new_n30252_, new_n30253_, new_n30254_, new_n30255_, new_n30256_,
    new_n30257_, new_n30258_, new_n30259_, new_n30260_, new_n30261_,
    new_n30262_, new_n30263_, new_n30264_, new_n30265_, new_n30266_,
    new_n30267_, new_n30268_, new_n30269_, new_n30270_, new_n30271_,
    new_n30272_, new_n30273_, new_n30274_, new_n30275_, new_n30276_,
    new_n30277_, new_n30278_, new_n30279_, new_n30280_, new_n30281_,
    new_n30282_, new_n30283_, new_n30284_, new_n30285_, new_n30286_,
    new_n30287_, new_n30288_, new_n30289_, new_n30290_, new_n30291_,
    new_n30292_, new_n30293_, new_n30294_, new_n30295_, new_n30296_,
    new_n30297_, new_n30298_, new_n30299_, new_n30300_, new_n30301_,
    new_n30302_, new_n30303_, new_n30304_, new_n30305_, new_n30306_,
    new_n30307_, new_n30308_, new_n30309_, new_n30310_, new_n30311_,
    new_n30312_, new_n30313_, new_n30314_, new_n30315_, new_n30316_,
    new_n30317_, new_n30318_, new_n30319_, new_n30320_, new_n30321_,
    new_n30322_, new_n30323_, new_n30324_, new_n30325_, new_n30326_,
    new_n30327_, new_n30328_, new_n30329_, new_n30330_, new_n30331_,
    new_n30332_, new_n30333_, new_n30334_, new_n30335_, new_n30336_,
    new_n30337_, new_n30338_, new_n30339_, new_n30340_, new_n30341_,
    new_n30342_, new_n30343_, new_n30344_, new_n30345_, new_n30346_,
    new_n30347_, new_n30348_, new_n30349_, new_n30350_, new_n30351_,
    new_n30352_, new_n30353_, new_n30354_, new_n30355_, new_n30356_,
    new_n30357_, new_n30358_, new_n30359_, new_n30360_, new_n30361_,
    new_n30362_, new_n30363_, new_n30364_, new_n30365_, new_n30366_,
    new_n30367_, new_n30368_, new_n30369_, new_n30370_, new_n30371_,
    new_n30372_, new_n30373_, new_n30374_, new_n30375_, new_n30376_,
    new_n30377_, new_n30378_, new_n30379_, new_n30380_, new_n30381_,
    new_n30382_, new_n30383_, new_n30384_, new_n30385_, new_n30386_,
    new_n30387_, new_n30388_, new_n30389_, new_n30390_, new_n30391_,
    new_n30392_, new_n30393_, new_n30394_, new_n30395_, new_n30396_,
    new_n30397_, new_n30398_, new_n30399_, new_n30400_, new_n30401_,
    new_n30402_, new_n30403_, new_n30404_, new_n30405_, new_n30406_,
    new_n30407_, new_n30408_, new_n30409_, new_n30410_, new_n30411_,
    new_n30412_, new_n30413_, new_n30414_, new_n30415_, new_n30416_,
    new_n30417_, new_n30418_, new_n30419_, new_n30420_, new_n30421_,
    new_n30422_, new_n30423_, new_n30424_, new_n30425_, new_n30426_,
    new_n30427_, new_n30428_, new_n30429_, new_n30430_, new_n30431_,
    new_n30432_, new_n30433_, new_n30434_, new_n30435_, new_n30436_,
    new_n30437_, new_n30438_, new_n30439_, new_n30440_, new_n30441_,
    new_n30442_, new_n30443_, new_n30444_, new_n30445_, new_n30446_,
    new_n30447_, new_n30448_, new_n30449_, new_n30450_, new_n30451_,
    new_n30452_, new_n30453_, new_n30454_, new_n30455_, new_n30456_,
    new_n30457_, new_n30458_, new_n30459_, new_n30460_, new_n30461_,
    new_n30462_, new_n30463_, new_n30464_, new_n30465_, new_n30466_,
    new_n30467_, new_n30468_, new_n30469_, new_n30470_, new_n30471_,
    new_n30472_, new_n30473_, new_n30474_, new_n30475_, new_n30476_,
    new_n30477_, new_n30478_, new_n30479_, new_n30480_, new_n30481_,
    new_n30482_, new_n30483_, new_n30484_, new_n30485_, new_n30486_,
    new_n30487_, new_n30488_, new_n30489_, new_n30490_, new_n30491_,
    new_n30492_, new_n30493_, new_n30494_, new_n30495_, new_n30496_,
    new_n30497_, new_n30498_, new_n30499_, new_n30500_, new_n30501_,
    new_n30502_, new_n30503_, new_n30504_, new_n30505_, new_n30506_,
    new_n30507_, new_n30508_, new_n30509_, new_n30510_, new_n30511_,
    new_n30512_, new_n30513_, new_n30514_, new_n30515_, new_n30516_,
    new_n30517_, new_n30518_, new_n30519_, new_n30520_, new_n30521_,
    new_n30522_, new_n30523_, new_n30524_, new_n30525_, new_n30526_,
    new_n30527_, new_n30528_, new_n30529_, new_n30530_, new_n30531_,
    new_n30532_, new_n30533_, new_n30534_, new_n30535_, new_n30536_,
    new_n30537_, new_n30538_, new_n30539_, new_n30540_, new_n30541_,
    new_n30542_, new_n30543_, new_n30544_, new_n30545_, new_n30546_,
    new_n30547_, new_n30548_, new_n30549_, new_n30550_, new_n30551_,
    new_n30552_, new_n30553_, new_n30554_, new_n30555_, new_n30556_,
    new_n30557_, new_n30558_, new_n30559_, new_n30560_, new_n30561_,
    new_n30562_, new_n30563_, new_n30564_, new_n30565_, new_n30566_,
    new_n30567_, new_n30568_, new_n30569_, new_n30570_, new_n30571_,
    new_n30572_, new_n30573_, new_n30574_, new_n30575_, new_n30576_,
    new_n30577_, new_n30578_, new_n30579_, new_n30580_, new_n30581_,
    new_n30582_, new_n30583_, new_n30584_, new_n30585_, new_n30586_,
    new_n30587_, new_n30588_, new_n30589_, new_n30590_, new_n30591_,
    new_n30592_, new_n30593_, new_n30594_, new_n30595_, new_n30596_,
    new_n30597_, new_n30598_, new_n30599_, new_n30600_, new_n30601_,
    new_n30602_, new_n30603_, new_n30604_, new_n30605_, new_n30606_,
    new_n30607_, new_n30608_, new_n30609_, new_n30610_, new_n30611_,
    new_n30612_, new_n30613_, new_n30614_, new_n30615_, new_n30616_,
    new_n30617_, new_n30618_, new_n30619_, new_n30620_, new_n30621_,
    new_n30622_, new_n30623_, new_n30624_, new_n30625_, new_n30626_,
    new_n30627_, new_n30628_, new_n30629_, new_n30630_, new_n30631_,
    new_n30632_, new_n30633_, new_n30634_, new_n30635_, new_n30636_,
    new_n30637_, new_n30638_, new_n30639_, new_n30640_, new_n30641_,
    new_n30642_, new_n30643_, new_n30644_, new_n30645_, new_n30646_,
    new_n30647_, new_n30648_, new_n30649_, new_n30650_, new_n30651_,
    new_n30652_, new_n30653_, new_n30654_, new_n30655_, new_n30656_,
    new_n30657_, new_n30658_, new_n30659_, new_n30660_, new_n30661_,
    new_n30662_, new_n30663_, new_n30664_, new_n30665_, new_n30666_,
    new_n30667_, new_n30668_, new_n30669_, new_n30670_, new_n30671_,
    new_n30672_, new_n30673_, new_n30674_, new_n30675_, new_n30676_,
    new_n30677_, new_n30678_, new_n30679_, new_n30680_, new_n30681_,
    new_n30682_, new_n30683_, new_n30684_, new_n30685_, new_n30686_,
    new_n30687_, new_n30688_, new_n30689_, new_n30690_, new_n30691_,
    new_n30692_, new_n30693_, new_n30694_, new_n30695_, new_n30696_,
    new_n30697_, new_n30698_, new_n30699_, new_n30700_, new_n30701_,
    new_n30702_, new_n30703_, new_n30704_, new_n30705_, new_n30706_,
    new_n30707_, new_n30708_, new_n30709_, new_n30710_, new_n30711_,
    new_n30712_, new_n30713_, new_n30714_, new_n30715_, new_n30716_,
    new_n30717_, new_n30718_, new_n30719_, new_n30720_, new_n30721_,
    new_n30722_, new_n30723_, new_n30724_, new_n30725_, new_n30726_,
    new_n30727_, new_n30728_, new_n30729_, new_n30730_, new_n30731_,
    new_n30732_, new_n30733_, new_n30734_, new_n30735_, new_n30736_,
    new_n30737_, new_n30738_, new_n30739_, new_n30740_, new_n30741_,
    new_n30742_, new_n30743_, new_n30744_, new_n30745_, new_n30746_,
    new_n30747_, new_n30748_, new_n30749_, new_n30750_, new_n30751_,
    new_n30752_, new_n30753_, new_n30754_, new_n30755_, new_n30756_,
    new_n30757_, new_n30758_, new_n30759_, new_n30760_, new_n30761_,
    new_n30762_, new_n30763_, new_n30764_, new_n30765_, new_n30766_,
    new_n30767_, new_n30768_, new_n30769_, new_n30770_, new_n30771_,
    new_n30772_, new_n30773_, new_n30774_, new_n30775_, new_n30776_,
    new_n30777_, new_n30778_, new_n30779_, new_n30780_, new_n30781_,
    new_n30782_, new_n30783_, new_n30784_, new_n30785_, new_n30786_,
    new_n30787_, new_n30788_, new_n30789_, new_n30790_, new_n30791_,
    new_n30792_, new_n30793_, new_n30794_, new_n30795_, new_n30796_,
    new_n30797_, new_n30798_, new_n30799_, new_n30800_, new_n30801_,
    new_n30802_, new_n30803_, new_n30804_, new_n30805_, new_n30806_,
    new_n30807_, new_n30808_, new_n30809_, new_n30810_, new_n30811_,
    new_n30812_, new_n30813_, new_n30814_, new_n30815_, new_n30816_,
    new_n30817_, new_n30818_, new_n30819_, new_n30820_, new_n30821_,
    new_n30822_, new_n30823_, new_n30824_, new_n30825_, new_n30826_,
    new_n30827_, new_n30828_, new_n30829_, new_n30830_, new_n30831_,
    new_n30832_, new_n30833_, new_n30834_, new_n30835_, new_n30836_,
    new_n30837_, new_n30838_, new_n30839_, new_n30840_, new_n30841_,
    new_n30842_, new_n30843_, new_n30844_, new_n30845_, new_n30846_,
    new_n30847_, new_n30848_, new_n30849_, new_n30850_, new_n30851_,
    new_n30852_, new_n30853_, new_n30854_, new_n30855_, new_n30856_,
    new_n30857_, new_n30858_, new_n30859_, new_n30860_, new_n30861_,
    new_n30862_, new_n30863_, new_n30864_, new_n30865_, new_n30866_,
    new_n30867_, new_n30868_, new_n30869_, new_n30870_, new_n30871_,
    new_n30872_, new_n30873_, new_n30874_, new_n30875_, new_n30876_,
    new_n30877_, new_n30878_, new_n30879_, new_n30880_, new_n30881_,
    new_n30882_, new_n30883_, new_n30884_, new_n30885_, new_n30886_,
    new_n30887_, new_n30888_, new_n30889_, new_n30890_, new_n30891_,
    new_n30892_, new_n30893_, new_n30894_, new_n30895_, new_n30896_,
    new_n30897_, new_n30898_, new_n30899_, new_n30900_, new_n30901_,
    new_n30902_, new_n30903_, new_n30904_, new_n30905_, new_n30906_,
    new_n30907_, new_n30908_, new_n30909_, new_n30910_, new_n30911_,
    new_n30912_, new_n30913_, new_n30914_, new_n30915_, new_n30916_,
    new_n30917_, new_n30918_, new_n30919_, new_n30920_, new_n30921_,
    new_n30922_, new_n30923_, new_n30924_, new_n30925_, new_n30926_,
    new_n30927_, new_n30928_, new_n30929_, new_n30930_, new_n30931_,
    new_n30932_, new_n30933_, new_n30934_, new_n30935_, new_n30936_,
    new_n30937_, new_n30938_, new_n30939_, new_n30940_, new_n30941_,
    new_n30942_, new_n30943_, new_n30944_, new_n30945_, new_n30946_,
    new_n30947_, new_n30948_, new_n30949_, new_n30950_, new_n30951_,
    new_n30952_, new_n30953_, new_n30954_, new_n30955_, new_n30956_,
    new_n30957_, new_n30958_, new_n30959_, new_n30960_, new_n30961_,
    new_n30962_, new_n30963_, new_n30964_, new_n30965_, new_n30966_,
    new_n30967_, new_n30968_, new_n30969_, new_n30970_, new_n30971_,
    new_n30972_, new_n30973_, new_n30974_, new_n30975_, new_n30976_,
    new_n30977_, new_n30978_, new_n30979_, new_n30980_, new_n30981_,
    new_n30982_, new_n30983_, new_n30984_, new_n30985_, new_n30986_,
    new_n30987_, new_n30988_, new_n30989_, new_n30990_, new_n30991_,
    new_n30992_, new_n30993_, new_n30994_, new_n30995_, new_n30996_,
    new_n30997_, new_n30998_, new_n30999_, new_n31000_, new_n31001_,
    new_n31002_, new_n31003_, new_n31004_, new_n31005_, new_n31006_,
    new_n31007_, new_n31008_, new_n31009_, new_n31010_, new_n31011_,
    new_n31012_, new_n31013_, new_n31014_, new_n31015_, new_n31016_,
    new_n31017_, new_n31018_, new_n31019_, new_n31020_, new_n31021_,
    new_n31022_, new_n31023_, new_n31024_, new_n31025_, new_n31026_,
    new_n31027_, new_n31028_, new_n31029_, new_n31030_, new_n31031_,
    new_n31032_, new_n31033_, new_n31034_, new_n31035_, new_n31036_,
    new_n31037_, new_n31038_, new_n31039_, new_n31040_, new_n31041_,
    new_n31042_, new_n31043_, new_n31044_, new_n31045_, new_n31046_,
    new_n31047_, new_n31048_, new_n31049_, new_n31050_, new_n31051_,
    new_n31052_, new_n31053_, new_n31054_, new_n31055_, new_n31056_,
    new_n31057_, new_n31058_, new_n31059_, new_n31060_, new_n31061_,
    new_n31062_, new_n31063_, new_n31064_, new_n31065_, new_n31066_,
    new_n31067_, new_n31068_, new_n31069_, new_n31070_, new_n31071_,
    new_n31072_, new_n31073_, new_n31074_, new_n31075_, new_n31076_,
    new_n31077_, new_n31078_, new_n31079_, new_n31080_, new_n31081_,
    new_n31082_, new_n31083_, new_n31084_, new_n31085_, new_n31086_,
    new_n31087_, new_n31088_, new_n31089_, new_n31090_, new_n31091_,
    new_n31092_, new_n31093_, new_n31094_, new_n31095_, new_n31096_,
    new_n31097_, new_n31098_, new_n31099_, new_n31100_, new_n31101_,
    new_n31102_, new_n31103_, new_n31104_, new_n31105_, new_n31106_,
    new_n31107_, new_n31108_, new_n31109_, new_n31110_, new_n31111_,
    new_n31112_, new_n31113_, new_n31114_, new_n31115_, new_n31116_,
    new_n31117_, new_n31118_, new_n31119_, new_n31120_, new_n31121_,
    new_n31122_, new_n31123_, new_n31124_, new_n31125_, new_n31126_,
    new_n31127_, new_n31128_, new_n31129_, new_n31130_, new_n31131_,
    new_n31132_, new_n31133_, new_n31134_, new_n31135_, new_n31136_,
    new_n31137_, new_n31138_, new_n31139_, new_n31140_, new_n31141_,
    new_n31142_, new_n31143_, new_n31144_, new_n31145_, new_n31146_,
    new_n31147_, new_n31148_, new_n31149_, new_n31150_, new_n31151_,
    new_n31152_, new_n31153_, new_n31154_, new_n31155_, new_n31156_,
    new_n31157_, new_n31158_, new_n31159_, new_n31160_, new_n31161_,
    new_n31162_, new_n31163_, new_n31164_, new_n31165_, new_n31166_,
    new_n31167_, new_n31168_, new_n31169_, new_n31170_, new_n31171_,
    new_n31172_, new_n31173_, new_n31174_, new_n31175_, new_n31176_,
    new_n31177_, new_n31178_, new_n31179_, new_n31180_, new_n31181_,
    new_n31182_, new_n31183_, new_n31184_, new_n31185_, new_n31186_,
    new_n31187_, new_n31188_, new_n31189_, new_n31190_, new_n31191_,
    new_n31192_, new_n31193_, new_n31194_, new_n31195_, new_n31196_,
    new_n31197_, new_n31198_, new_n31199_, new_n31200_, new_n31201_,
    new_n31202_, new_n31203_, new_n31204_, new_n31205_, new_n31206_,
    new_n31207_, new_n31208_, new_n31209_, new_n31210_, new_n31211_,
    new_n31212_, new_n31213_, new_n31214_, new_n31215_, new_n31216_,
    new_n31217_, new_n31218_, new_n31219_, new_n31220_, new_n31221_,
    new_n31222_, new_n31223_, new_n31224_, new_n31225_, new_n31226_,
    new_n31227_, new_n31228_, new_n31229_, new_n31230_, new_n31231_,
    new_n31232_, new_n31233_, new_n31234_, new_n31235_, new_n31236_,
    new_n31237_, new_n31238_, new_n31239_, new_n31240_, new_n31241_,
    new_n31242_, new_n31243_, new_n31244_, new_n31245_, new_n31246_,
    new_n31247_, new_n31248_, new_n31249_, new_n31250_, new_n31251_,
    new_n31252_, new_n31253_, new_n31254_, new_n31255_, new_n31256_,
    new_n31257_, new_n31258_, new_n31259_, new_n31260_, new_n31261_,
    new_n31262_, new_n31263_, new_n31264_, new_n31265_, new_n31266_,
    new_n31267_, new_n31268_, new_n31269_, new_n31270_, new_n31271_,
    new_n31272_, new_n31273_, new_n31274_, new_n31275_, new_n31276_,
    new_n31277_, new_n31278_, new_n31279_, new_n31280_, new_n31281_,
    new_n31282_, new_n31283_, new_n31284_, new_n31285_, new_n31286_,
    new_n31287_, new_n31288_, new_n31289_, new_n31290_, new_n31291_,
    new_n31292_, new_n31293_, new_n31294_, new_n31295_, new_n31296_,
    new_n31297_, new_n31298_, new_n31299_, new_n31300_, new_n31301_,
    new_n31302_, new_n31303_, new_n31304_, new_n31305_, new_n31306_,
    new_n31307_, new_n31308_, new_n31309_, new_n31310_, new_n31311_,
    new_n31312_, new_n31313_, new_n31314_, new_n31315_, new_n31316_,
    new_n31317_, new_n31318_, new_n31319_, new_n31320_, new_n31321_,
    new_n31322_, new_n31323_, new_n31324_, new_n31325_, new_n31326_,
    new_n31327_, new_n31328_, new_n31329_, new_n31330_, new_n31331_,
    new_n31332_, new_n31333_, new_n31334_, new_n31335_, new_n31336_,
    new_n31337_, new_n31338_, new_n31339_, new_n31340_, new_n31341_,
    new_n31342_, new_n31343_, new_n31344_, new_n31345_, new_n31346_,
    new_n31347_, new_n31348_, new_n31349_, new_n31350_, new_n31351_,
    new_n31352_, new_n31353_, new_n31354_, new_n31355_, new_n31356_,
    new_n31357_, new_n31358_, new_n31359_, new_n31360_, new_n31361_,
    new_n31362_, new_n31363_, new_n31364_, new_n31365_, new_n31366_,
    new_n31367_, new_n31368_, new_n31369_, new_n31370_, new_n31371_,
    new_n31372_, new_n31373_, new_n31374_, new_n31375_, new_n31376_,
    new_n31377_, new_n31378_, new_n31379_, new_n31380_, new_n31381_,
    new_n31382_, new_n31383_, new_n31384_, new_n31385_, new_n31386_,
    new_n31387_, new_n31388_, new_n31389_, new_n31390_, new_n31391_,
    new_n31392_, new_n31393_, new_n31394_, new_n31395_, new_n31396_,
    new_n31397_, new_n31398_, new_n31399_, new_n31400_, new_n31401_,
    new_n31402_, new_n31403_, new_n31404_, new_n31405_, new_n31406_,
    new_n31407_, new_n31408_, new_n31409_, new_n31410_, new_n31411_,
    new_n31412_, new_n31413_, new_n31414_, new_n31415_, new_n31416_,
    new_n31417_, new_n31418_, new_n31419_, new_n31420_, new_n31421_,
    new_n31422_, new_n31423_, new_n31424_, new_n31425_, new_n31426_,
    new_n31427_, new_n31428_, new_n31429_, new_n31430_, new_n31431_,
    new_n31432_, new_n31433_, new_n31434_, new_n31435_, new_n31436_,
    new_n31437_, new_n31438_, new_n31439_, new_n31440_, new_n31441_,
    new_n31442_, new_n31443_, new_n31444_, new_n31445_, new_n31446_,
    new_n31447_, new_n31448_, new_n31449_, new_n31450_, new_n31451_,
    new_n31452_, new_n31453_, new_n31454_, new_n31455_, new_n31456_,
    new_n31457_, new_n31458_, new_n31459_, new_n31460_, new_n31461_,
    new_n31462_, new_n31463_, new_n31464_, new_n31465_, new_n31466_,
    new_n31467_, new_n31468_, new_n31469_, new_n31470_, new_n31471_,
    new_n31472_, new_n31473_, new_n31474_, new_n31475_, new_n31476_,
    new_n31477_, new_n31478_, new_n31479_, new_n31480_, new_n31481_,
    new_n31482_, new_n31483_, new_n31484_, new_n31485_, new_n31486_,
    new_n31487_, new_n31488_, new_n31489_, new_n31490_, new_n31491_,
    new_n31492_, new_n31493_, new_n31494_, new_n31495_, new_n31496_,
    new_n31497_, new_n31498_, new_n31499_, new_n31500_, new_n31501_,
    new_n31502_, new_n31503_, new_n31504_, new_n31505_, new_n31506_,
    new_n31507_, new_n31508_, new_n31509_, new_n31510_, new_n31511_,
    new_n31512_, new_n31513_, new_n31514_, new_n31515_, new_n31516_,
    new_n31517_, new_n31518_, new_n31519_, new_n31520_, new_n31521_,
    new_n31522_, new_n31523_, new_n31524_, new_n31525_, new_n31526_,
    new_n31527_, new_n31528_, new_n31529_, new_n31530_, new_n31531_,
    new_n31532_, new_n31533_, new_n31534_, new_n31535_, new_n31536_,
    new_n31537_, new_n31538_, new_n31539_, new_n31540_, new_n31541_,
    new_n31542_, new_n31543_, new_n31544_, new_n31545_, new_n31546_,
    new_n31547_, new_n31548_, new_n31549_, new_n31550_, new_n31551_,
    new_n31552_, new_n31553_, new_n31554_, new_n31555_, new_n31556_,
    new_n31557_, new_n31558_, new_n31559_, new_n31560_, new_n31561_,
    new_n31562_, new_n31563_, new_n31564_, new_n31565_, new_n31566_,
    new_n31567_, new_n31568_, new_n31569_, new_n31570_, new_n31571_,
    new_n31572_, new_n31573_, new_n31574_, new_n31575_, new_n31576_,
    new_n31577_, new_n31578_, new_n31579_, new_n31580_, new_n31581_,
    new_n31582_, new_n31583_, new_n31584_, new_n31585_, new_n31586_,
    new_n31587_, new_n31588_, new_n31589_, new_n31590_, new_n31591_,
    new_n31592_, new_n31593_, new_n31594_, new_n31595_, new_n31596_,
    new_n31597_, new_n31598_, new_n31599_, new_n31600_, new_n31601_,
    new_n31602_, new_n31603_, new_n31604_, new_n31605_, new_n31606_,
    new_n31607_, new_n31608_, new_n31609_, new_n31610_, new_n31611_,
    new_n31612_, new_n31613_, new_n31614_, new_n31615_, new_n31616_,
    new_n31617_, new_n31618_, new_n31619_, new_n31620_, new_n31621_,
    new_n31622_, new_n31623_, new_n31624_, new_n31625_, new_n31626_,
    new_n31627_, new_n31628_, new_n31629_, new_n31630_, new_n31631_,
    new_n31632_, new_n31633_, new_n31634_, new_n31635_, new_n31636_,
    new_n31637_, new_n31638_, new_n31639_, new_n31640_, new_n31641_,
    new_n31642_, new_n31643_, new_n31644_, new_n31645_, new_n31646_,
    new_n31647_, new_n31648_, new_n31649_, new_n31650_, new_n31651_,
    new_n31652_, new_n31653_, new_n31654_, new_n31655_, new_n31656_,
    new_n31657_, new_n31658_, new_n31659_, new_n31660_, new_n31661_,
    new_n31662_, new_n31663_, new_n31664_, new_n31665_, new_n31666_,
    new_n31667_, new_n31668_, new_n31669_, new_n31670_, new_n31671_,
    new_n31672_, new_n31673_, new_n31674_, new_n31675_, new_n31676_,
    new_n31677_, new_n31678_, new_n31679_, new_n31680_, new_n31681_,
    new_n31682_, new_n31683_, new_n31684_, new_n31685_, new_n31686_,
    new_n31687_, new_n31688_, new_n31689_, new_n31690_, new_n31691_,
    new_n31692_, new_n31693_, new_n31694_, new_n31695_, new_n31696_,
    new_n31697_, new_n31698_, new_n31699_, new_n31700_, new_n31701_,
    new_n31702_, new_n31703_, new_n31704_, new_n31705_, new_n31706_,
    new_n31707_, new_n31708_, new_n31709_, new_n31710_, new_n31711_,
    new_n31712_, new_n31713_, new_n31714_, new_n31715_, new_n31716_,
    new_n31717_, new_n31718_, new_n31719_, new_n31720_, new_n31721_,
    new_n31722_, new_n31723_, new_n31724_, new_n31725_, new_n31726_,
    new_n31727_, new_n31728_, new_n31729_, new_n31730_, new_n31731_,
    new_n31732_, new_n31733_, new_n31734_, new_n31735_, new_n31736_,
    new_n31737_, new_n31738_, new_n31739_, new_n31740_, new_n31741_,
    new_n31742_, new_n31743_, new_n31744_, new_n31745_, new_n31746_,
    new_n31747_, new_n31748_, new_n31749_, new_n31750_, new_n31751_,
    new_n31752_, new_n31753_, new_n31754_, new_n31755_, new_n31756_,
    new_n31757_, new_n31758_, new_n31759_, new_n31760_, new_n31761_,
    new_n31762_, new_n31763_, new_n31764_, new_n31765_, new_n31766_,
    new_n31767_, new_n31768_, new_n31769_, new_n31770_, new_n31771_,
    new_n31772_, new_n31773_, new_n31774_, new_n31775_, new_n31776_,
    new_n31777_, new_n31778_, new_n31779_, new_n31780_, new_n31781_,
    new_n31782_, new_n31783_, new_n31784_, new_n31785_, new_n31786_,
    new_n31787_, new_n31788_, new_n31789_, new_n31790_, new_n31791_,
    new_n31792_, new_n31793_, new_n31794_, new_n31795_, new_n31796_,
    new_n31797_, new_n31798_, new_n31799_, new_n31800_, new_n31801_,
    new_n31802_, new_n31803_, new_n31804_, new_n31805_, new_n31806_,
    new_n31807_, new_n31808_, new_n31809_, new_n31810_, new_n31811_,
    new_n31812_, new_n31813_, new_n31814_, new_n31815_, new_n31816_,
    new_n31817_, new_n31818_, new_n31819_, new_n31820_, new_n31821_,
    new_n31822_, new_n31823_, new_n31824_, new_n31825_, new_n31826_,
    new_n31827_, new_n31828_, new_n31829_, new_n31830_, new_n31831_,
    new_n31832_, new_n31833_, new_n31834_, new_n31835_, new_n31836_,
    new_n31837_, new_n31838_, new_n31839_, new_n31840_, new_n31841_,
    new_n31842_, new_n31843_, new_n31844_, new_n31845_, new_n31846_,
    new_n31847_, new_n31848_, new_n31849_, new_n31850_, new_n31851_,
    new_n31852_, new_n31853_, new_n31854_, new_n31855_, new_n31856_,
    new_n31857_, new_n31858_, new_n31859_, new_n31860_, new_n31861_,
    new_n31862_, new_n31863_, new_n31864_, new_n31865_, new_n31866_,
    new_n31867_, new_n31868_, new_n31869_, new_n31870_, new_n31871_,
    new_n31872_, new_n31873_, new_n31874_, new_n31875_, new_n31876_,
    new_n31877_, new_n31878_, new_n31879_, new_n31880_, new_n31881_,
    new_n31882_, new_n31883_, new_n31884_, new_n31885_, new_n31886_,
    new_n31887_, new_n31888_, new_n31889_, new_n31890_, new_n31891_,
    new_n31892_, new_n31893_, new_n31894_, new_n31895_, new_n31896_,
    new_n31897_, new_n31898_, new_n31899_, new_n31900_, new_n31901_,
    new_n31902_, new_n31903_, new_n31904_, new_n31905_, new_n31906_,
    new_n31907_, new_n31908_, new_n31909_, new_n31910_, new_n31911_,
    new_n31912_, new_n31913_, new_n31914_, new_n31915_, new_n31916_,
    new_n31917_, new_n31918_, new_n31919_, new_n31920_, new_n31921_,
    new_n31922_, new_n31923_, new_n31924_, new_n31925_, new_n31926_,
    new_n31927_, new_n31928_, new_n31929_, new_n31930_, new_n31931_,
    new_n31932_, new_n31933_, new_n31934_, new_n31935_, new_n31936_,
    new_n31937_, new_n31938_, new_n31939_, new_n31940_, new_n31941_,
    new_n31942_, new_n31943_, new_n31944_, new_n31945_, new_n31946_,
    new_n31947_, new_n31948_, new_n31949_, new_n31950_, new_n31951_,
    new_n31952_, new_n31953_, new_n31954_, new_n31955_, new_n31956_,
    new_n31957_, new_n31958_, new_n31959_, new_n31960_, new_n31961_,
    new_n31962_, new_n31963_, new_n31964_, new_n31965_, new_n31966_,
    new_n31967_, new_n31968_, new_n31969_, new_n31970_, new_n31971_,
    new_n31972_, new_n31973_, new_n31974_, new_n31975_, new_n31976_,
    new_n31977_, new_n31978_, new_n31979_, new_n31980_, new_n31981_,
    new_n31982_, new_n31983_, new_n31984_, new_n31985_, new_n31986_,
    new_n31987_, new_n31988_, new_n31989_, new_n31990_, new_n31991_,
    new_n31992_, new_n31993_, new_n31994_, new_n31995_, new_n31996_,
    new_n31997_, new_n31998_, new_n31999_, new_n32000_, new_n32001_,
    new_n32002_, new_n32003_, new_n32004_, new_n32005_, new_n32006_,
    new_n32007_, new_n32008_, new_n32009_, new_n32010_, new_n32011_,
    new_n32012_, new_n32013_, new_n32014_, new_n32015_, new_n32016_,
    new_n32017_, new_n32018_, new_n32019_, new_n32020_, new_n32021_,
    new_n32022_, new_n32023_, new_n32024_, new_n32025_, new_n32026_,
    new_n32027_, new_n32028_, new_n32029_, new_n32030_, new_n32031_,
    new_n32032_, new_n32033_, new_n32034_, new_n32035_, new_n32036_,
    new_n32037_, new_n32038_, new_n32039_, new_n32040_, new_n32041_,
    new_n32042_, new_n32043_, new_n32044_, new_n32045_, new_n32046_,
    new_n32047_, new_n32048_, new_n32049_, new_n32050_, new_n32051_,
    new_n32052_, new_n32053_, new_n32054_, new_n32055_, new_n32056_,
    new_n32057_, new_n32058_, new_n32059_, new_n32060_, new_n32061_,
    new_n32062_, new_n32063_, new_n32064_, new_n32065_, new_n32066_,
    new_n32067_, new_n32068_, new_n32069_, new_n32070_, new_n32071_,
    new_n32072_, new_n32073_, new_n32074_, new_n32075_, new_n32076_,
    new_n32077_, new_n32078_, new_n32079_, new_n32080_, new_n32081_,
    new_n32082_, new_n32083_, new_n32084_, new_n32085_, new_n32086_,
    new_n32087_, new_n32088_, new_n32089_, new_n32090_, new_n32091_,
    new_n32092_, new_n32093_, new_n32094_, new_n32095_, new_n32096_,
    new_n32097_, new_n32098_, new_n32099_, new_n32100_, new_n32101_,
    new_n32102_, new_n32103_, new_n32104_, new_n32105_, new_n32106_,
    new_n32107_, new_n32108_, new_n32109_, new_n32110_, new_n32111_,
    new_n32112_, new_n32113_, new_n32114_, new_n32115_, new_n32116_,
    new_n32117_, new_n32118_, new_n32119_, new_n32120_, new_n32121_,
    new_n32122_, new_n32123_, new_n32124_, new_n32125_, new_n32126_,
    new_n32127_, new_n32128_, new_n32129_, new_n32130_, new_n32131_,
    new_n32132_, new_n32133_, new_n32134_, new_n32135_, new_n32136_,
    new_n32137_, new_n32138_, new_n32139_, new_n32140_, new_n32141_,
    new_n32142_, new_n32143_, new_n32144_, new_n32145_, new_n32146_,
    new_n32147_, new_n32148_, new_n32149_, new_n32150_, new_n32151_,
    new_n32152_, new_n32153_, new_n32154_, new_n32155_, new_n32156_,
    new_n32157_, new_n32158_, new_n32159_, new_n32160_, new_n32161_,
    new_n32162_, new_n32163_, new_n32164_, new_n32165_, new_n32166_,
    new_n32167_, new_n32168_, new_n32169_, new_n32170_, new_n32171_,
    new_n32172_, new_n32173_, new_n32174_, new_n32175_, new_n32176_,
    new_n32177_, new_n32178_, new_n32179_, new_n32180_, new_n32181_,
    new_n32182_, new_n32183_, new_n32184_, new_n32185_, new_n32186_,
    new_n32187_, new_n32188_, new_n32189_, new_n32190_, new_n32191_,
    new_n32192_, new_n32193_, new_n32194_, new_n32195_, new_n32196_,
    new_n32197_, new_n32198_, new_n32199_, new_n32200_, new_n32201_,
    new_n32202_, new_n32203_, new_n32204_, new_n32205_, new_n32206_,
    new_n32207_, new_n32208_, new_n32209_, new_n32210_, new_n32211_,
    new_n32212_, new_n32213_, new_n32214_, new_n32215_, new_n32216_,
    new_n32217_, new_n32218_, new_n32219_, new_n32220_, new_n32221_,
    new_n32222_, new_n32223_, new_n32224_, new_n32225_, new_n32226_,
    new_n32227_, new_n32228_, new_n32229_, new_n32230_, new_n32231_,
    new_n32232_, new_n32233_, new_n32234_, new_n32235_, new_n32236_,
    new_n32237_, new_n32238_, new_n32239_, new_n32240_, new_n32241_,
    new_n32242_, new_n32243_, new_n32244_, new_n32245_, new_n32246_,
    new_n32247_, new_n32248_, new_n32249_, new_n32250_, new_n32251_,
    new_n32252_, new_n32253_, new_n32254_, new_n32255_, new_n32256_,
    new_n32257_, new_n32258_, new_n32259_, new_n32260_, new_n32261_,
    new_n32262_, new_n32263_, new_n32264_, new_n32265_, new_n32266_,
    new_n32267_, new_n32268_, new_n32269_, new_n32270_, new_n32271_,
    new_n32272_, new_n32273_, new_n32274_, new_n32275_, new_n32276_,
    new_n32277_, new_n32278_, new_n32279_, new_n32280_, new_n32281_,
    new_n32282_, new_n32283_, new_n32284_, new_n32285_, new_n32286_,
    new_n32287_, new_n32288_, new_n32289_, new_n32290_, new_n32291_,
    new_n32292_, new_n32293_, new_n32294_, new_n32295_, new_n32296_,
    new_n32297_, new_n32298_, new_n32299_, new_n32300_, new_n32301_,
    new_n32302_, new_n32303_, new_n32304_, new_n32305_, new_n32306_,
    new_n32307_, new_n32308_, new_n32309_, new_n32310_, new_n32311_,
    new_n32312_, new_n32313_, new_n32314_, new_n32315_, new_n32316_,
    new_n32317_, new_n32318_, new_n32319_, new_n32320_, new_n32321_,
    new_n32322_, new_n32323_, new_n32324_, new_n32325_, new_n32326_,
    new_n32327_, new_n32328_, new_n32329_, new_n32330_, new_n32331_,
    new_n32332_, new_n32333_, new_n32334_, new_n32335_, new_n32336_,
    new_n32337_, new_n32338_, new_n32339_, new_n32340_, new_n32341_,
    new_n32342_, new_n32343_, new_n32344_, new_n32345_, new_n32346_,
    new_n32347_, new_n32348_, new_n32349_, new_n32350_, new_n32351_,
    new_n32352_, new_n32353_, new_n32354_, new_n32355_, new_n32356_,
    new_n32357_, new_n32358_, new_n32359_, new_n32360_, new_n32361_,
    new_n32362_, new_n32363_, new_n32364_, new_n32365_, new_n32366_,
    new_n32367_, new_n32368_, new_n32369_, new_n32370_, new_n32371_,
    new_n32372_, new_n32373_, new_n32374_, new_n32375_, new_n32376_,
    new_n32377_, new_n32378_, new_n32379_, new_n32380_, new_n32381_,
    new_n32382_, new_n32383_, new_n32384_, new_n32385_, new_n32386_,
    new_n32387_, new_n32388_, new_n32389_, new_n32390_, new_n32391_,
    new_n32392_, new_n32393_, new_n32394_, new_n32395_, new_n32396_,
    new_n32397_, new_n32398_, new_n32399_, new_n32400_, new_n32401_,
    new_n32402_, new_n32403_, new_n32404_, new_n32405_, new_n32406_,
    new_n32407_, new_n32408_, new_n32409_, new_n32410_, new_n32411_,
    new_n32412_, new_n32413_, new_n32414_, new_n32415_, new_n32416_,
    new_n32417_, new_n32418_, new_n32419_, new_n32420_, new_n32421_,
    new_n32422_, new_n32423_, new_n32424_, new_n32425_, new_n32426_,
    new_n32427_, new_n32428_, new_n32429_, new_n32430_, new_n32431_,
    new_n32432_, new_n32433_, new_n32434_, new_n32435_, new_n32436_,
    new_n32437_, new_n32438_, new_n32439_, new_n32440_, new_n32441_,
    new_n32442_, new_n32443_, new_n32444_, new_n32445_, new_n32446_,
    new_n32447_, new_n32448_, new_n32449_, new_n32450_, new_n32451_,
    new_n32452_, new_n32453_, new_n32454_, new_n32455_, new_n32456_,
    new_n32457_, new_n32458_, new_n32459_, new_n32460_, new_n32461_,
    new_n32462_, new_n32463_, new_n32464_, new_n32465_, new_n32466_,
    new_n32467_, new_n32468_, new_n32469_, new_n32470_, new_n32471_,
    new_n32472_, new_n32473_, new_n32474_, new_n32475_, new_n32476_,
    new_n32477_, new_n32478_, new_n32479_, new_n32480_, new_n32481_,
    new_n32482_, new_n32483_, new_n32484_, new_n32485_, new_n32486_,
    new_n32487_, new_n32488_, new_n32489_, new_n32490_, new_n32491_,
    new_n32492_, new_n32493_, new_n32494_, new_n32495_, new_n32496_,
    new_n32497_, new_n32498_, new_n32499_, new_n32500_, new_n32501_,
    new_n32502_, new_n32503_, new_n32504_, new_n32505_, new_n32506_,
    new_n32507_, new_n32508_, new_n32509_, new_n32510_, new_n32511_,
    new_n32512_, new_n32513_, new_n32514_, new_n32515_, new_n32516_,
    new_n32517_, new_n32518_, new_n32519_, new_n32520_, new_n32521_,
    new_n32522_, new_n32523_, new_n32524_, new_n32525_, new_n32526_,
    new_n32527_, new_n32528_, new_n32529_, new_n32530_, new_n32531_,
    new_n32532_, new_n32533_, new_n32534_, new_n32535_, new_n32536_,
    new_n32537_, new_n32538_, new_n32539_, new_n32540_, new_n32541_,
    new_n32542_, new_n32543_, new_n32544_, new_n32545_, new_n32546_,
    new_n32547_, new_n32548_, new_n32549_, new_n32550_, new_n32551_,
    new_n32552_, new_n32553_, new_n32554_, new_n32555_, new_n32556_,
    new_n32557_, new_n32558_, new_n32559_, new_n32560_, new_n32561_,
    new_n32562_, new_n32563_, new_n32564_, new_n32565_, new_n32566_,
    new_n32567_, new_n32568_, new_n32569_, new_n32570_, new_n32571_,
    new_n32572_, new_n32573_, new_n32574_, new_n32575_, new_n32576_,
    new_n32577_, new_n32578_, new_n32579_, new_n32580_, new_n32581_,
    new_n32582_, new_n32583_, new_n32584_, new_n32585_, new_n32586_,
    new_n32587_, new_n32588_, new_n32589_, new_n32590_, new_n32591_,
    new_n32592_, new_n32593_, new_n32594_, new_n32595_, new_n32596_,
    new_n32597_, new_n32598_, new_n32599_, new_n32600_, new_n32601_,
    new_n32602_, new_n32603_, new_n32604_, new_n32605_, new_n32606_,
    new_n32607_, new_n32608_, new_n32609_, new_n32610_, new_n32611_,
    new_n32612_, new_n32613_, new_n32614_, new_n32615_, new_n32616_,
    new_n32617_, new_n32618_, new_n32619_, new_n32620_, new_n32621_,
    new_n32622_, new_n32623_, new_n32624_, new_n32625_, new_n32626_,
    new_n32627_, new_n32628_, new_n32629_, new_n32630_, new_n32631_,
    new_n32632_, new_n32633_, new_n32634_, new_n32635_, new_n32636_,
    new_n32637_, new_n32638_, new_n32639_, new_n32640_, new_n32641_,
    new_n32642_, new_n32643_, new_n32644_, new_n32645_, new_n32646_,
    new_n32647_, new_n32648_, new_n32649_, new_n32650_, new_n32651_,
    new_n32652_, new_n32653_, new_n32654_, new_n32655_, new_n32656_,
    new_n32657_, new_n32658_, new_n32659_, new_n32660_, new_n32661_,
    new_n32662_, new_n32663_, new_n32664_, new_n32665_, new_n32666_,
    new_n32667_, new_n32668_, new_n32669_, new_n32670_, new_n32671_,
    new_n32672_, new_n32673_, new_n32674_, new_n32675_, new_n32676_,
    new_n32677_, new_n32678_, new_n32679_, new_n32680_, new_n32681_,
    new_n32682_, new_n32683_, new_n32684_, new_n32685_, new_n32686_,
    new_n32687_, new_n32688_, new_n32689_, new_n32690_, new_n32691_,
    new_n32692_, new_n32693_, new_n32694_, new_n32695_, new_n32696_,
    new_n32697_, new_n32698_, new_n32699_, new_n32700_, new_n32701_,
    new_n32702_, new_n32703_, new_n32704_, new_n32705_, new_n32706_,
    new_n32707_, new_n32708_, new_n32709_, new_n32710_, new_n32711_,
    new_n32712_, new_n32713_, new_n32714_, new_n32715_, new_n32716_,
    new_n32717_, new_n32718_, new_n32719_, new_n32720_, new_n32721_,
    new_n32722_, new_n32723_, new_n32724_, new_n32725_, new_n32726_,
    new_n32727_, new_n32728_, new_n32729_, new_n32730_, new_n32731_,
    new_n32732_, new_n32733_, new_n32734_, new_n32735_, new_n32736_,
    new_n32737_, new_n32738_, new_n32739_, new_n32740_, new_n32741_,
    new_n32742_, new_n32743_, new_n32744_, new_n32745_, new_n32746_,
    new_n32747_, new_n32748_, new_n32749_, new_n32750_, new_n32751_,
    new_n32752_, new_n32753_, new_n32754_, new_n32755_, new_n32756_,
    new_n32757_, new_n32758_, new_n32759_, new_n32760_, new_n32761_,
    new_n32762_, new_n32763_, new_n32764_, new_n32765_, new_n32766_,
    new_n32767_, new_n32768_, new_n32769_, new_n32770_, new_n32771_,
    new_n32772_, new_n32773_, new_n32774_, new_n32775_, new_n32776_,
    new_n32777_, new_n32778_, new_n32779_, new_n32780_, new_n32781_,
    new_n32782_, new_n32783_, new_n32784_, new_n32785_, new_n32786_,
    new_n32787_, new_n32788_, new_n32789_, new_n32790_, new_n32791_,
    new_n32792_, new_n32793_, new_n32794_, new_n32795_, new_n32796_,
    new_n32797_, new_n32798_, new_n32799_, new_n32800_, new_n32801_,
    new_n32802_, new_n32803_, new_n32804_, new_n32805_, new_n32806_,
    new_n32807_, new_n32808_, new_n32809_, new_n32810_, new_n32811_,
    new_n32812_, new_n32813_, new_n32814_, new_n32815_, new_n32816_,
    new_n32817_, new_n32818_, new_n32819_, new_n32820_, new_n32821_,
    new_n32822_, new_n32823_, new_n32824_, new_n32825_, new_n32826_,
    new_n32827_, new_n32828_, new_n32829_, new_n32830_, new_n32831_,
    new_n32832_, new_n32833_, new_n32834_, new_n32835_, new_n32836_,
    new_n32837_, new_n32838_, new_n32839_, new_n32840_, new_n32841_,
    new_n32842_, new_n32843_, new_n32844_, new_n32845_, new_n32846_,
    new_n32847_, new_n32848_, new_n32849_, new_n32850_, new_n32851_,
    new_n32852_, new_n32853_, new_n32854_, new_n32855_, new_n32856_,
    new_n32857_, new_n32858_, new_n32859_, new_n32860_, new_n32861_,
    new_n32862_, new_n32863_, new_n32864_, new_n32865_, new_n32866_,
    new_n32867_, new_n32868_, new_n32869_, new_n32870_, new_n32871_,
    new_n32872_, new_n32873_, new_n32874_, new_n32875_, new_n32876_,
    new_n32877_, new_n32878_, new_n32879_, new_n32880_, new_n32881_,
    new_n32882_, new_n32883_, new_n32884_, new_n32885_, new_n32886_,
    new_n32887_, new_n32888_, new_n32889_, new_n32890_, new_n32891_,
    new_n32892_, new_n32893_, new_n32894_, new_n32895_, new_n32896_,
    new_n32897_, new_n32898_, new_n32899_, new_n32900_, new_n32901_,
    new_n32902_, new_n32903_, new_n32904_, new_n32905_, new_n32906_,
    new_n32907_, new_n32908_, new_n32909_, new_n32910_, new_n32911_,
    new_n32912_, new_n32913_, new_n32914_, new_n32915_, new_n32916_,
    new_n32917_, new_n32918_, new_n32919_, new_n32920_, new_n32921_,
    new_n32922_, new_n32923_, new_n32924_, new_n32925_, new_n32926_,
    new_n32927_, new_n32928_, new_n32929_, new_n32930_, new_n32931_,
    new_n32932_, new_n32933_, new_n32934_, new_n32935_, new_n32936_,
    new_n32937_, new_n32938_, new_n32939_, new_n32940_, new_n32941_,
    new_n32942_, new_n32943_, new_n32944_, new_n32945_, new_n32946_,
    new_n32947_, new_n32948_, new_n32949_, new_n32950_, new_n32951_,
    new_n32952_, new_n32953_, new_n32954_, new_n32955_, new_n32956_,
    new_n32957_, new_n32958_, new_n32959_, new_n32960_, new_n32961_,
    new_n32962_, new_n32963_, new_n32964_, new_n32965_, new_n32966_,
    new_n32967_, new_n32968_, new_n32969_, new_n32970_, new_n32971_,
    new_n32972_, new_n32973_, new_n32974_, new_n32975_, new_n32976_,
    new_n32977_, new_n32978_, new_n32979_, new_n32980_, new_n32981_,
    new_n32982_, new_n32983_, new_n32984_, new_n32985_, new_n32986_,
    new_n32987_, new_n32988_, new_n32989_, new_n32990_, new_n32991_,
    new_n32992_, new_n32993_, new_n32994_, new_n32995_, new_n32996_,
    new_n32997_, new_n32998_, new_n32999_, new_n33000_, new_n33001_,
    new_n33002_, new_n33003_, new_n33004_, new_n33005_, new_n33006_,
    new_n33007_, new_n33008_, new_n33009_, new_n33010_, new_n33011_,
    new_n33012_, new_n33013_, new_n33014_, new_n33015_, new_n33016_,
    new_n33017_, new_n33018_, new_n33019_, new_n33020_, new_n33021_,
    new_n33022_, new_n33023_, new_n33024_, new_n33025_, new_n33026_,
    new_n33027_, new_n33028_, new_n33029_, new_n33030_, new_n33031_,
    new_n33032_, new_n33033_, new_n33034_, new_n33035_, new_n33036_,
    new_n33037_, new_n33038_, new_n33039_, new_n33040_, new_n33041_,
    new_n33042_, new_n33043_, new_n33044_, new_n33045_, new_n33046_,
    new_n33047_, new_n33048_, new_n33049_, new_n33050_, new_n33051_,
    new_n33052_, new_n33053_, new_n33054_, new_n33055_, new_n33056_,
    new_n33057_, new_n33058_, new_n33059_, new_n33060_, new_n33061_,
    new_n33062_, new_n33063_, new_n33064_, new_n33065_, new_n33066_,
    new_n33067_, new_n33068_, new_n33069_, new_n33070_, new_n33071_,
    new_n33072_, new_n33073_, new_n33074_, new_n33075_, new_n33076_,
    new_n33077_, new_n33078_, new_n33079_, new_n33080_, new_n33081_,
    new_n33082_, new_n33083_, new_n33084_, new_n33085_, new_n33086_,
    new_n33087_, new_n33088_, new_n33089_, new_n33090_, new_n33091_,
    new_n33092_, new_n33093_, new_n33094_, new_n33095_, new_n33096_,
    new_n33097_, new_n33098_, new_n33099_, new_n33100_, new_n33101_,
    new_n33102_, new_n33103_, new_n33104_, new_n33105_, new_n33106_,
    new_n33107_, new_n33108_, new_n33109_, new_n33110_, new_n33111_,
    new_n33112_, new_n33113_, new_n33114_, new_n33115_, new_n33116_,
    new_n33117_, new_n33118_, new_n33119_, new_n33120_, new_n33121_,
    new_n33122_, new_n33123_, new_n33124_, new_n33125_, new_n33126_,
    new_n33127_, new_n33128_, new_n33129_, new_n33130_, new_n33131_,
    new_n33132_, new_n33133_, new_n33134_, new_n33135_, new_n33136_,
    new_n33137_, new_n33138_, new_n33139_, new_n33140_, new_n33141_,
    new_n33142_, new_n33143_, new_n33144_, new_n33145_, new_n33146_,
    new_n33147_, new_n33148_, new_n33149_, new_n33150_, new_n33151_,
    new_n33152_, new_n33153_, new_n33154_, new_n33155_, new_n33156_,
    new_n33157_, new_n33158_, new_n33159_, new_n33160_, new_n33161_,
    new_n33162_, new_n33163_, new_n33164_, new_n33165_, new_n33166_,
    new_n33167_, new_n33168_, new_n33169_, new_n33170_, new_n33171_,
    new_n33172_, new_n33173_, new_n33174_, new_n33175_, new_n33176_,
    new_n33177_, new_n33178_, new_n33179_, new_n33180_, new_n33181_,
    new_n33182_, new_n33183_, new_n33184_, new_n33185_, new_n33186_,
    new_n33187_, new_n33188_, new_n33189_, new_n33190_, new_n33191_,
    new_n33192_, new_n33193_, new_n33194_, new_n33195_, new_n33196_,
    new_n33197_, new_n33198_, new_n33199_, new_n33200_, new_n33201_,
    new_n33202_, new_n33203_, new_n33204_, new_n33205_, new_n33206_,
    new_n33207_, new_n33208_, new_n33209_, new_n33210_, new_n33211_,
    new_n33212_, new_n33213_, new_n33214_, new_n33215_, new_n33216_,
    new_n33217_, new_n33218_, new_n33219_, new_n33220_, new_n33221_,
    new_n33222_, new_n33223_, new_n33224_, new_n33225_, new_n33226_,
    new_n33227_, new_n33228_, new_n33229_, new_n33230_, new_n33231_,
    new_n33232_, new_n33233_, new_n33234_, new_n33235_, new_n33236_,
    new_n33237_, new_n33238_, new_n33239_, new_n33240_, new_n33241_,
    new_n33242_, new_n33243_, new_n33244_, new_n33245_, new_n33246_,
    new_n33247_, new_n33248_, new_n33249_, new_n33250_, new_n33251_,
    new_n33252_, new_n33253_, new_n33254_, new_n33255_, new_n33256_,
    new_n33257_, new_n33258_, new_n33259_, new_n33260_, new_n33261_,
    new_n33262_, new_n33263_, new_n33264_, new_n33265_, new_n33266_,
    new_n33267_, new_n33268_, new_n33269_, new_n33270_, new_n33271_,
    new_n33272_, new_n33273_, new_n33274_, new_n33275_, new_n33276_,
    new_n33277_, new_n33278_, new_n33279_, new_n33280_, new_n33281_,
    new_n33282_, new_n33283_, new_n33284_, new_n33285_, new_n33286_,
    new_n33287_, new_n33288_, new_n33289_, new_n33290_, new_n33291_,
    new_n33292_, new_n33293_, new_n33294_, new_n33295_, new_n33296_,
    new_n33297_, new_n33298_, new_n33299_, new_n33300_, new_n33301_,
    new_n33302_, new_n33303_, new_n33304_, new_n33305_, new_n33306_,
    new_n33307_, new_n33308_, new_n33309_, new_n33310_, new_n33311_,
    new_n33312_, new_n33313_, new_n33314_, new_n33315_, new_n33316_,
    new_n33317_, new_n33318_, new_n33319_, new_n33320_, new_n33321_,
    new_n33322_, new_n33323_, new_n33324_, new_n33325_, new_n33326_,
    new_n33327_, new_n33328_, new_n33329_, new_n33330_, new_n33331_,
    new_n33332_, new_n33333_, new_n33334_, new_n33335_, new_n33336_,
    new_n33337_, new_n33338_, new_n33339_, new_n33340_, new_n33341_,
    new_n33342_, new_n33343_, new_n33344_, new_n33345_, new_n33346_,
    new_n33347_, new_n33348_, new_n33349_, new_n33350_, new_n33351_,
    new_n33352_, new_n33353_, new_n33354_, new_n33355_, new_n33356_,
    new_n33357_, new_n33358_, new_n33359_, new_n33360_, new_n33361_,
    new_n33362_, new_n33363_, new_n33364_, new_n33365_, new_n33366_,
    new_n33367_, new_n33368_, new_n33369_, new_n33370_, new_n33371_,
    new_n33372_, new_n33373_, new_n33374_, new_n33375_, new_n33376_,
    new_n33377_, new_n33378_, new_n33379_, new_n33380_, new_n33381_,
    new_n33382_, new_n33383_, new_n33384_, new_n33385_, new_n33386_,
    new_n33387_, new_n33388_, new_n33389_, new_n33390_, new_n33391_,
    new_n33392_, new_n33393_, new_n33394_, new_n33395_, new_n33396_,
    new_n33397_, new_n33398_, new_n33399_, new_n33400_, new_n33401_,
    new_n33402_, new_n33403_, new_n33404_, new_n33405_, new_n33406_,
    new_n33407_, new_n33408_, new_n33409_, new_n33410_, new_n33411_,
    new_n33412_, new_n33413_, new_n33414_, new_n33415_, new_n33416_,
    new_n33417_, new_n33418_, new_n33419_, new_n33420_, new_n33421_,
    new_n33422_, new_n33423_, new_n33424_, new_n33425_, new_n33426_,
    new_n33427_, new_n33428_, new_n33429_, new_n33430_, new_n33431_,
    new_n33432_, new_n33433_, new_n33434_, new_n33435_, new_n33436_,
    new_n33437_, new_n33438_, new_n33439_, new_n33440_, new_n33441_,
    new_n33442_, new_n33443_, new_n33444_, new_n33445_, new_n33446_,
    new_n33447_, new_n33448_, new_n33449_, new_n33450_, new_n33451_,
    new_n33452_, new_n33453_, new_n33454_, new_n33455_, new_n33456_,
    new_n33457_, new_n33458_, new_n33459_, new_n33460_, new_n33461_,
    new_n33462_, new_n33463_, new_n33464_, new_n33465_, new_n33466_,
    new_n33467_, new_n33468_, new_n33469_, new_n33470_, new_n33471_,
    new_n33472_, new_n33473_, new_n33474_, new_n33475_, new_n33476_,
    new_n33477_, new_n33478_, new_n33479_, new_n33480_, new_n33481_,
    new_n33482_, new_n33483_, new_n33484_, new_n33485_, new_n33486_,
    new_n33487_, new_n33488_, new_n33489_, new_n33490_, new_n33491_,
    new_n33492_, new_n33493_, new_n33494_, new_n33495_, new_n33496_,
    new_n33497_, new_n33498_, new_n33499_, new_n33500_, new_n33501_,
    new_n33502_, new_n33503_, new_n33504_, new_n33505_, new_n33506_,
    new_n33507_, new_n33508_, new_n33509_, new_n33510_, new_n33511_,
    new_n33512_, new_n33513_, new_n33514_, new_n33515_, new_n33516_,
    new_n33517_, new_n33518_, new_n33519_, new_n33520_, new_n33521_,
    new_n33522_, new_n33523_, new_n33524_, new_n33525_, new_n33526_,
    new_n33527_, new_n33528_, new_n33529_, new_n33530_, new_n33531_,
    new_n33532_, new_n33533_, new_n33534_, new_n33535_, new_n33536_,
    new_n33537_, new_n33538_, new_n33539_, new_n33540_, new_n33541_,
    new_n33542_, new_n33543_, new_n33544_, new_n33545_, new_n33546_,
    new_n33547_, new_n33548_, new_n33549_, new_n33550_, new_n33551_,
    new_n33552_, new_n33553_, new_n33554_, new_n33555_, new_n33556_,
    new_n33557_, new_n33558_, new_n33559_, new_n33560_, new_n33561_,
    new_n33562_, new_n33563_, new_n33564_, new_n33565_, new_n33566_,
    new_n33567_, new_n33568_, new_n33569_, new_n33570_, new_n33571_,
    new_n33572_, new_n33573_, new_n33574_, new_n33575_, new_n33576_,
    new_n33577_, new_n33578_, new_n33579_, new_n33580_, new_n33581_,
    new_n33582_, new_n33583_, new_n33584_, new_n33585_, new_n33586_,
    new_n33587_, new_n33588_, new_n33589_, new_n33590_, new_n33591_,
    new_n33592_, new_n33593_, new_n33594_, new_n33595_, new_n33596_,
    new_n33597_, new_n33598_, new_n33599_, new_n33600_, new_n33601_,
    new_n33602_, new_n33603_, new_n33604_, new_n33605_, new_n33606_,
    new_n33607_, new_n33608_, new_n33609_, new_n33610_, new_n33611_,
    new_n33612_, new_n33613_, new_n33614_, new_n33615_, new_n33616_,
    new_n33617_, new_n33618_, new_n33619_, new_n33620_, new_n33621_,
    new_n33622_, new_n33623_, new_n33624_, new_n33625_, new_n33626_,
    new_n33627_, new_n33628_, new_n33629_, new_n33630_, new_n33631_,
    new_n33632_, new_n33633_, new_n33634_, new_n33635_, new_n33636_,
    new_n33637_, new_n33638_, new_n33639_, new_n33640_, new_n33641_,
    new_n33642_, new_n33643_, new_n33644_, new_n33645_, new_n33646_,
    new_n33647_, new_n33648_, new_n33649_, new_n33650_, new_n33651_,
    new_n33652_, new_n33653_, new_n33654_, new_n33655_, new_n33656_,
    new_n33657_, new_n33658_, new_n33659_, new_n33660_, new_n33661_,
    new_n33662_, new_n33663_, new_n33664_, new_n33665_, new_n33666_,
    new_n33667_, new_n33668_, new_n33669_, new_n33670_, new_n33671_,
    new_n33672_, new_n33673_, new_n33674_, new_n33675_, new_n33676_,
    new_n33677_, new_n33678_, new_n33679_, new_n33680_, new_n33681_,
    new_n33682_, new_n33683_, new_n33684_, new_n33685_, new_n33686_,
    new_n33687_, new_n33688_, new_n33689_, new_n33690_, new_n33691_,
    new_n33692_, new_n33693_, new_n33694_, new_n33695_, new_n33696_,
    new_n33697_, new_n33698_, new_n33699_, new_n33700_, new_n33701_,
    new_n33702_, new_n33703_, new_n33704_, new_n33705_, new_n33706_,
    new_n33707_, new_n33708_, new_n33709_, new_n33710_, new_n33711_,
    new_n33712_, new_n33713_, new_n33714_, new_n33715_, new_n33716_,
    new_n33717_, new_n33718_, new_n33719_, new_n33720_, new_n33721_,
    new_n33722_, new_n33723_, new_n33724_, new_n33725_, new_n33726_,
    new_n33727_, new_n33728_, new_n33729_, new_n33730_, new_n33731_,
    new_n33732_, new_n33733_, new_n33734_, new_n33735_, new_n33736_,
    new_n33737_, new_n33738_, new_n33739_, new_n33740_, new_n33741_,
    new_n33742_;
  assign new_n2966_ = ~new_n9273_ | ~new_n9347_;
  assign new_n2967_ = ~pi1231 | ~new_n9348_;
  assign new_n2968_ = ~new_n9264_ | ~new_n9329_;
  assign new_n2969_ = new_n3012_ & po0164;
  assign new_n2970_ = pi0999 & new_n3139_ & new_n3140_ & pi0993;
  assign new_n2971_ = pi0104 & pi0037;
  assign new_n2972_ = pi0105 & pi0036;
  assign new_n2973_ = pi0102 & pi0103;
  assign po0161 = ~po0164 | ~new_n2970_ | ~new_n21008_;
  assign po0163 = ~new_n3142_ | ~po0162 | ~new_n3141_ | ~pi0550;
  assign po0164 = ~pi1448 | ~new_n21018_ | ~new_n3143_ | ~pi1442 | ~new_n3145_;
  assign po0162 = ~new_n21007_ | ~new_n2970_;
  assign po0128 = ~new_n3244_ | ~new_n3245_ | ~new_n3246_;
  assign po0127 = ~new_n3241_ | ~new_n3242_ | ~new_n3243_;
  assign po0126 = ~new_n3238_ | ~new_n3239_ | ~new_n3240_;
  assign po0125 = ~new_n3235_ | ~new_n3236_ | ~new_n3237_;
  assign po0124 = ~new_n3232_ | ~new_n3233_ | ~new_n3234_;
  assign po0123 = ~new_n3229_ | ~new_n3230_ | ~new_n3231_;
  assign po0122 = ~new_n3226_ | ~new_n3227_ | ~new_n3228_;
  assign po0121 = ~new_n3223_ | ~new_n3224_ | ~new_n3225_;
  assign po0120 = ~new_n3220_ | ~new_n3221_ | ~new_n3222_;
  assign po0119 = ~new_n3217_ | ~new_n3218_ | ~new_n3219_;
  assign po0118 = ~new_n3214_ | ~new_n3215_ | ~new_n3216_;
  assign po0117 = ~new_n3211_ | ~new_n3212_ | ~new_n3213_;
  assign po0116 = ~new_n3208_ | ~new_n3209_ | ~new_n3210_;
  assign po0115 = ~new_n3205_ | ~new_n3206_ | ~new_n3207_;
  assign po0114 = ~new_n3202_ | ~new_n3203_ | ~new_n3204_;
  assign po0113 = ~new_n3199_ | ~new_n3200_ | ~new_n3201_;
  assign po0112 = ~new_n3196_ | ~new_n3197_ | ~new_n3198_;
  assign po0111 = ~new_n3193_ | ~new_n3194_ | ~new_n3195_;
  assign po0110 = ~new_n3190_ | ~new_n3191_ | ~new_n3192_;
  assign po0109 = ~new_n3187_ | ~new_n3188_ | ~new_n3189_;
  assign po0108 = ~new_n3184_ | ~new_n3185_ | ~new_n3186_;
  assign po0107 = ~new_n3181_ | ~new_n3182_ | ~new_n3183_;
  assign po0106 = ~new_n3178_ | ~new_n3179_ | ~new_n3180_;
  assign po0105 = ~new_n3175_ | ~new_n3176_ | ~new_n3177_;
  assign po0104 = ~new_n3172_ | ~new_n3173_ | ~new_n3174_;
  assign po0103 = ~new_n3169_ | ~new_n3170_ | ~new_n3171_;
  assign po0102 = ~new_n3166_ | ~new_n3167_ | ~new_n3168_;
  assign po0101 = ~new_n3163_ | ~new_n3164_ | ~new_n3165_;
  assign po0100 = ~new_n3160_ | ~new_n3161_ | ~new_n3162_;
  assign po0099 = ~new_n3157_ | ~new_n3158_ | ~new_n3159_;
  assign po0098 = ~new_n3154_ | ~new_n3155_ | ~new_n3156_;
  assign po0097 = ~new_n3151_ | ~new_n3152_ | ~new_n3153_;
  assign new_n3010_ = ~new_n21018_;
  assign new_n3011_ = ~new_n21008_;
  assign new_n3012_ = ~po0164 | ~new_n3149_;
  assign po0129 = ~new_n3248_ | ~new_n3247_;
  assign po0130 = ~new_n3250_ | ~new_n3249_;
  assign po0131 = ~new_n3252_ | ~new_n3251_;
  assign po0132 = ~new_n3254_ | ~new_n3253_;
  assign po0133 = ~new_n3256_ | ~new_n3255_;
  assign po0134 = ~new_n3258_ | ~new_n3257_;
  assign po0135 = ~new_n3260_ | ~new_n3259_;
  assign po0136 = ~new_n3262_ | ~new_n3261_;
  assign po0137 = ~new_n3264_ | ~new_n3263_;
  assign po0138 = ~new_n3266_ | ~new_n3265_;
  assign po0139 = ~new_n3268_ | ~new_n3267_;
  assign po0140 = ~new_n3270_ | ~new_n3269_;
  assign po0141 = ~new_n3272_ | ~new_n3271_;
  assign po0142 = ~new_n3274_ | ~new_n3273_;
  assign po0143 = ~new_n3276_ | ~new_n3275_;
  assign po0144 = ~new_n3278_ | ~new_n3277_;
  assign po0145 = ~new_n3280_ | ~new_n3279_;
  assign po0146 = ~new_n3282_ | ~new_n3281_;
  assign po0147 = ~new_n3284_ | ~new_n3283_;
  assign po0148 = ~new_n3286_ | ~new_n3285_;
  assign po0149 = ~new_n3288_ | ~new_n3287_;
  assign po0150 = ~new_n3290_ | ~new_n3289_;
  assign po0151 = ~new_n3292_ | ~new_n3291_;
  assign po0152 = ~new_n3294_ | ~new_n3293_;
  assign po0153 = ~new_n3296_ | ~new_n3295_;
  assign po0154 = ~new_n3298_ | ~new_n3297_;
  assign po0155 = ~new_n3300_ | ~new_n3299_;
  assign po0156 = ~new_n3302_ | ~new_n3301_;
  assign po0157 = ~new_n3304_ | ~new_n3303_;
  assign po0158 = ~new_n3306_ | ~new_n3305_;
  assign po0159 = ~new_n3308_ | ~new_n3307_;
  assign po0160 = ~new_n3310_ | ~new_n3309_;
  assign new_n3045_ = ~new_n3312_ | ~new_n3311_;
  assign new_n3046_ = ~new_n3314_ | ~new_n3313_;
  assign new_n3047_ = ~new_n3316_ | ~new_n3315_;
  assign new_n3048_ = ~new_n3318_ | ~new_n3317_;
  assign new_n3049_ = ~new_n3320_ | ~new_n3319_;
  assign new_n3050_ = ~new_n3322_ | ~new_n3321_;
  assign new_n3051_ = ~new_n3324_ | ~new_n3323_;
  assign new_n3052_ = ~new_n3326_ | ~new_n3325_;
  assign new_n3053_ = ~new_n3328_ | ~new_n3327_;
  assign new_n3054_ = ~new_n3330_ | ~new_n3329_;
  assign new_n3055_ = ~new_n3332_ | ~new_n3331_;
  assign new_n3056_ = ~new_n3334_ | ~new_n3333_;
  assign new_n3057_ = ~new_n3336_ | ~new_n3335_;
  assign new_n3058_ = ~new_n3338_ | ~new_n3337_;
  assign new_n3059_ = ~new_n3340_ | ~new_n3339_;
  assign new_n3060_ = ~new_n3342_ | ~new_n3341_;
  assign new_n3061_ = ~new_n3344_ | ~new_n3343_;
  assign new_n3062_ = ~new_n3346_ | ~new_n3345_;
  assign new_n3063_ = ~new_n3348_ | ~new_n3347_;
  assign new_n3064_ = ~new_n3350_ | ~new_n3349_;
  assign new_n3065_ = ~new_n3352_ | ~new_n3351_;
  assign new_n3066_ = ~new_n3354_ | ~new_n3353_;
  assign new_n3067_ = ~new_n3356_ | ~new_n3355_;
  assign new_n3068_ = ~new_n3358_ | ~new_n3357_;
  assign new_n3069_ = ~new_n3360_ | ~new_n3359_;
  assign new_n3070_ = ~new_n3362_ | ~new_n3361_;
  assign new_n3071_ = ~new_n3364_ | ~new_n3363_;
  assign new_n3072_ = ~new_n3366_ | ~new_n3365_;
  assign new_n3073_ = ~new_n3368_ | ~new_n3367_;
  assign new_n3074_ = ~new_n3370_ | ~new_n3369_;
  assign new_n3075_ = ~new_n3372_ | ~new_n3371_;
  assign new_n3076_ = ~new_n3374_ | ~new_n3373_;
  assign new_n3077_ = ~new_n3376_ | ~new_n3375_;
  assign new_n3078_ = ~new_n3378_ | ~new_n3377_;
  assign new_n3079_ = ~new_n3380_ | ~new_n3379_;
  assign new_n3080_ = ~new_n3382_ | ~new_n3381_;
  assign new_n3081_ = ~new_n3384_ | ~new_n3383_;
  assign new_n3082_ = ~new_n3386_ | ~new_n3385_;
  assign new_n3083_ = ~new_n3388_ | ~new_n3387_;
  assign new_n3084_ = ~new_n3390_ | ~new_n3389_;
  assign new_n3085_ = ~new_n3392_ | ~new_n3391_;
  assign new_n3086_ = ~new_n3394_ | ~new_n3393_;
  assign new_n3087_ = ~new_n3396_ | ~new_n3395_;
  assign new_n3088_ = ~new_n3398_ | ~new_n3397_;
  assign new_n3089_ = ~new_n3400_ | ~new_n3399_;
  assign new_n3090_ = ~new_n3402_ | ~new_n3401_;
  assign new_n3091_ = ~new_n3404_ | ~new_n3403_;
  assign new_n3092_ = ~new_n3406_ | ~new_n3405_;
  assign new_n3093_ = ~new_n3408_ | ~new_n3407_;
  assign new_n3094_ = ~new_n3410_ | ~new_n3409_;
  assign new_n3095_ = ~new_n3412_ | ~new_n3411_;
  assign new_n3096_ = ~new_n3414_ | ~new_n3413_;
  assign new_n3097_ = ~new_n3416_ | ~new_n3415_;
  assign new_n3098_ = ~new_n3418_ | ~new_n3417_;
  assign new_n3099_ = ~new_n3420_ | ~new_n3419_;
  assign new_n3100_ = ~new_n3422_ | ~new_n3421_;
  assign new_n3101_ = ~new_n3424_ | ~new_n3423_;
  assign new_n3102_ = ~new_n3426_ | ~new_n3425_;
  assign new_n3103_ = ~new_n3428_ | ~new_n3427_;
  assign new_n3104_ = ~new_n3430_ | ~new_n3429_;
  assign new_n3105_ = ~new_n3432_ | ~new_n3431_;
  assign new_n3106_ = ~new_n3434_ | ~new_n3433_;
  assign new_n3107_ = ~new_n3436_ | ~new_n3435_;
  assign new_n3108_ = ~new_n3438_ | ~new_n3437_;
  assign po0082 = ~new_n3440_ | ~new_n3439_;
  assign po0083 = ~new_n3442_ | ~new_n3441_;
  assign po0084 = ~new_n3444_ | ~new_n3443_;
  assign po0085 = ~new_n3446_ | ~new_n3445_;
  assign po0086 = ~new_n3448_ | ~new_n3447_;
  assign po0087 = ~new_n3450_ | ~new_n3449_;
  assign po0088 = ~new_n3452_ | ~new_n3451_;
  assign po0089 = ~new_n3454_ | ~new_n3453_;
  assign po0062 = ~new_n3456_ | ~new_n3455_;
  assign po0063 = ~new_n3458_ | ~new_n3457_;
  assign po0064 = ~new_n3460_ | ~new_n3459_;
  assign po0065 = ~new_n3462_ | ~new_n3461_;
  assign po0066 = ~new_n3464_ | ~new_n3463_;
  assign po0067 = ~new_n3466_ | ~new_n3465_;
  assign po0068 = ~new_n3468_ | ~new_n3467_;
  assign po0069 = ~new_n3470_ | ~new_n3469_;
  assign po0070 = ~new_n3472_ | ~new_n3471_;
  assign po0071 = ~new_n3474_ | ~new_n3473_;
  assign po0090 = ~new_n3476_ | ~new_n3475_;
  assign po0072 = ~new_n3478_ | ~new_n3477_;
  assign po0073 = ~new_n3480_ | ~new_n3479_;
  assign po0074 = ~new_n3482_ | ~new_n3481_;
  assign po0075 = ~new_n3484_ | ~new_n3483_;
  assign po0076 = ~new_n3486_ | ~new_n3485_;
  assign po0077 = ~new_n3488_ | ~new_n3487_;
  assign po0078 = ~new_n3490_ | ~new_n3489_;
  assign po0079 = ~new_n3492_ | ~new_n3491_;
  assign po0080 = ~new_n3494_ | ~new_n3493_;
  assign po0081 = ~new_n3496_ | ~new_n3495_;
  assign po0091 = ~new_n3498_ | ~new_n3497_;
  assign new_n3139_ = ~pi1001 & ~pi0558 & ~pi0557 & ~pi0556;
  assign new_n3140_ = ~pi0998 & ~pi0555;
  assign new_n3141_ = ~pi0109 & ~pi0108 & ~pi0552 & ~pi0544 & ~pi0549;
  assign new_n3142_ = ~pi0106 & ~pi0107;
  assign new_n3143_ = ~pi1004 & ~pi1006 & ~pi1447 & ~pi1007 & ~pi1450;
  assign new_n3144_ = ~new_n21028_ | ~new_n21003_ | ~new_n21005_;
  assign new_n3145_ = ~pi1005;
  assign new_n3146_ = ~new_n3144_;
  assign new_n3147_ = ~po0164;
  assign new_n3148_ = ~po0162;
  assign new_n3149_ = ~new_n21008_ | ~new_n2970_;
  assign new_n3150_ = ~new_n3012_;
  assign new_n3151_ = ~pi0861 | ~new_n2969_;
  assign new_n3152_ = ~pi1310 | ~new_n3147_;
  assign new_n3153_ = ~pi0038 | ~new_n3150_;
  assign new_n3154_ = ~pi0862 | ~new_n2969_;
  assign new_n3155_ = ~pi1311 | ~new_n3147_;
  assign new_n3156_ = ~pi0039 | ~new_n3150_;
  assign new_n3157_ = ~pi0863 | ~new_n2969_;
  assign new_n3158_ = ~pi1312 | ~new_n3147_;
  assign new_n3159_ = ~pi0040 | ~new_n3150_;
  assign new_n3160_ = ~pi0864 | ~new_n2969_;
  assign new_n3161_ = ~pi1313 | ~new_n3147_;
  assign new_n3162_ = ~pi0041 | ~new_n3150_;
  assign new_n3163_ = ~pi0865 | ~new_n2969_;
  assign new_n3164_ = ~pi1314 | ~new_n3147_;
  assign new_n3165_ = ~pi0042 | ~new_n3150_;
  assign new_n3166_ = ~pi0866 | ~new_n2969_;
  assign new_n3167_ = ~pi1315 | ~new_n3147_;
  assign new_n3168_ = ~pi0043 | ~new_n3150_;
  assign new_n3169_ = ~pi0867 | ~new_n2969_;
  assign new_n3170_ = ~pi1316 | ~new_n3147_;
  assign new_n3171_ = ~pi0044 | ~new_n3150_;
  assign new_n3172_ = ~pi0868 | ~new_n2969_;
  assign new_n3173_ = ~pi1317 | ~new_n3147_;
  assign new_n3174_ = ~pi0045 | ~new_n3150_;
  assign new_n3175_ = ~pi0869 | ~new_n2969_;
  assign new_n3176_ = ~pi1318 | ~new_n3147_;
  assign new_n3177_ = ~pi0046 | ~new_n3150_;
  assign new_n3178_ = ~pi0870 | ~new_n2969_;
  assign new_n3179_ = ~pi1319 | ~new_n3147_;
  assign new_n3180_ = ~pi0047 | ~new_n3150_;
  assign new_n3181_ = ~pi0871 | ~new_n2969_;
  assign new_n3182_ = ~pi1320 | ~new_n3147_;
  assign new_n3183_ = ~pi0048 | ~new_n3150_;
  assign new_n3184_ = ~pi0872 | ~new_n2969_;
  assign new_n3185_ = ~pi1321 | ~new_n3147_;
  assign new_n3186_ = ~pi0049 | ~new_n3150_;
  assign new_n3187_ = ~pi0873 | ~new_n2969_;
  assign new_n3188_ = ~pi1322 | ~new_n3147_;
  assign new_n3189_ = ~pi0050 | ~new_n3150_;
  assign new_n3190_ = ~pi0874 | ~new_n2969_;
  assign new_n3191_ = ~pi1323 | ~new_n3147_;
  assign new_n3192_ = ~pi0051 | ~new_n3150_;
  assign new_n3193_ = ~pi0875 | ~new_n2969_;
  assign new_n3194_ = ~pi1324 | ~new_n3147_;
  assign new_n3195_ = ~pi0052 | ~new_n3150_;
  assign new_n3196_ = ~pi0876 | ~new_n2969_;
  assign new_n3197_ = ~pi1325 | ~new_n3147_;
  assign new_n3198_ = ~pi0053 | ~new_n3150_;
  assign new_n3199_ = ~pi0877 | ~new_n2969_;
  assign new_n3200_ = ~pi1326 | ~new_n3147_;
  assign new_n3201_ = ~pi0054 | ~new_n3150_;
  assign new_n3202_ = ~pi0878 | ~new_n2969_;
  assign new_n3203_ = ~pi1327 | ~new_n3147_;
  assign new_n3204_ = ~pi0055 | ~new_n3150_;
  assign new_n3205_ = ~pi0879 | ~new_n2969_;
  assign new_n3206_ = ~pi1328 | ~new_n3147_;
  assign new_n3207_ = ~pi0056 | ~new_n3150_;
  assign new_n3208_ = ~pi0880 | ~new_n2969_;
  assign new_n3209_ = ~pi1329 | ~new_n3147_;
  assign new_n3210_ = ~pi0057 | ~new_n3150_;
  assign new_n3211_ = ~pi0881 | ~new_n2969_;
  assign new_n3212_ = ~pi1330 | ~new_n3147_;
  assign new_n3213_ = ~pi0058 | ~new_n3150_;
  assign new_n3214_ = ~pi0882 | ~new_n2969_;
  assign new_n3215_ = ~pi1331 | ~new_n3147_;
  assign new_n3216_ = ~pi0059 | ~new_n3150_;
  assign new_n3217_ = ~pi0883 | ~new_n2969_;
  assign new_n3218_ = ~pi1332 | ~new_n3147_;
  assign new_n3219_ = ~pi0060 | ~new_n3150_;
  assign new_n3220_ = ~pi0884 | ~new_n2969_;
  assign new_n3221_ = ~pi1333 | ~new_n3147_;
  assign new_n3222_ = ~pi0061 | ~new_n3150_;
  assign new_n3223_ = ~pi0885 | ~new_n2969_;
  assign new_n3224_ = ~pi1334 | ~new_n3147_;
  assign new_n3225_ = ~pi0062 | ~new_n3150_;
  assign new_n3226_ = ~pi0886 | ~new_n2969_;
  assign new_n3227_ = ~pi1335 | ~new_n3147_;
  assign new_n3228_ = ~pi0063 | ~new_n3150_;
  assign new_n3229_ = ~pi0887 | ~new_n2969_;
  assign new_n3230_ = ~pi1336 | ~new_n3147_;
  assign new_n3231_ = ~pi0064 | ~new_n3150_;
  assign new_n3232_ = ~pi0888 | ~new_n2969_;
  assign new_n3233_ = ~pi1337 | ~new_n3147_;
  assign new_n3234_ = ~pi0065 | ~new_n3150_;
  assign new_n3235_ = ~pi0889 | ~new_n2969_;
  assign new_n3236_ = ~pi1338 | ~new_n3147_;
  assign new_n3237_ = ~pi0066 | ~new_n3150_;
  assign new_n3238_ = ~pi0890 | ~new_n2969_;
  assign new_n3239_ = ~pi1339 | ~new_n3147_;
  assign new_n3240_ = ~pi0067 | ~new_n3150_;
  assign new_n3241_ = ~pi0891 | ~new_n2969_;
  assign new_n3242_ = ~pi1340 | ~new_n3147_;
  assign new_n3243_ = ~pi0068 | ~new_n3150_;
  assign new_n3244_ = ~pi0892 | ~new_n2969_;
  assign new_n3245_ = ~pi1341 | ~new_n3147_;
  assign new_n3246_ = ~pi0069 | ~new_n3150_;
  assign new_n3247_ = ~pi0070 | ~po0162;
  assign new_n3248_ = ~pi0861 | ~new_n3148_;
  assign new_n3249_ = ~pi0071 | ~po0162;
  assign new_n3250_ = ~pi0862 | ~new_n3148_;
  assign new_n3251_ = ~pi0072 | ~po0162;
  assign new_n3252_ = ~pi0863 | ~new_n3148_;
  assign new_n3253_ = ~pi0073 | ~po0162;
  assign new_n3254_ = ~pi0864 | ~new_n3148_;
  assign new_n3255_ = ~pi0074 | ~po0162;
  assign new_n3256_ = ~pi0865 | ~new_n3148_;
  assign new_n3257_ = ~pi0075 | ~po0162;
  assign new_n3258_ = ~pi0866 | ~new_n3148_;
  assign new_n3259_ = ~pi0076 | ~po0162;
  assign new_n3260_ = ~pi0867 | ~new_n3148_;
  assign new_n3261_ = ~pi0077 | ~po0162;
  assign new_n3262_ = ~pi0868 | ~new_n3148_;
  assign new_n3263_ = ~pi0078 | ~po0162;
  assign new_n3264_ = ~pi0869 | ~new_n3148_;
  assign new_n3265_ = ~pi0079 | ~po0162;
  assign new_n3266_ = ~pi0870 | ~new_n3148_;
  assign new_n3267_ = ~pi0080 | ~po0162;
  assign new_n3268_ = ~pi0871 | ~new_n3148_;
  assign new_n3269_ = ~pi0081 | ~po0162;
  assign new_n3270_ = ~pi0872 | ~new_n3148_;
  assign new_n3271_ = ~pi0082 | ~po0162;
  assign new_n3272_ = ~pi0873 | ~new_n3148_;
  assign new_n3273_ = ~pi0083 | ~po0162;
  assign new_n3274_ = ~pi0874 | ~new_n3148_;
  assign new_n3275_ = ~pi0084 | ~po0162;
  assign new_n3276_ = ~pi0875 | ~new_n3148_;
  assign new_n3277_ = ~pi0085 | ~po0162;
  assign new_n3278_ = ~pi0876 | ~new_n3148_;
  assign new_n3279_ = ~pi0086 | ~po0162;
  assign new_n3280_ = ~pi0877 | ~new_n3148_;
  assign new_n3281_ = ~pi0087 | ~po0162;
  assign new_n3282_ = ~pi0878 | ~new_n3148_;
  assign new_n3283_ = ~pi0088 | ~po0162;
  assign new_n3284_ = ~pi0879 | ~new_n3148_;
  assign new_n3285_ = ~pi0089 | ~po0162;
  assign new_n3286_ = ~pi0880 | ~new_n3148_;
  assign new_n3287_ = ~pi0090 | ~po0162;
  assign new_n3288_ = ~pi0881 | ~new_n3148_;
  assign new_n3289_ = ~pi0091 | ~po0162;
  assign new_n3290_ = ~pi0882 | ~new_n3148_;
  assign new_n3291_ = ~pi0092 | ~po0162;
  assign new_n3292_ = ~pi0883 | ~new_n3148_;
  assign new_n3293_ = ~pi0093 | ~po0162;
  assign new_n3294_ = ~pi0884 | ~new_n3148_;
  assign new_n3295_ = ~pi0094 | ~po0162;
  assign new_n3296_ = ~pi0885 | ~new_n3148_;
  assign new_n3297_ = ~pi0095 | ~po0162;
  assign new_n3298_ = ~pi0886 | ~new_n3148_;
  assign new_n3299_ = ~pi0096 | ~po0162;
  assign new_n3300_ = ~pi0887 | ~new_n3148_;
  assign new_n3301_ = ~pi0097 | ~po0162;
  assign new_n3302_ = ~pi0888 | ~new_n3148_;
  assign new_n3303_ = ~pi0098 | ~po0162;
  assign new_n3304_ = ~pi0889 | ~new_n3148_;
  assign new_n3305_ = ~pi0099 | ~po0162;
  assign new_n3306_ = ~pi0890 | ~new_n3148_;
  assign new_n3307_ = ~pi0100 | ~po0162;
  assign new_n3308_ = ~pi0891 | ~new_n3148_;
  assign new_n3309_ = ~pi0101 | ~po0162;
  assign new_n3310_ = ~pi0892 | ~new_n3148_;
  assign new_n3311_ = ~pi0079 | ~new_n3011_;
  assign new_n3312_ = ~pi0047 | ~new_n21008_;
  assign new_n3313_ = ~pi0078 | ~new_n3011_;
  assign new_n3314_ = ~pi0046 | ~new_n21008_;
  assign new_n3315_ = ~pi0077 | ~new_n3011_;
  assign new_n3316_ = ~pi0045 | ~new_n21008_;
  assign new_n3317_ = ~pi0076 | ~new_n3011_;
  assign new_n3318_ = ~pi0044 | ~new_n21008_;
  assign new_n3319_ = ~pi0075 | ~new_n3011_;
  assign new_n3320_ = ~pi0043 | ~new_n21008_;
  assign new_n3321_ = ~pi0074 | ~new_n3011_;
  assign new_n3322_ = ~pi0042 | ~new_n21008_;
  assign new_n3323_ = ~pi0073 | ~new_n3011_;
  assign new_n3324_ = ~pi0041 | ~new_n21008_;
  assign new_n3325_ = ~pi0101 | ~new_n3011_;
  assign new_n3326_ = ~pi0069 | ~new_n21008_;
  assign new_n3327_ = ~pi0100 | ~new_n3011_;
  assign new_n3328_ = ~pi0068 | ~new_n21008_;
  assign new_n3329_ = ~pi0072 | ~new_n3011_;
  assign new_n3330_ = ~pi0040 | ~new_n21008_;
  assign new_n3331_ = ~pi0099 | ~new_n3011_;
  assign new_n3332_ = ~pi0067 | ~new_n21008_;
  assign new_n3333_ = ~pi0098 | ~new_n3011_;
  assign new_n3334_ = ~pi0066 | ~new_n21008_;
  assign new_n3335_ = ~pi0097 | ~new_n3011_;
  assign new_n3336_ = ~pi0065 | ~new_n21008_;
  assign new_n3337_ = ~pi0096 | ~new_n3011_;
  assign new_n3338_ = ~pi0064 | ~new_n21008_;
  assign new_n3339_ = ~pi0095 | ~new_n3011_;
  assign new_n3340_ = ~pi0063 | ~new_n21008_;
  assign new_n3341_ = ~pi0094 | ~new_n3011_;
  assign new_n3342_ = ~pi0062 | ~new_n21008_;
  assign new_n3343_ = ~pi0093 | ~new_n3011_;
  assign new_n3344_ = ~pi0061 | ~new_n21008_;
  assign new_n3345_ = ~pi0092 | ~new_n3011_;
  assign new_n3346_ = ~pi0060 | ~new_n21008_;
  assign new_n3347_ = ~pi0091 | ~new_n3011_;
  assign new_n3348_ = ~pi0059 | ~new_n21008_;
  assign new_n3349_ = ~pi0090 | ~new_n3011_;
  assign new_n3350_ = ~pi0058 | ~new_n21008_;
  assign new_n3351_ = ~pi0071 | ~new_n3011_;
  assign new_n3352_ = ~pi0039 | ~new_n21008_;
  assign new_n3353_ = ~pi0089 | ~new_n3011_;
  assign new_n3354_ = ~pi0057 | ~new_n21008_;
  assign new_n3355_ = ~pi0088 | ~new_n3011_;
  assign new_n3356_ = ~pi0056 | ~new_n21008_;
  assign new_n3357_ = ~pi0087 | ~new_n3011_;
  assign new_n3358_ = ~pi0055 | ~new_n21008_;
  assign new_n3359_ = ~pi0086 | ~new_n3011_;
  assign new_n3360_ = ~pi0054 | ~new_n21008_;
  assign new_n3361_ = ~pi0085 | ~new_n3011_;
  assign new_n3362_ = ~pi0053 | ~new_n21008_;
  assign new_n3363_ = ~pi0084 | ~new_n3011_;
  assign new_n3364_ = ~pi0052 | ~new_n21008_;
  assign new_n3365_ = ~pi0083 | ~new_n3011_;
  assign new_n3366_ = ~pi0051 | ~new_n21008_;
  assign new_n3367_ = ~pi0082 | ~new_n3011_;
  assign new_n3368_ = ~pi0050 | ~new_n21008_;
  assign new_n3369_ = ~pi0081 | ~new_n3011_;
  assign new_n3370_ = ~pi0049 | ~new_n21008_;
  assign new_n3371_ = ~pi0080 | ~new_n3011_;
  assign new_n3372_ = ~pi0048 | ~new_n21008_;
  assign new_n3373_ = ~pi0070 | ~new_n3011_;
  assign new_n3374_ = ~pi0038 | ~new_n21008_;
  assign new_n3375_ = ~pi0023 | ~new_n3010_;
  assign new_n3376_ = ~pi0047 | ~new_n21018_;
  assign new_n3377_ = ~pi0024 | ~new_n3010_;
  assign new_n3378_ = ~pi0046 | ~new_n21018_;
  assign new_n3379_ = ~pi0025 | ~new_n3010_;
  assign new_n3380_ = ~pi0045 | ~new_n21018_;
  assign new_n3381_ = ~pi0026 | ~new_n3010_;
  assign new_n3382_ = ~pi0044 | ~new_n21018_;
  assign new_n3383_ = ~pi0027 | ~new_n3010_;
  assign new_n3384_ = ~pi0043 | ~new_n21018_;
  assign new_n3385_ = ~pi0028 | ~new_n3010_;
  assign new_n3386_ = ~pi0042 | ~new_n21018_;
  assign new_n3387_ = ~pi0029 | ~new_n3010_;
  assign new_n3388_ = ~pi0041 | ~new_n21018_;
  assign new_n3389_ = ~pi0001 | ~new_n3010_;
  assign new_n3390_ = ~pi0069 | ~new_n21018_;
  assign new_n3391_ = ~pi0002 | ~new_n3010_;
  assign new_n3392_ = ~pi0068 | ~new_n21018_;
  assign new_n3393_ = ~pi0030 | ~new_n3010_;
  assign new_n3394_ = ~pi0040 | ~new_n21018_;
  assign new_n3395_ = ~pi0003 | ~new_n3010_;
  assign new_n3396_ = ~pi0067 | ~new_n21018_;
  assign new_n3397_ = ~pi0004 | ~new_n3010_;
  assign new_n3398_ = ~pi0066 | ~new_n21018_;
  assign new_n3399_ = ~pi0005 | ~new_n3010_;
  assign new_n3400_ = ~pi0065 | ~new_n21018_;
  assign new_n3401_ = ~pi0006 | ~new_n3010_;
  assign new_n3402_ = ~pi0064 | ~new_n21018_;
  assign new_n3403_ = ~pi0007 | ~new_n3010_;
  assign new_n3404_ = ~pi0063 | ~new_n21018_;
  assign new_n3405_ = ~pi0008 | ~new_n3010_;
  assign new_n3406_ = ~pi0062 | ~new_n21018_;
  assign new_n3407_ = ~pi0009 | ~new_n3010_;
  assign new_n3408_ = ~pi0061 | ~new_n21018_;
  assign new_n3409_ = ~pi0010 | ~new_n3010_;
  assign new_n3410_ = ~pi0060 | ~new_n21018_;
  assign new_n3411_ = ~pi0011 | ~new_n3010_;
  assign new_n3412_ = ~pi0059 | ~new_n21018_;
  assign new_n3413_ = ~pi0012 | ~new_n3010_;
  assign new_n3414_ = ~pi0058 | ~new_n21018_;
  assign new_n3415_ = ~pi0031 | ~new_n3010_;
  assign new_n3416_ = ~pi0039 | ~new_n21018_;
  assign new_n3417_ = ~pi0013 | ~new_n3010_;
  assign new_n3418_ = ~pi0057 | ~new_n21018_;
  assign new_n3419_ = ~pi0014 | ~new_n3010_;
  assign new_n3420_ = ~pi0056 | ~new_n21018_;
  assign new_n3421_ = ~pi0015 | ~new_n3010_;
  assign new_n3422_ = ~pi0055 | ~new_n21018_;
  assign new_n3423_ = ~pi0016 | ~new_n3010_;
  assign new_n3424_ = ~pi0054 | ~new_n21018_;
  assign new_n3425_ = ~pi0017 | ~new_n3010_;
  assign new_n3426_ = ~pi0053 | ~new_n21018_;
  assign new_n3427_ = ~pi0018 | ~new_n3010_;
  assign new_n3428_ = ~pi0052 | ~new_n21018_;
  assign new_n3429_ = ~pi0019 | ~new_n3010_;
  assign new_n3430_ = ~pi0051 | ~new_n21018_;
  assign new_n3431_ = ~pi0020 | ~new_n3010_;
  assign new_n3432_ = ~pi0050 | ~new_n21018_;
  assign new_n3433_ = ~pi0021 | ~new_n3010_;
  assign new_n3434_ = ~pi0049 | ~new_n21018_;
  assign new_n3435_ = ~pi0022 | ~new_n3010_;
  assign new_n3436_ = ~pi0048 | ~new_n21018_;
  assign new_n3437_ = ~pi0032 | ~new_n3010_;
  assign new_n3438_ = ~pi0038 | ~new_n21018_;
  assign new_n3439_ = ~pi0579 | ~new_n3144_;
  assign new_n3440_ = ~pi0130 | ~new_n3146_;
  assign new_n3441_ = ~pi0580 | ~new_n3144_;
  assign new_n3442_ = ~pi0131 | ~new_n3146_;
  assign new_n3443_ = ~pi0581 | ~new_n3144_;
  assign new_n3444_ = ~pi0132 | ~new_n3146_;
  assign new_n3445_ = ~pi0582 | ~new_n3144_;
  assign new_n3446_ = ~pi0133 | ~new_n3146_;
  assign new_n3447_ = ~pi0583 | ~new_n3144_;
  assign new_n3448_ = ~pi0134 | ~new_n3146_;
  assign new_n3449_ = ~pi0584 | ~new_n3144_;
  assign new_n3450_ = ~pi0135 | ~new_n3146_;
  assign new_n3451_ = ~pi0585 | ~new_n3144_;
  assign new_n3452_ = ~pi0136 | ~new_n3146_;
  assign new_n3453_ = ~pi0586 | ~new_n3144_;
  assign new_n3454_ = ~pi0137 | ~new_n3146_;
  assign new_n3455_ = ~pi0559 | ~new_n3144_;
  assign new_n3456_ = ~pi0110 | ~new_n3146_;
  assign new_n3457_ = ~pi0560 | ~new_n3144_;
  assign new_n3458_ = ~pi0111 | ~new_n3146_;
  assign new_n3459_ = ~pi0561 | ~new_n3144_;
  assign new_n3460_ = ~pi0112 | ~new_n3146_;
  assign new_n3461_ = ~pi0562 | ~new_n3144_;
  assign new_n3462_ = ~pi0113 | ~new_n3146_;
  assign new_n3463_ = ~pi0563 | ~new_n3144_;
  assign new_n3464_ = ~pi0114 | ~new_n3146_;
  assign new_n3465_ = ~pi0564 | ~new_n3144_;
  assign new_n3466_ = ~pi0115 | ~new_n3146_;
  assign new_n3467_ = ~pi0565 | ~new_n3144_;
  assign new_n3468_ = ~pi0116 | ~new_n3146_;
  assign new_n3469_ = ~pi0566 | ~new_n3144_;
  assign new_n3470_ = ~pi0117 | ~new_n3146_;
  assign new_n3471_ = ~pi0567 | ~new_n3144_;
  assign new_n3472_ = ~pi0118 | ~new_n3146_;
  assign new_n3473_ = ~pi0568 | ~new_n3144_;
  assign new_n3474_ = ~pi0119 | ~new_n3146_;
  assign new_n3475_ = ~pi0587 | ~new_n3144_;
  assign new_n3476_ = ~pi0138 | ~new_n3146_;
  assign new_n3477_ = ~pi0569 | ~new_n3144_;
  assign new_n3478_ = ~pi0120 | ~new_n3146_;
  assign new_n3479_ = ~pi0570 | ~new_n3144_;
  assign new_n3480_ = ~pi0121 | ~new_n3146_;
  assign new_n3481_ = ~pi0571 | ~new_n3144_;
  assign new_n3482_ = ~pi0122 | ~new_n3146_;
  assign new_n3483_ = ~pi0572 | ~new_n3144_;
  assign new_n3484_ = ~pi0123 | ~new_n3146_;
  assign new_n3485_ = ~pi0573 | ~new_n3144_;
  assign new_n3486_ = ~pi0124 | ~new_n3146_;
  assign new_n3487_ = ~pi0574 | ~new_n3144_;
  assign new_n3488_ = ~pi0125 | ~new_n3146_;
  assign new_n3489_ = ~pi0575 | ~new_n3144_;
  assign new_n3490_ = ~pi0126 | ~new_n3146_;
  assign new_n3491_ = ~pi0576 | ~new_n3144_;
  assign new_n3492_ = ~pi0127 | ~new_n3146_;
  assign new_n3493_ = ~pi0577 | ~new_n3144_;
  assign new_n3494_ = ~pi0128 | ~new_n3146_;
  assign new_n3495_ = ~pi0578 | ~new_n3144_;
  assign new_n3496_ = ~pi0129 | ~new_n3146_;
  assign new_n3497_ = ~pi0588 | ~new_n3144_;
  assign new_n3498_ = ~pi0139 | ~new_n3146_;
  assign new_n3499_ = ~pi1240 | ~new_n9330_;
  assign new_n3500_ = ~new_n9282_ | ~new_n9365_;
  assign new_n3501_ = ~pi1222 | ~new_n9366_;
  assign new_n3502_ = ~new_n9277_ | ~new_n9355_;
  assign new_n3503_ = ~pi1227 | ~new_n9356_;
  assign new_n3504_ = ~new_n9268_ | ~new_n9337_;
  assign new_n3505_ = ~pi1236 | ~new_n9338_;
  assign new_n3506_ = ~new_n9261_ | ~new_n9323_;
  assign new_n3507_ = ~pi1243 | ~new_n9324_;
  assign new_n3508_ = ~new_n2971_ & ~pi0547;
  assign new_n3509_ = new_n4510_ & new_n3605_;
  assign new_n3510_ = new_n4844_ & new_n5481_;
  assign new_n3511_ = new_n4845_ & new_n5481_;
  assign new_n3512_ = new_n4511_ & new_n3509_;
  assign new_n3513_ = new_n5479_ & new_n3607_;
  assign new_n3514_ = new_n4846_ & new_n5497_;
  assign new_n3515_ = new_n5480_ & new_n3618_;
  assign new_n3516_ = new_n5452_ & new_n3618_;
  assign new_n3517_ = new_n5453_ & new_n3618_;
  assign new_n3518_ = new_n4847_ & new_n5497_;
  assign new_n3519_ = new_n6598_ & new_n6591_;
  assign new_n3520_ = new_n6548_ & new_n4360_;
  assign new_n3521_ = new_n6497_ & new_n4357_;
  assign new_n3522_ = new_n6446_ & new_n4354_;
  assign new_n3523_ = new_n6395_ & new_n6388_;
  assign new_n3524_ = new_n6345_ & new_n4349_;
  assign new_n3525_ = new_n6293_ & new_n4345_;
  assign new_n3526_ = new_n6241_ & new_n4341_;
  assign new_n3527_ = new_n6192_ & new_n6184_;
  assign new_n3528_ = new_n6141_ & new_n4332_;
  assign new_n3529_ = new_n6089_ & new_n4328_;
  assign new_n3530_ = new_n6037_ & new_n4324_;
  assign new_n3531_ = new_n5985_ & new_n5977_;
  assign new_n3532_ = new_n5934_ & new_n4316_;
  assign new_n3533_ = new_n5882_ & new_n4308_;
  assign new_n3534_ = new_n5830_ & new_n4302_;
  assign new_n3535_ = new_n5478_ & new_n5468_;
  assign new_n3536_ = pi0176 & new_n4416_;
  assign new_n3537_ = new_n5468_ & pi0175;
  assign new_n3538_ = new_n5107_ & new_n4405_;
  assign new_n3539_ = new_n3536_ & new_n5452_;
  assign new_n3540_ = new_n3536_ & new_n5453_;
  assign new_n3541_ = pi0177 & new_n4416_;
  assign new_n3542_ = pi0177 & new_n4405_;
  assign new_n3543_ = new_n5109_ & new_n4405_;
  assign new_n3544_ = new_n5108_ & new_n4405_;
  assign new_n3545_ = new_n5510_ & new_n4405_;
  assign new_n3546_ = new_n5509_ & pi0178;
  assign new_n3547_ = new_n5466_ & new_n4374_;
  assign new_n3548_ = new_n3539_ & new_n5449_;
  assign new_n3549_ = new_n3784_ & new_n3517_;
  assign new_n3550_ = new_n3538_ & new_n3784_;
  assign new_n3551_ = new_n3517_ & new_n4397_;
  assign new_n3552_ = new_n3538_ & new_n4397_;
  assign new_n3553_ = new_n3542_ & pi0547;
  assign new_n3554_ = new_n3542_ & new_n3787_;
  assign new_n3555_ = new_n5465_ & new_n5729_;
  assign new_n3556_ = new_n5466_ & new_n5729_;
  assign new_n3557_ = pi0175 & new_n4416_;
  assign new_n3558_ = new_n4404_ & new_n4246_;
  assign new_n3559_ = new_n3541_ & new_n4414_;
  assign new_n3560_ = new_n3540_ & new_n4413_;
  assign new_n3561_ = new_n8251_ & new_n3540_;
  assign new_n3562_ = new_n5467_ & new_n4260_;
  assign new_n3563_ = new_n5467_ & new_n5661_;
  assign new_n3564_ = new_n5465_ & new_n4374_;
  assign new_n3565_ = pi0178 & new_n4407_;
  assign new_n3566_ = new_n4407_ & new_n4277_;
  assign new_n3567_ = new_n5466_ & new_n5764_;
  assign new_n3568_ = new_n5695_ & new_n4374_ & new_n4263_;
  assign new_n3569_ = pi0070 & new_n5468_;
  assign new_n3570_ = pi0071 & new_n5468_;
  assign new_n3571_ = pi0072 & new_n5468_;
  assign new_n3572_ = pi0073 & new_n5468_;
  assign new_n3573_ = pi0074 & new_n5468_;
  assign new_n3574_ = pi0075 & new_n5468_;
  assign new_n3575_ = pi0076 & new_n5468_;
  assign new_n3576_ = pi0077 & new_n5468_;
  assign new_n3577_ = pi0094 & new_n3535_;
  assign new_n3578_ = pi0086 & new_n3535_;
  assign new_n3579_ = pi0095 & new_n3535_;
  assign new_n3580_ = pi0087 & new_n3535_;
  assign new_n3581_ = pi0096 & new_n3535_;
  assign new_n3582_ = pi0088 & new_n3535_;
  assign new_n3583_ = pi0097 & new_n3535_;
  assign new_n3584_ = pi0089 & new_n3535_;
  assign new_n3585_ = pi0098 & new_n3535_;
  assign new_n3586_ = pi0090 & new_n3535_;
  assign new_n3587_ = pi0099 & new_n3535_;
  assign new_n3588_ = pi0091 & new_n3535_;
  assign new_n3589_ = pi0100 & new_n3535_;
  assign new_n3590_ = pi0092 & new_n3535_;
  assign new_n3591_ = pi0101 & new_n3535_;
  assign new_n3592_ = pi0093 & new_n3535_;
  assign new_n3593_ = new_n3537_ & new_n4264_;
  assign new_n3594_ = new_n3537_ & new_n4260_;
  assign new_n3595_ = new_n3537_ & new_n4257_;
  assign new_n3596_ = new_n3537_ & new_n4263_;
  assign new_n3597_ = new_n3537_ & new_n4258_;
  assign new_n3598_ = new_n3537_ & new_n4266_;
  assign new_n3599_ = new_n3537_ & new_n4230_;
  assign new_n3600_ = new_n3547_ & new_n4230_;
  assign new_n3601_ = new_n3537_ & new_n4374_;
  assign new_n3602_ = new_n3547_ & new_n4269_;
  assign new_n3603_ = new_n3565_ & new_n4264_;
  assign new_n3604_ = new_n3547_ & new_n5746_;
  assign new_n3605_ = new_n5500_ & new_n5678_;
  assign new_n3606_ = new_n4816_ & new_n5507_;
  assign new_n3607_ = new_n3568_ & new_n5764_ & new_n4258_;
  assign new_n3608_ = new_n3568_ & new_n3619_ & new_n5678_;
  assign new_n3609_ = pi0176 & pi0177;
  assign new_n3610_ = new_n3536_ & new_n5479_;
  assign new_n3611_ = new_n3536_ & new_n5480_;
  assign new_n3612_ = new_n5712_ & new_n5763_;
  assign new_n3613_ = new_n4425_ & new_n4295_;
  assign new_n3614_ = new_n5808_ & new_n4425_;
  assign new_n3615_ = new_n9118_ & new_n4295_;
  assign new_n3616_ = new_n9118_ & new_n5808_;
  assign new_n3617_ = new_n5729_ & new_n5678_;
  assign new_n3618_ = new_n3568_ & new_n3605_;
  assign new_n3619_ = new_n5746_ & new_n5763_;
  assign new_n3620_ = pi0308 & pi0309;
  assign new_n3621_ = new_n3620_ & new_n5488_;
  assign new_n3622_ = pi0310 & new_n4249_;
  assign new_n3623_ = new_n3620_ & new_n3622_;
  assign new_n3624_ = pi0311 & new_n4250_;
  assign new_n3625_ = new_n3620_ & new_n3624_;
  assign new_n3626_ = new_n3620_ & new_n5623_;
  assign new_n3627_ = pi0308 & new_n5624_;
  assign new_n3628_ = new_n3622_ & new_n4253_;
  assign new_n3629_ = new_n3628_ & pi0308;
  assign new_n3630_ = new_n3624_ & new_n4253_;
  assign new_n3631_ = new_n3630_ & pi0308;
  assign new_n3632_ = pi0308 & new_n5625_;
  assign new_n3633_ = new_n5626_ & new_n3622_;
  assign new_n3634_ = new_n5626_ & new_n3624_;
  assign new_n3635_ = new_n5626_ & new_n5623_;
  assign new_n3636_ = new_n5624_ & new_n4256_;
  assign new_n3637_ = ~pi0308 & ~pi0309;
  assign new_n3638_ = new_n3622_ & new_n3637_;
  assign new_n3639_ = new_n3624_ & new_n3637_;
  assign new_n3640_ = new_n5625_ & new_n4256_;
  assign new_n3641_ = new_n5812_ & new_n4426_;
  assign new_n3642_ = new_n4427_ & new_n4338_;
  assign new_n3643_ = new_n4426_ & new_n4298_;
  assign new_n3644_ = new_n5813_ & new_n3643_;
  assign new_n3645_ = new_n4246_ & new_n5471_;
  assign new_n3646_ = pi0316 & new_n4312_;
  assign new_n3647_ = new_n5800_ & new_n3643_;
  assign new_n3648_ = pi0314 & new_n4284_;
  assign new_n3649_ = new_n5802_ & new_n4284_;
  assign new_n3650_ = new_n5801_ & new_n3643_;
  assign new_n3651_ = new_n5802_ & pi0316;
  assign new_n3652_ = new_n5799_ & new_n4284_;
  assign new_n3653_ = new_n3652_ & new_n3643_;
  assign new_n3654_ = new_n9124_ & new_n4338_;
  assign new_n3655_ = new_n5814_ & new_n5813_;
  assign new_n3656_ = new_n5814_ & new_n5800_;
  assign new_n3657_ = ~pi0316 & ~pi0314;
  assign new_n3658_ = new_n5814_ & new_n5801_;
  assign new_n3659_ = new_n5814_ & new_n3652_;
  assign new_n3660_ = new_n5816_ & new_n4427_;
  assign new_n3661_ = new_n5800_ & new_n3641_;
  assign new_n3662_ = new_n5801_ & new_n3641_;
  assign new_n3663_ = new_n3652_ & new_n3641_;
  assign new_n3664_ = new_n5816_ & new_n9124_;
  assign new_n3665_ = new_n9121_ & new_n5812_;
  assign new_n3666_ = new_n3665_ & new_n5813_;
  assign new_n3667_ = new_n3665_ & new_n5800_;
  assign new_n3668_ = new_n3665_ & new_n5801_;
  assign new_n3669_ = new_n3665_ & new_n3652_;
  assign new_n3670_ = new_n4374_ & new_n4372_;
  assign new_n3671_ = new_n6641_ & new_n9126_ & new_n9125_;
  assign new_n3672_ = new_n6649_ & new_n6648_;
  assign new_n3673_ = new_n4402_ & new_n6682_;
  assign new_n3674_ = new_n4824_ & new_n6678_;
  assign new_n3675_ = pi0311 & new_n4384_;
  assign new_n3676_ = new_n6699_ & new_n6704_;
  assign new_n3677_ = new_n3676_ & new_n3675_;
  assign new_n3678_ = new_n4249_ & new_n4384_;
  assign new_n3679_ = new_n3676_ & new_n3678_;
  assign new_n3680_ = new_n6714_ & pi0311;
  assign new_n3681_ = new_n3676_ & new_n3680_;
  assign new_n3682_ = new_n6714_ & new_n4249_;
  assign new_n3683_ = new_n3676_ & new_n3682_;
  assign new_n3684_ = new_n6699_ & new_n4381_;
  assign new_n3685_ = new_n3684_ & new_n3675_;
  assign new_n3686_ = new_n3684_ & new_n3678_;
  assign new_n3687_ = new_n3684_ & new_n3680_;
  assign new_n3688_ = new_n3684_ & new_n3682_;
  assign new_n3689_ = new_n6704_ & new_n4421_;
  assign new_n3690_ = new_n3689_ & new_n3675_;
  assign new_n3691_ = new_n3689_ & new_n3678_;
  assign new_n3692_ = new_n3689_ & new_n3680_;
  assign new_n3693_ = new_n3689_ & new_n3682_;
  assign new_n3694_ = new_n4421_ & new_n4381_;
  assign new_n3695_ = new_n3675_ & new_n3694_;
  assign new_n3696_ = new_n3678_ & new_n3694_;
  assign new_n3697_ = new_n3680_ & new_n3694_;
  assign new_n3698_ = new_n3682_ & new_n3694_;
  assign new_n3699_ = new_n4428_ & new_n4422_;
  assign new_n3700_ = new_n3699_ & new_n3624_;
  assign new_n3701_ = new_n3699_ & new_n5623_;
  assign new_n3702_ = new_n3699_ & new_n5488_;
  assign new_n3703_ = new_n3699_ & new_n3622_;
  assign new_n3704_ = new_n9190_ & new_n4422_;
  assign new_n3705_ = new_n3704_ & new_n3624_;
  assign new_n3706_ = new_n3704_ & new_n5623_;
  assign new_n3707_ = new_n3704_ & new_n5488_;
  assign new_n3708_ = new_n3704_ & new_n3622_;
  assign new_n3709_ = new_n8672_ & new_n4428_;
  assign new_n3710_ = new_n3709_ & new_n3624_;
  assign new_n3711_ = new_n3709_ & new_n5623_;
  assign new_n3712_ = new_n3709_ & new_n5488_;
  assign new_n3713_ = new_n3709_ & new_n3622_;
  assign new_n3714_ = new_n8672_ & new_n9190_;
  assign new_n3715_ = new_n3714_ & new_n3624_;
  assign new_n3716_ = new_n3714_ & new_n5623_;
  assign new_n3717_ = new_n3714_ & new_n5488_;
  assign new_n3718_ = new_n3714_ & new_n3622_;
  assign new_n3719_ = new_n9193_ & new_n5447_;
  assign new_n3720_ = new_n3719_ & new_n3678_;
  assign new_n3721_ = new_n3719_ & new_n3675_;
  assign new_n3722_ = new_n3719_ & new_n3682_;
  assign new_n3723_ = new_n3719_ & new_n3680_;
  assign new_n3724_ = new_n9193_ & new_n4423_;
  assign new_n3725_ = new_n3724_ & new_n3678_;
  assign new_n3726_ = new_n3724_ & new_n3675_;
  assign new_n3727_ = new_n3724_ & new_n3682_;
  assign new_n3728_ = new_n3724_ & new_n3680_;
  assign new_n3729_ = new_n5447_ & new_n4429_;
  assign new_n3730_ = new_n3729_ & new_n3678_;
  assign new_n3731_ = new_n3729_ & new_n3675_;
  assign new_n3732_ = new_n3729_ & new_n3682_;
  assign new_n3733_ = new_n3729_ & new_n3680_;
  assign new_n3734_ = new_n4429_ & new_n4423_;
  assign new_n3735_ = new_n3734_ & new_n3678_;
  assign new_n3736_ = new_n3734_ & new_n3675_;
  assign new_n3737_ = new_n3734_ & new_n3682_;
  assign new_n3738_ = new_n3734_ & new_n3680_;
  assign new_n3739_ = new_n8931_ & new_n5624_;
  assign new_n3740_ = new_n8931_ & new_n3628_;
  assign new_n3741_ = new_n8931_ & new_n3630_;
  assign new_n3742_ = new_n8931_ & new_n5625_;
  assign new_n3743_ = new_n8931_ & pi0309;
  assign new_n3744_ = new_n3743_ & new_n5488_;
  assign new_n3745_ = new_n3743_ & new_n3622_;
  assign new_n3746_ = new_n3743_ & new_n3624_;
  assign new_n3747_ = new_n3743_ & new_n5623_;
  assign new_n3748_ = new_n5624_ & new_n4424_;
  assign new_n3749_ = new_n3628_ & new_n4424_;
  assign new_n3750_ = new_n3630_ & new_n4424_;
  assign new_n3751_ = new_n5625_ & new_n4424_;
  assign new_n3752_ = pi0309 & new_n4424_;
  assign new_n3753_ = new_n3752_ & new_n5488_;
  assign new_n3754_ = new_n3752_ & new_n3622_;
  assign new_n3755_ = new_n3752_ & new_n3624_;
  assign new_n3756_ = new_n3752_ & new_n5623_;
  assign new_n3757_ = new_n3548_ & new_n3508_;
  assign new_n3758_ = pi0507 & new_n3560_;
  assign new_n3759_ = new_n8514_ & new_n5289_ & new_n8515_ & new_n8516_;
  assign new_n3760_ = new_n9103_ & new_n9102_;
  assign new_n3761_ = ~new_n5370_ | ~new_n5368_ | ~new_n5369_ | ~new_n5371_;
  assign new_n3762_ = ~new_n5366_ | ~new_n5364_ | ~new_n5365_ | ~new_n5367_;
  assign new_n3763_ = ~new_n5362_ | ~new_n5360_ | ~new_n5361_ | ~new_n5363_;
  assign new_n3764_ = ~new_n5358_ | ~new_n5356_ | ~new_n5357_ | ~new_n5359_;
  assign new_n3765_ = ~new_n5354_ | ~new_n5352_ | ~new_n5353_ | ~new_n5355_;
  assign new_n3766_ = ~new_n5350_ | ~new_n5348_ | ~new_n5349_ | ~new_n5351_;
  assign new_n3767_ = ~new_n5346_ | ~new_n5344_ | ~new_n5345_ | ~new_n5347_;
  assign new_n3768_ = ~new_n5342_ | ~new_n5340_ | ~new_n5341_ | ~new_n5343_;
  assign new_n3769_ = ~new_n5434_ | ~new_n5432_ | ~new_n5433_ | ~new_n5435_;
  assign new_n3770_ = ~new_n5430_ | ~new_n5428_ | ~new_n5429_ | ~new_n5431_;
  assign new_n3771_ = ~new_n5426_ | ~new_n5424_ | ~new_n5425_ | ~new_n5427_;
  assign new_n3772_ = ~new_n5422_ | ~new_n5420_ | ~new_n5421_ | ~new_n5423_;
  assign new_n3773_ = ~new_n5418_ | ~new_n5416_ | ~new_n5417_ | ~new_n5419_;
  assign new_n3774_ = ~new_n5414_ | ~new_n5412_ | ~new_n5413_ | ~new_n5415_;
  assign new_n3775_ = ~new_n5410_ | ~new_n5408_ | ~new_n5409_ | ~new_n5411_;
  assign new_n3776_ = ~new_n5406_ | ~new_n5404_ | ~new_n5405_ | ~new_n5407_;
  assign new_n3777_ = ~new_n5338_ | ~new_n5336_ | ~new_n5337_ | ~new_n5339_;
  assign new_n3778_ = ~new_n5334_ | ~new_n5332_ | ~new_n5333_ | ~new_n5335_;
  assign new_n3779_ = ~new_n5330_ | ~new_n5328_ | ~new_n5329_ | ~new_n5331_;
  assign new_n3780_ = ~new_n5326_ | ~new_n5324_ | ~new_n5325_ | ~new_n5327_;
  assign new_n3781_ = ~new_n5322_ | ~new_n5320_ | ~new_n5321_ | ~new_n5323_;
  assign new_n3782_ = ~new_n5318_ | ~new_n5316_ | ~new_n5317_ | ~new_n5319_;
  assign new_n3783_ = ~new_n5314_ | ~new_n5312_ | ~new_n5313_ | ~new_n5315_;
  assign new_n3784_ = ~new_n5310_ | ~new_n5308_ | ~new_n5309_ | ~new_n5311_;
  assign new_n3785_ = pi0307 & new_n4363_;
  assign new_n3786_ = ~new_n2971_;
  assign new_n3787_ = ~pi0547;
  assign new_n3788_ = pi0308 & new_n4363_;
  assign po0611 = ~new_n9093_ | ~new_n8539_;
  assign po0610 = ~new_n8538_ | ~new_n8537_;
  assign po0608 = ~new_n5491_ | ~new_n9181_ | ~new_n9180_;
  assign po0606 = ~new_n5491_ | ~new_n9177_ | ~new_n9176_;
  assign po0604 = ~new_n8526_ | ~new_n8525_;
  assign po0601 = ~new_n5483_ | ~new_n9169_ | ~new_n9168_;
  assign po0599 = ~new_n5483_ | ~new_n9159_ | ~new_n9158_;
  assign po0598 = new_n8513_ & new_n9063_;
  assign po0597 = ~new_n8508_ | ~new_n5286_ | ~new_n8510_ | ~new_n5285_ | ~new_n8507_;
  assign po0596 = ~new_n8500_ | ~new_n5283_ | ~new_n8502_ | ~new_n5282_ | ~new_n8499_;
  assign po0595 = ~new_n8492_ | ~new_n5280_ | ~new_n8494_ | ~new_n5279_ | ~new_n8491_;
  assign po0594 = ~new_n8484_ | ~new_n5277_ | ~new_n8486_ | ~new_n5276_ | ~new_n8483_;
  assign po0593 = ~new_n8476_ | ~new_n5274_ | ~new_n8478_ | ~new_n5273_ | ~new_n8475_;
  assign po0592 = ~new_n8468_ | ~new_n5271_ | ~new_n8470_ | ~new_n5270_ | ~new_n8467_;
  assign po0591 = ~new_n8460_ | ~new_n5268_ | ~new_n8462_ | ~new_n5267_ | ~new_n8459_;
  assign po0590 = ~new_n8452_ | ~new_n5265_ | ~new_n8454_ | ~new_n5264_ | ~new_n8451_;
  assign po0589 = ~new_n8444_ | ~new_n5262_ | ~new_n8446_ | ~new_n5261_ | ~new_n8443_;
  assign po0588 = ~new_n8436_ | ~new_n5259_ | ~new_n8438_ | ~new_n5258_ | ~new_n8435_;
  assign po0587 = ~new_n8428_ | ~new_n5256_ | ~new_n8430_ | ~new_n5255_ | ~new_n8427_;
  assign po0586 = ~new_n8420_ | ~new_n5253_ | ~new_n8422_ | ~new_n5252_ | ~new_n8419_;
  assign po0585 = ~new_n8412_ | ~new_n5250_ | ~new_n8414_ | ~new_n5249_ | ~new_n8411_;
  assign po0584 = ~new_n8404_ | ~new_n5247_ | ~new_n8406_ | ~new_n5246_ | ~new_n8403_;
  assign po0583 = ~new_n8396_ | ~new_n5244_ | ~new_n8398_ | ~new_n5243_ | ~new_n8395_;
  assign po0582 = ~new_n8388_ | ~new_n5241_ | ~new_n8390_ | ~new_n5240_ | ~new_n8387_;
  assign po0581 = ~new_n8380_ | ~new_n5238_ | ~new_n8382_ | ~new_n5237_ | ~new_n8379_;
  assign po0580 = ~new_n8372_ | ~new_n5235_ | ~new_n8374_ | ~new_n5234_ | ~new_n8371_;
  assign po0579 = ~new_n8364_ | ~new_n5232_ | ~new_n8366_ | ~new_n5231_ | ~new_n8363_;
  assign po0578 = ~new_n8356_ | ~new_n5229_ | ~new_n8358_ | ~new_n5228_ | ~new_n8355_;
  assign po0577 = ~new_n8348_ | ~new_n5226_ | ~new_n8350_ | ~new_n5225_ | ~new_n8347_;
  assign po0576 = ~new_n8340_ | ~new_n5223_ | ~new_n8342_ | ~new_n5222_ | ~new_n8339_;
  assign po0575 = ~new_n8332_ | ~new_n5220_ | ~new_n8334_ | ~new_n5219_ | ~new_n8331_;
  assign po0574 = ~new_n8324_ | ~new_n5217_ | ~new_n8326_ | ~new_n5216_ | ~new_n8323_;
  assign po0573 = ~new_n8316_ | ~new_n5214_ | ~new_n8318_ | ~new_n5213_ | ~new_n8315_;
  assign po0572 = ~new_n5212_ | ~new_n5210_;
  assign po0571 = ~new_n5207_ | ~new_n5205_;
  assign po0570 = ~new_n8285_ | ~new_n5201_ | ~new_n8289_ | ~new_n8288_ | ~new_n5199_;
  assign po0569 = ~new_n8275_ | ~new_n5197_ | ~new_n8279_ | ~new_n8278_ | ~new_n5195_;
  assign po0568 = ~new_n8265_ | ~new_n5193_ | ~new_n8269_ | ~new_n8268_ | ~new_n5191_;
  assign po0567 = ~new_n8255_ | ~new_n5189_ | ~new_n8259_ | ~new_n8258_ | ~new_n5187_;
  assign po0566 = ~new_n8248_ | ~new_n8247_;
  assign po0565 = ~new_n8245_ | ~new_n8246_ | ~new_n8244_;
  assign po0564 = ~new_n8242_ | ~new_n8243_ | ~new_n8241_;
  assign po0563 = ~new_n8239_ | ~new_n8240_ | ~new_n8238_;
  assign po0562 = ~new_n8236_ | ~new_n8237_ | ~new_n8235_;
  assign po0561 = ~new_n8233_ | ~new_n8234_ | ~new_n8232_;
  assign po0560 = ~new_n8230_ | ~new_n8231_ | ~new_n8229_;
  assign po0559 = ~new_n8227_ | ~new_n8228_ | ~new_n8226_;
  assign po0558 = ~new_n8224_ | ~new_n8225_ | ~new_n8223_;
  assign po0557 = ~new_n8221_ | ~new_n8222_ | ~new_n8220_;
  assign po0556 = ~new_n8218_ | ~new_n8219_ | ~new_n8217_;
  assign po0555 = ~new_n8215_ | ~new_n8216_ | ~new_n8214_;
  assign po0554 = ~new_n8212_ | ~new_n8213_ | ~new_n8211_;
  assign po0553 = ~new_n8209_ | ~new_n8210_ | ~new_n8208_;
  assign po0552 = ~new_n8206_ | ~new_n8207_ | ~new_n8205_;
  assign po0551 = ~new_n8203_ | ~new_n8204_ | ~new_n8202_;
  assign po0550 = ~new_n8200_ | ~new_n8201_ | ~new_n8199_;
  assign po0549 = ~new_n8197_ | ~new_n8198_ | ~new_n8196_;
  assign po0548 = ~new_n8194_ | ~new_n8195_ | ~new_n8193_;
  assign po0547 = ~new_n8191_ | ~new_n8192_ | ~new_n8190_;
  assign po0546 = ~new_n8188_ | ~new_n8189_ | ~new_n8187_;
  assign po0545 = ~new_n8185_ | ~new_n8186_ | ~new_n8184_;
  assign po0544 = ~new_n8183_ | ~new_n8182_ | ~new_n8181_;
  assign po0543 = ~new_n8180_ | ~new_n8179_ | ~new_n8178_;
  assign po0542 = ~new_n8177_ | ~new_n8176_ | ~new_n8175_;
  assign po0541 = ~new_n8174_ | ~new_n8173_ | ~new_n8172_;
  assign po0540 = ~new_n8171_ | ~new_n8170_ | ~new_n8169_;
  assign po0539 = ~new_n8168_ | ~new_n8167_ | ~new_n8166_;
  assign po0538 = ~new_n8165_ | ~new_n8164_ | ~new_n8163_;
  assign po0537 = ~new_n8162_ | ~new_n8161_ | ~new_n8160_;
  assign po0536 = ~new_n8159_ | ~new_n8158_ | ~new_n8157_;
  assign po0535 = ~new_n8156_ | ~new_n8155_ | ~new_n8154_;
  assign po0534 = ~new_n8150_ | ~new_n8151_ | ~new_n8149_;
  assign po0533 = ~new_n8145_ | ~new_n8147_ | ~new_n8146_ | ~new_n8148_ | ~new_n8144_;
  assign po0532 = ~new_n8140_ | ~new_n8142_ | ~new_n8141_ | ~new_n8143_ | ~new_n8139_;
  assign po0531 = ~new_n8135_ | ~new_n8137_ | ~new_n8136_ | ~new_n8138_ | ~new_n8134_;
  assign po0530 = ~new_n8129_ | ~new_n8132_ | ~new_n5185_ | ~new_n8130_;
  assign po0529 = ~new_n8124_ | ~new_n8127_ | ~new_n5184_ | ~new_n8125_;
  assign po0528 = ~new_n8119_ | ~new_n8122_ | ~new_n5183_ | ~new_n8120_;
  assign po0527 = ~new_n8114_ | ~new_n8117_ | ~new_n5182_ | ~new_n8115_;
  assign po0526 = ~new_n8109_ | ~new_n8112_ | ~new_n5181_ | ~new_n8110_;
  assign po0525 = ~new_n8104_ | ~new_n8107_ | ~new_n5180_ | ~new_n8105_;
  assign po0524 = ~new_n8099_ | ~new_n8102_ | ~new_n5179_ | ~new_n8100_;
  assign po0523 = ~new_n8094_ | ~new_n8097_ | ~new_n5178_ | ~new_n8095_;
  assign po0522 = ~new_n8089_ | ~new_n8092_ | ~new_n5177_ | ~new_n8090_;
  assign po0521 = ~new_n8084_ | ~new_n8087_ | ~new_n5176_ | ~new_n8085_;
  assign po0520 = ~new_n8079_ | ~new_n8082_ | ~new_n5175_ | ~new_n8080_;
  assign po0519 = ~new_n8074_ | ~new_n8077_ | ~new_n5174_ | ~new_n8075_;
  assign po0518 = ~new_n8072_ | ~new_n8070_ | ~new_n5173_;
  assign po0517 = ~new_n8068_ | ~new_n8066_ | ~new_n5172_;
  assign po0516 = ~new_n8064_ | ~new_n8062_ | ~new_n5171_;
  assign po0515 = ~new_n5170_ | ~new_n8059_ | ~new_n8058_;
  assign po0514 = ~new_n5169_ | ~new_n8055_ | ~new_n8054_;
  assign po0513 = ~new_n5168_ | ~new_n8051_ | ~new_n8050_;
  assign po0512 = ~new_n5167_ | ~new_n8047_ | ~new_n8046_;
  assign po0511 = ~new_n5166_ | ~new_n8043_ | ~new_n8042_;
  assign po0510 = ~new_n5165_ | ~new_n8039_ | ~new_n8038_;
  assign po0509 = ~new_n5164_ | ~new_n8035_ | ~new_n8034_;
  assign po0508 = ~new_n5163_ | ~new_n8031_ | ~new_n8030_;
  assign po0507 = ~new_n5162_ | ~new_n8027_ | ~new_n8026_;
  assign po0506 = ~new_n5161_ | ~new_n8023_ | ~new_n8022_;
  assign po0505 = ~new_n5160_ | ~new_n8019_ | ~new_n8018_;
  assign po0504 = ~new_n5159_ | ~new_n8015_ | ~new_n8014_;
  assign po0503 = ~new_n5158_ | ~new_n8011_ | ~new_n8010_;
  assign po0502 = pi0443 & new_n7915_;
  assign po0501 = ~new_n5157_ | ~new_n8006_;
  assign po0500 = ~new_n5156_ | ~new_n8003_;
  assign po0499 = ~new_n5155_ | ~new_n8000_;
  assign po0498 = ~new_n5154_ | ~new_n7997_;
  assign po0497 = ~new_n5153_ | ~new_n7994_;
  assign po0496 = ~new_n5152_ | ~new_n7991_;
  assign po0495 = ~new_n5151_ | ~new_n7988_;
  assign po0494 = ~new_n5150_ | ~new_n7985_;
  assign po0493 = ~new_n5149_ | ~new_n7982_;
  assign po0492 = ~new_n5148_ | ~new_n7979_;
  assign po0491 = ~new_n5147_ | ~new_n7976_;
  assign po0490 = ~new_n5146_ | ~new_n7973_;
  assign po0489 = ~new_n5145_ | ~new_n7970_;
  assign po0488 = ~new_n5144_ | ~new_n7967_;
  assign po0487 = ~new_n5143_ | ~new_n7964_;
  assign po0486 = ~new_n7963_ | ~new_n7962_ | ~new_n7961_;
  assign po0485 = ~new_n7960_ | ~new_n7959_ | ~new_n7958_;
  assign po0484 = ~new_n7957_ | ~new_n7956_ | ~new_n7955_;
  assign po0483 = ~new_n7954_ | ~new_n7953_ | ~new_n7952_;
  assign po0482 = ~new_n7951_ | ~new_n7950_ | ~new_n7949_;
  assign po0481 = ~new_n7948_ | ~new_n7947_ | ~new_n7946_;
  assign po0480 = ~new_n7945_ | ~new_n7944_ | ~new_n7943_;
  assign po0479 = ~new_n7942_ | ~new_n7941_ | ~new_n7940_;
  assign po0478 = ~new_n7939_ | ~new_n7938_ | ~new_n7937_;
  assign po0477 = ~new_n7936_ | ~new_n7935_ | ~new_n7934_;
  assign po0476 = ~new_n7933_ | ~new_n7932_ | ~new_n7931_;
  assign po0475 = ~new_n7930_ | ~new_n7929_ | ~new_n7928_;
  assign po0474 = ~new_n7927_ | ~new_n7926_ | ~new_n7925_;
  assign po0473 = ~new_n7924_ | ~new_n7923_ | ~new_n7922_;
  assign po0472 = ~new_n7921_ | ~new_n7920_ | ~new_n7919_;
  assign po0471 = ~new_n7918_ | ~new_n7917_ | ~new_n7916_;
  assign po0470 = ~new_n7912_ | ~new_n7911_ | ~new_n7910_;
  assign po0469 = ~new_n7909_ | ~new_n7908_ | ~new_n7907_;
  assign po0468 = ~new_n7906_ | ~new_n7905_ | ~new_n7904_;
  assign po0467 = ~new_n7903_ | ~new_n7902_ | ~new_n7901_;
  assign po0466 = ~new_n7900_ | ~new_n7899_ | ~new_n7898_;
  assign po0465 = ~new_n7897_ | ~new_n7896_ | ~new_n7895_;
  assign po0464 = ~new_n7894_ | ~new_n7893_ | ~new_n7892_;
  assign po0463 = ~new_n7891_ | ~new_n7890_ | ~new_n7889_;
  assign po0462 = ~new_n7888_ | ~new_n7887_ | ~new_n7886_;
  assign po0461 = ~new_n7885_ | ~new_n7884_ | ~new_n7883_;
  assign po0460 = ~new_n7882_ | ~new_n7881_ | ~new_n7880_;
  assign po0459 = ~new_n7879_ | ~new_n7878_ | ~new_n7877_;
  assign po0458 = ~new_n7876_ | ~new_n7875_ | ~new_n7874_;
  assign po0457 = ~new_n7873_ | ~new_n7872_ | ~new_n7871_;
  assign po0456 = ~new_n7870_ | ~new_n7869_ | ~new_n7868_;
  assign po0455 = ~new_n7867_ | ~new_n7866_ | ~new_n7865_;
  assign po0454 = ~new_n7864_ | ~new_n7863_ | ~new_n7862_;
  assign po0453 = ~new_n7861_ | ~new_n7860_ | ~new_n7859_;
  assign po0452 = ~new_n7858_ | ~new_n7857_ | ~new_n7856_;
  assign po0451 = ~new_n7855_ | ~new_n7854_ | ~new_n7853_;
  assign po0450 = ~new_n7852_ | ~new_n7851_ | ~new_n7850_;
  assign po0449 = ~new_n7849_ | ~new_n7848_ | ~new_n7847_;
  assign po0448 = ~new_n7846_ | ~new_n7845_ | ~new_n7844_;
  assign po0447 = ~new_n7843_ | ~new_n7842_ | ~new_n7841_;
  assign po0446 = ~new_n7840_ | ~new_n7839_ | ~new_n7838_;
  assign po0445 = ~new_n7837_ | ~new_n7836_ | ~new_n7835_;
  assign po0444 = ~new_n7834_ | ~new_n7833_ | ~new_n7832_;
  assign po0443 = ~new_n7831_ | ~new_n7830_ | ~new_n7829_;
  assign po0442 = ~new_n7828_ | ~new_n7827_ | ~new_n7826_;
  assign po0441 = ~new_n7825_ | ~new_n7824_ | ~new_n7823_;
  assign po0440 = ~new_n7822_ | ~new_n7821_ | ~new_n7820_;
  assign po0439 = ~new_n7812_ | ~new_n5141_ | ~new_n7809_ | ~new_n7811_ | ~new_n7810_;
  assign po0438 = ~new_n7804_ | ~new_n5140_ | ~new_n7801_ | ~new_n7802_ | ~new_n7803_;
  assign po0437 = ~new_n7796_ | ~new_n5139_ | ~new_n7793_ | ~new_n7794_ | ~new_n7795_;
  assign po0436 = ~new_n7788_ | ~new_n5138_ | ~new_n7785_ | ~new_n7786_ | ~new_n7787_;
  assign po0435 = ~new_n7778_ | ~new_n5137_ | ~new_n7779_ | ~new_n7777_ | ~new_n7780_;
  assign po0434 = ~new_n7770_ | ~new_n5136_ | ~new_n7771_ | ~new_n7769_ | ~new_n7772_;
  assign po0433 = ~new_n7762_ | ~new_n5135_ | ~new_n7763_ | ~new_n7761_ | ~new_n7764_;
  assign po0432 = ~new_n7754_ | ~new_n5134_ | ~new_n7755_ | ~new_n7753_ | ~new_n7756_;
  assign po0431 = ~new_n7746_ | ~new_n5133_ | ~new_n7747_ | ~new_n7748_ | ~new_n7745_;
  assign po0430 = ~new_n7738_ | ~new_n5132_ | ~new_n7739_ | ~new_n7740_ | ~new_n7737_;
  assign po0429 = ~new_n7730_ | ~new_n7732_ | ~new_n5131_ | ~new_n7731_ | ~new_n7729_;
  assign po0428 = ~new_n7722_ | ~new_n7724_ | ~new_n5130_ | ~new_n7723_ | ~new_n7721_;
  assign po0427 = ~new_n7714_ | ~new_n5129_ | ~new_n7716_ | ~new_n7715_ | ~new_n7713_;
  assign po0426 = ~new_n7706_ | ~new_n5128_ | ~new_n7708_ | ~new_n7707_ | ~new_n7705_;
  assign po0425 = ~new_n7698_ | ~new_n5127_ | ~new_n7700_ | ~new_n7699_ | ~new_n7697_;
  assign po0424 = ~new_n7690_ | ~new_n5126_ | ~new_n7692_ | ~new_n7691_ | ~new_n7689_;
  assign po0423 = ~new_n7682_ | ~new_n5125_ | ~new_n7683_ | ~new_n7684_ | ~new_n7681_;
  assign po0422 = ~new_n7674_ | ~new_n5124_ | ~new_n7675_ | ~new_n7676_ | ~new_n7673_;
  assign po0421 = ~new_n7666_ | ~new_n5123_ | ~new_n7667_ | ~new_n7668_ | ~new_n7665_;
  assign po0420 = ~new_n7658_ | ~new_n5122_ | ~new_n7659_ | ~new_n7660_ | ~new_n7657_;
  assign po0419 = ~new_n7650_ | ~new_n5121_ | ~new_n7652_ | ~new_n7651_ | ~new_n7649_;
  assign po0418 = ~new_n7642_ | ~new_n5120_ | ~new_n7644_ | ~new_n7643_ | ~new_n7641_;
  assign po0417 = ~new_n7634_ | ~new_n5119_ | ~new_n7635_ | ~new_n7636_ | ~new_n7633_;
  assign po0416 = ~new_n7626_ | ~new_n5118_ | ~new_n7627_ | ~new_n7628_ | ~new_n7625_;
  assign po0415 = ~new_n7618_ | ~new_n5117_ | ~new_n7619_ | ~new_n7620_ | ~new_n7617_;
  assign po0414 = ~new_n7610_ | ~new_n5116_ | ~new_n7611_ | ~new_n7612_ | ~new_n7609_;
  assign po0413 = ~new_n7602_ | ~new_n5115_ | ~new_n7603_ | ~new_n7604_ | ~new_n7601_;
  assign po0412 = ~new_n7594_ | ~new_n5114_ | ~new_n7596_ | ~new_n7595_ | ~new_n7593_;
  assign po0411 = ~new_n7588_ | ~new_n5113_ | ~new_n7585_ | ~new_n7586_ | ~new_n7587_;
  assign po0410 = ~new_n7580_ | ~new_n5112_ | ~new_n7577_ | ~new_n7578_ | ~new_n7579_;
  assign po0409 = ~new_n7572_ | ~new_n5111_ | ~new_n7569_ | ~new_n7570_ | ~new_n7571_;
  assign po0408 = ~new_n7564_ | ~new_n5110_ | ~new_n7561_ | ~new_n7562_ | ~new_n7563_;
  assign po0407 = new_n7552_ & new_n9062_;
  assign po0406 = ~new_n7530_ | ~new_n7531_ | ~new_n7529_;
  assign po0405 = ~new_n7506_ | ~new_n7507_ | ~new_n7505_;
  assign po0404 = ~new_n7482_ | ~new_n7483_ | ~new_n7481_;
  assign po0403 = ~new_n7458_ | ~new_n7459_ | ~new_n7457_;
  assign po0402 = ~new_n7434_ | ~new_n7435_ | ~new_n7433_;
  assign po0401 = ~new_n5049_ | ~new_n7410_;
  assign po0400 = ~new_n5039_ | ~new_n7386_;
  assign po0399 = ~new_n5029_ | ~new_n7362_;
  assign po0398 = ~new_n5019_ | ~new_n7338_;
  assign po0397 = ~new_n5009_ | ~new_n7314_;
  assign po0396 = ~new_n5001_ | ~new_n7290_;
  assign po0395 = ~new_n7266_ | ~new_n7267_ | ~new_n7265_;
  assign po0394 = ~new_n7242_ | ~new_n7243_ | ~new_n7241_;
  assign po0393 = ~new_n7218_ | ~new_n7219_ | ~new_n7217_;
  assign po0392 = ~new_n7194_ | ~new_n7195_ | ~new_n7193_;
  assign po0391 = ~new_n4967_ | ~new_n7170_;
  assign po0390 = ~new_n4959_ | ~new_n7146_;
  assign po0389 = ~new_n7122_ | ~new_n7123_ | ~new_n7121_;
  assign po0388 = ~new_n7098_ | ~new_n7099_ | ~new_n7097_;
  assign po0387 = ~new_n7074_ | ~new_n7075_ | ~new_n7073_;
  assign po0386 = ~new_n7050_ | ~new_n7051_ | ~new_n7049_;
  assign po0385 = ~new_n7026_ | ~new_n7027_ | ~new_n7025_;
  assign po0384 = ~new_n7002_ | ~new_n7003_ | ~new_n7001_;
  assign po0383 = ~new_n6978_ | ~new_n6979_ | ~new_n6977_;
  assign po0382 = ~new_n6954_ | ~new_n6955_ | ~new_n6953_;
  assign po0381 = ~new_n6930_ | ~new_n6931_ | ~new_n6929_;
  assign po0380 = ~new_n6906_ | ~new_n6907_ | ~new_n6905_;
  assign po0379 = ~new_n6882_ | ~new_n6883_ | ~new_n6881_;
  assign po0378 = ~new_n6858_ | ~new_n6859_ | ~new_n6857_;
  assign po0377 = ~new_n6834_ | ~new_n6835_ | ~new_n6833_;
  assign po0376 = ~new_n6811_ | ~new_n6810_ | ~new_n6809_;
  assign po0375 = ~new_n6772_ | ~new_n6771_;
  assign po0374 = ~new_n6766_ | ~new_n6765_;
  assign po0373 = ~new_n6755_ | ~new_n6754_;
  assign po0372 = ~new_n6747_ | ~new_n6746_;
  assign po0371 = pi0312 & new_n6735_;
  assign po0365 = ~new_n4807_ | ~new_n6638_;
  assign po0364 = ~new_n4805_ | ~new_n6633_;
  assign po0363 = ~new_n4803_ | ~new_n6628_;
  assign po0362 = ~new_n4801_ | ~new_n6623_;
  assign po0361 = ~new_n4799_ | ~new_n6618_;
  assign po0360 = ~new_n4797_ | ~new_n6613_;
  assign po0359 = ~new_n4795_ | ~new_n6608_;
  assign po0358 = ~new_n4793_ | ~new_n6603_;
  assign po0357 = ~new_n4789_ | ~new_n6588_;
  assign po0356 = ~new_n4787_ | ~new_n6583_;
  assign po0355 = ~new_n4785_ | ~new_n6578_;
  assign po0354 = ~new_n4783_ | ~new_n6573_;
  assign po0353 = ~new_n4781_ | ~new_n6568_;
  assign po0352 = ~new_n4779_ | ~new_n6563_;
  assign po0351 = ~new_n4777_ | ~new_n6558_;
  assign po0350 = ~new_n4775_ | ~new_n6553_;
  assign po0349 = ~new_n4771_ | ~new_n6537_;
  assign po0348 = ~new_n4769_ | ~new_n6532_;
  assign po0347 = ~new_n4767_ | ~new_n6527_;
  assign po0346 = ~new_n4765_ | ~new_n6522_;
  assign po0345 = ~new_n4763_ | ~new_n6517_;
  assign po0344 = ~new_n4761_ | ~new_n6512_;
  assign po0343 = ~new_n4759_ | ~new_n6507_;
  assign po0342 = ~new_n4757_ | ~new_n6502_;
  assign po0341 = ~new_n4754_ | ~new_n6486_;
  assign po0340 = ~new_n4752_ | ~new_n6481_;
  assign po0339 = ~new_n4750_ | ~new_n6476_;
  assign po0338 = ~new_n4748_ | ~new_n6471_;
  assign po0337 = ~new_n4746_ | ~new_n6466_;
  assign po0336 = ~new_n4744_ | ~new_n6461_;
  assign po0335 = ~new_n4742_ | ~new_n6456_;
  assign po0334 = ~new_n4740_ | ~new_n6451_;
  assign po0333 = ~new_n4736_ | ~new_n6435_;
  assign po0332 = ~new_n4734_ | ~new_n6430_;
  assign po0331 = ~new_n4732_ | ~new_n6425_;
  assign po0330 = ~new_n4730_ | ~new_n6420_;
  assign po0329 = ~new_n4728_ | ~new_n6415_;
  assign po0328 = ~new_n4726_ | ~new_n6410_;
  assign po0327 = ~new_n4724_ | ~new_n6405_;
  assign po0326 = ~new_n4722_ | ~new_n6400_;
  assign po0325 = ~new_n6384_ | ~new_n6385_ | ~new_n4718_;
  assign po0324 = ~new_n6379_ | ~new_n6380_ | ~new_n4716_;
  assign po0323 = ~new_n6374_ | ~new_n6375_ | ~new_n4714_;
  assign po0322 = ~new_n6369_ | ~new_n6370_ | ~new_n4712_;
  assign po0321 = ~new_n6364_ | ~new_n6365_ | ~new_n4710_;
  assign po0320 = ~new_n6359_ | ~new_n6360_ | ~new_n4708_;
  assign po0319 = ~new_n6354_ | ~new_n6355_ | ~new_n4706_;
  assign po0318 = ~new_n6349_ | ~new_n6350_ | ~new_n4704_;
  assign po0317 = ~new_n6332_ | ~new_n6333_ | ~new_n4700_;
  assign po0316 = ~new_n6327_ | ~new_n6328_ | ~new_n4698_;
  assign po0315 = ~new_n6322_ | ~new_n6323_ | ~new_n4696_;
  assign po0314 = ~new_n6317_ | ~new_n6318_ | ~new_n4694_;
  assign po0313 = ~new_n6312_ | ~new_n6313_ | ~new_n4692_;
  assign po0312 = ~new_n6307_ | ~new_n6308_ | ~new_n4690_;
  assign po0311 = ~new_n6302_ | ~new_n6303_ | ~new_n4688_;
  assign po0310 = ~new_n6297_ | ~new_n6298_ | ~new_n4686_;
  assign po0309 = ~new_n6280_ | ~new_n6281_ | ~new_n4682_;
  assign po0308 = ~new_n6275_ | ~new_n6276_ | ~new_n4680_;
  assign po0307 = ~new_n6270_ | ~new_n6271_ | ~new_n4678_;
  assign po0306 = ~new_n6265_ | ~new_n6266_ | ~new_n4676_;
  assign po0305 = ~new_n6260_ | ~new_n6261_ | ~new_n4674_;
  assign po0304 = ~new_n6255_ | ~new_n6256_ | ~new_n4672_;
  assign po0303 = ~new_n6250_ | ~new_n6251_ | ~new_n4670_;
  assign po0302 = ~new_n6245_ | ~new_n6246_ | ~new_n4668_;
  assign po0301 = ~new_n6231_ | ~new_n6232_ | ~new_n4665_;
  assign po0300 = ~new_n6226_ | ~new_n6227_ | ~new_n4663_;
  assign po0299 = ~new_n6221_ | ~new_n6222_ | ~new_n4661_;
  assign po0298 = ~new_n6216_ | ~new_n6217_ | ~new_n4659_;
  assign po0297 = ~new_n6211_ | ~new_n6212_ | ~new_n4657_;
  assign po0296 = ~new_n6206_ | ~new_n6207_ | ~new_n4655_;
  assign po0295 = ~new_n6201_ | ~new_n6202_ | ~new_n4653_;
  assign po0294 = ~new_n6196_ | ~new_n6197_ | ~new_n4651_;
  assign po0293 = ~new_n6180_ | ~new_n6181_ | ~new_n4648_;
  assign po0292 = ~new_n6175_ | ~new_n6176_ | ~new_n4646_;
  assign po0291 = ~new_n6170_ | ~new_n6171_ | ~new_n4644_;
  assign po0290 = ~new_n6165_ | ~new_n6166_ | ~new_n4642_;
  assign po0289 = ~new_n6160_ | ~new_n6161_ | ~new_n4640_;
  assign po0288 = ~new_n6155_ | ~new_n6156_ | ~new_n4638_;
  assign po0287 = ~new_n6150_ | ~new_n6151_ | ~new_n4636_;
  assign po0286 = ~new_n6145_ | ~new_n6146_ | ~new_n4634_;
  assign po0285 = ~new_n6128_ | ~new_n6129_ | ~new_n4630_;
  assign po0284 = ~new_n6123_ | ~new_n6124_ | ~new_n4628_;
  assign po0283 = ~new_n6118_ | ~new_n6119_ | ~new_n4626_;
  assign po0282 = ~new_n6113_ | ~new_n6114_ | ~new_n4624_;
  assign po0281 = ~new_n6108_ | ~new_n6109_ | ~new_n4622_;
  assign po0280 = ~new_n6103_ | ~new_n6104_ | ~new_n4620_;
  assign po0279 = ~new_n6098_ | ~new_n6099_ | ~new_n4618_;
  assign po0278 = ~new_n6093_ | ~new_n6094_ | ~new_n4616_;
  assign po0277 = ~new_n6076_ | ~new_n6077_ | ~new_n4612_;
  assign po0276 = ~new_n6071_ | ~new_n6072_ | ~new_n4610_;
  assign po0275 = ~new_n6066_ | ~new_n6067_ | ~new_n4608_;
  assign po0274 = ~new_n6061_ | ~new_n6062_ | ~new_n4606_;
  assign po0273 = ~new_n6056_ | ~new_n6057_ | ~new_n4604_;
  assign po0272 = ~new_n6051_ | ~new_n6052_ | ~new_n4602_;
  assign po0271 = ~new_n6046_ | ~new_n6047_ | ~new_n4600_;
  assign po0270 = ~new_n6041_ | ~new_n6042_ | ~new_n4598_;
  assign po0269 = ~new_n6024_ | ~new_n6025_ | ~new_n4595_;
  assign po0268 = ~new_n6019_ | ~new_n6020_ | ~new_n4593_;
  assign po0267 = ~new_n6014_ | ~new_n6015_ | ~new_n4591_;
  assign po0266 = ~new_n6009_ | ~new_n6010_ | ~new_n4589_;
  assign po0265 = ~new_n6004_ | ~new_n6005_ | ~new_n4587_;
  assign po0264 = ~new_n5999_ | ~new_n6000_ | ~new_n4585_;
  assign po0263 = ~new_n5994_ | ~new_n5995_ | ~new_n4583_;
  assign po0262 = ~new_n5989_ | ~new_n5990_ | ~new_n4581_;
  assign po0261 = ~new_n5973_ | ~new_n5974_ | ~new_n4577_;
  assign po0260 = ~new_n5968_ | ~new_n5969_ | ~new_n4575_;
  assign po0259 = ~new_n5963_ | ~new_n5964_ | ~new_n4573_;
  assign po0258 = ~new_n5958_ | ~new_n5959_ | ~new_n4571_;
  assign po0257 = ~new_n5953_ | ~new_n5954_ | ~new_n4569_;
  assign po0256 = ~new_n5948_ | ~new_n5949_ | ~new_n4567_;
  assign po0255 = ~new_n5943_ | ~new_n5944_ | ~new_n4565_;
  assign po0254 = ~new_n5938_ | ~new_n5939_ | ~new_n4563_;
  assign po0253 = ~new_n5921_ | ~new_n5922_ | ~new_n4559_;
  assign po0252 = ~new_n5916_ | ~new_n5917_ | ~new_n4557_;
  assign po0251 = ~new_n5911_ | ~new_n5912_ | ~new_n4555_;
  assign po0250 = ~new_n5906_ | ~new_n5907_ | ~new_n4553_;
  assign po0249 = ~new_n5901_ | ~new_n5902_ | ~new_n4551_;
  assign po0248 = ~new_n5896_ | ~new_n5897_ | ~new_n4549_;
  assign po0247 = ~new_n5891_ | ~new_n5892_ | ~new_n4547_;
  assign po0246 = ~new_n5886_ | ~new_n5887_ | ~new_n4545_;
  assign po0245 = ~new_n5869_ | ~new_n5870_ | ~new_n4541_;
  assign po0244 = ~new_n5864_ | ~new_n5865_ | ~new_n4539_;
  assign po0243 = ~new_n5859_ | ~new_n5860_ | ~new_n4537_;
  assign po0242 = ~new_n5854_ | ~new_n5855_ | ~new_n4535_;
  assign po0241 = ~new_n5849_ | ~new_n5850_ | ~new_n4533_;
  assign po0240 = ~new_n5844_ | ~new_n5845_ | ~new_n4531_;
  assign po0239 = ~new_n5839_ | ~new_n5840_ | ~new_n4529_;
  assign po0238 = ~new_n5834_ | ~new_n5835_ | ~new_n4527_;
  assign po0237 = ~new_n4523_ | ~new_n9115_ | ~new_n9114_;
  assign po0236 = ~new_n5791_ | ~new_n5485_ | ~new_n5790_ | ~new_n5792_;
  assign po0235 = ~new_n4519_ | ~new_n5788_;
  assign po0233 = pi0174 & new_n9093_;
  assign po0232 = pi0173 & new_n9093_;
  assign po0231 = pi0172 & new_n9093_;
  assign po0230 = pi0171 & new_n9093_;
  assign po0229 = pi0170 & new_n9093_;
  assign po0228 = pi0169 & new_n9093_;
  assign po0227 = pi0168 & new_n9093_;
  assign po0226 = pi0167 & new_n9093_;
  assign po0225 = pi0166 & new_n9093_;
  assign po0224 = pi0165 & new_n9093_;
  assign po0223 = pi0164 & new_n9093_;
  assign po0222 = pi0163 & new_n9093_;
  assign po0221 = pi0162 & new_n9093_;
  assign po0220 = pi0161 & new_n9093_;
  assign po0219 = pi0160 & new_n9093_;
  assign po0218 = pi0159 & new_n9093_;
  assign po0217 = pi0158 & new_n9093_;
  assign po0216 = pi0157 & new_n9093_;
  assign po0215 = pi0156 & new_n9093_;
  assign po0214 = pi0155 & new_n9093_;
  assign po0213 = pi0154 & new_n9093_;
  assign po0212 = pi0153 & new_n9093_;
  assign po0211 = pi0152 & new_n9093_;
  assign po0210 = pi0151 & new_n9093_;
  assign po0209 = pi0150 & new_n9093_;
  assign po0208 = pi0149 & new_n9093_;
  assign po0207 = pi0148 & new_n9093_;
  assign po0206 = pi0147 & new_n9093_;
  assign po0205 = pi0146 & new_n9093_;
  assign po0204 = pi0145 & new_n9093_;
  assign po0201 = ~new_n5619_ | ~new_n9090_ | ~new_n9089_;
  assign po0200 = ~new_n4467_ | ~new_n9088_ | ~new_n9087_;
  assign po0199 = ~new_n4466_ | ~new_n5613_;
  assign po0198 = ~new_n5600_ | ~new_n5599_ | ~new_n5598_;
  assign po0197 = ~new_n5597_ | ~new_n5596_ | ~new_n5595_;
  assign po0196 = ~new_n5594_ | ~new_n5593_ | ~new_n5592_;
  assign po0195 = ~new_n5591_ | ~new_n5590_ | ~new_n5589_;
  assign po0194 = ~new_n5588_ | ~new_n5587_ | ~new_n5586_;
  assign po0193 = ~new_n5585_ | ~new_n5584_ | ~new_n5583_;
  assign po0192 = ~new_n5582_ | ~new_n5581_ | ~new_n5580_;
  assign po0191 = ~new_n5579_ | ~new_n5578_ | ~new_n5577_;
  assign po0190 = ~new_n5576_ | ~new_n5575_ | ~new_n5574_;
  assign po0189 = ~new_n5573_ | ~new_n5572_ | ~new_n5571_;
  assign po0188 = ~new_n5570_ | ~new_n5569_ | ~new_n5568_;
  assign po0187 = ~new_n5567_ | ~new_n5566_ | ~new_n5565_;
  assign po0186 = ~new_n5564_ | ~new_n5563_ | ~new_n5562_;
  assign po0185 = ~new_n5561_ | ~new_n5560_ | ~new_n5559_;
  assign po0184 = ~new_n5558_ | ~new_n5557_ | ~new_n5556_;
  assign po0183 = ~new_n5555_ | ~new_n5554_ | ~new_n5553_;
  assign po0182 = ~new_n5552_ | ~new_n5551_ | ~new_n5550_;
  assign po0181 = ~new_n5549_ | ~new_n5548_ | ~new_n5547_;
  assign po0180 = ~new_n5546_ | ~new_n5545_ | ~new_n5544_;
  assign po0179 = ~new_n5543_ | ~new_n5542_ | ~new_n5541_;
  assign po0178 = ~new_n5540_ | ~new_n5539_ | ~new_n5538_;
  assign po0177 = ~new_n5537_ | ~new_n5536_ | ~new_n5535_;
  assign po0176 = ~new_n5534_ | ~new_n5533_ | ~new_n5532_;
  assign po0175 = ~new_n5531_ | ~new_n5530_ | ~new_n5529_;
  assign po0174 = ~new_n5528_ | ~new_n5527_ | ~new_n5526_;
  assign po0173 = ~new_n5525_ | ~new_n5524_ | ~new_n5523_;
  assign po0172 = ~new_n5522_ | ~new_n5521_ | ~new_n5520_;
  assign po0171 = ~new_n5519_ | ~new_n5518_ | ~new_n5517_;
  assign po0170 = ~new_n5516_ | ~new_n5515_ | ~new_n5514_;
  assign po0169 = ~new_n5513_ | ~new_n5512_ | ~new_n5511_;
  assign new_n4218_ = ~new_n5402_ | ~new_n5400_ | ~new_n5401_ | ~new_n5403_;
  assign new_n4219_ = ~new_n5398_ | ~new_n5396_ | ~new_n5397_ | ~new_n5399_;
  assign new_n4220_ = ~new_n5394_ | ~new_n5392_ | ~new_n5393_ | ~new_n5395_;
  assign new_n4221_ = ~new_n5390_ | ~new_n5388_ | ~new_n5389_ | ~new_n5391_;
  assign new_n4222_ = ~new_n5386_ | ~new_n5384_ | ~new_n5385_ | ~new_n5387_;
  assign new_n4223_ = ~new_n5382_ | ~new_n5380_ | ~new_n5381_ | ~new_n5383_;
  assign new_n4224_ = ~new_n5378_ | ~new_n5376_ | ~new_n5377_ | ~new_n5379_;
  assign new_n4225_ = ~new_n5374_ | ~new_n5372_ | ~new_n5373_ | ~new_n5375_;
  assign new_n4226_ = ~new_n3613_ | ~new_n5798_;
  assign new_n4227_ = ~new_n3615_ | ~new_n5798_;
  assign new_n4228_ = ~new_n3614_ | ~new_n5798_;
  assign new_n4229_ = ~new_n3616_ | ~new_n5798_;
  assign new_n4230_ = ~new_n4502_ | ~new_n4499_ | ~new_n4500_ | ~new_n4503_ | ~new_n4501_;
  assign new_n4231_ = ~pi0548;
  assign new_n4232_ = ~pi0141;
  assign new_n4233_ = ~pi0141 | ~new_n4241_;
  assign new_n4234_ = ~new_n5464_ | ~new_n4235_;
  assign new_n4235_ = ~pi0140;
  assign new_n4236_ = ~pi0140 | ~new_n5464_;
  assign new_n4237_ = ~pi0509;
  assign new_n4238_ = ~pi0141 | ~new_n4235_;
  assign new_n4239_ = pi0141 | pi0140;
  assign new_n4240_ = ~pi0033;
  assign new_n4241_ = ~pi0142;
  assign new_n4242_ = ~pi0142 | ~new_n4243_;
  assign new_n4243_ = ~pi0548 | ~new_n4240_;
  assign new_n4244_ = pi0033 | pi0548;
  assign new_n4245_ = ~pi0177;
  assign new_n4246_ = ~pi0176;
  assign new_n4247_ = pi0310 | pi0311;
  assign new_n4248_ = ~new_n5623_ | ~new_n4253_;
  assign new_n4249_ = ~pi0311;
  assign new_n4250_ = ~pi0310;
  assign new_n4251_ = ~pi0310 | ~pi0311;
  assign new_n4252_ = ~new_n5488_ | ~new_n4253_;
  assign new_n4253_ = ~pi0309;
  assign new_n4254_ = ~pi0309 | ~new_n4256_;
  assign new_n4255_ = ~new_n5626_ | ~new_n5488_;
  assign new_n4256_ = ~pi0308;
  assign new_n4257_ = ~new_n4497_ | ~new_n4494_ | ~new_n4495_ | ~new_n4498_ | ~new_n4496_;
  assign new_n4258_ = ~new_n4482_ | ~new_n4479_ | ~new_n4480_ | ~new_n4483_ | ~new_n4481_;
  assign new_n4259_ = ~new_n4230_ | ~new_n4266_;
  assign new_n4260_ = ~new_n4477_ | ~new_n4474_ | ~new_n4475_ | ~new_n4478_ | ~new_n4476_;
  assign new_n4261_ = ~new_n5622_ | ~new_n4241_;
  assign new_n4262_ = ~new_n5449_ | ~new_n3786_;
  assign new_n4263_ = ~new_n4487_ | ~new_n4484_ | ~new_n4485_ | ~new_n4488_ | ~new_n4486_;
  assign new_n4264_ = ~new_n4472_ | ~new_n4469_ | ~new_n4470_ | ~new_n4473_ | ~new_n4471_;
  assign new_n4265_ = ~new_n3509_ | ~new_n5644_;
  assign new_n4266_ = ~new_n4507_ | ~new_n4504_ | ~new_n4505_ | ~new_n4508_ | ~new_n4506_;
  assign new_n4267_ = ~new_n4260_ | ~new_n4264_;
  assign new_n4268_ = ~new_n5661_ | ~new_n4264_;
  assign new_n4269_ = ~new_n5763_ | ~new_n4266_;
  assign new_n4270_ = ~new_n5644_ | ~new_n5661_;
  assign new_n4271_ = ~new_n3607_ | ~new_n5453_;
  assign new_n4272_ = ~new_n3608_ | ~new_n5453_;
  assign new_n4273_ = ~new_n3608_ | ~new_n5452_;
  assign new_n4274_ = ~new_n5644_ | ~new_n4260_;
  assign new_n4275_ = ~new_n4512_ | ~new_n3509_;
  assign new_n4276_ = ~new_n9105_ | ~new_n23632_ | ~new_n5469_ | ~new_n4418_ | ~new_n9104_;
  assign new_n4277_ = ~pi0178;
  assign new_n4278_ = ~pi0178 | ~new_n5785_;
  assign new_n4279_ = pi0175 | pi0177;
  assign new_n4280_ = ~pi0176 | ~new_n4245_;
  assign new_n4281_ = pi0176 | pi0177;
  assign new_n4282_ = ~new_n23871_ | ~pi0175;
  assign new_n4283_ = ~new_n5822_ | ~new_n4277_;
  assign new_n4284_ = ~pi0316;
  assign new_n4285_ = ~pi0315;
  assign new_n4286_ = ~pi0315 | ~pi0316;
  assign new_n4287_ = ~pi0314;
  assign new_n4288_ = ~pi0314 | ~new_n5804_;
  assign new_n4289_ = ~pi0313;
  assign new_n4290_ = ~pi0313 | ~new_n5805_;
  assign new_n4291_ = pi0175 | pi0176;
  assign new_n4292_ = ~new_n5451_ | ~pi0547;
  assign new_n4293_ = ~new_n4309_ | ~new_n5797_;
  assign new_n4294_ = ~new_n4293_ | ~new_n4284_;
  assign new_n4295_ = ~new_n4336_ | ~new_n5807_;
  assign new_n4296_ = ~pi0316 | ~new_n4297_;
  assign new_n4297_ = ~new_n4306_ | ~new_n4314_;
  assign new_n4298_ = ~new_n5487_ | ~new_n5811_;
  assign new_n4299_ = ~new_n4312_ | ~new_n4284_;
  assign new_n4300_ = ~new_n5803_ | ~new_n3642_;
  assign new_n4301_ = ~new_n4300_ | ~new_n5823_;
  assign new_n4302_ = ~new_n4290_ | ~new_n5819_;
  assign new_n4303_ = ~new_n4542_ | ~new_n3648_;
  assign new_n4304_ = ~new_n4297_ | ~new_n4284_;
  assign new_n4305_ = ~new_n3646_ | ~new_n3642_;
  assign new_n4306_ = ~pi0316 | ~new_n4293_;
  assign new_n4307_ = ~new_n4305_ | ~new_n5875_;
  assign new_n4308_ = ~new_n4303_ | ~new_n5873_;
  assign new_n4309_ = ~pi0316 | ~new_n4285_;
  assign new_n4310_ = ~new_n4560_ | ~new_n5796_;
  assign new_n4311_ = ~new_n5799_ | ~pi0316;
  assign new_n4312_ = ~new_n4304_ | ~new_n4311_;
  assign new_n4313_ = ~new_n3649_ | ~new_n3642_;
  assign new_n4314_ = ~new_n5798_ | ~new_n4284_;
  assign new_n4315_ = ~new_n4313_ | ~new_n5927_;
  assign new_n4316_ = ~new_n4310_ | ~new_n5925_;
  assign new_n4317_ = ~new_n4578_ | ~new_n3648_;
  assign new_n4318_ = ~new_n3651_ | ~new_n3642_;
  assign new_n4319_ = ~new_n4318_ | ~new_n5978_;
  assign new_n4320_ = ~new_n5804_ | ~pi0313 | ~new_n4287_;
  assign new_n4321_ = ~new_n9121_ | ~new_n4298_;
  assign new_n4322_ = ~new_n3654_ | ~new_n5803_;
  assign new_n4323_ = ~new_n4322_ | ~new_n6030_;
  assign new_n4324_ = ~new_n4320_ | ~new_n6028_;
  assign new_n4325_ = ~new_n4613_ | ~new_n3657_;
  assign new_n4326_ = ~new_n3654_ | ~new_n3646_;
  assign new_n4327_ = ~new_n4326_ | ~new_n6082_;
  assign new_n4328_ = ~new_n4325_ | ~new_n6080_;
  assign new_n4329_ = ~new_n4631_ | ~new_n5796_;
  assign new_n4330_ = ~new_n3654_ | ~new_n3649_;
  assign new_n4331_ = ~new_n4330_ | ~new_n6134_;
  assign new_n4332_ = ~new_n4329_ | ~new_n6132_;
  assign new_n4333_ = ~new_n3657_ | ~pi0313 | ~new_n4285_;
  assign new_n4334_ = ~new_n3654_ | ~new_n3651_;
  assign new_n4335_ = ~new_n4334_ | ~new_n6185_;
  assign new_n4336_ = ~new_n5805_ | ~new_n4289_;
  assign new_n4337_ = ~new_n3641_ | ~new_n5813_;
  assign new_n4338_ = ~new_n4524_ | ~new_n4337_;
  assign new_n4339_ = ~new_n3660_ | ~new_n5803_;
  assign new_n4340_ = ~new_n4339_ | ~new_n4337_;
  assign new_n4341_ = ~new_n4336_ | ~new_n5487_;
  assign new_n4342_ = ~new_n4683_ | ~new_n3648_;
  assign new_n4343_ = ~new_n3660_ | ~new_n3646_;
  assign new_n4344_ = ~new_n4343_ | ~new_n6286_;
  assign new_n4345_ = ~new_n4342_ | ~new_n6284_;
  assign new_n4346_ = ~new_n4701_ | ~new_n5796_;
  assign new_n4347_ = ~new_n3660_ | ~new_n3649_;
  assign new_n4348_ = ~new_n4347_ | ~new_n6338_;
  assign new_n4349_ = ~new_n4346_ | ~new_n6336_;
  assign new_n4350_ = ~new_n4719_ | ~new_n3648_;
  assign new_n4351_ = ~new_n3660_ | ~new_n3651_;
  assign new_n4352_ = ~new_n4737_ | ~new_n5804_;
  assign new_n4353_ = ~new_n3664_ | ~new_n5803_;
  assign new_n4354_ = ~new_n4352_ | ~new_n6438_;
  assign new_n4355_ = ~new_n3657_ | ~pi0315 | ~new_n4289_;
  assign new_n4356_ = ~new_n3664_ | ~new_n3646_;
  assign new_n4357_ = ~new_n4355_ | ~new_n6489_;
  assign new_n4358_ = ~new_n4772_ | ~new_n5796_;
  assign new_n4359_ = ~new_n3664_ | ~new_n3649_;
  assign new_n4360_ = ~new_n4358_ | ~new_n6540_;
  assign new_n4361_ = ~new_n4790_ | ~new_n3657_;
  assign new_n4362_ = ~new_n3664_ | ~new_n3651_;
  assign new_n4363_ = ~pi0545;
  assign new_n4364_ = ~new_n5695_ | ~new_n4258_;
  assign new_n4365_ = ~new_n3670_ | ~new_n4269_;
  assign new_n4366_ = ~new_n27144_;
  assign new_n4367_ = ~new_n22221_;
  assign new_n4368_ = ~new_n21854_;
  assign new_n4369_ = ~new_n25105_;
  assign new_n4370_ = ~new_n27146_;
  assign new_n4371_ = ~new_n21624_;
  assign new_n4372_ = ~new_n5746_ | ~new_n4230_;
  assign new_n4373_ = ~new_n3606_ | ~new_n5479_;
  assign new_n4374_ = ~new_n4492_ | ~new_n4489_ | ~new_n4490_ | ~new_n4493_ | ~new_n4491_;
  assign new_n4375_ = ~new_n4818_ | ~new_n3617_;
  assign new_n4376_ = ~new_n4823_ | ~new_n9132_ | ~new_n9131_;
  assign new_n4377_ = ~new_n6680_ | ~new_n4378_ | ~new_n4275_;
  assign new_n4378_ = ~new_n5470_ | ~new_n4374_;
  assign new_n4379_ = ~pi0308 | ~new_n6659_;
  assign new_n4380_ = ~pi0308 | ~new_n6661_;
  assign new_n4381_ = ~new_n4252_ | ~new_n4383_;
  assign new_n4382_ = ~new_n4830_ | ~new_n3673_;
  assign new_n4383_ = ~pi0309 | ~new_n4251_;
  assign new_n4384_ = ~new_n4247_ | ~new_n4251_;
  assign new_n4385_ = ~new_n5506_ | ~new_n5479_ | ~new_n4374_;
  assign new_n4386_ = ~new_n3674_ | ~new_n4399_;
  assign new_n4387_ = ~new_n4271_ | ~new_n6715_;
  assign new_n4388_ = ~new_n23877_;
  assign new_n4389_ = ~new_n6734_ | ~new_n5486_ | ~new_n4283_;
  assign new_n4390_ = ~new_n4291_ | ~new_n4279_;
  assign new_n4391_ = ~new_n5450_ | ~new_n4257_ | ~new_n4260_;
  assign new_n4392_ = ~new_n5661_ | ~new_n4257_ | ~new_n3786_;
  assign new_n4393_ = ~new_n23443_;
  assign new_n4394_ = ~new_n22636_;
  assign new_n4395_ = ~new_n5451_ | ~new_n4245_;
  assign new_n4396_ = ~pi0508;
  assign new_n4397_ = ~new_n3784_;
  assign new_n4398_ = ~new_n4817_ | ~new_n3606_;
  assign new_n4399_ = ~new_n3617_ | ~new_n5470_;
  assign new_n4400_ = ~new_n5508_ | ~new_n5678_;
  assign new_n4401_ = ~new_n5508_ | ~new_n4258_;
  assign new_n4402_ = ~new_n4820_ | ~new_n4819_ | ~new_n3605_;
  assign new_n4403_ = ~pi0176 | ~new_n4404_;
  assign new_n4404_ = ~new_n5492_ | ~new_n6786_;
  assign new_n4405_ = ~new_n7559_ | ~new_n7558_;
  assign new_n4406_ = ~new_n3546_ | ~new_n7819_;
  assign new_n4407_ = ~new_n7914_ | ~new_n7913_;
  assign new_n4408_ = ~new_n3546_ | ~new_n8009_;
  assign new_n4409_ = ~new_n3546_ | ~new_n8153_;
  assign new_n4410_ = ~new_n6646_ | ~new_n6645_;
  assign new_n4411_ = ~new_n6643_ | ~new_n6642_;
  assign new_n4412_ = ~pi0507;
  assign new_n4413_ = pi0547 | new_n2971_;
  assign new_n4414_ = ~new_n22288_;
  assign new_n4415_ = ~new_n22288_ | ~new_n3541_;
  assign new_n4416_ = ~new_n5186_ | ~new_n5490_;
  assign new_n4417_ = ~new_n5300_ | ~new_n5294_ | ~new_n5297_ | ~new_n5304_;
  assign new_n4418_ = ~new_n5438_ | ~new_n3618_ | ~new_n4264_;
  assign new_n4419_ = ~pi0551;
  assign new_n4420_ = ~pi0553;
  assign new_n4421_ = ~new_n4255_ | ~new_n4380_;
  assign new_n4422_ = ~new_n4379_ | ~new_n8671_;
  assign new_n4423_ = ~new_n5445_ | ~new_n4248_;
  assign new_n4424_ = ~new_n4254_ | ~new_n8930_;
  assign new_n4425_ = ~new_n9117_ | ~new_n9116_;
  assign new_n4426_ = ~new_n9120_ | ~new_n9119_;
  assign new_n4427_ = ~new_n9123_ | ~new_n9122_;
  assign new_n4428_ = ~new_n9189_ | ~new_n9188_;
  assign new_n4429_ = ~new_n9192_ | ~new_n9191_;
  assign po0165 = ~new_n9077_ | ~new_n9076_;
  assign po0166 = ~new_n9079_ | ~new_n9078_;
  assign po0167 = ~new_n9081_ | ~new_n9080_;
  assign po0168 = ~new_n9083_ | ~new_n9082_;
  assign new_n4434_ = ~new_n9092_ | ~new_n9091_;
  assign new_n4435_ = new_n4239_ & new_n5442_;
  assign po0202 = ~new_n9095_ | ~new_n9094_;
  assign po0203 = ~new_n9097_ | ~new_n9096_;
  assign po0234 = ~new_n9111_ | ~new_n9110_;
  assign new_n4439_ = new_n4808_ & new_n3512_;
  assign po0366 = ~new_n9128_ | ~new_n9127_;
  assign po0367 = ~new_n9136_ | ~new_n9135_;
  assign new_n4442_ = ~new_n9143_ | ~new_n9142_;
  assign new_n4443_ = ~new_n9140_ | ~new_n9139_;
  assign po0368 = ~new_n9146_ | ~new_n9145_;
  assign po0369 = ~new_n9148_ | ~new_n9147_;
  assign po0370 = ~new_n9152_ | ~new_n9151_;
  assign new_n4447_ = ~pi0144 & ~pi0509;
  assign po0600 = ~new_n9167_ | ~new_n9166_;
  assign po0602 = ~new_n9171_ | ~new_n9170_;
  assign po0603 = ~new_n9173_ | ~new_n9172_;
  assign po0605 = ~new_n9175_ | ~new_n9174_;
  assign po0607 = ~new_n9179_ | ~new_n9178_;
  assign po0609 = ~new_n9183_ | ~new_n9182_;
  assign po0612 = ~new_n9185_ | ~new_n9184_;
  assign po0613 = ~new_n9187_ | ~new_n9186_;
  assign new_n4456_ = ~new_n9195_ | ~new_n9194_;
  assign new_n4457_ = ~new_n9197_ | ~new_n9196_;
  assign new_n4458_ = ~new_n9199_ | ~new_n9198_;
  assign new_n4459_ = new_n27131_ & new_n3512_;
  assign new_n4460_ = ~new_n9201_ | ~new_n9200_;
  assign new_n4461_ = ~new_n9203_ | ~new_n9202_;
  assign new_n4462_ = ~new_n9205_ | ~new_n9204_;
  assign new_n4463_ = ~new_n9207_ | ~new_n9206_;
  assign new_n4464_ = ~new_n9209_ | ~new_n9208_;
  assign new_n4465_ = pi0142 & new_n5603_;
  assign new_n4466_ = new_n5612_ & new_n4236_;
  assign new_n4467_ = new_n5614_ & new_n4234_;
  assign new_n4468_ = pi0548 & pi0142;
  assign new_n4469_ = new_n5630_ & new_n5628_ & new_n5629_ & new_n5631_;
  assign new_n4470_ = new_n5634_ & new_n5632_ & new_n5633_ & new_n5635_;
  assign new_n4471_ = new_n5637_ & new_n5636_;
  assign new_n4472_ = new_n5639_ & new_n5638_;
  assign new_n4473_ = new_n5642_ & new_n5640_ & new_n5641_ & new_n5643_;
  assign new_n4474_ = new_n5647_ & new_n5645_ & new_n5646_ & new_n5648_;
  assign new_n4475_ = new_n5651_ & new_n5649_ & new_n5650_ & new_n5652_;
  assign new_n4476_ = new_n5654_ & new_n5653_;
  assign new_n4477_ = new_n5656_ & new_n5655_;
  assign new_n4478_ = new_n5659_ & new_n5657_ & new_n5658_ & new_n5660_;
  assign new_n4479_ = new_n5664_ & new_n5662_ & new_n5663_ & new_n5665_;
  assign new_n4480_ = new_n5668_ & new_n5666_ & new_n5667_ & new_n5669_;
  assign new_n4481_ = new_n5671_ & new_n5670_;
  assign new_n4482_ = new_n5673_ & new_n5672_;
  assign new_n4483_ = new_n5676_ & new_n5674_ & new_n5675_ & new_n5677_;
  assign new_n4484_ = new_n5698_ & new_n5696_ & new_n5697_ & new_n5699_;
  assign new_n4485_ = new_n5702_ & new_n5700_ & new_n5701_ & new_n5703_;
  assign new_n4486_ = new_n5705_ & new_n5704_;
  assign new_n4487_ = new_n5707_ & new_n5706_;
  assign new_n4488_ = new_n5710_ & new_n5708_ & new_n5709_ & new_n5711_;
  assign new_n4489_ = new_n5715_ & new_n5713_ & new_n5714_ & new_n5716_;
  assign new_n4490_ = new_n5719_ & new_n5717_ & new_n5718_ & new_n5720_;
  assign new_n4491_ = new_n5722_ & new_n5721_;
  assign new_n4492_ = new_n5724_ & new_n5723_;
  assign new_n4493_ = new_n5727_ & new_n5725_ & new_n5726_ & new_n5728_;
  assign new_n4494_ = new_n5681_ & new_n5679_ & new_n5680_ & new_n5682_;
  assign new_n4495_ = new_n5685_ & new_n5683_ & new_n5684_ & new_n5686_;
  assign new_n4496_ = new_n5688_ & new_n5687_;
  assign new_n4497_ = new_n5690_ & new_n5689_;
  assign new_n4498_ = new_n5693_ & new_n5691_ & new_n5692_ & new_n5694_;
  assign new_n4499_ = new_n5749_ & new_n5747_ & new_n5748_ & new_n5750_;
  assign new_n4500_ = new_n5753_ & new_n5751_ & new_n5752_ & new_n5754_;
  assign new_n4501_ = new_n5756_ & new_n5755_;
  assign new_n4502_ = new_n5758_ & new_n5757_;
  assign new_n4503_ = new_n5761_ & new_n5759_ & new_n5760_ & new_n5762_;
  assign new_n4504_ = new_n5732_ & new_n5730_ & new_n5731_ & new_n5733_;
  assign new_n4505_ = new_n5736_ & new_n5734_ & new_n5735_ & new_n5737_;
  assign new_n4506_ = new_n5739_ & new_n5738_;
  assign new_n4507_ = new_n5741_ & new_n5740_;
  assign new_n4508_ = new_n5744_ & new_n5742_ & new_n5743_ & new_n5745_;
  assign new_n4509_ = new_n3508_ & new_n5449_;
  assign new_n4510_ = new_n5712_ & new_n4374_;
  assign new_n4511_ = new_n5479_ & new_n4257_;
  assign new_n4512_ = new_n5480_ & new_n4257_;
  assign new_n4513_ = new_n5767_ & new_n5765_ & new_n5766_ & new_n5768_;
  assign new_n4514_ = new_n5771_ & new_n5769_ & new_n5770_ & new_n5772_;
  assign new_n4515_ = new_n5695_ & new_n3786_;
  assign new_n4516_ = new_n4374_ & new_n4263_ & new_n4264_;
  assign new_n4517_ = new_n5777_ & new_n4391_ & new_n4392_;
  assign new_n4518_ = new_n5782_ & new_n4245_;
  assign new_n4519_ = new_n5787_ & new_n4280_;
  assign new_n4520_ = new_n5496_ & new_n3786_;
  assign new_n4521_ = pi0175 & pi0178;
  assign new_n4522_ = new_n5494_ & new_n5484_;
  assign new_n4523_ = new_n4522_ & new_n5795_;
  assign new_n4524_ = new_n4321_ & new_n5815_;
  assign new_n4525_ = new_n5827_ & new_n5468_;
  assign new_n4526_ = new_n5832_ & new_n5831_;
  assign new_n4527_ = new_n4526_ & new_n5833_;
  assign new_n4528_ = new_n5837_ & new_n5836_;
  assign new_n4529_ = new_n4528_ & new_n5838_;
  assign new_n4530_ = new_n5842_ & new_n5841_;
  assign new_n4531_ = new_n4530_ & new_n5843_;
  assign new_n4532_ = new_n5847_ & new_n5846_;
  assign new_n4533_ = new_n4532_ & new_n5848_;
  assign new_n4534_ = new_n5852_ & new_n5851_;
  assign new_n4535_ = new_n4534_ & new_n5853_;
  assign new_n4536_ = new_n5857_ & new_n5856_;
  assign new_n4537_ = new_n4536_ & new_n5858_;
  assign new_n4538_ = new_n5862_ & new_n5861_;
  assign new_n4539_ = new_n4538_ & new_n5863_;
  assign new_n4540_ = new_n5867_ & new_n5866_;
  assign new_n4541_ = new_n4540_ & new_n5868_;
  assign new_n4542_ = pi0313 & pi0315;
  assign new_n4543_ = new_n5879_ & new_n5468_;
  assign new_n4544_ = new_n5884_ & new_n5883_;
  assign new_n4545_ = new_n4544_ & new_n5885_;
  assign new_n4546_ = new_n5889_ & new_n5888_;
  assign new_n4547_ = new_n4546_ & new_n5890_;
  assign new_n4548_ = new_n5894_ & new_n5893_;
  assign new_n4549_ = new_n4548_ & new_n5895_;
  assign new_n4550_ = new_n5899_ & new_n5898_;
  assign new_n4551_ = new_n4550_ & new_n5900_;
  assign new_n4552_ = new_n5904_ & new_n5903_;
  assign new_n4553_ = new_n4552_ & new_n5905_;
  assign new_n4554_ = new_n5909_ & new_n5908_;
  assign new_n4555_ = new_n4554_ & new_n5910_;
  assign new_n4556_ = new_n5914_ & new_n5913_;
  assign new_n4557_ = new_n4556_ & new_n5915_;
  assign new_n4558_ = new_n5919_ & new_n5918_;
  assign new_n4559_ = new_n4558_ & new_n5920_;
  assign new_n4560_ = pi0313 & pi0314;
  assign new_n4561_ = new_n5931_ & new_n5468_;
  assign new_n4562_ = new_n5936_ & new_n5935_;
  assign new_n4563_ = new_n4562_ & new_n5937_;
  assign new_n4564_ = new_n5941_ & new_n5940_;
  assign new_n4565_ = new_n4564_ & new_n5942_;
  assign new_n4566_ = new_n5946_ & new_n5945_;
  assign new_n4567_ = new_n4566_ & new_n5947_;
  assign new_n4568_ = new_n5951_ & new_n5950_;
  assign new_n4569_ = new_n4568_ & new_n5952_;
  assign new_n4570_ = new_n5956_ & new_n5955_;
  assign new_n4571_ = new_n4570_ & new_n5957_;
  assign new_n4572_ = new_n5961_ & new_n5960_;
  assign new_n4573_ = new_n4572_ & new_n5962_;
  assign new_n4574_ = new_n5966_ & new_n5965_;
  assign new_n4575_ = new_n4574_ & new_n5967_;
  assign new_n4576_ = new_n5971_ & new_n5970_;
  assign new_n4577_ = new_n4576_ & new_n5972_;
  assign new_n4578_ = pi0313 & new_n4285_;
  assign new_n4579_ = new_n5982_ & new_n5468_;
  assign new_n4580_ = new_n5987_ & new_n5986_;
  assign new_n4581_ = new_n4580_ & new_n5988_;
  assign new_n4582_ = new_n5992_ & new_n5991_;
  assign new_n4583_ = new_n4582_ & new_n5993_;
  assign new_n4584_ = new_n5997_ & new_n5996_;
  assign new_n4585_ = new_n4584_ & new_n5998_;
  assign new_n4586_ = new_n6002_ & new_n6001_;
  assign new_n4587_ = new_n4586_ & new_n6003_;
  assign new_n4588_ = new_n6007_ & new_n6006_;
  assign new_n4589_ = new_n4588_ & new_n6008_;
  assign new_n4590_ = new_n6012_ & new_n6011_;
  assign new_n4591_ = new_n4590_ & new_n6013_;
  assign new_n4592_ = new_n6017_ & new_n6016_;
  assign new_n4593_ = new_n4592_ & new_n6018_;
  assign new_n4594_ = new_n6022_ & new_n6021_;
  assign new_n4595_ = new_n4594_ & new_n6023_;
  assign new_n4596_ = new_n6034_ & new_n5468_;
  assign new_n4597_ = new_n6039_ & new_n6038_;
  assign new_n4598_ = new_n4597_ & new_n6040_;
  assign new_n4599_ = new_n6044_ & new_n6043_;
  assign new_n4600_ = new_n4599_ & new_n6045_;
  assign new_n4601_ = new_n6049_ & new_n6048_;
  assign new_n4602_ = new_n4601_ & new_n6050_;
  assign new_n4603_ = new_n6054_ & new_n6053_;
  assign new_n4604_ = new_n4603_ & new_n6055_;
  assign new_n4605_ = new_n6059_ & new_n6058_;
  assign new_n4606_ = new_n4605_ & new_n6060_;
  assign new_n4607_ = new_n6064_ & new_n6063_;
  assign new_n4608_ = new_n4607_ & new_n6065_;
  assign new_n4609_ = new_n6069_ & new_n6068_;
  assign new_n4610_ = new_n4609_ & new_n6070_;
  assign new_n4611_ = new_n6074_ & new_n6073_;
  assign new_n4612_ = new_n4611_ & new_n6075_;
  assign new_n4613_ = pi0313 & pi0315;
  assign new_n4614_ = new_n6086_ & new_n5468_;
  assign new_n4615_ = new_n6091_ & new_n6090_;
  assign new_n4616_ = new_n4615_ & new_n6092_;
  assign new_n4617_ = new_n6096_ & new_n6095_;
  assign new_n4618_ = new_n4617_ & new_n6097_;
  assign new_n4619_ = new_n6101_ & new_n6100_;
  assign new_n4620_ = new_n4619_ & new_n6102_;
  assign new_n4621_ = new_n6106_ & new_n6105_;
  assign new_n4622_ = new_n4621_ & new_n6107_;
  assign new_n4623_ = new_n6111_ & new_n6110_;
  assign new_n4624_ = new_n4623_ & new_n6112_;
  assign new_n4625_ = new_n6116_ & new_n6115_;
  assign new_n4626_ = new_n4625_ & new_n6117_;
  assign new_n4627_ = new_n6121_ & new_n6120_;
  assign new_n4628_ = new_n4627_ & new_n6122_;
  assign new_n4629_ = new_n6126_ & new_n6125_;
  assign new_n4630_ = new_n4629_ & new_n6127_;
  assign new_n4631_ = pi0313 & new_n4287_;
  assign new_n4632_ = new_n6138_ & new_n5468_;
  assign new_n4633_ = new_n6143_ & new_n6142_;
  assign new_n4634_ = new_n4633_ & new_n6144_;
  assign new_n4635_ = new_n6148_ & new_n6147_;
  assign new_n4636_ = new_n4635_ & new_n6149_;
  assign new_n4637_ = new_n6153_ & new_n6152_;
  assign new_n4638_ = new_n4637_ & new_n6154_;
  assign new_n4639_ = new_n6158_ & new_n6157_;
  assign new_n4640_ = new_n4639_ & new_n6159_;
  assign new_n4641_ = new_n6163_ & new_n6162_;
  assign new_n4642_ = new_n4641_ & new_n6164_;
  assign new_n4643_ = new_n6168_ & new_n6167_;
  assign new_n4644_ = new_n4643_ & new_n6169_;
  assign new_n4645_ = new_n6173_ & new_n6172_;
  assign new_n4646_ = new_n4645_ & new_n6174_;
  assign new_n4647_ = new_n6178_ & new_n6177_;
  assign new_n4648_ = new_n4647_ & new_n6179_;
  assign new_n4649_ = new_n6189_ & new_n5468_;
  assign new_n4650_ = new_n6194_ & new_n6193_;
  assign new_n4651_ = new_n4650_ & new_n6195_;
  assign new_n4652_ = new_n6199_ & new_n6198_;
  assign new_n4653_ = new_n4652_ & new_n6200_;
  assign new_n4654_ = new_n6204_ & new_n6203_;
  assign new_n4655_ = new_n4654_ & new_n6205_;
  assign new_n4656_ = new_n6209_ & new_n6208_;
  assign new_n4657_ = new_n4656_ & new_n6210_;
  assign new_n4658_ = new_n6214_ & new_n6213_;
  assign new_n4659_ = new_n4658_ & new_n6215_;
  assign new_n4660_ = new_n6219_ & new_n6218_;
  assign new_n4661_ = new_n4660_ & new_n6220_;
  assign new_n4662_ = new_n6224_ & new_n6223_;
  assign new_n4663_ = new_n4662_ & new_n6225_;
  assign new_n4664_ = new_n6229_ & new_n6228_;
  assign new_n4665_ = new_n4664_ & new_n6230_;
  assign new_n4666_ = new_n6238_ & new_n5468_;
  assign new_n4667_ = new_n6243_ & new_n6242_;
  assign new_n4668_ = new_n4667_ & new_n6244_;
  assign new_n4669_ = new_n6248_ & new_n6247_;
  assign new_n4670_ = new_n4669_ & new_n6249_;
  assign new_n4671_ = new_n6253_ & new_n6252_;
  assign new_n4672_ = new_n4671_ & new_n6254_;
  assign new_n4673_ = new_n6258_ & new_n6257_;
  assign new_n4674_ = new_n4673_ & new_n6259_;
  assign new_n4675_ = new_n6263_ & new_n6262_;
  assign new_n4676_ = new_n4675_ & new_n6264_;
  assign new_n4677_ = new_n6268_ & new_n6267_;
  assign new_n4678_ = new_n4677_ & new_n6269_;
  assign new_n4679_ = new_n6273_ & new_n6272_;
  assign new_n4680_ = new_n4679_ & new_n6274_;
  assign new_n4681_ = new_n6278_ & new_n6277_;
  assign new_n4682_ = new_n4681_ & new_n6279_;
  assign new_n4683_ = pi0315 & new_n4289_;
  assign new_n4684_ = new_n6290_ & new_n5468_;
  assign new_n4685_ = new_n6295_ & new_n6294_;
  assign new_n4686_ = new_n4685_ & new_n6296_;
  assign new_n4687_ = new_n6300_ & new_n6299_;
  assign new_n4688_ = new_n4687_ & new_n6301_;
  assign new_n4689_ = new_n6305_ & new_n6304_;
  assign new_n4690_ = new_n4689_ & new_n6306_;
  assign new_n4691_ = new_n6310_ & new_n6309_;
  assign new_n4692_ = new_n4691_ & new_n6311_;
  assign new_n4693_ = new_n6315_ & new_n6314_;
  assign new_n4694_ = new_n4693_ & new_n6316_;
  assign new_n4695_ = new_n6320_ & new_n6319_;
  assign new_n4696_ = new_n4695_ & new_n6321_;
  assign new_n4697_ = new_n6325_ & new_n6324_;
  assign new_n4698_ = new_n4697_ & new_n6326_;
  assign new_n4699_ = new_n6330_ & new_n6329_;
  assign new_n4700_ = new_n4699_ & new_n6331_;
  assign new_n4701_ = pi0314 & new_n4289_;
  assign new_n4702_ = new_n6342_ & new_n5468_;
  assign new_n4703_ = new_n6347_ & new_n6346_;
  assign new_n4704_ = new_n4703_ & new_n6348_;
  assign new_n4705_ = new_n6352_ & new_n6351_;
  assign new_n4706_ = new_n4705_ & new_n6353_;
  assign new_n4707_ = new_n6357_ & new_n6356_;
  assign new_n4708_ = new_n4707_ & new_n6358_;
  assign new_n4709_ = new_n6362_ & new_n6361_;
  assign new_n4710_ = new_n4709_ & new_n6363_;
  assign new_n4711_ = new_n6367_ & new_n6366_;
  assign new_n4712_ = new_n4711_ & new_n6368_;
  assign new_n4713_ = new_n6372_ & new_n6371_;
  assign new_n4714_ = new_n4713_ & new_n6373_;
  assign new_n4715_ = new_n6377_ & new_n6376_;
  assign new_n4716_ = new_n4715_ & new_n6378_;
  assign new_n4717_ = new_n6382_ & new_n6381_;
  assign new_n4718_ = new_n4717_ & new_n6383_;
  assign new_n4719_ = ~pi0313 & ~pi0315;
  assign new_n4720_ = new_n6393_ & new_n5468_;
  assign new_n4721_ = new_n6399_ & new_n6397_ & new_n6396_;
  assign new_n4722_ = new_n4721_ & new_n6398_;
  assign new_n4723_ = new_n6404_ & new_n6402_ & new_n6401_;
  assign new_n4724_ = new_n4723_ & new_n6403_;
  assign new_n4725_ = new_n6409_ & new_n6407_ & new_n6406_;
  assign new_n4726_ = new_n4725_ & new_n6408_;
  assign new_n4727_ = new_n6414_ & new_n6412_ & new_n6411_;
  assign new_n4728_ = new_n4727_ & new_n6413_;
  assign new_n4729_ = new_n6419_ & new_n6417_ & new_n6416_;
  assign new_n4730_ = new_n4729_ & new_n6418_;
  assign new_n4731_ = new_n6424_ & new_n6422_ & new_n6421_;
  assign new_n4732_ = new_n4731_ & new_n6423_;
  assign new_n4733_ = new_n6429_ & new_n6427_ & new_n6426_;
  assign new_n4734_ = new_n4733_ & new_n6428_;
  assign new_n4735_ = new_n6434_ & new_n6432_ & new_n6431_;
  assign new_n4736_ = new_n4735_ & new_n6433_;
  assign new_n4737_ = ~pi0314 & ~pi0313;
  assign new_n4738_ = new_n6444_ & new_n5468_;
  assign new_n4739_ = new_n6450_ & new_n6448_ & new_n6447_;
  assign new_n4740_ = new_n4739_ & new_n6449_;
  assign new_n4741_ = new_n6455_ & new_n6453_ & new_n6452_;
  assign new_n4742_ = new_n4741_ & new_n6454_;
  assign new_n4743_ = new_n6460_ & new_n6458_ & new_n6457_;
  assign new_n4744_ = new_n4743_ & new_n6459_;
  assign new_n4745_ = new_n6465_ & new_n6463_ & new_n6462_;
  assign new_n4746_ = new_n4745_ & new_n6464_;
  assign new_n4747_ = new_n6470_ & new_n6468_ & new_n6467_;
  assign new_n4748_ = new_n4747_ & new_n6469_;
  assign new_n4749_ = new_n6475_ & new_n6473_ & new_n6472_;
  assign new_n4750_ = new_n4749_ & new_n6474_;
  assign new_n4751_ = new_n6480_ & new_n6478_ & new_n6477_;
  assign new_n4752_ = new_n4751_ & new_n6479_;
  assign new_n4753_ = new_n6485_ & new_n6483_ & new_n6482_;
  assign new_n4754_ = new_n4753_ & new_n6484_;
  assign new_n4755_ = new_n6495_ & new_n5468_;
  assign new_n4756_ = new_n6501_ & new_n6499_ & new_n6498_;
  assign new_n4757_ = new_n4756_ & new_n6500_;
  assign new_n4758_ = new_n6506_ & new_n6504_ & new_n6503_;
  assign new_n4759_ = new_n4758_ & new_n6505_;
  assign new_n4760_ = new_n6511_ & new_n6509_ & new_n6508_;
  assign new_n4761_ = new_n4760_ & new_n6510_;
  assign new_n4762_ = new_n6516_ & new_n6514_ & new_n6513_;
  assign new_n4763_ = new_n4762_ & new_n6515_;
  assign new_n4764_ = new_n6521_ & new_n6519_ & new_n6518_;
  assign new_n4765_ = new_n4764_ & new_n6520_;
  assign new_n4766_ = new_n6526_ & new_n6524_ & new_n6523_;
  assign new_n4767_ = new_n4766_ & new_n6525_;
  assign new_n4768_ = new_n6531_ & new_n6529_ & new_n6528_;
  assign new_n4769_ = new_n4768_ & new_n6530_;
  assign new_n4770_ = new_n6536_ & new_n6534_ & new_n6533_;
  assign new_n4771_ = new_n4770_ & new_n6535_;
  assign new_n4772_ = ~pi0314 & ~pi0313;
  assign new_n4773_ = new_n6546_ & new_n5468_;
  assign new_n4774_ = new_n6552_ & new_n6550_ & new_n6549_;
  assign new_n4775_ = new_n4774_ & new_n6551_;
  assign new_n4776_ = new_n6557_ & new_n6555_ & new_n6554_;
  assign new_n4777_ = new_n4776_ & new_n6556_;
  assign new_n4778_ = new_n6562_ & new_n6560_ & new_n6559_;
  assign new_n4779_ = new_n4778_ & new_n6561_;
  assign new_n4780_ = new_n6567_ & new_n6565_ & new_n6564_;
  assign new_n4781_ = new_n4780_ & new_n6566_;
  assign new_n4782_ = new_n6572_ & new_n6570_ & new_n6569_;
  assign new_n4783_ = new_n4782_ & new_n6571_;
  assign new_n4784_ = new_n6577_ & new_n6575_ & new_n6574_;
  assign new_n4785_ = new_n4784_ & new_n6576_;
  assign new_n4786_ = new_n6582_ & new_n6580_ & new_n6579_;
  assign new_n4787_ = new_n4786_ & new_n6581_;
  assign new_n4788_ = new_n6587_ & new_n6585_ & new_n6584_;
  assign new_n4789_ = new_n4788_ & new_n6586_;
  assign new_n4790_ = ~pi0313 & ~pi0315;
  assign new_n4791_ = new_n6596_ & new_n5468_;
  assign new_n4792_ = new_n6602_ & new_n6600_ & new_n6599_;
  assign new_n4793_ = new_n4792_ & new_n6601_;
  assign new_n4794_ = new_n6607_ & new_n6605_ & new_n6604_;
  assign new_n4795_ = new_n4794_ & new_n6606_;
  assign new_n4796_ = new_n6612_ & new_n6610_ & new_n6609_;
  assign new_n4797_ = new_n4796_ & new_n6611_;
  assign new_n4798_ = new_n6617_ & new_n6615_ & new_n6614_;
  assign new_n4799_ = new_n4798_ & new_n6616_;
  assign new_n4800_ = new_n6622_ & new_n6620_ & new_n6619_;
  assign new_n4801_ = new_n4800_ & new_n6621_;
  assign new_n4802_ = new_n6627_ & new_n6625_ & new_n6624_;
  assign new_n4803_ = new_n4802_ & new_n6626_;
  assign new_n4804_ = new_n6632_ & new_n6630_ & new_n6629_;
  assign new_n4805_ = new_n4804_ & new_n6631_;
  assign new_n4806_ = new_n6637_ & new_n6635_ & new_n6634_;
  assign new_n4807_ = new_n4806_ & new_n6636_;
  assign new_n4808_ = new_n5496_ & new_n27131_;
  assign new_n4809_ = pi0545 & pi0178;
  assign new_n4810_ = new_n5678_ & new_n4260_;
  assign new_n4811_ = new_n4263_ & new_n4274_;
  assign new_n4812_ = new_n6651_ & new_n5489_;
  assign new_n4813_ = new_n4812_ & new_n6650_;
  assign new_n4814_ = new_n6654_ & new_n5486_;
  assign new_n4815_ = new_n6658_ & new_n6657_;
  assign new_n4816_ = new_n5712_ & new_n5695_;
  assign new_n4817_ = new_n3617_ & new_n5453_;
  assign new_n4818_ = new_n5746_ & new_n4257_;
  assign new_n4819_ = new_n5712_ & new_n4257_;
  assign new_n4820_ = new_n5729_ & new_n5480_;
  assign new_n4821_ = new_n6664_ & new_n6667_ & new_n6666_;
  assign new_n4822_ = new_n6676_ & new_n6675_ & new_n5495_;
  assign new_n4823_ = new_n9133_ & new_n4822_ & new_n6677_ & new_n9134_;
  assign new_n4824_ = new_n3673_ & new_n6684_ & new_n4398_;
  assign new_n4825_ = pi0310 & new_n5626_;
  assign new_n4826_ = pi0308 & new_n4249_;
  assign new_n4827_ = new_n4275_ & new_n4272_ & new_n4273_;
  assign new_n4828_ = new_n4827_ & new_n4401_ & new_n4400_;
  assign new_n4829_ = new_n5661_ & new_n3612_;
  assign new_n4830_ = new_n6689_ & new_n6688_;
  assign new_n4831_ = new_n6694_ & new_n6692_;
  assign new_n4832_ = new_n4831_ & new_n4833_ & new_n6695_;
  assign new_n4833_ = new_n6696_ & new_n6697_;
  assign new_n4834_ = new_n6708_ & new_n6706_;
  assign new_n4835_ = new_n4834_ & new_n6707_;
  assign new_n4836_ = new_n6711_ & new_n6710_;
  assign new_n4837_ = new_n4838_ & new_n6718_;
  assign new_n4838_ = new_n6721_ & new_n6720_;
  assign new_n4839_ = new_n6724_ & new_n6723_;
  assign new_n4840_ = new_n6732_ & new_n6730_;
  assign new_n4841_ = new_n6743_ & new_n6744_;
  assign new_n4842_ = new_n6750_ & new_n6748_;
  assign new_n4843_ = new_n6782_ & new_n6781_ & new_n5489_;
  assign new_n4844_ = new_n3612_ & new_n5452_;
  assign new_n4845_ = new_n3612_ & new_n5479_;
  assign new_n4846_ = new_n5764_ & new_n5712_;
  assign new_n4847_ = new_n3612_ & new_n5746_;
  assign new_n4848_ = new_n6792_ & new_n6791_;
  assign new_n4849_ = new_n6794_ & new_n6788_ & new_n6789_ & new_n4850_ & new_n6793_;
  assign new_n4850_ = new_n4851_ & new_n6797_;
  assign new_n4851_ = new_n6795_ & new_n6796_;
  assign new_n4852_ = new_n6799_ & new_n6801_ & new_n6802_ & new_n6800_ & new_n6798_;
  assign new_n4853_ = new_n6804_ & new_n6806_ & new_n6807_ & new_n6803_ & new_n6805_;
  assign new_n4854_ = new_n4853_ & new_n4852_;
  assign new_n4855_ = new_n6816_ & new_n6815_;
  assign new_n4856_ = new_n6817_ & new_n6813_ & new_n4857_ & new_n6818_;
  assign new_n4857_ = new_n4858_ & new_n6821_;
  assign new_n4858_ = new_n6819_ & new_n6820_;
  assign new_n4859_ = new_n6823_ & new_n6825_ & new_n6826_ & new_n6824_ & new_n6822_;
  assign new_n4860_ = new_n6827_ & new_n6829_ & new_n6828_ & new_n6830_;
  assign new_n4861_ = new_n6831_ & new_n4860_ & new_n4859_;
  assign new_n4862_ = new_n4863_ & new_n6837_;
  assign new_n4863_ = new_n6840_ & new_n6839_;
  assign new_n4864_ = new_n4865_ & new_n6845_;
  assign new_n4865_ = new_n6843_ & new_n6844_;
  assign new_n4866_ = new_n4864_ & new_n6842_ & new_n6841_;
  assign new_n4867_ = new_n6847_ & new_n6849_ & new_n6850_ & new_n6848_ & new_n6846_;
  assign new_n4868_ = new_n6851_ & new_n6853_ & new_n6852_ & new_n6854_;
  assign new_n4869_ = new_n6855_ & new_n4868_ & new_n4867_;
  assign new_n4870_ = new_n6861_ & new_n6860_;
  assign new_n4871_ = new_n6864_ & new_n6863_;
  assign new_n4872_ = new_n4873_ & new_n6869_;
  assign new_n4873_ = new_n6867_ & new_n6868_;
  assign new_n4874_ = new_n4872_ & new_n6866_ & new_n6865_;
  assign new_n4875_ = new_n6871_ & new_n6873_ & new_n6874_ & new_n6872_ & new_n6870_;
  assign new_n4876_ = new_n6875_ & new_n6877_ & new_n6876_ & new_n6878_;
  assign new_n4877_ = new_n6879_ & new_n4876_ & new_n4875_;
  assign new_n4878_ = new_n4879_ & new_n6885_;
  assign new_n4879_ = new_n6888_ & new_n6887_;
  assign new_n4880_ = new_n4881_ & new_n6893_;
  assign new_n4881_ = new_n6891_ & new_n6892_;
  assign new_n4882_ = new_n4880_ & new_n6890_ & new_n6889_;
  assign new_n4883_ = new_n6895_ & new_n6897_ & new_n6898_ & new_n6896_ & new_n6894_;
  assign new_n4884_ = new_n6899_ & new_n6901_ & new_n6900_ & new_n6902_;
  assign new_n4885_ = new_n6903_ & new_n4884_ & new_n4883_;
  assign new_n4886_ = new_n4887_ & new_n6908_;
  assign new_n4887_ = new_n6912_ & new_n6911_;
  assign new_n4888_ = new_n4889_ & new_n6917_;
  assign new_n4889_ = new_n6915_ & new_n6916_;
  assign new_n4890_ = new_n4888_ & new_n6914_ & new_n6913_;
  assign new_n4891_ = new_n6919_ & new_n6921_ & new_n6922_ & new_n6920_ & new_n6918_;
  assign new_n4892_ = new_n6923_ & new_n6925_ & new_n6924_ & new_n6926_;
  assign new_n4893_ = new_n6927_ & new_n4892_ & new_n4891_;
  assign new_n4894_ = new_n4895_ & new_n6932_;
  assign new_n4895_ = new_n6936_ & new_n6935_;
  assign new_n4896_ = new_n4897_ & new_n6941_;
  assign new_n4897_ = new_n6939_ & new_n6940_;
  assign new_n4898_ = new_n4896_ & new_n6938_ & new_n6937_;
  assign new_n4899_ = new_n6943_ & new_n6945_ & new_n6946_ & new_n6944_ & new_n6942_;
  assign new_n4900_ = new_n6947_ & new_n6949_ & new_n6948_ & new_n6950_;
  assign new_n4901_ = new_n6951_ & new_n4900_ & new_n4899_;
  assign new_n4902_ = new_n4903_ & new_n6956_;
  assign new_n4903_ = new_n6960_ & new_n6959_;
  assign new_n4904_ = new_n4905_ & new_n6965_;
  assign new_n4905_ = new_n6963_ & new_n6964_;
  assign new_n4906_ = new_n4904_ & new_n6962_ & new_n6961_;
  assign new_n4907_ = new_n6967_ & new_n6969_ & new_n6970_ & new_n6968_ & new_n6966_;
  assign new_n4908_ = new_n6971_ & new_n6973_ & new_n6972_ & new_n6974_;
  assign new_n4909_ = new_n6975_ & new_n4908_ & new_n4907_;
  assign new_n4910_ = new_n4911_ & new_n6980_;
  assign new_n4911_ = new_n6984_ & new_n6983_;
  assign new_n4912_ = new_n6987_ & new_n6989_ & new_n6988_;
  assign new_n4913_ = new_n4912_ & new_n6986_ & new_n6985_;
  assign new_n4914_ = new_n6991_ & new_n6993_ & new_n6994_ & new_n6992_ & new_n6990_;
  assign new_n4915_ = new_n6997_ & new_n6995_ & new_n6996_ & new_n6998_;
  assign new_n4916_ = new_n6999_ & new_n4915_ & new_n4914_;
  assign new_n4917_ = new_n4918_ & new_n7004_;
  assign new_n4918_ = new_n7008_ & new_n7007_;
  assign new_n4919_ = new_n7013_ & new_n7012_;
  assign new_n4920_ = new_n7009_ & new_n4919_ & new_n7011_ & new_n7010_;
  assign new_n4921_ = new_n7015_ & new_n7017_ & new_n7018_ & new_n7016_ & new_n7014_;
  assign new_n4922_ = new_n7021_ & new_n7019_ & new_n7020_ & new_n7022_;
  assign new_n4923_ = new_n7023_ & new_n4922_ & new_n4921_;
  assign new_n4924_ = new_n4925_ & new_n7029_;
  assign new_n4925_ = new_n7032_ & new_n7031_;
  assign new_n4926_ = new_n7037_ & new_n7036_;
  assign new_n4927_ = new_n7033_ & new_n4926_ & new_n7035_ & new_n7034_;
  assign new_n4928_ = new_n7039_ & new_n7041_ & new_n7042_ & new_n7040_ & new_n7038_;
  assign new_n4929_ = new_n7045_ & new_n7043_ & new_n7044_ & new_n7046_;
  assign new_n4930_ = new_n7047_ & new_n4929_ & new_n4928_;
  assign new_n4931_ = new_n4932_ & new_n7053_;
  assign new_n4932_ = new_n7056_ & new_n7055_;
  assign new_n4933_ = new_n7061_ & new_n7060_;
  assign new_n4934_ = new_n7057_ & new_n4933_ & new_n7059_ & new_n7058_;
  assign new_n4935_ = new_n7063_ & new_n7065_ & new_n7066_ & new_n7064_ & new_n7062_;
  assign new_n4936_ = new_n7069_ & new_n7067_ & new_n7068_ & new_n7070_;
  assign new_n4937_ = new_n7071_ & new_n4936_ & new_n4935_;
  assign new_n4938_ = new_n4939_ & new_n7076_;
  assign new_n4939_ = new_n7080_ & new_n7079_;
  assign new_n4940_ = new_n7085_ & new_n7084_;
  assign new_n4941_ = new_n7081_ & new_n4940_ & new_n7083_ & new_n7082_;
  assign new_n4942_ = new_n7087_ & new_n7089_ & new_n7090_ & new_n7088_ & new_n7086_;
  assign new_n4943_ = new_n7093_ & new_n7091_ & new_n7092_ & new_n7094_;
  assign new_n4944_ = new_n7095_ & new_n4943_ & new_n4942_;
  assign new_n4945_ = new_n4946_ & new_n7100_;
  assign new_n4946_ = new_n7104_ & new_n7103_;
  assign new_n4947_ = new_n7109_ & new_n7108_;
  assign new_n4948_ = new_n7105_ & new_n4947_ & new_n7107_ & new_n7106_;
  assign new_n4949_ = new_n7111_ & new_n7113_ & new_n7114_ & new_n7112_ & new_n7110_;
  assign new_n4950_ = new_n7117_ & new_n7115_ & new_n7116_ & new_n7118_;
  assign new_n4951_ = new_n7119_ & new_n4950_ & new_n4949_;
  assign new_n4952_ = new_n7128_ & new_n7127_;
  assign new_n4953_ = new_n7133_ & new_n7132_;
  assign new_n4954_ = new_n7129_ & new_n4953_ & new_n7131_ & new_n7130_;
  assign new_n4955_ = new_n4952_ & new_n7124_ & new_n7125_ & new_n4954_ & new_n7126_;
  assign new_n4956_ = new_n7135_ & new_n7137_ & new_n7138_ & new_n7136_ & new_n7134_;
  assign new_n4957_ = new_n7141_ & new_n7139_ & new_n7140_ & new_n7142_;
  assign new_n4958_ = new_n7143_ & new_n4957_ & new_n4956_;
  assign new_n4959_ = new_n7147_ & new_n7145_;
  assign new_n4960_ = new_n7152_ & new_n7151_;
  assign new_n4961_ = new_n7157_ & new_n7156_;
  assign new_n4962_ = new_n7153_ & new_n4961_ & new_n7155_ & new_n7154_;
  assign new_n4963_ = new_n4960_ & new_n7148_ & new_n7149_ & new_n4962_ & new_n7150_;
  assign new_n4964_ = new_n7159_ & new_n7161_ & new_n7162_ & new_n7160_ & new_n7158_;
  assign new_n4965_ = new_n7165_ & new_n7163_ & new_n7164_ & new_n7166_;
  assign new_n4966_ = new_n7167_ & new_n4965_ & new_n4964_;
  assign new_n4967_ = new_n7171_ & new_n7169_;
  assign new_n4968_ = new_n4969_ & new_n7173_;
  assign new_n4969_ = new_n7176_ & new_n7175_;
  assign new_n4970_ = new_n7181_ & new_n7180_;
  assign new_n4971_ = new_n7177_ & new_n4970_ & new_n7179_ & new_n7178_;
  assign new_n4972_ = new_n7183_ & new_n7185_ & new_n7186_ & new_n7184_ & new_n7182_;
  assign new_n4973_ = new_n7189_ & new_n7187_ & new_n7188_ & new_n7190_;
  assign new_n4974_ = new_n7191_ & new_n4973_ & new_n4972_;
  assign new_n4975_ = new_n7200_ & new_n7199_;
  assign new_n4976_ = new_n7202_ & new_n7197_ & new_n4977_ & new_n7203_ & new_n7201_;
  assign new_n4977_ = new_n7205_ & new_n7204_;
  assign new_n4978_ = new_n7207_ & new_n7209_ & new_n7210_ & new_n7208_ & new_n7206_;
  assign new_n4979_ = new_n7213_ & new_n7211_ & new_n7212_ & new_n7214_;
  assign new_n4980_ = new_n7215_ & new_n4979_ & new_n4978_;
  assign new_n4981_ = new_n4982_ & new_n7221_;
  assign new_n4982_ = new_n7224_ & new_n7223_;
  assign new_n4983_ = new_n7229_ & new_n7228_;
  assign new_n4984_ = new_n7225_ & new_n4983_ & new_n7227_ & new_n7226_;
  assign new_n4985_ = new_n7231_ & new_n7233_ & new_n7234_ & new_n7232_ & new_n7230_;
  assign new_n4986_ = new_n7237_ & new_n7235_ & new_n7236_ & new_n7238_;
  assign new_n4987_ = new_n7239_ & new_n4986_ & new_n4985_;
  assign new_n4988_ = new_n7248_ & new_n7247_;
  assign new_n4989_ = new_n7250_ & new_n7245_ & new_n4990_ & new_n7251_ & new_n7249_;
  assign new_n4990_ = new_n7253_ & new_n7252_;
  assign new_n4991_ = new_n7255_ & new_n7257_ & new_n7258_ & new_n7256_ & new_n7254_;
  assign new_n4992_ = new_n7261_ & new_n7259_ & new_n7260_ & new_n7262_;
  assign new_n4993_ = new_n7263_ & new_n4992_ & new_n4991_;
  assign new_n4994_ = new_n7272_ & new_n7271_;
  assign new_n4995_ = new_n7277_ & new_n7276_;
  assign new_n4996_ = new_n7273_ & new_n4995_ & new_n7275_ & new_n7274_;
  assign new_n4997_ = new_n7270_ & new_n5000_ & new_n7268_ & new_n4996_ & new_n4994_;
  assign new_n4998_ = new_n7279_ & new_n7281_ & new_n7282_ & new_n7280_ & new_n7278_;
  assign new_n4999_ = new_n7285_ & new_n7283_ & new_n7284_ & new_n7286_;
  assign new_n5000_ = new_n7287_ & new_n4999_ & new_n4998_;
  assign new_n5001_ = new_n7291_ & new_n7289_;
  assign new_n5002_ = new_n7296_ & new_n7295_;
  assign new_n5003_ = new_n7301_ & new_n7300_;
  assign new_n5004_ = new_n7297_ & new_n5003_ & new_n7299_ & new_n7298_;
  assign new_n5005_ = new_n7294_ & new_n5008_ & new_n7292_ & new_n5004_ & new_n5002_;
  assign new_n5006_ = new_n7303_ & new_n7305_ & new_n7306_ & new_n7304_ & new_n7302_;
  assign new_n5007_ = new_n7309_ & new_n7307_ & new_n7308_ & new_n7310_;
  assign new_n5008_ = new_n7311_ & new_n5006_ & new_n5007_;
  assign new_n5009_ = new_n7315_ & new_n7313_;
  assign new_n5010_ = new_n7320_ & new_n7319_;
  assign new_n5011_ = new_n7325_ & new_n7324_;
  assign new_n5012_ = new_n7321_ & new_n5011_ & new_n7323_ & new_n7322_;
  assign new_n5013_ = new_n7317_ & new_n7316_ & new_n5012_ & new_n5010_ & new_n7318_;
  assign new_n5014_ = new_n7328_ & new_n7327_ & new_n7326_;
  assign new_n5015_ = new_n7330_ & new_n7329_;
  assign new_n5016_ = new_n7333_ & new_n7332_ & new_n7331_;
  assign new_n5017_ = new_n7335_ & new_n7334_;
  assign new_n5018_ = new_n5014_ & new_n5017_ & new_n5016_ & new_n5015_;
  assign new_n5019_ = new_n7339_ & new_n7337_;
  assign new_n5020_ = new_n7344_ & new_n7343_;
  assign new_n5021_ = new_n7349_ & new_n7348_;
  assign new_n5022_ = new_n7345_ & new_n5021_ & new_n7347_ & new_n7346_;
  assign new_n5023_ = new_n7341_ & new_n7340_ & new_n5022_ & new_n5020_ & new_n7342_;
  assign new_n5024_ = new_n7352_ & new_n7351_ & new_n7350_;
  assign new_n5025_ = new_n7354_ & new_n7353_;
  assign new_n5026_ = new_n7357_ & new_n7356_ & new_n7355_;
  assign new_n5027_ = new_n7359_ & new_n7358_;
  assign new_n5028_ = new_n5024_ & new_n5027_ & new_n5026_ & new_n5025_;
  assign new_n5029_ = new_n7363_ & new_n7361_;
  assign new_n5030_ = new_n7368_ & new_n7367_;
  assign new_n5031_ = new_n7373_ & new_n7372_;
  assign new_n5032_ = new_n7369_ & new_n5031_ & new_n7371_ & new_n7370_;
  assign new_n5033_ = new_n7365_ & new_n5032_ & new_n7364_ & new_n5030_ & new_n7366_;
  assign new_n5034_ = new_n7376_ & new_n7375_ & new_n7374_;
  assign new_n5035_ = new_n7378_ & new_n7377_;
  assign new_n5036_ = new_n7381_ & new_n7380_ & new_n7379_;
  assign new_n5037_ = new_n7383_ & new_n7382_;
  assign new_n5038_ = new_n5034_ & new_n5036_ & new_n5037_ & new_n5035_;
  assign new_n5039_ = new_n7387_ & new_n7385_;
  assign new_n5040_ = new_n7392_ & new_n7391_;
  assign new_n5041_ = new_n7397_ & new_n7396_;
  assign new_n5042_ = new_n7393_ & new_n5041_ & new_n7395_ & new_n7394_;
  assign new_n5043_ = new_n7389_ & new_n5042_ & new_n5040_ & new_n7388_ & new_n7390_;
  assign new_n5044_ = new_n7400_ & new_n7399_ & new_n7398_;
  assign new_n5045_ = new_n7402_ & new_n7401_;
  assign new_n5046_ = new_n7405_ & new_n7404_ & new_n7403_;
  assign new_n5047_ = new_n7407_ & new_n7406_;
  assign new_n5048_ = new_n5044_ & new_n5046_ & new_n5047_ & new_n5045_;
  assign new_n5049_ = new_n7411_ & new_n7409_;
  assign new_n5050_ = new_n7413_ & new_n7412_;
  assign new_n5051_ = new_n7416_ & new_n7415_;
  assign new_n5052_ = new_n7421_ & new_n7420_;
  assign new_n5053_ = new_n7417_ & new_n5052_ & new_n7419_ & new_n7418_;
  assign new_n5054_ = new_n7424_ & new_n7423_ & new_n7422_;
  assign new_n5055_ = new_n7426_ & new_n7425_;
  assign new_n5056_ = new_n7429_ & new_n7428_ & new_n7427_;
  assign new_n5057_ = new_n7431_ & new_n7430_;
  assign new_n5058_ = new_n5054_ & new_n5056_ & new_n5057_ & new_n5055_;
  assign new_n5059_ = new_n7437_ & new_n7436_;
  assign new_n5060_ = new_n7440_ & new_n7439_;
  assign new_n5061_ = new_n7445_ & new_n7444_;
  assign new_n5062_ = new_n7441_ & new_n5061_ & new_n7443_ & new_n7442_;
  assign new_n5063_ = new_n7448_ & new_n7447_ & new_n7446_;
  assign new_n5064_ = new_n7450_ & new_n7449_;
  assign new_n5065_ = new_n7453_ & new_n7452_ & new_n7451_;
  assign new_n5066_ = new_n7455_ & new_n7454_;
  assign new_n5067_ = new_n5063_ & new_n5065_ & new_n5066_ & new_n5064_;
  assign new_n5068_ = new_n7461_ & new_n7460_;
  assign new_n5069_ = new_n7464_ & new_n7463_;
  assign new_n5070_ = new_n7469_ & new_n7468_;
  assign new_n5071_ = new_n7465_ & new_n5070_ & new_n7467_ & new_n7466_;
  assign new_n5072_ = new_n7472_ & new_n7471_ & new_n7470_;
  assign new_n5073_ = new_n7474_ & new_n7473_;
  assign new_n5074_ = new_n7477_ & new_n7476_ & new_n7475_;
  assign new_n5075_ = new_n7479_ & new_n7478_;
  assign new_n5076_ = new_n5072_ & new_n5074_ & new_n5075_ & new_n5073_;
  assign new_n5077_ = new_n7485_ & new_n7484_;
  assign new_n5078_ = new_n7488_ & new_n7487_;
  assign new_n5079_ = new_n7493_ & new_n7492_;
  assign new_n5080_ = new_n7489_ & new_n5079_ & new_n7491_ & new_n7490_;
  assign new_n5081_ = new_n7496_ & new_n7495_ & new_n7494_;
  assign new_n5082_ = new_n7498_ & new_n7497_;
  assign new_n5083_ = new_n7501_ & new_n7500_ & new_n7499_;
  assign new_n5084_ = new_n7503_ & new_n7502_;
  assign new_n5085_ = new_n5081_ & new_n5083_ & new_n5084_ & new_n5082_;
  assign new_n5086_ = new_n7509_ & new_n7508_;
  assign new_n5087_ = new_n7512_ & new_n7511_;
  assign new_n5088_ = new_n7517_ & new_n7516_;
  assign new_n5089_ = new_n7513_ & new_n5088_ & new_n7515_ & new_n7514_;
  assign new_n5090_ = new_n7520_ & new_n7519_ & new_n7518_;
  assign new_n5091_ = new_n7522_ & new_n7521_;
  assign new_n5092_ = new_n7525_ & new_n7524_ & new_n7523_;
  assign new_n5093_ = new_n7527_ & new_n7526_;
  assign new_n5094_ = new_n5090_ & new_n5092_ & new_n5093_ & new_n5091_;
  assign new_n5095_ = new_n7554_ & new_n4403_;
  assign new_n5096_ = new_n7533_ & new_n7532_;
  assign new_n5097_ = new_n7536_ & new_n7535_;
  assign new_n5098_ = new_n5097_ & new_n7537_;
  assign new_n5099_ = new_n7540_ & new_n7542_ & new_n7541_;
  assign new_n5100_ = new_n5099_ & new_n7539_ & new_n7538_;
  assign new_n5101_ = new_n7534_ & new_n5100_ & new_n5098_ & new_n5096_;
  assign new_n5102_ = new_n7545_ & new_n7544_ & new_n7543_;
  assign new_n5103_ = new_n7547_ & new_n7546_;
  assign new_n5104_ = new_n5103_ & new_n5102_ & new_n7548_;
  assign new_n5105_ = new_n7550_ & new_n7549_;
  assign new_n5106_ = new_n7554_ & new_n5104_ & new_n5105_ & new_n7551_ & new_n7553_;
  assign new_n5107_ = pi0178 & new_n4260_;
  assign new_n5108_ = pi0176 & new_n4277_;
  assign new_n5109_ = new_n5661_ & pi0178;
  assign new_n5110_ = new_n7567_ & new_n7565_ & new_n7566_ & new_n7568_;
  assign new_n5111_ = new_n7575_ & new_n7573_ & new_n7574_ & new_n7576_;
  assign new_n5112_ = new_n7581_ & new_n7583_ & new_n7584_ & new_n7582_;
  assign new_n5113_ = new_n7589_ & new_n7591_ & new_n7592_ & new_n7590_;
  assign new_n5114_ = new_n7597_ & new_n7599_ & new_n7600_ & new_n7598_;
  assign new_n5115_ = new_n7605_ & new_n7607_ & new_n7608_ & new_n7606_;
  assign new_n5116_ = new_n7613_ & new_n7615_ & new_n7616_ & new_n7614_;
  assign new_n5117_ = new_n7621_ & new_n7623_ & new_n7624_ & new_n7622_;
  assign new_n5118_ = new_n7629_ & new_n7631_ & new_n7632_ & new_n7630_;
  assign new_n5119_ = new_n7637_ & new_n7639_ & new_n7640_ & new_n7638_;
  assign new_n5120_ = new_n7645_ & new_n7647_ & new_n7648_ & new_n7646_;
  assign new_n5121_ = new_n7653_ & new_n7655_ & new_n7656_ & new_n7654_;
  assign new_n5122_ = new_n7661_ & new_n7663_ & new_n7662_ & new_n7664_;
  assign new_n5123_ = new_n7669_ & new_n7671_ & new_n7670_ & new_n7672_;
  assign new_n5124_ = new_n7677_ & new_n7679_ & new_n7678_ & new_n7680_;
  assign new_n5125_ = new_n7685_ & new_n7687_ & new_n7686_ & new_n7688_;
  assign new_n5126_ = new_n7693_ & new_n7695_ & new_n7694_ & new_n7696_;
  assign new_n5127_ = new_n7701_ & new_n7703_ & new_n7702_ & new_n7704_;
  assign new_n5128_ = new_n7709_ & new_n7711_ & new_n7710_ & new_n7712_;
  assign new_n5129_ = new_n7717_ & new_n7719_ & new_n7718_ & new_n7720_;
  assign new_n5130_ = new_n7725_ & new_n7727_ & new_n7726_ & new_n7728_;
  assign new_n5131_ = new_n7733_ & new_n7735_ & new_n7734_ & new_n7736_;
  assign new_n5132_ = new_n7741_ & new_n7743_ & new_n7742_ & new_n7744_;
  assign new_n5133_ = new_n7749_ & new_n7751_ & new_n7750_ & new_n7752_;
  assign new_n5134_ = new_n7757_ & new_n7759_ & new_n7758_ & new_n7760_;
  assign new_n5135_ = new_n7765_ & new_n7767_ & new_n7766_ & new_n7768_;
  assign new_n5136_ = new_n7775_ & new_n7773_ & new_n7774_ & new_n7776_;
  assign new_n5137_ = new_n7783_ & new_n7781_ & new_n7782_ & new_n7784_;
  assign new_n5138_ = new_n7791_ & new_n7789_ & new_n7790_ & new_n7792_;
  assign new_n5139_ = new_n7797_ & new_n7798_ & new_n7799_ & new_n7800_;
  assign new_n5140_ = new_n7805_ & new_n7806_ & new_n7807_ & new_n7808_;
  assign new_n5141_ = new_n7813_ & new_n7814_ & new_n7815_ & new_n7816_;
  assign new_n5142_ = new_n5449_ & new_n3546_;
  assign new_n5143_ = new_n7965_ & new_n7966_;
  assign new_n5144_ = new_n7968_ & new_n7969_;
  assign new_n5145_ = new_n7971_ & new_n7972_;
  assign new_n5146_ = new_n7974_ & new_n7975_;
  assign new_n5147_ = new_n7977_ & new_n7978_;
  assign new_n5148_ = new_n7980_ & new_n7981_;
  assign new_n5149_ = new_n7983_ & new_n7984_;
  assign new_n5150_ = new_n7986_ & new_n7987_;
  assign new_n5151_ = new_n7989_ & new_n7990_;
  assign new_n5152_ = new_n7992_ & new_n7993_;
  assign new_n5153_ = new_n7995_ & new_n7996_;
  assign new_n5154_ = new_n7998_ & new_n7999_;
  assign new_n5155_ = new_n8001_ & new_n8002_;
  assign new_n5156_ = new_n8004_ & new_n8005_;
  assign new_n5157_ = new_n8007_ & new_n8008_;
  assign new_n5158_ = new_n8013_ & new_n8012_;
  assign new_n5159_ = new_n8017_ & new_n8016_;
  assign new_n5160_ = new_n8021_ & new_n8020_;
  assign new_n5161_ = new_n8025_ & new_n8024_;
  assign new_n5162_ = new_n8029_ & new_n8028_;
  assign new_n5163_ = new_n8033_ & new_n8032_;
  assign new_n5164_ = new_n8037_ & new_n8036_;
  assign new_n5165_ = new_n8041_ & new_n8040_;
  assign new_n5166_ = new_n8045_ & new_n8044_;
  assign new_n5167_ = new_n8049_ & new_n8048_;
  assign new_n5168_ = new_n8053_ & new_n8052_;
  assign new_n5169_ = new_n8057_ & new_n8056_;
  assign new_n5170_ = new_n8061_ & new_n8060_;
  assign new_n5171_ = new_n8063_ & new_n8065_;
  assign new_n5172_ = new_n8067_ & new_n8069_;
  assign new_n5173_ = new_n8071_ & new_n8073_;
  assign new_n5174_ = new_n8078_ & new_n8076_;
  assign new_n5175_ = new_n8083_ & new_n8081_;
  assign new_n5176_ = new_n8088_ & new_n8086_;
  assign new_n5177_ = new_n8093_ & new_n8091_;
  assign new_n5178_ = new_n8098_ & new_n8096_;
  assign new_n5179_ = new_n8103_ & new_n8101_;
  assign new_n5180_ = new_n8108_ & new_n8106_;
  assign new_n5181_ = new_n8113_ & new_n8111_;
  assign new_n5182_ = new_n8118_ & new_n8116_;
  assign new_n5183_ = new_n8123_ & new_n8121_;
  assign new_n5184_ = new_n8128_ & new_n8126_;
  assign new_n5185_ = new_n8133_ & new_n8131_;
  assign new_n5186_ = new_n5492_ & new_n5485_ & new_n5484_;
  assign new_n5187_ = new_n5188_ & new_n8254_ & new_n8253_;
  assign new_n5188_ = new_n8257_ & new_n8256_;
  assign new_n5189_ = new_n5190_ & new_n8260_;
  assign new_n5190_ = new_n8262_ & new_n8261_;
  assign new_n5191_ = new_n5192_ & new_n8264_ & new_n8263_;
  assign new_n5192_ = new_n8267_ & new_n8266_;
  assign new_n5193_ = new_n5194_ & new_n8270_;
  assign new_n5194_ = new_n8272_ & new_n8271_;
  assign new_n5195_ = new_n5196_ & new_n8274_ & new_n8273_;
  assign new_n5196_ = new_n8277_ & new_n8276_;
  assign new_n5197_ = new_n5198_ & new_n8280_;
  assign new_n5198_ = new_n8282_ & new_n8281_;
  assign new_n5199_ = new_n5200_ & new_n8284_ & new_n8283_;
  assign new_n5200_ = new_n8287_ & new_n8286_;
  assign new_n5201_ = new_n5202_ & new_n8290_;
  assign new_n5202_ = new_n8292_ & new_n8291_;
  assign new_n5203_ = new_n8294_ & new_n8293_ & new_n5472_;
  assign new_n5204_ = new_n8296_ & new_n8297_;
  assign new_n5205_ = new_n5206_ & new_n8300_;
  assign new_n5206_ = new_n8302_ & new_n8301_;
  assign new_n5207_ = new_n5204_ & new_n8299_ & new_n8298_ & new_n5203_ & new_n8295_;
  assign new_n5208_ = new_n8304_ & new_n8303_ & new_n5472_;
  assign new_n5209_ = new_n8306_ & new_n8307_;
  assign new_n5210_ = new_n5211_ & new_n8310_;
  assign new_n5211_ = new_n8312_ & new_n8311_;
  assign new_n5212_ = new_n5209_ & new_n8309_ & new_n8308_ & new_n5208_ & new_n8305_;
  assign new_n5213_ = new_n8314_ & new_n8313_ & new_n5472_;
  assign new_n5214_ = new_n5215_ & new_n8317_;
  assign new_n5215_ = new_n8320_ & new_n8319_;
  assign new_n5216_ = new_n8322_ & new_n8321_ & new_n5472_;
  assign new_n5217_ = new_n5218_ & new_n8325_;
  assign new_n5218_ = new_n8328_ & new_n8327_;
  assign new_n5219_ = new_n8330_ & new_n8329_ & new_n5472_;
  assign new_n5220_ = new_n5221_ & new_n8333_;
  assign new_n5221_ = new_n8336_ & new_n8335_;
  assign new_n5222_ = new_n8338_ & new_n8337_ & new_n5472_;
  assign new_n5223_ = new_n5224_ & new_n8341_;
  assign new_n5224_ = new_n8344_ & new_n8343_;
  assign new_n5225_ = new_n8346_ & new_n8345_ & new_n5472_;
  assign new_n5226_ = new_n5227_ & new_n8349_;
  assign new_n5227_ = new_n8352_ & new_n8351_;
  assign new_n5228_ = new_n8354_ & new_n8353_ & new_n5472_;
  assign new_n5229_ = new_n5230_ & new_n8357_;
  assign new_n5230_ = new_n8360_ & new_n8359_;
  assign new_n5231_ = new_n8362_ & new_n8361_ & new_n5472_;
  assign new_n5232_ = new_n5233_ & new_n8365_;
  assign new_n5233_ = new_n8368_ & new_n8367_;
  assign new_n5234_ = new_n8370_ & new_n8369_ & new_n5472_;
  assign new_n5235_ = new_n5236_ & new_n8373_;
  assign new_n5236_ = new_n8376_ & new_n8375_;
  assign new_n5237_ = new_n8378_ & new_n8377_ & new_n5472_;
  assign new_n5238_ = new_n5239_ & new_n8381_;
  assign new_n5239_ = new_n8384_ & new_n8383_;
  assign new_n5240_ = new_n8386_ & new_n8385_ & new_n5472_;
  assign new_n5241_ = new_n5242_ & new_n8389_;
  assign new_n5242_ = new_n8392_ & new_n8391_;
  assign new_n5243_ = new_n8394_ & new_n8393_ & new_n5472_;
  assign new_n5244_ = new_n5245_ & new_n8397_;
  assign new_n5245_ = new_n8400_ & new_n8399_;
  assign new_n5246_ = new_n8402_ & new_n8401_ & new_n5472_;
  assign new_n5247_ = new_n5248_ & new_n8405_;
  assign new_n5248_ = new_n8408_ & new_n8407_;
  assign new_n5249_ = new_n8410_ & new_n8409_ & new_n5472_;
  assign new_n5250_ = new_n5251_ & new_n8413_;
  assign new_n5251_ = new_n8416_ & new_n8415_;
  assign new_n5252_ = new_n8418_ & new_n8417_ & new_n5472_;
  assign new_n5253_ = new_n5254_ & new_n8421_;
  assign new_n5254_ = new_n8424_ & new_n8423_;
  assign new_n5255_ = new_n8426_ & new_n8425_;
  assign new_n5256_ = new_n5257_ & new_n8429_;
  assign new_n5257_ = new_n8432_ & new_n8431_;
  assign new_n5258_ = new_n8434_ & new_n8433_;
  assign new_n5259_ = new_n5260_ & new_n8437_;
  assign new_n5260_ = new_n8440_ & new_n8439_;
  assign new_n5261_ = new_n8442_ & new_n8441_;
  assign new_n5262_ = new_n5263_ & new_n8445_;
  assign new_n5263_ = new_n8448_ & new_n8447_;
  assign new_n5264_ = new_n8450_ & new_n8449_;
  assign new_n5265_ = new_n5266_ & new_n8453_;
  assign new_n5266_ = new_n8456_ & new_n8455_;
  assign new_n5267_ = new_n8458_ & new_n8457_;
  assign new_n5268_ = new_n5269_ & new_n8461_;
  assign new_n5269_ = new_n8464_ & new_n8463_;
  assign new_n5270_ = new_n8466_ & new_n8465_;
  assign new_n5271_ = new_n5272_ & new_n8469_;
  assign new_n5272_ = new_n8472_ & new_n8471_;
  assign new_n5273_ = new_n8474_ & new_n8473_;
  assign new_n5274_ = new_n5275_ & new_n8477_;
  assign new_n5275_ = new_n8480_ & new_n8479_;
  assign new_n5276_ = new_n8482_ & new_n8481_;
  assign new_n5277_ = new_n5278_ & new_n8485_;
  assign new_n5278_ = new_n8488_ & new_n8487_;
  assign new_n5279_ = new_n8490_ & new_n8489_;
  assign new_n5280_ = new_n5281_ & new_n8493_;
  assign new_n5281_ = new_n8496_ & new_n8495_;
  assign new_n5282_ = new_n8498_ & new_n8497_;
  assign new_n5283_ = new_n5284_ & new_n8501_;
  assign new_n5284_ = new_n8504_ & new_n8503_;
  assign new_n5285_ = new_n8506_ & new_n8505_;
  assign new_n5286_ = new_n5287_ & new_n8509_;
  assign new_n5287_ = new_n8512_ & new_n8511_;
  assign new_n5288_ = new_n8520_ & new_n8521_;
  assign new_n5289_ = new_n5288_ & new_n8517_;
  assign new_n5290_ = new_n8518_ & new_n4415_;
  assign new_n5291_ = ~new_n22088_ & ~new_n8519_;
  assign new_n5292_ = ~pi0146 & ~pi0145 & ~pi0148 & ~pi0147;
  assign new_n5293_ = ~pi0150 & ~pi0149 & ~pi0152 & ~pi0151;
  assign new_n5294_ = new_n5293_ & new_n5292_;
  assign new_n5295_ = ~pi0154 & ~pi0153 & ~pi0156 & ~pi0155;
  assign new_n5296_ = ~pi0158 & ~pi0157 & ~pi0160 & ~pi0159;
  assign new_n5297_ = new_n5296_ & new_n5295_;
  assign new_n5298_ = ~pi0162 & ~pi0161 & ~pi0164 & ~pi0163;
  assign new_n5299_ = ~pi0166 & ~pi0165 & ~pi0168 & ~pi0167;
  assign new_n5300_ = new_n5299_ & new_n5298_;
  assign new_n5301_ = ~pi0169 & ~pi0170;
  assign new_n5302_ = ~pi0171 & ~pi0172;
  assign new_n5303_ = ~pi0173 & ~pi0174;
  assign new_n5304_ = new_n8522_ & new_n5301_ & new_n5302_ & new_n5303_;
  assign new_n5305_ = ~pi0143 & ~pi0144 & ~pi0508;
  assign new_n5306_ = new_n8531_ & new_n3786_;
  assign new_n5307_ = new_n8529_ & new_n4291_;
  assign new_n5308_ = new_n8545_ & new_n8543_ & new_n8544_ & new_n8546_;
  assign new_n5309_ = new_n8549_ & new_n8547_ & new_n8548_ & new_n8550_;
  assign new_n5310_ = new_n8553_ & new_n8551_ & new_n8552_ & new_n8554_;
  assign new_n5311_ = new_n8557_ & new_n8555_ & new_n8556_ & new_n8558_;
  assign new_n5312_ = new_n8561_ & new_n8559_ & new_n8560_ & new_n8562_;
  assign new_n5313_ = new_n8565_ & new_n8563_ & new_n8564_ & new_n8566_;
  assign new_n5314_ = new_n8569_ & new_n8567_ & new_n8568_ & new_n8570_;
  assign new_n5315_ = new_n8573_ & new_n8571_ & new_n8572_ & new_n8574_;
  assign new_n5316_ = new_n8577_ & new_n8575_ & new_n8576_ & new_n8578_;
  assign new_n5317_ = new_n8581_ & new_n8579_ & new_n8580_ & new_n8582_;
  assign new_n5318_ = new_n8585_ & new_n8583_ & new_n8584_ & new_n8586_;
  assign new_n5319_ = new_n8589_ & new_n8587_ & new_n8588_ & new_n8590_;
  assign new_n5320_ = new_n8593_ & new_n8591_ & new_n8592_ & new_n8594_;
  assign new_n5321_ = new_n8597_ & new_n8595_ & new_n8596_ & new_n8598_;
  assign new_n5322_ = new_n8601_ & new_n8599_ & new_n8600_ & new_n8602_;
  assign new_n5323_ = new_n8605_ & new_n8603_ & new_n8604_ & new_n8606_;
  assign new_n5324_ = new_n8609_ & new_n8607_ & new_n8608_ & new_n8610_;
  assign new_n5325_ = new_n8613_ & new_n8611_ & new_n8612_ & new_n8614_;
  assign new_n5326_ = new_n8617_ & new_n8615_ & new_n8616_ & new_n8618_;
  assign new_n5327_ = new_n8621_ & new_n8619_ & new_n8620_ & new_n8622_;
  assign new_n5328_ = new_n8625_ & new_n8623_ & new_n8624_ & new_n8626_;
  assign new_n5329_ = new_n8629_ & new_n8627_ & new_n8628_ & new_n8630_;
  assign new_n5330_ = new_n8633_ & new_n8631_ & new_n8632_ & new_n8634_;
  assign new_n5331_ = new_n8637_ & new_n8635_ & new_n8636_ & new_n8638_;
  assign new_n5332_ = new_n8641_ & new_n8639_ & new_n8640_ & new_n8642_;
  assign new_n5333_ = new_n8645_ & new_n8643_ & new_n8644_ & new_n8646_;
  assign new_n5334_ = new_n8649_ & new_n8647_ & new_n8648_ & new_n8650_;
  assign new_n5335_ = new_n8653_ & new_n8651_ & new_n8652_ & new_n8654_;
  assign new_n5336_ = new_n8657_ & new_n8655_ & new_n8656_ & new_n8658_;
  assign new_n5337_ = new_n8661_ & new_n8659_ & new_n8660_ & new_n8662_;
  assign new_n5338_ = new_n8665_ & new_n8663_ & new_n8664_ & new_n8666_;
  assign new_n5339_ = new_n8669_ & new_n8667_ & new_n8668_ & new_n8670_;
  assign new_n5340_ = new_n8675_ & new_n8673_ & new_n8674_ & new_n8676_;
  assign new_n5341_ = new_n8679_ & new_n8677_ & new_n8678_ & new_n8680_;
  assign new_n5342_ = new_n8683_ & new_n8681_ & new_n8682_ & new_n8684_;
  assign new_n5343_ = new_n8687_ & new_n8685_ & new_n8686_ & new_n8688_;
  assign new_n5344_ = new_n8691_ & new_n8689_ & new_n8690_ & new_n8692_;
  assign new_n5345_ = new_n8695_ & new_n8693_ & new_n8694_ & new_n8696_;
  assign new_n5346_ = new_n8699_ & new_n8697_ & new_n8698_ & new_n8700_;
  assign new_n5347_ = new_n8703_ & new_n8701_ & new_n8702_ & new_n8704_;
  assign new_n5348_ = new_n8707_ & new_n8705_ & new_n8706_ & new_n8708_;
  assign new_n5349_ = new_n8711_ & new_n8709_ & new_n8710_ & new_n8712_;
  assign new_n5350_ = new_n8715_ & new_n8713_ & new_n8714_ & new_n8716_;
  assign new_n5351_ = new_n8719_ & new_n8717_ & new_n8718_ & new_n8720_;
  assign new_n5352_ = new_n8723_ & new_n8721_ & new_n8722_ & new_n8724_;
  assign new_n5353_ = new_n8727_ & new_n8725_ & new_n8726_ & new_n8728_;
  assign new_n5354_ = new_n8731_ & new_n8729_ & new_n8730_ & new_n8732_;
  assign new_n5355_ = new_n8735_ & new_n8733_ & new_n8734_ & new_n8736_;
  assign new_n5356_ = new_n8739_ & new_n8737_ & new_n8738_ & new_n8740_;
  assign new_n5357_ = new_n8743_ & new_n8741_ & new_n8742_ & new_n8744_;
  assign new_n5358_ = new_n8747_ & new_n8745_ & new_n8746_ & new_n8748_;
  assign new_n5359_ = new_n8751_ & new_n8749_ & new_n8750_ & new_n8752_;
  assign new_n5360_ = new_n8755_ & new_n8753_ & new_n8754_ & new_n8756_;
  assign new_n5361_ = new_n8759_ & new_n8757_ & new_n8758_ & new_n8760_;
  assign new_n5362_ = new_n8763_ & new_n8761_ & new_n8762_ & new_n8764_;
  assign new_n5363_ = new_n8767_ & new_n8765_ & new_n8766_ & new_n8768_;
  assign new_n5364_ = new_n8771_ & new_n8769_ & new_n8770_ & new_n8772_;
  assign new_n5365_ = new_n8775_ & new_n8773_ & new_n8774_ & new_n8776_;
  assign new_n5366_ = new_n8779_ & new_n8777_ & new_n8778_ & new_n8780_;
  assign new_n5367_ = new_n8783_ & new_n8781_ & new_n8782_ & new_n8784_;
  assign new_n5368_ = new_n8787_ & new_n8785_ & new_n8786_ & new_n8788_;
  assign new_n5369_ = new_n8791_ & new_n8789_ & new_n8790_ & new_n8792_;
  assign new_n5370_ = new_n8795_ & new_n8793_ & new_n8794_ & new_n8796_;
  assign new_n5371_ = new_n8799_ & new_n8797_ & new_n8798_ & new_n8800_;
  assign new_n5372_ = new_n8804_ & new_n8802_ & new_n8803_ & new_n8805_;
  assign new_n5373_ = new_n8808_ & new_n8806_ & new_n8807_ & new_n8809_;
  assign new_n5374_ = new_n8812_ & new_n8810_ & new_n8811_ & new_n8813_;
  assign new_n5375_ = new_n8816_ & new_n8814_ & new_n8815_ & new_n8817_;
  assign new_n5376_ = new_n8820_ & new_n8818_ & new_n8819_ & new_n8821_;
  assign new_n5377_ = new_n8824_ & new_n8822_ & new_n8823_ & new_n8825_;
  assign new_n5378_ = new_n8828_ & new_n8826_ & new_n8827_ & new_n8829_;
  assign new_n5379_ = new_n8832_ & new_n8830_ & new_n8831_ & new_n8833_;
  assign new_n5380_ = new_n8836_ & new_n8834_ & new_n8835_ & new_n8837_;
  assign new_n5381_ = new_n8840_ & new_n8838_ & new_n8839_ & new_n8841_;
  assign new_n5382_ = new_n8844_ & new_n8842_ & new_n8843_ & new_n8845_;
  assign new_n5383_ = new_n8848_ & new_n8846_ & new_n8847_ & new_n8849_;
  assign new_n5384_ = new_n8852_ & new_n8850_ & new_n8851_ & new_n8853_;
  assign new_n5385_ = new_n8856_ & new_n8854_ & new_n8855_ & new_n8857_;
  assign new_n5386_ = new_n8860_ & new_n8858_ & new_n8859_ & new_n8861_;
  assign new_n5387_ = new_n8864_ & new_n8862_ & new_n8863_ & new_n8865_;
  assign new_n5388_ = new_n8868_ & new_n8866_ & new_n8867_ & new_n8869_;
  assign new_n5389_ = new_n8872_ & new_n8870_ & new_n8871_ & new_n8873_;
  assign new_n5390_ = new_n8876_ & new_n8874_ & new_n8875_ & new_n8877_;
  assign new_n5391_ = new_n8880_ & new_n8878_ & new_n8879_ & new_n8881_;
  assign new_n5392_ = new_n8884_ & new_n8882_ & new_n8883_ & new_n8885_;
  assign new_n5393_ = new_n8888_ & new_n8886_ & new_n8887_ & new_n8889_;
  assign new_n5394_ = new_n8892_ & new_n8890_ & new_n8891_ & new_n8893_;
  assign new_n5395_ = new_n8896_ & new_n8894_ & new_n8895_ & new_n8897_;
  assign new_n5396_ = new_n8900_ & new_n8898_ & new_n8899_ & new_n8901_;
  assign new_n5397_ = new_n8904_ & new_n8902_ & new_n8903_ & new_n8905_;
  assign new_n5398_ = new_n8908_ & new_n8906_ & new_n8907_ & new_n8909_;
  assign new_n5399_ = new_n8912_ & new_n8910_ & new_n8911_ & new_n8913_;
  assign new_n5400_ = new_n8916_ & new_n8914_ & new_n8915_ & new_n8917_;
  assign new_n5401_ = new_n8920_ & new_n8918_ & new_n8919_ & new_n8921_;
  assign new_n5402_ = new_n8924_ & new_n8922_ & new_n8923_ & new_n8925_;
  assign new_n5403_ = new_n8928_ & new_n8926_ & new_n8927_ & new_n8929_;
  assign new_n5404_ = new_n8934_ & new_n8932_ & new_n8933_ & new_n8935_;
  assign new_n5405_ = new_n8938_ & new_n8936_ & new_n8937_ & new_n8939_;
  assign new_n5406_ = new_n8942_ & new_n8940_ & new_n8941_ & new_n8943_;
  assign new_n5407_ = new_n8946_ & new_n8944_ & new_n8945_ & new_n8947_;
  assign new_n5408_ = new_n8950_ & new_n8948_ & new_n8949_ & new_n8951_;
  assign new_n5409_ = new_n8954_ & new_n8952_ & new_n8953_ & new_n8955_;
  assign new_n5410_ = new_n8958_ & new_n8956_ & new_n8957_ & new_n8959_;
  assign new_n5411_ = new_n8962_ & new_n8960_ & new_n8961_ & new_n8963_;
  assign new_n5412_ = new_n8966_ & new_n8964_ & new_n8965_ & new_n8967_;
  assign new_n5413_ = new_n8970_ & new_n8968_ & new_n8969_ & new_n8971_;
  assign new_n5414_ = new_n8974_ & new_n8972_ & new_n8973_ & new_n8975_;
  assign new_n5415_ = new_n8978_ & new_n8976_ & new_n8977_ & new_n8979_;
  assign new_n5416_ = new_n8982_ & new_n8980_ & new_n8981_ & new_n8983_;
  assign new_n5417_ = new_n8986_ & new_n8984_ & new_n8985_ & new_n8987_;
  assign new_n5418_ = new_n8990_ & new_n8988_ & new_n8989_ & new_n8991_;
  assign new_n5419_ = new_n8994_ & new_n8992_ & new_n8993_ & new_n8995_;
  assign new_n5420_ = new_n8998_ & new_n8996_ & new_n8997_ & new_n8999_;
  assign new_n5421_ = new_n9002_ & new_n9000_ & new_n9001_ & new_n9003_;
  assign new_n5422_ = new_n9006_ & new_n9004_ & new_n9005_ & new_n9007_;
  assign new_n5423_ = new_n9010_ & new_n9008_ & new_n9009_ & new_n9011_;
  assign new_n5424_ = new_n9014_ & new_n9012_ & new_n9013_ & new_n9015_;
  assign new_n5425_ = new_n9018_ & new_n9016_ & new_n9017_ & new_n9019_;
  assign new_n5426_ = new_n9022_ & new_n9020_ & new_n9021_ & new_n9023_;
  assign new_n5427_ = new_n9026_ & new_n9024_ & new_n9025_ & new_n9027_;
  assign new_n5428_ = new_n9030_ & new_n9028_ & new_n9029_ & new_n9031_;
  assign new_n5429_ = new_n9034_ & new_n9032_ & new_n9033_ & new_n9035_;
  assign new_n5430_ = new_n9038_ & new_n9036_ & new_n9037_ & new_n9039_;
  assign new_n5431_ = new_n9042_ & new_n9040_ & new_n9041_ & new_n9043_;
  assign new_n5432_ = new_n9046_ & new_n9044_ & new_n9045_ & new_n9047_;
  assign new_n5433_ = new_n9050_ & new_n9048_ & new_n9049_ & new_n9051_;
  assign new_n5434_ = new_n9054_ & new_n9052_ & new_n9053_ & new_n9055_;
  assign new_n5435_ = new_n9058_ & new_n9056_ & new_n9057_ & new_n9059_;
  assign new_n5436_ = new_n9099_ & new_n9098_;
  assign new_n5437_ = ~new_n4517_ | ~new_n3760_;
  assign new_n5438_ = new_n9107_ & new_n9106_;
  assign new_n5439_ = ~new_n4814_ | ~new_n6653_;
  assign new_n5440_ = ~pi0348;
  assign new_n5441_ = ~new_n3546_ | ~new_n5437_;
  assign new_n5442_ = ~pi0035;
  assign new_n5443_ = ~new_n5307_ | ~new_n5490_;
  assign new_n5444_ = ~new_n5490_ | ~new_n4395_;
  assign new_n5445_ = ~pi0309 | ~new_n4247_;
  assign new_n5446_ = ~new_n4813_ | ~new_n3671_ | ~new_n3672_;
  assign new_n5447_ = ~new_n4423_;
  assign new_n5448_ = ~pi0033 | ~new_n3786_;
  assign new_n5449_ = ~new_n4261_;
  assign new_n5450_ = ~new_n4262_;
  assign new_n5451_ = ~new_n4291_;
  assign new_n5452_ = ~new_n4268_;
  assign new_n5453_ = ~new_n4267_;
  assign new_n5454_ = ~new_n4398_;
  assign new_n5455_ = ~new_n4399_;
  assign new_n5456_ = ~new_n4400_;
  assign new_n5457_ = ~new_n4401_;
  assign new_n5458_ = ~new_n4275_;
  assign new_n5459_ = ~new_n4273_;
  assign new_n5460_ = ~new_n4272_;
  assign new_n5461_ = ~new_n4271_;
  assign new_n5462_ = ~new_n4402_;
  assign new_n5463_ = ~new_n4417_;
  assign new_n5464_ = ~new_n4233_;
  assign new_n5465_ = ~new_n4409_;
  assign new_n5466_ = ~new_n4408_;
  assign new_n5467_ = ~new_n4406_;
  assign new_n5468_ = ~new_n4283_;
  assign new_n5469_ = ~new_n22894_;
  assign new_n5470_ = ~new_n4373_;
  assign new_n5471_ = ~new_n5451_ | ~new_n3787_;
  assign new_n5472_ = ~new_n5503_ | ~new_n4416_;
  assign new_n5473_ = ~new_n3539_ | ~new_n4261_;
  assign new_n5474_ = ~new_n4403_;
  assign new_n5475_ = ~new_n4415_;
  assign new_n5476_ = ~new_n4236_;
  assign new_n5477_ = ~new_n4234_;
  assign new_n5478_ = ~new_n4292_;
  assign new_n5479_ = ~new_n4270_;
  assign new_n5480_ = ~new_n4274_;
  assign new_n5481_ = ~new_n4375_;
  assign new_n5482_ = ~new_n4337_;
  assign new_n5483_ = ~new_n5305_ | ~new_n5463_;
  assign new_n5484_ = ~new_n4521_ | ~new_n5510_;
  assign new_n5485_ = ~new_n4277_ | ~new_n3787_ | ~new_n4246_ | ~pi0177;
  assign new_n5486_ = ~new_n4809_ | ~new_n3609_;
  assign new_n5487_ = ~new_n3614_ | ~new_n5809_;
  assign new_n5488_ = ~new_n4251_;
  assign new_n5489_ = ~new_n5506_ | ~new_n4269_;
  assign new_n5490_ = ~new_n3546_ | ~new_n8249_;
  assign new_n5491_ = ~new_n5608_ | ~new_n4241_;
  assign new_n5492_ = ~new_n5503_ | ~new_n4277_;
  assign new_n5493_ = ~new_n3609_ | ~new_n4388_;
  assign new_n5494_ = ~new_n2971_ | ~new_n4246_ | ~pi0178;
  assign new_n5495_ = ~new_n4810_ | ~new_n5764_;
  assign new_n5496_ = ~new_n4279_;
  assign new_n5497_ = ~new_n4385_;
  assign new_n5498_ = ~new_n4306_;
  assign new_n5499_ = ~new_n4314_;
  assign new_n5500_ = ~new_n4259_;
  assign new_n5501_ = ~new_n4282_;
  assign new_n5502_ = ~new_n4238_;
  assign new_n5503_ = ~new_n4395_;
  assign new_n5504_ = ~new_n4392_;
  assign new_n5505_ = ~new_n4391_;
  assign new_n5506_ = ~new_n4364_;
  assign new_n5507_ = ~new_n4372_;
  assign new_n5508_ = ~new_n4378_;
  assign new_n5509_ = ~new_n4280_;
  assign new_n5510_ = ~new_n4281_;
  assign new_n5511_ = ~pi0539 | ~new_n5477_;
  assign new_n5512_ = ~pi0538 | ~new_n5476_;
  assign new_n5513_ = ~pi0110 | ~new_n4233_;
  assign new_n5514_ = ~pi0538 | ~new_n5477_;
  assign new_n5515_ = ~pi0537 | ~new_n5476_;
  assign new_n5516_ = ~pi0111 | ~new_n4233_;
  assign new_n5517_ = ~pi0537 | ~new_n5477_;
  assign new_n5518_ = ~pi0536 | ~new_n5476_;
  assign new_n5519_ = ~pi0112 | ~new_n4233_;
  assign new_n5520_ = ~pi0536 | ~new_n5477_;
  assign new_n5521_ = ~pi0535 | ~new_n5476_;
  assign new_n5522_ = ~pi0113 | ~new_n4233_;
  assign new_n5523_ = ~pi0535 | ~new_n5477_;
  assign new_n5524_ = ~pi0534 | ~new_n5476_;
  assign new_n5525_ = ~pi0114 | ~new_n4233_;
  assign new_n5526_ = ~pi0534 | ~new_n5477_;
  assign new_n5527_ = ~pi0533 | ~new_n5476_;
  assign new_n5528_ = ~pi0115 | ~new_n4233_;
  assign new_n5529_ = ~pi0533 | ~new_n5477_;
  assign new_n5530_ = ~pi0532 | ~new_n5476_;
  assign new_n5531_ = ~pi0116 | ~new_n4233_;
  assign new_n5532_ = ~pi0532 | ~new_n5477_;
  assign new_n5533_ = ~pi0531 | ~new_n5476_;
  assign new_n5534_ = ~pi0117 | ~new_n4233_;
  assign new_n5535_ = ~pi0531 | ~new_n5477_;
  assign new_n5536_ = ~pi0530 | ~new_n5476_;
  assign new_n5537_ = ~pi0118 | ~new_n4233_;
  assign new_n5538_ = ~pi0530 | ~new_n5477_;
  assign new_n5539_ = ~pi0529 | ~new_n5476_;
  assign new_n5540_ = ~pi0119 | ~new_n4233_;
  assign new_n5541_ = ~pi0529 | ~new_n5477_;
  assign new_n5542_ = ~pi0528 | ~new_n5476_;
  assign new_n5543_ = ~pi0120 | ~new_n4233_;
  assign new_n5544_ = ~pi0528 | ~new_n5477_;
  assign new_n5545_ = ~pi0527 | ~new_n5476_;
  assign new_n5546_ = ~pi0121 | ~new_n4233_;
  assign new_n5547_ = ~pi0527 | ~new_n5477_;
  assign new_n5548_ = ~pi0526 | ~new_n5476_;
  assign new_n5549_ = ~pi0122 | ~new_n4233_;
  assign new_n5550_ = ~pi0526 | ~new_n5477_;
  assign new_n5551_ = ~pi0525 | ~new_n5476_;
  assign new_n5552_ = ~pi0123 | ~new_n4233_;
  assign new_n5553_ = ~pi0525 | ~new_n5477_;
  assign new_n5554_ = ~pi0524 | ~new_n5476_;
  assign new_n5555_ = ~pi0124 | ~new_n4233_;
  assign new_n5556_ = ~pi0524 | ~new_n5477_;
  assign new_n5557_ = ~pi0523 | ~new_n5476_;
  assign new_n5558_ = ~pi0125 | ~new_n4233_;
  assign new_n5559_ = ~pi0523 | ~new_n5477_;
  assign new_n5560_ = ~pi0522 | ~new_n5476_;
  assign new_n5561_ = ~pi0126 | ~new_n4233_;
  assign new_n5562_ = ~pi0522 | ~new_n5477_;
  assign new_n5563_ = ~pi0521 | ~new_n5476_;
  assign new_n5564_ = ~pi0127 | ~new_n4233_;
  assign new_n5565_ = ~pi0521 | ~new_n5477_;
  assign new_n5566_ = ~pi0520 | ~new_n5476_;
  assign new_n5567_ = ~pi0128 | ~new_n4233_;
  assign new_n5568_ = ~pi0520 | ~new_n5477_;
  assign new_n5569_ = ~pi0519 | ~new_n5476_;
  assign new_n5570_ = ~pi0129 | ~new_n4233_;
  assign new_n5571_ = ~pi0519 | ~new_n5477_;
  assign new_n5572_ = ~pi0518 | ~new_n5476_;
  assign new_n5573_ = ~pi0130 | ~new_n4233_;
  assign new_n5574_ = ~pi0518 | ~new_n5477_;
  assign new_n5575_ = ~pi0517 | ~new_n5476_;
  assign new_n5576_ = ~pi0131 | ~new_n4233_;
  assign new_n5577_ = ~pi0517 | ~new_n5477_;
  assign new_n5578_ = ~pi0516 | ~new_n5476_;
  assign new_n5579_ = ~pi0132 | ~new_n4233_;
  assign new_n5580_ = ~pi0516 | ~new_n5477_;
  assign new_n5581_ = ~pi0515 | ~new_n5476_;
  assign new_n5582_ = ~pi0133 | ~new_n4233_;
  assign new_n5583_ = ~pi0515 | ~new_n5477_;
  assign new_n5584_ = ~pi0514 | ~new_n5476_;
  assign new_n5585_ = ~pi0134 | ~new_n4233_;
  assign new_n5586_ = ~pi0514 | ~new_n5477_;
  assign new_n5587_ = ~pi0513 | ~new_n5476_;
  assign new_n5588_ = ~pi0135 | ~new_n4233_;
  assign new_n5589_ = ~pi0513 | ~new_n5477_;
  assign new_n5590_ = ~pi0512 | ~new_n5476_;
  assign new_n5591_ = ~pi0136 | ~new_n4233_;
  assign new_n5592_ = ~pi0512 | ~new_n5477_;
  assign new_n5593_ = ~pi0511 | ~new_n5476_;
  assign new_n5594_ = ~pi0137 | ~new_n4233_;
  assign new_n5595_ = ~pi0511 | ~new_n5477_;
  assign new_n5596_ = ~pi0510 | ~new_n5476_;
  assign new_n5597_ = ~pi0138 | ~new_n4233_;
  assign new_n5598_ = ~pi0510 | ~new_n5477_;
  assign new_n5599_ = ~pi0509 | ~new_n5476_;
  assign new_n5600_ = ~pi0139 | ~new_n4233_;
  assign new_n5601_ = ~new_n4243_;
  assign new_n5602_ = ~new_n5601_ | ~new_n3786_;
  assign new_n5603_ = ~pi0034 | ~new_n5502_;
  assign new_n5604_ = ~new_n4244_;
  assign new_n5605_ = ~new_n5604_ | ~new_n3786_;
  assign new_n5606_ = pi0142 | pi0034;
  assign new_n5607_ = ~new_n9069_ | ~new_n9068_ | ~new_n5606_;
  assign new_n5608_ = ~new_n4239_;
  assign new_n5609_ = ~new_n5502_ | ~new_n4244_ | ~new_n2971_;
  assign new_n5610_ = ~new_n5608_ | ~pi0033 | ~new_n4231_;
  assign new_n5611_ = ~new_n5609_ | ~new_n5610_;
  assign new_n5612_ = ~new_n4465_ | ~new_n5611_;
  assign new_n5613_ = ~pi0140 | ~new_n5607_;
  assign new_n5614_ = ~new_n5464_ | ~new_n2971_;
  assign new_n5615_ = ~new_n4468_ | ~new_n9071_;
  assign new_n5616_ = ~pi0140 | ~new_n4243_;
  assign new_n5617_ = ~pi0034 | ~new_n4241_;
  assign new_n5618_ = ~new_n5617_ | ~new_n5616_;
  assign new_n5619_ = ~new_n5618_ | ~new_n4232_;
  assign new_n5620_ = ~new_n5442_ | ~new_n4239_;
  assign new_n5621_ = ~pi0140 | ~new_n4232_;
  assign new_n5622_ = ~new_n4238_ | ~new_n5621_;
  assign new_n5623_ = ~new_n4247_;
  assign new_n5624_ = ~new_n4252_;
  assign new_n5625_ = ~new_n4248_;
  assign new_n5626_ = ~new_n4254_;
  assign new_n5627_ = ~new_n4255_;
  assign new_n5628_ = ~pi0306 | ~new_n3640_;
  assign new_n5629_ = ~pi0298 | ~new_n3639_;
  assign new_n5630_ = ~pi0290 | ~new_n3638_;
  assign new_n5631_ = ~pi0282 | ~new_n3636_;
  assign new_n5632_ = ~pi0274 | ~new_n3635_;
  assign new_n5633_ = ~pi0266 | ~new_n3634_;
  assign new_n5634_ = ~pi0258 | ~new_n3633_;
  assign new_n5635_ = ~pi0250 | ~new_n5627_;
  assign new_n5636_ = ~pi0242 | ~new_n3632_;
  assign new_n5637_ = ~pi0234 | ~new_n3631_;
  assign new_n5638_ = ~pi0226 | ~new_n3629_;
  assign new_n5639_ = ~pi0218 | ~new_n3627_;
  assign new_n5640_ = ~pi0210 | ~new_n3626_;
  assign new_n5641_ = ~pi0202 | ~new_n3625_;
  assign new_n5642_ = ~pi0194 | ~new_n3623_;
  assign new_n5643_ = ~pi0186 | ~new_n3621_;
  assign new_n5644_ = ~new_n4264_;
  assign new_n5645_ = ~pi0305 | ~new_n3640_;
  assign new_n5646_ = ~pi0297 | ~new_n3639_;
  assign new_n5647_ = ~pi0289 | ~new_n3638_;
  assign new_n5648_ = ~pi0281 | ~new_n3636_;
  assign new_n5649_ = ~pi0273 | ~new_n3635_;
  assign new_n5650_ = ~pi0265 | ~new_n3634_;
  assign new_n5651_ = ~pi0257 | ~new_n3633_;
  assign new_n5652_ = ~pi0249 | ~new_n5627_;
  assign new_n5653_ = ~pi0241 | ~new_n3632_;
  assign new_n5654_ = ~pi0233 | ~new_n3631_;
  assign new_n5655_ = ~pi0225 | ~new_n3629_;
  assign new_n5656_ = ~pi0217 | ~new_n3627_;
  assign new_n5657_ = ~pi0209 | ~new_n3626_;
  assign new_n5658_ = ~pi0201 | ~new_n3625_;
  assign new_n5659_ = ~pi0193 | ~new_n3623_;
  assign new_n5660_ = ~pi0185 | ~new_n3621_;
  assign new_n5661_ = ~new_n4260_;
  assign new_n5662_ = ~pi0302 | ~new_n3640_;
  assign new_n5663_ = ~pi0294 | ~new_n3639_;
  assign new_n5664_ = ~pi0286 | ~new_n3638_;
  assign new_n5665_ = ~pi0278 | ~new_n3636_;
  assign new_n5666_ = ~pi0270 | ~new_n3635_;
  assign new_n5667_ = ~pi0262 | ~new_n3634_;
  assign new_n5668_ = ~pi0254 | ~new_n3633_;
  assign new_n5669_ = ~pi0246 | ~new_n5627_;
  assign new_n5670_ = ~pi0238 | ~new_n3632_;
  assign new_n5671_ = ~pi0230 | ~new_n3631_;
  assign new_n5672_ = ~pi0222 | ~new_n3629_;
  assign new_n5673_ = ~pi0214 | ~new_n3627_;
  assign new_n5674_ = ~pi0206 | ~new_n3626_;
  assign new_n5675_ = ~pi0198 | ~new_n3625_;
  assign new_n5676_ = ~pi0190 | ~new_n3623_;
  assign new_n5677_ = ~pi0182 | ~new_n3621_;
  assign new_n5678_ = ~new_n4258_;
  assign new_n5679_ = ~pi0304 | ~new_n3640_;
  assign new_n5680_ = ~pi0296 | ~new_n3639_;
  assign new_n5681_ = ~pi0288 | ~new_n3638_;
  assign new_n5682_ = ~pi0280 | ~new_n3636_;
  assign new_n5683_ = ~pi0272 | ~new_n3635_;
  assign new_n5684_ = ~pi0264 | ~new_n3634_;
  assign new_n5685_ = ~pi0256 | ~new_n3633_;
  assign new_n5686_ = ~pi0248 | ~new_n5627_;
  assign new_n5687_ = ~pi0240 | ~new_n3632_;
  assign new_n5688_ = ~pi0232 | ~new_n3631_;
  assign new_n5689_ = ~pi0224 | ~new_n3629_;
  assign new_n5690_ = ~pi0216 | ~new_n3627_;
  assign new_n5691_ = ~pi0208 | ~new_n3626_;
  assign new_n5692_ = ~pi0200 | ~new_n3625_;
  assign new_n5693_ = ~pi0192 | ~new_n3623_;
  assign new_n5694_ = ~pi0184 | ~new_n3621_;
  assign new_n5695_ = ~new_n4257_;
  assign new_n5696_ = ~pi0303 | ~new_n3640_;
  assign new_n5697_ = ~pi0295 | ~new_n3639_;
  assign new_n5698_ = ~pi0287 | ~new_n3638_;
  assign new_n5699_ = ~pi0279 | ~new_n3636_;
  assign new_n5700_ = ~pi0271 | ~new_n3635_;
  assign new_n5701_ = ~pi0263 | ~new_n3634_;
  assign new_n5702_ = ~pi0255 | ~new_n3633_;
  assign new_n5703_ = ~pi0247 | ~new_n5627_;
  assign new_n5704_ = ~pi0239 | ~new_n3632_;
  assign new_n5705_ = ~pi0231 | ~new_n3631_;
  assign new_n5706_ = ~pi0223 | ~new_n3629_;
  assign new_n5707_ = ~pi0215 | ~new_n3627_;
  assign new_n5708_ = ~pi0207 | ~new_n3626_;
  assign new_n5709_ = ~pi0199 | ~new_n3625_;
  assign new_n5710_ = ~pi0191 | ~new_n3623_;
  assign new_n5711_ = ~pi0183 | ~new_n3621_;
  assign new_n5712_ = ~new_n4263_;
  assign new_n5713_ = ~pi0299 | ~new_n3640_;
  assign new_n5714_ = ~pi0291 | ~new_n3639_;
  assign new_n5715_ = ~pi0283 | ~new_n3638_;
  assign new_n5716_ = ~pi0275 | ~new_n3636_;
  assign new_n5717_ = ~pi0267 | ~new_n3635_;
  assign new_n5718_ = ~pi0259 | ~new_n3634_;
  assign new_n5719_ = ~pi0251 | ~new_n3633_;
  assign new_n5720_ = ~pi0243 | ~new_n5627_;
  assign new_n5721_ = ~pi0235 | ~new_n3632_;
  assign new_n5722_ = ~pi0227 | ~new_n3631_;
  assign new_n5723_ = ~pi0219 | ~new_n3629_;
  assign new_n5724_ = ~pi0211 | ~new_n3627_;
  assign new_n5725_ = ~pi0203 | ~new_n3626_;
  assign new_n5726_ = ~pi0195 | ~new_n3625_;
  assign new_n5727_ = ~pi0187 | ~new_n3623_;
  assign new_n5728_ = ~pi0179 | ~new_n3621_;
  assign new_n5729_ = ~new_n4374_;
  assign new_n5730_ = ~pi0301 | ~new_n3640_;
  assign new_n5731_ = ~pi0293 | ~new_n3639_;
  assign new_n5732_ = ~pi0285 | ~new_n3638_;
  assign new_n5733_ = ~pi0277 | ~new_n3636_;
  assign new_n5734_ = ~pi0269 | ~new_n3635_;
  assign new_n5735_ = ~pi0261 | ~new_n3634_;
  assign new_n5736_ = ~pi0253 | ~new_n3633_;
  assign new_n5737_ = ~pi0245 | ~new_n5627_;
  assign new_n5738_ = ~pi0237 | ~new_n3632_;
  assign new_n5739_ = ~pi0229 | ~new_n3631_;
  assign new_n5740_ = ~pi0221 | ~new_n3629_;
  assign new_n5741_ = ~pi0213 | ~new_n3627_;
  assign new_n5742_ = ~pi0205 | ~new_n3626_;
  assign new_n5743_ = ~pi0197 | ~new_n3625_;
  assign new_n5744_ = ~pi0189 | ~new_n3623_;
  assign new_n5745_ = ~pi0181 | ~new_n3621_;
  assign new_n5746_ = ~new_n4266_;
  assign new_n5747_ = ~pi0300 | ~new_n3640_;
  assign new_n5748_ = ~pi0292 | ~new_n3639_;
  assign new_n5749_ = ~pi0284 | ~new_n3638_;
  assign new_n5750_ = ~pi0276 | ~new_n3636_;
  assign new_n5751_ = ~pi0268 | ~new_n3635_;
  assign new_n5752_ = ~pi0260 | ~new_n3634_;
  assign new_n5753_ = ~pi0252 | ~new_n3633_;
  assign new_n5754_ = ~pi0244 | ~new_n5627_;
  assign new_n5755_ = ~pi0236 | ~new_n3632_;
  assign new_n5756_ = ~pi0228 | ~new_n3631_;
  assign new_n5757_ = ~pi0220 | ~new_n3629_;
  assign new_n5758_ = ~pi0212 | ~new_n3627_;
  assign new_n5759_ = ~pi0204 | ~new_n3626_;
  assign new_n5760_ = ~pi0196 | ~new_n3625_;
  assign new_n5761_ = ~pi0188 | ~new_n3623_;
  assign new_n5762_ = ~pi0180 | ~new_n3621_;
  assign new_n5763_ = ~new_n4230_;
  assign new_n5764_ = ~new_n4269_;
  assign new_n5765_ = ~new_n3517_ | ~new_n4394_;
  assign new_n5766_ = ~new_n3516_ | ~new_n4393_;
  assign new_n5767_ = ~new_n3513_ | ~new_n4368_;
  assign new_n5768_ = ~new_n5461_ | ~new_n4371_;
  assign new_n5769_ = ~new_n5460_ | ~new_n4366_;
  assign new_n5770_ = ~new_n5459_ | ~new_n4369_;
  assign new_n5771_ = ~new_n3512_ | ~new_n4367_;
  assign new_n5772_ = ~new_n5458_ | ~new_n4370_;
  assign new_n5773_ = ~new_n4514_ | ~new_n4513_;
  assign new_n5774_ = ~new_n3619_ | ~new_n9100_ | ~new_n9101_ | ~new_n4516_ | ~new_n5678_;
  assign new_n5775_ = ~new_n4265_;
  assign new_n5776_ = ~new_n5436_ | ~new_n5775_;
  assign new_n5777_ = ~new_n4515_ | ~new_n9072_;
  assign new_n5778_ = ~new_n5437_;
  assign new_n5779_ = ~new_n4418_;
  assign new_n5780_ = pi0546 | pi0545;
  assign new_n5781_ = ~new_n4276_;
  assign new_n5782_ = ~new_n4509_ | ~new_n5459_;
  assign new_n5783_ = ~new_n4518_ | ~new_n5781_;
  assign new_n5784_ = ~pi0177 | ~new_n2971_;
  assign new_n5785_ = ~pi0176 | ~new_n9109_ | ~new_n9108_;
  assign new_n5786_ = ~new_n4278_;
  assign new_n5787_ = ~pi0177 | ~new_n9113_ | ~new_n9112_;
  assign new_n5788_ = ~pi0176 | ~new_n4278_;
  assign new_n5789_ = ~new_n5785_ | ~new_n5494_;
  assign new_n5790_ = ~new_n4520_ | ~new_n5786_;
  assign new_n5791_ = ~pi0177 | ~new_n5789_;
  assign new_n5792_ = ~new_n3546_ | ~new_n5785_;
  assign new_n5793_ = ~new_n5501_ | ~new_n5510_;
  assign new_n5794_ = ~new_n5785_ | ~new_n5493_;
  assign new_n5795_ = ~new_n3546_ | ~new_n4276_;
  assign new_n5796_ = ~new_n4309_;
  assign new_n5797_ = ~pi0315 | ~new_n4284_;
  assign new_n5798_ = ~new_n4293_;
  assign new_n5799_ = ~new_n4297_;
  assign new_n5800_ = ~new_n4304_;
  assign new_n5801_ = ~new_n4311_;
  assign new_n5802_ = ~new_n4312_;
  assign new_n5803_ = ~new_n4299_;
  assign new_n5804_ = ~new_n4286_;
  assign new_n5805_ = ~new_n4288_;
  assign new_n5806_ = ~new_n4336_;
  assign new_n5807_ = ~pi0313 | ~new_n4288_;
  assign new_n5808_ = ~new_n4295_;
  assign new_n5809_ = ~new_n4294_;
  assign new_n5810_ = ~new_n5809_ | ~new_n4425_;
  assign new_n5811_ = ~new_n5810_ | ~new_n4295_;
  assign new_n5812_ = ~new_n4298_;
  assign new_n5813_ = ~new_n4296_;
  assign new_n5814_ = ~new_n4321_;
  assign new_n5815_ = ~new_n4296_ | ~new_n4298_;
  assign new_n5816_ = ~new_n4338_;
  assign new_n5817_ = ~new_n4300_;
  assign new_n5818_ = ~new_n4290_;
  assign new_n5819_ = ~new_n3613_ | ~new_n5809_;
  assign new_n5820_ = ~new_n4302_;
  assign new_n5821_ = ~pi0177 | ~new_n4246_;
  assign new_n5822_ = ~new_n4282_ | ~new_n4280_ | ~new_n5821_;
  assign new_n5823_ = ~new_n5813_ | ~new_n3643_;
  assign new_n5824_ = ~new_n4301_;
  assign new_n5825_ = ~new_n3645_ | ~new_n4301_;
  assign new_n5826_ = ~new_n5820_ | ~new_n5825_;
  assign new_n5827_ = ~pi0175 | ~new_n4290_;
  assign new_n5828_ = ~new_n4525_ | ~new_n5826_;
  assign new_n5829_ = ~new_n5824_ | ~new_n5478_;
  assign new_n5830_ = ~new_n3645_ | ~new_n5829_;
  assign new_n5831_ = ~new_n3601_ | ~new_n5818_;
  assign new_n5832_ = ~new_n3592_ | ~new_n3644_;
  assign new_n5833_ = ~new_n3591_ | ~new_n5817_;
  assign new_n5834_ = ~new_n3534_ | ~new_n3576_;
  assign new_n5835_ = ~pi0179 | ~new_n5828_;
  assign new_n5836_ = ~new_n3599_ | ~new_n5818_;
  assign new_n5837_ = ~new_n3590_ | ~new_n3644_;
  assign new_n5838_ = ~new_n3589_ | ~new_n5817_;
  assign new_n5839_ = ~new_n3575_ | ~new_n3534_;
  assign new_n5840_ = ~pi0180 | ~new_n5828_;
  assign new_n5841_ = ~new_n3598_ | ~new_n5818_;
  assign new_n5842_ = ~new_n3588_ | ~new_n3644_;
  assign new_n5843_ = ~new_n3587_ | ~new_n5817_;
  assign new_n5844_ = ~new_n3574_ | ~new_n3534_;
  assign new_n5845_ = ~pi0181 | ~new_n5828_;
  assign new_n5846_ = ~new_n3597_ | ~new_n5818_;
  assign new_n5847_ = ~new_n3586_ | ~new_n3644_;
  assign new_n5848_ = ~new_n3585_ | ~new_n5817_;
  assign new_n5849_ = ~new_n3573_ | ~new_n3534_;
  assign new_n5850_ = ~pi0182 | ~new_n5828_;
  assign new_n5851_ = ~new_n3596_ | ~new_n5818_;
  assign new_n5852_ = ~new_n3584_ | ~new_n3644_;
  assign new_n5853_ = ~new_n3583_ | ~new_n5817_;
  assign new_n5854_ = ~new_n3572_ | ~new_n3534_;
  assign new_n5855_ = ~pi0183 | ~new_n5828_;
  assign new_n5856_ = ~new_n3595_ | ~new_n5818_;
  assign new_n5857_ = ~new_n3582_ | ~new_n3644_;
  assign new_n5858_ = ~new_n3581_ | ~new_n5817_;
  assign new_n5859_ = ~new_n3571_ | ~new_n3534_;
  assign new_n5860_ = ~pi0184 | ~new_n5828_;
  assign new_n5861_ = ~new_n3594_ | ~new_n5818_;
  assign new_n5862_ = ~new_n3580_ | ~new_n3644_;
  assign new_n5863_ = ~new_n3579_ | ~new_n5817_;
  assign new_n5864_ = ~new_n3570_ | ~new_n3534_;
  assign new_n5865_ = ~pi0185 | ~new_n5828_;
  assign new_n5866_ = ~new_n3593_ | ~new_n5818_;
  assign new_n5867_ = ~new_n3578_ | ~new_n3644_;
  assign new_n5868_ = ~new_n3577_ | ~new_n5817_;
  assign new_n5869_ = ~new_n3569_ | ~new_n3534_;
  assign new_n5870_ = ~pi0186 | ~new_n5828_;
  assign new_n5871_ = ~new_n4305_;
  assign new_n5872_ = ~new_n4303_;
  assign new_n5873_ = ~new_n5498_ | ~new_n3613_;
  assign new_n5874_ = ~new_n4308_;
  assign new_n5875_ = ~new_n5800_ | ~new_n3643_;
  assign new_n5876_ = ~new_n4307_;
  assign new_n5877_ = ~new_n3645_ | ~new_n4307_;
  assign new_n5878_ = ~new_n5874_ | ~new_n5877_;
  assign new_n5879_ = ~pi0175 | ~new_n4303_;
  assign new_n5880_ = ~new_n4543_ | ~new_n5878_;
  assign new_n5881_ = ~new_n5876_ | ~new_n5478_;
  assign new_n5882_ = ~new_n3645_ | ~new_n5881_;
  assign new_n5883_ = ~new_n5872_ | ~new_n3601_;
  assign new_n5884_ = ~new_n3647_ | ~new_n3592_;
  assign new_n5885_ = ~new_n5871_ | ~new_n3591_;
  assign new_n5886_ = ~new_n3533_ | ~new_n3576_;
  assign new_n5887_ = ~pi0187 | ~new_n5880_;
  assign new_n5888_ = ~new_n5872_ | ~new_n3599_;
  assign new_n5889_ = ~new_n3647_ | ~new_n3590_;
  assign new_n5890_ = ~new_n5871_ | ~new_n3589_;
  assign new_n5891_ = ~new_n3533_ | ~new_n3575_;
  assign new_n5892_ = ~pi0188 | ~new_n5880_;
  assign new_n5893_ = ~new_n5872_ | ~new_n3598_;
  assign new_n5894_ = ~new_n3647_ | ~new_n3588_;
  assign new_n5895_ = ~new_n5871_ | ~new_n3587_;
  assign new_n5896_ = ~new_n3533_ | ~new_n3574_;
  assign new_n5897_ = ~pi0189 | ~new_n5880_;
  assign new_n5898_ = ~new_n5872_ | ~new_n3597_;
  assign new_n5899_ = ~new_n3647_ | ~new_n3586_;
  assign new_n5900_ = ~new_n5871_ | ~new_n3585_;
  assign new_n5901_ = ~new_n3533_ | ~new_n3573_;
  assign new_n5902_ = ~pi0190 | ~new_n5880_;
  assign new_n5903_ = ~new_n5872_ | ~new_n3596_;
  assign new_n5904_ = ~new_n3647_ | ~new_n3584_;
  assign new_n5905_ = ~new_n5871_ | ~new_n3583_;
  assign new_n5906_ = ~new_n3533_ | ~new_n3572_;
  assign new_n5907_ = ~pi0191 | ~new_n5880_;
  assign new_n5908_ = ~new_n5872_ | ~new_n3595_;
  assign new_n5909_ = ~new_n3647_ | ~new_n3582_;
  assign new_n5910_ = ~new_n5871_ | ~new_n3581_;
  assign new_n5911_ = ~new_n3533_ | ~new_n3571_;
  assign new_n5912_ = ~pi0192 | ~new_n5880_;
  assign new_n5913_ = ~new_n5872_ | ~new_n3594_;
  assign new_n5914_ = ~new_n3647_ | ~new_n3580_;
  assign new_n5915_ = ~new_n5871_ | ~new_n3579_;
  assign new_n5916_ = ~new_n3533_ | ~new_n3570_;
  assign new_n5917_ = ~pi0193 | ~new_n5880_;
  assign new_n5918_ = ~new_n5872_ | ~new_n3593_;
  assign new_n5919_ = ~new_n3647_ | ~new_n3578_;
  assign new_n5920_ = ~new_n5871_ | ~new_n3577_;
  assign new_n5921_ = ~new_n3533_ | ~new_n3569_;
  assign new_n5922_ = ~pi0194 | ~new_n5880_;
  assign new_n5923_ = ~new_n4313_;
  assign new_n5924_ = ~new_n4310_;
  assign new_n5925_ = ~new_n5499_ | ~new_n3613_;
  assign new_n5926_ = ~new_n4316_;
  assign new_n5927_ = ~new_n5801_ | ~new_n3643_;
  assign new_n5928_ = ~new_n4315_;
  assign new_n5929_ = ~new_n3645_ | ~new_n4315_;
  assign new_n5930_ = ~new_n5926_ | ~new_n5929_;
  assign new_n5931_ = ~pi0175 | ~new_n4310_;
  assign new_n5932_ = ~new_n4561_ | ~new_n5930_;
  assign new_n5933_ = ~new_n5928_ | ~new_n5478_;
  assign new_n5934_ = ~new_n3645_ | ~new_n5933_;
  assign new_n5935_ = ~new_n5924_ | ~new_n3601_;
  assign new_n5936_ = ~new_n3650_ | ~new_n3592_;
  assign new_n5937_ = ~new_n5923_ | ~new_n3591_;
  assign new_n5938_ = ~new_n3532_ | ~new_n3576_;
  assign new_n5939_ = ~pi0195 | ~new_n5932_;
  assign new_n5940_ = ~new_n5924_ | ~new_n3599_;
  assign new_n5941_ = ~new_n3650_ | ~new_n3590_;
  assign new_n5942_ = ~new_n5923_ | ~new_n3589_;
  assign new_n5943_ = ~new_n3532_ | ~new_n3575_;
  assign new_n5944_ = ~pi0196 | ~new_n5932_;
  assign new_n5945_ = ~new_n5924_ | ~new_n3598_;
  assign new_n5946_ = ~new_n3650_ | ~new_n3588_;
  assign new_n5947_ = ~new_n5923_ | ~new_n3587_;
  assign new_n5948_ = ~new_n3532_ | ~new_n3574_;
  assign new_n5949_ = ~pi0197 | ~new_n5932_;
  assign new_n5950_ = ~new_n5924_ | ~new_n3597_;
  assign new_n5951_ = ~new_n3650_ | ~new_n3586_;
  assign new_n5952_ = ~new_n5923_ | ~new_n3585_;
  assign new_n5953_ = ~new_n3532_ | ~new_n3573_;
  assign new_n5954_ = ~pi0198 | ~new_n5932_;
  assign new_n5955_ = ~new_n5924_ | ~new_n3596_;
  assign new_n5956_ = ~new_n3650_ | ~new_n3584_;
  assign new_n5957_ = ~new_n5923_ | ~new_n3583_;
  assign new_n5958_ = ~new_n3532_ | ~new_n3572_;
  assign new_n5959_ = ~pi0199 | ~new_n5932_;
  assign new_n5960_ = ~new_n5924_ | ~new_n3595_;
  assign new_n5961_ = ~new_n3650_ | ~new_n3582_;
  assign new_n5962_ = ~new_n5923_ | ~new_n3581_;
  assign new_n5963_ = ~new_n3532_ | ~new_n3571_;
  assign new_n5964_ = ~pi0200 | ~new_n5932_;
  assign new_n5965_ = ~new_n5924_ | ~new_n3594_;
  assign new_n5966_ = ~new_n3650_ | ~new_n3580_;
  assign new_n5967_ = ~new_n5923_ | ~new_n3579_;
  assign new_n5968_ = ~new_n3532_ | ~new_n3570_;
  assign new_n5969_ = ~pi0201 | ~new_n5932_;
  assign new_n5970_ = ~new_n5924_ | ~new_n3593_;
  assign new_n5971_ = ~new_n3650_ | ~new_n3578_;
  assign new_n5972_ = ~new_n5923_ | ~new_n3577_;
  assign new_n5973_ = ~new_n3532_ | ~new_n3569_;
  assign new_n5974_ = ~pi0202 | ~new_n5932_;
  assign new_n5975_ = ~new_n4318_;
  assign new_n5976_ = ~new_n4317_;
  assign new_n5977_ = ~new_n4226_;
  assign new_n5978_ = ~new_n3652_ | ~new_n3643_;
  assign new_n5979_ = ~new_n4319_;
  assign new_n5980_ = ~new_n3645_ | ~new_n4319_;
  assign new_n5981_ = ~new_n5980_ | ~new_n4226_;
  assign new_n5982_ = ~pi0175 | ~new_n4317_;
  assign new_n5983_ = ~new_n4579_ | ~new_n5981_;
  assign new_n5984_ = ~new_n5979_ | ~new_n5478_;
  assign new_n5985_ = ~new_n3645_ | ~new_n5984_;
  assign new_n5986_ = ~new_n5976_ | ~new_n3601_;
  assign new_n5987_ = ~new_n3653_ | ~new_n3592_;
  assign new_n5988_ = ~new_n5975_ | ~new_n3591_;
  assign new_n5989_ = ~new_n3531_ | ~new_n3576_;
  assign new_n5990_ = ~pi0203 | ~new_n5983_;
  assign new_n5991_ = ~new_n5976_ | ~new_n3599_;
  assign new_n5992_ = ~new_n3653_ | ~new_n3590_;
  assign new_n5993_ = ~new_n5975_ | ~new_n3589_;
  assign new_n5994_ = ~new_n3531_ | ~new_n3575_;
  assign new_n5995_ = ~pi0204 | ~new_n5983_;
  assign new_n5996_ = ~new_n5976_ | ~new_n3598_;
  assign new_n5997_ = ~new_n3653_ | ~new_n3588_;
  assign new_n5998_ = ~new_n5975_ | ~new_n3587_;
  assign new_n5999_ = ~new_n3531_ | ~new_n3574_;
  assign new_n6000_ = ~pi0205 | ~new_n5983_;
  assign new_n6001_ = ~new_n5976_ | ~new_n3597_;
  assign new_n6002_ = ~new_n3653_ | ~new_n3586_;
  assign new_n6003_ = ~new_n5975_ | ~new_n3585_;
  assign new_n6004_ = ~new_n3531_ | ~new_n3573_;
  assign new_n6005_ = ~pi0206 | ~new_n5983_;
  assign new_n6006_ = ~new_n5976_ | ~new_n3596_;
  assign new_n6007_ = ~new_n3653_ | ~new_n3584_;
  assign new_n6008_ = ~new_n5975_ | ~new_n3583_;
  assign new_n6009_ = ~new_n3531_ | ~new_n3572_;
  assign new_n6010_ = ~pi0207 | ~new_n5983_;
  assign new_n6011_ = ~new_n5976_ | ~new_n3595_;
  assign new_n6012_ = ~new_n3653_ | ~new_n3582_;
  assign new_n6013_ = ~new_n5975_ | ~new_n3581_;
  assign new_n6014_ = ~new_n3531_ | ~new_n3571_;
  assign new_n6015_ = ~pi0208 | ~new_n5983_;
  assign new_n6016_ = ~new_n5976_ | ~new_n3594_;
  assign new_n6017_ = ~new_n3653_ | ~new_n3580_;
  assign new_n6018_ = ~new_n5975_ | ~new_n3579_;
  assign new_n6019_ = ~new_n3531_ | ~new_n3570_;
  assign new_n6020_ = ~pi0209 | ~new_n5983_;
  assign new_n6021_ = ~new_n5976_ | ~new_n3593_;
  assign new_n6022_ = ~new_n3653_ | ~new_n3578_;
  assign new_n6023_ = ~new_n5975_ | ~new_n3577_;
  assign new_n6024_ = ~new_n3531_ | ~new_n3569_;
  assign new_n6025_ = ~pi0210 | ~new_n5983_;
  assign new_n6026_ = ~new_n4322_;
  assign new_n6027_ = ~new_n4320_;
  assign new_n6028_ = ~new_n3615_ | ~new_n5809_;
  assign new_n6029_ = ~new_n4324_;
  assign new_n6030_ = ~new_n5814_ | ~new_n5813_;
  assign new_n6031_ = ~new_n4323_;
  assign new_n6032_ = ~new_n3645_ | ~new_n4323_;
  assign new_n6033_ = ~new_n6029_ | ~new_n6032_;
  assign new_n6034_ = ~pi0175 | ~new_n4320_;
  assign new_n6035_ = ~new_n4596_ | ~new_n6033_;
  assign new_n6036_ = ~new_n6031_ | ~new_n5478_;
  assign new_n6037_ = ~new_n3645_ | ~new_n6036_;
  assign new_n6038_ = ~new_n6027_ | ~new_n3601_;
  assign new_n6039_ = ~new_n3655_ | ~new_n3592_;
  assign new_n6040_ = ~new_n6026_ | ~new_n3591_;
  assign new_n6041_ = ~new_n3530_ | ~new_n3576_;
  assign new_n6042_ = ~pi0211 | ~new_n6035_;
  assign new_n6043_ = ~new_n6027_ | ~new_n3599_;
  assign new_n6044_ = ~new_n3655_ | ~new_n3590_;
  assign new_n6045_ = ~new_n6026_ | ~new_n3589_;
  assign new_n6046_ = ~new_n3530_ | ~new_n3575_;
  assign new_n6047_ = ~pi0212 | ~new_n6035_;
  assign new_n6048_ = ~new_n6027_ | ~new_n3598_;
  assign new_n6049_ = ~new_n3655_ | ~new_n3588_;
  assign new_n6050_ = ~new_n6026_ | ~new_n3587_;
  assign new_n6051_ = ~new_n3530_ | ~new_n3574_;
  assign new_n6052_ = ~pi0213 | ~new_n6035_;
  assign new_n6053_ = ~new_n6027_ | ~new_n3597_;
  assign new_n6054_ = ~new_n3655_ | ~new_n3586_;
  assign new_n6055_ = ~new_n6026_ | ~new_n3585_;
  assign new_n6056_ = ~new_n3530_ | ~new_n3573_;
  assign new_n6057_ = ~pi0214 | ~new_n6035_;
  assign new_n6058_ = ~new_n6027_ | ~new_n3596_;
  assign new_n6059_ = ~new_n3655_ | ~new_n3584_;
  assign new_n6060_ = ~new_n6026_ | ~new_n3583_;
  assign new_n6061_ = ~new_n3530_ | ~new_n3572_;
  assign new_n6062_ = ~pi0215 | ~new_n6035_;
  assign new_n6063_ = ~new_n6027_ | ~new_n3595_;
  assign new_n6064_ = ~new_n3655_ | ~new_n3582_;
  assign new_n6065_ = ~new_n6026_ | ~new_n3581_;
  assign new_n6066_ = ~new_n3530_ | ~new_n3571_;
  assign new_n6067_ = ~pi0216 | ~new_n6035_;
  assign new_n6068_ = ~new_n6027_ | ~new_n3594_;
  assign new_n6069_ = ~new_n3655_ | ~new_n3580_;
  assign new_n6070_ = ~new_n6026_ | ~new_n3579_;
  assign new_n6071_ = ~new_n3530_ | ~new_n3570_;
  assign new_n6072_ = ~pi0217 | ~new_n6035_;
  assign new_n6073_ = ~new_n6027_ | ~new_n3593_;
  assign new_n6074_ = ~new_n3655_ | ~new_n3578_;
  assign new_n6075_ = ~new_n6026_ | ~new_n3577_;
  assign new_n6076_ = ~new_n3530_ | ~new_n3569_;
  assign new_n6077_ = ~pi0218 | ~new_n6035_;
  assign new_n6078_ = ~new_n4326_;
  assign new_n6079_ = ~new_n4325_;
  assign new_n6080_ = ~new_n3615_ | ~new_n5498_;
  assign new_n6081_ = ~new_n4328_;
  assign new_n6082_ = ~new_n5814_ | ~new_n5800_;
  assign new_n6083_ = ~new_n4327_;
  assign new_n6084_ = ~new_n3645_ | ~new_n4327_;
  assign new_n6085_ = ~new_n6081_ | ~new_n6084_;
  assign new_n6086_ = ~pi0175 | ~new_n4325_;
  assign new_n6087_ = ~new_n4614_ | ~new_n6085_;
  assign new_n6088_ = ~new_n6083_ | ~new_n5478_;
  assign new_n6089_ = ~new_n3645_ | ~new_n6088_;
  assign new_n6090_ = ~new_n6079_ | ~new_n3601_;
  assign new_n6091_ = ~new_n3656_ | ~new_n3592_;
  assign new_n6092_ = ~new_n6078_ | ~new_n3591_;
  assign new_n6093_ = ~new_n3529_ | ~new_n3576_;
  assign new_n6094_ = ~pi0219 | ~new_n6087_;
  assign new_n6095_ = ~new_n6079_ | ~new_n3599_;
  assign new_n6096_ = ~new_n3656_ | ~new_n3590_;
  assign new_n6097_ = ~new_n6078_ | ~new_n3589_;
  assign new_n6098_ = ~new_n3529_ | ~new_n3575_;
  assign new_n6099_ = ~pi0220 | ~new_n6087_;
  assign new_n6100_ = ~new_n6079_ | ~new_n3598_;
  assign new_n6101_ = ~new_n3656_ | ~new_n3588_;
  assign new_n6102_ = ~new_n6078_ | ~new_n3587_;
  assign new_n6103_ = ~new_n3529_ | ~new_n3574_;
  assign new_n6104_ = ~pi0221 | ~new_n6087_;
  assign new_n6105_ = ~new_n6079_ | ~new_n3597_;
  assign new_n6106_ = ~new_n3656_ | ~new_n3586_;
  assign new_n6107_ = ~new_n6078_ | ~new_n3585_;
  assign new_n6108_ = ~new_n3529_ | ~new_n3573_;
  assign new_n6109_ = ~pi0222 | ~new_n6087_;
  assign new_n6110_ = ~new_n6079_ | ~new_n3596_;
  assign new_n6111_ = ~new_n3656_ | ~new_n3584_;
  assign new_n6112_ = ~new_n6078_ | ~new_n3583_;
  assign new_n6113_ = ~new_n3529_ | ~new_n3572_;
  assign new_n6114_ = ~pi0223 | ~new_n6087_;
  assign new_n6115_ = ~new_n6079_ | ~new_n3595_;
  assign new_n6116_ = ~new_n3656_ | ~new_n3582_;
  assign new_n6117_ = ~new_n6078_ | ~new_n3581_;
  assign new_n6118_ = ~new_n3529_ | ~new_n3571_;
  assign new_n6119_ = ~pi0224 | ~new_n6087_;
  assign new_n6120_ = ~new_n6079_ | ~new_n3594_;
  assign new_n6121_ = ~new_n3656_ | ~new_n3580_;
  assign new_n6122_ = ~new_n6078_ | ~new_n3579_;
  assign new_n6123_ = ~new_n3529_ | ~new_n3570_;
  assign new_n6124_ = ~pi0225 | ~new_n6087_;
  assign new_n6125_ = ~new_n6079_ | ~new_n3593_;
  assign new_n6126_ = ~new_n3656_ | ~new_n3578_;
  assign new_n6127_ = ~new_n6078_ | ~new_n3577_;
  assign new_n6128_ = ~new_n3529_ | ~new_n3569_;
  assign new_n6129_ = ~pi0226 | ~new_n6087_;
  assign new_n6130_ = ~new_n4330_;
  assign new_n6131_ = ~new_n4329_;
  assign new_n6132_ = ~new_n3615_ | ~new_n5499_;
  assign new_n6133_ = ~new_n4332_;
  assign new_n6134_ = ~new_n5814_ | ~new_n5801_;
  assign new_n6135_ = ~new_n4331_;
  assign new_n6136_ = ~new_n3645_ | ~new_n4331_;
  assign new_n6137_ = ~new_n6133_ | ~new_n6136_;
  assign new_n6138_ = ~pi0175 | ~new_n4329_;
  assign new_n6139_ = ~new_n4632_ | ~new_n6137_;
  assign new_n6140_ = ~new_n6135_ | ~new_n5478_;
  assign new_n6141_ = ~new_n3645_ | ~new_n6140_;
  assign new_n6142_ = ~new_n6131_ | ~new_n3601_;
  assign new_n6143_ = ~new_n3658_ | ~new_n3592_;
  assign new_n6144_ = ~new_n6130_ | ~new_n3591_;
  assign new_n6145_ = ~new_n3528_ | ~new_n3576_;
  assign new_n6146_ = ~pi0227 | ~new_n6139_;
  assign new_n6147_ = ~new_n6131_ | ~new_n3599_;
  assign new_n6148_ = ~new_n3658_ | ~new_n3590_;
  assign new_n6149_ = ~new_n6130_ | ~new_n3589_;
  assign new_n6150_ = ~new_n3528_ | ~new_n3575_;
  assign new_n6151_ = ~pi0228 | ~new_n6139_;
  assign new_n6152_ = ~new_n6131_ | ~new_n3598_;
  assign new_n6153_ = ~new_n3658_ | ~new_n3588_;
  assign new_n6154_ = ~new_n6130_ | ~new_n3587_;
  assign new_n6155_ = ~new_n3528_ | ~new_n3574_;
  assign new_n6156_ = ~pi0229 | ~new_n6139_;
  assign new_n6157_ = ~new_n6131_ | ~new_n3597_;
  assign new_n6158_ = ~new_n3658_ | ~new_n3586_;
  assign new_n6159_ = ~new_n6130_ | ~new_n3585_;
  assign new_n6160_ = ~new_n3528_ | ~new_n3573_;
  assign new_n6161_ = ~pi0230 | ~new_n6139_;
  assign new_n6162_ = ~new_n6131_ | ~new_n3596_;
  assign new_n6163_ = ~new_n3658_ | ~new_n3584_;
  assign new_n6164_ = ~new_n6130_ | ~new_n3583_;
  assign new_n6165_ = ~new_n3528_ | ~new_n3572_;
  assign new_n6166_ = ~pi0231 | ~new_n6139_;
  assign new_n6167_ = ~new_n6131_ | ~new_n3595_;
  assign new_n6168_ = ~new_n3658_ | ~new_n3582_;
  assign new_n6169_ = ~new_n6130_ | ~new_n3581_;
  assign new_n6170_ = ~new_n3528_ | ~new_n3571_;
  assign new_n6171_ = ~pi0232 | ~new_n6139_;
  assign new_n6172_ = ~new_n6131_ | ~new_n3594_;
  assign new_n6173_ = ~new_n3658_ | ~new_n3580_;
  assign new_n6174_ = ~new_n6130_ | ~new_n3579_;
  assign new_n6175_ = ~new_n3528_ | ~new_n3570_;
  assign new_n6176_ = ~pi0233 | ~new_n6139_;
  assign new_n6177_ = ~new_n6131_ | ~new_n3593_;
  assign new_n6178_ = ~new_n3658_ | ~new_n3578_;
  assign new_n6179_ = ~new_n6130_ | ~new_n3577_;
  assign new_n6180_ = ~new_n3528_ | ~new_n3569_;
  assign new_n6181_ = ~pi0234 | ~new_n6139_;
  assign new_n6182_ = ~new_n4334_;
  assign new_n6183_ = ~new_n4333_;
  assign new_n6184_ = ~new_n4227_;
  assign new_n6185_ = ~new_n5814_ | ~new_n3652_;
  assign new_n6186_ = ~new_n4335_;
  assign new_n6187_ = ~new_n3645_ | ~new_n4335_;
  assign new_n6188_ = ~new_n6187_ | ~new_n4227_;
  assign new_n6189_ = ~pi0175 | ~new_n4333_;
  assign new_n6190_ = ~new_n4649_ | ~new_n6188_;
  assign new_n6191_ = ~new_n6186_ | ~new_n5478_;
  assign new_n6192_ = ~new_n3645_ | ~new_n6191_;
  assign new_n6193_ = ~new_n6183_ | ~new_n3601_;
  assign new_n6194_ = ~new_n3659_ | ~new_n3592_;
  assign new_n6195_ = ~new_n6182_ | ~new_n3591_;
  assign new_n6196_ = ~new_n3527_ | ~new_n3576_;
  assign new_n6197_ = ~pi0235 | ~new_n6190_;
  assign new_n6198_ = ~new_n6183_ | ~new_n3599_;
  assign new_n6199_ = ~new_n3659_ | ~new_n3590_;
  assign new_n6200_ = ~new_n6182_ | ~new_n3589_;
  assign new_n6201_ = ~new_n3527_ | ~new_n3575_;
  assign new_n6202_ = ~pi0236 | ~new_n6190_;
  assign new_n6203_ = ~new_n6183_ | ~new_n3598_;
  assign new_n6204_ = ~new_n3659_ | ~new_n3588_;
  assign new_n6205_ = ~new_n6182_ | ~new_n3587_;
  assign new_n6206_ = ~new_n3527_ | ~new_n3574_;
  assign new_n6207_ = ~pi0237 | ~new_n6190_;
  assign new_n6208_ = ~new_n6183_ | ~new_n3597_;
  assign new_n6209_ = ~new_n3659_ | ~new_n3586_;
  assign new_n6210_ = ~new_n6182_ | ~new_n3585_;
  assign new_n6211_ = ~new_n3527_ | ~new_n3573_;
  assign new_n6212_ = ~pi0238 | ~new_n6190_;
  assign new_n6213_ = ~new_n6183_ | ~new_n3596_;
  assign new_n6214_ = ~new_n3659_ | ~new_n3584_;
  assign new_n6215_ = ~new_n6182_ | ~new_n3583_;
  assign new_n6216_ = ~new_n3527_ | ~new_n3572_;
  assign new_n6217_ = ~pi0239 | ~new_n6190_;
  assign new_n6218_ = ~new_n6183_ | ~new_n3595_;
  assign new_n6219_ = ~new_n3659_ | ~new_n3582_;
  assign new_n6220_ = ~new_n6182_ | ~new_n3581_;
  assign new_n6221_ = ~new_n3527_ | ~new_n3571_;
  assign new_n6222_ = ~pi0240 | ~new_n6190_;
  assign new_n6223_ = ~new_n6183_ | ~new_n3594_;
  assign new_n6224_ = ~new_n3659_ | ~new_n3580_;
  assign new_n6225_ = ~new_n6182_ | ~new_n3579_;
  assign new_n6226_ = ~new_n3527_ | ~new_n3570_;
  assign new_n6227_ = ~pi0241 | ~new_n6190_;
  assign new_n6228_ = ~new_n6183_ | ~new_n3593_;
  assign new_n6229_ = ~new_n3659_ | ~new_n3578_;
  assign new_n6230_ = ~new_n6182_ | ~new_n3577_;
  assign new_n6231_ = ~new_n3527_ | ~new_n3569_;
  assign new_n6232_ = ~pi0242 | ~new_n6190_;
  assign new_n6233_ = ~new_n4339_;
  assign new_n6234_ = ~new_n4341_;
  assign new_n6235_ = ~new_n4340_;
  assign new_n6236_ = ~new_n3645_ | ~new_n4340_;
  assign new_n6237_ = ~new_n6234_ | ~new_n6236_;
  assign new_n6238_ = ~pi0175 | ~new_n4336_;
  assign new_n6239_ = ~new_n4666_ | ~new_n6237_;
  assign new_n6240_ = ~new_n6235_ | ~new_n5478_;
  assign new_n6241_ = ~new_n3645_ | ~new_n6240_;
  assign new_n6242_ = ~new_n5806_ | ~new_n3601_;
  assign new_n6243_ = ~new_n5482_ | ~new_n3592_;
  assign new_n6244_ = ~new_n6233_ | ~new_n3591_;
  assign new_n6245_ = ~new_n3526_ | ~new_n3576_;
  assign new_n6246_ = ~pi0243 | ~new_n6239_;
  assign new_n6247_ = ~new_n5806_ | ~new_n3599_;
  assign new_n6248_ = ~new_n5482_ | ~new_n3590_;
  assign new_n6249_ = ~new_n6233_ | ~new_n3589_;
  assign new_n6250_ = ~new_n3526_ | ~new_n3575_;
  assign new_n6251_ = ~pi0244 | ~new_n6239_;
  assign new_n6252_ = ~new_n5806_ | ~new_n3598_;
  assign new_n6253_ = ~new_n5482_ | ~new_n3588_;
  assign new_n6254_ = ~new_n6233_ | ~new_n3587_;
  assign new_n6255_ = ~new_n3526_ | ~new_n3574_;
  assign new_n6256_ = ~pi0245 | ~new_n6239_;
  assign new_n6257_ = ~new_n5806_ | ~new_n3597_;
  assign new_n6258_ = ~new_n5482_ | ~new_n3586_;
  assign new_n6259_ = ~new_n6233_ | ~new_n3585_;
  assign new_n6260_ = ~new_n3526_ | ~new_n3573_;
  assign new_n6261_ = ~pi0246 | ~new_n6239_;
  assign new_n6262_ = ~new_n5806_ | ~new_n3596_;
  assign new_n6263_ = ~new_n5482_ | ~new_n3584_;
  assign new_n6264_ = ~new_n6233_ | ~new_n3583_;
  assign new_n6265_ = ~new_n3526_ | ~new_n3572_;
  assign new_n6266_ = ~pi0247 | ~new_n6239_;
  assign new_n6267_ = ~new_n5806_ | ~new_n3595_;
  assign new_n6268_ = ~new_n5482_ | ~new_n3582_;
  assign new_n6269_ = ~new_n6233_ | ~new_n3581_;
  assign new_n6270_ = ~new_n3526_ | ~new_n3571_;
  assign new_n6271_ = ~pi0248 | ~new_n6239_;
  assign new_n6272_ = ~new_n5806_ | ~new_n3594_;
  assign new_n6273_ = ~new_n5482_ | ~new_n3580_;
  assign new_n6274_ = ~new_n6233_ | ~new_n3579_;
  assign new_n6275_ = ~new_n3526_ | ~new_n3570_;
  assign new_n6276_ = ~pi0249 | ~new_n6239_;
  assign new_n6277_ = ~new_n5806_ | ~new_n3593_;
  assign new_n6278_ = ~new_n5482_ | ~new_n3578_;
  assign new_n6279_ = ~new_n6233_ | ~new_n3577_;
  assign new_n6280_ = ~new_n3526_ | ~new_n3569_;
  assign new_n6281_ = ~pi0250 | ~new_n6239_;
  assign new_n6282_ = ~new_n4343_;
  assign new_n6283_ = ~new_n4342_;
  assign new_n6284_ = ~new_n5498_ | ~new_n3614_;
  assign new_n6285_ = ~new_n4345_;
  assign new_n6286_ = ~new_n5800_ | ~new_n3641_;
  assign new_n6287_ = ~new_n4344_;
  assign new_n6288_ = ~new_n3645_ | ~new_n4344_;
  assign new_n6289_ = ~new_n6285_ | ~new_n6288_;
  assign new_n6290_ = ~pi0175 | ~new_n4342_;
  assign new_n6291_ = ~new_n4684_ | ~new_n6289_;
  assign new_n6292_ = ~new_n6287_ | ~new_n5478_;
  assign new_n6293_ = ~new_n3645_ | ~new_n6292_;
  assign new_n6294_ = ~new_n6283_ | ~new_n3601_;
  assign new_n6295_ = ~new_n3661_ | ~new_n3592_;
  assign new_n6296_ = ~new_n6282_ | ~new_n3591_;
  assign new_n6297_ = ~new_n3525_ | ~new_n3576_;
  assign new_n6298_ = ~pi0251 | ~new_n6291_;
  assign new_n6299_ = ~new_n6283_ | ~new_n3599_;
  assign new_n6300_ = ~new_n3661_ | ~new_n3590_;
  assign new_n6301_ = ~new_n6282_ | ~new_n3589_;
  assign new_n6302_ = ~new_n3525_ | ~new_n3575_;
  assign new_n6303_ = ~pi0252 | ~new_n6291_;
  assign new_n6304_ = ~new_n6283_ | ~new_n3598_;
  assign new_n6305_ = ~new_n3661_ | ~new_n3588_;
  assign new_n6306_ = ~new_n6282_ | ~new_n3587_;
  assign new_n6307_ = ~new_n3525_ | ~new_n3574_;
  assign new_n6308_ = ~pi0253 | ~new_n6291_;
  assign new_n6309_ = ~new_n6283_ | ~new_n3597_;
  assign new_n6310_ = ~new_n3661_ | ~new_n3586_;
  assign new_n6311_ = ~new_n6282_ | ~new_n3585_;
  assign new_n6312_ = ~new_n3525_ | ~new_n3573_;
  assign new_n6313_ = ~pi0254 | ~new_n6291_;
  assign new_n6314_ = ~new_n6283_ | ~new_n3596_;
  assign new_n6315_ = ~new_n3661_ | ~new_n3584_;
  assign new_n6316_ = ~new_n6282_ | ~new_n3583_;
  assign new_n6317_ = ~new_n3525_ | ~new_n3572_;
  assign new_n6318_ = ~pi0255 | ~new_n6291_;
  assign new_n6319_ = ~new_n6283_ | ~new_n3595_;
  assign new_n6320_ = ~new_n3661_ | ~new_n3582_;
  assign new_n6321_ = ~new_n6282_ | ~new_n3581_;
  assign new_n6322_ = ~new_n3525_ | ~new_n3571_;
  assign new_n6323_ = ~pi0256 | ~new_n6291_;
  assign new_n6324_ = ~new_n6283_ | ~new_n3594_;
  assign new_n6325_ = ~new_n3661_ | ~new_n3580_;
  assign new_n6326_ = ~new_n6282_ | ~new_n3579_;
  assign new_n6327_ = ~new_n3525_ | ~new_n3570_;
  assign new_n6328_ = ~pi0257 | ~new_n6291_;
  assign new_n6329_ = ~new_n6283_ | ~new_n3593_;
  assign new_n6330_ = ~new_n3661_ | ~new_n3578_;
  assign new_n6331_ = ~new_n6282_ | ~new_n3577_;
  assign new_n6332_ = ~new_n3525_ | ~new_n3569_;
  assign new_n6333_ = ~pi0258 | ~new_n6291_;
  assign new_n6334_ = ~new_n4347_;
  assign new_n6335_ = ~new_n4346_;
  assign new_n6336_ = ~new_n5499_ | ~new_n3614_;
  assign new_n6337_ = ~new_n4349_;
  assign new_n6338_ = ~new_n5801_ | ~new_n3641_;
  assign new_n6339_ = ~new_n4348_;
  assign new_n6340_ = ~new_n3645_ | ~new_n4348_;
  assign new_n6341_ = ~new_n6337_ | ~new_n6340_;
  assign new_n6342_ = ~pi0175 | ~new_n4346_;
  assign new_n6343_ = ~new_n4702_ | ~new_n6341_;
  assign new_n6344_ = ~new_n6339_ | ~new_n5478_;
  assign new_n6345_ = ~new_n3645_ | ~new_n6344_;
  assign new_n6346_ = ~new_n6335_ | ~new_n3601_;
  assign new_n6347_ = ~new_n3662_ | ~new_n3592_;
  assign new_n6348_ = ~new_n6334_ | ~new_n3591_;
  assign new_n6349_ = ~new_n3524_ | ~new_n3576_;
  assign new_n6350_ = ~pi0259 | ~new_n6343_;
  assign new_n6351_ = ~new_n6335_ | ~new_n3599_;
  assign new_n6352_ = ~new_n3662_ | ~new_n3590_;
  assign new_n6353_ = ~new_n6334_ | ~new_n3589_;
  assign new_n6354_ = ~new_n3524_ | ~new_n3575_;
  assign new_n6355_ = ~pi0260 | ~new_n6343_;
  assign new_n6356_ = ~new_n6335_ | ~new_n3598_;
  assign new_n6357_ = ~new_n3662_ | ~new_n3588_;
  assign new_n6358_ = ~new_n6334_ | ~new_n3587_;
  assign new_n6359_ = ~new_n3524_ | ~new_n3574_;
  assign new_n6360_ = ~pi0261 | ~new_n6343_;
  assign new_n6361_ = ~new_n6335_ | ~new_n3597_;
  assign new_n6362_ = ~new_n3662_ | ~new_n3586_;
  assign new_n6363_ = ~new_n6334_ | ~new_n3585_;
  assign new_n6364_ = ~new_n3524_ | ~new_n3573_;
  assign new_n6365_ = ~pi0262 | ~new_n6343_;
  assign new_n6366_ = ~new_n6335_ | ~new_n3596_;
  assign new_n6367_ = ~new_n3662_ | ~new_n3584_;
  assign new_n6368_ = ~new_n6334_ | ~new_n3583_;
  assign new_n6369_ = ~new_n3524_ | ~new_n3572_;
  assign new_n6370_ = ~pi0263 | ~new_n6343_;
  assign new_n6371_ = ~new_n6335_ | ~new_n3595_;
  assign new_n6372_ = ~new_n3662_ | ~new_n3582_;
  assign new_n6373_ = ~new_n6334_ | ~new_n3581_;
  assign new_n6374_ = ~new_n3524_ | ~new_n3571_;
  assign new_n6375_ = ~pi0264 | ~new_n6343_;
  assign new_n6376_ = ~new_n6335_ | ~new_n3594_;
  assign new_n6377_ = ~new_n3662_ | ~new_n3580_;
  assign new_n6378_ = ~new_n6334_ | ~new_n3579_;
  assign new_n6379_ = ~new_n3524_ | ~new_n3570_;
  assign new_n6380_ = ~pi0265 | ~new_n6343_;
  assign new_n6381_ = ~new_n6335_ | ~new_n3593_;
  assign new_n6382_ = ~new_n3662_ | ~new_n3578_;
  assign new_n6383_ = ~new_n6334_ | ~new_n3577_;
  assign new_n6384_ = ~new_n3524_ | ~new_n3569_;
  assign new_n6385_ = ~pi0266 | ~new_n6343_;
  assign new_n6386_ = ~new_n4351_;
  assign new_n6387_ = ~new_n4350_;
  assign new_n6388_ = ~new_n4228_;
  assign new_n6389_ = ~new_n3652_ | ~new_n3641_;
  assign new_n6390_ = ~new_n4351_ | ~new_n6389_;
  assign new_n6391_ = ~new_n3645_ | ~new_n6390_;
  assign new_n6392_ = ~new_n6391_ | ~new_n4228_;
  assign new_n6393_ = ~pi0175 | ~new_n4350_;
  assign new_n6394_ = ~new_n4720_ | ~new_n6392_;
  assign new_n6395_ = ~new_n3645_ | ~new_n4292_;
  assign new_n6396_ = ~new_n6387_ | ~new_n3601_;
  assign new_n6397_ = ~new_n3663_ | ~new_n3592_;
  assign new_n6398_ = ~new_n6386_ | ~new_n3591_;
  assign new_n6399_ = ~new_n3523_ | ~new_n3576_;
  assign new_n6400_ = ~pi0267 | ~new_n6394_;
  assign new_n6401_ = ~new_n6387_ | ~new_n3599_;
  assign new_n6402_ = ~new_n3663_ | ~new_n3590_;
  assign new_n6403_ = ~new_n6386_ | ~new_n3589_;
  assign new_n6404_ = ~new_n3523_ | ~new_n3575_;
  assign new_n6405_ = ~pi0268 | ~new_n6394_;
  assign new_n6406_ = ~new_n6387_ | ~new_n3598_;
  assign new_n6407_ = ~new_n3663_ | ~new_n3588_;
  assign new_n6408_ = ~new_n6386_ | ~new_n3587_;
  assign new_n6409_ = ~new_n3523_ | ~new_n3574_;
  assign new_n6410_ = ~pi0269 | ~new_n6394_;
  assign new_n6411_ = ~new_n6387_ | ~new_n3597_;
  assign new_n6412_ = ~new_n3663_ | ~new_n3586_;
  assign new_n6413_ = ~new_n6386_ | ~new_n3585_;
  assign new_n6414_ = ~new_n3523_ | ~new_n3573_;
  assign new_n6415_ = ~pi0270 | ~new_n6394_;
  assign new_n6416_ = ~new_n6387_ | ~new_n3596_;
  assign new_n6417_ = ~new_n3663_ | ~new_n3584_;
  assign new_n6418_ = ~new_n6386_ | ~new_n3583_;
  assign new_n6419_ = ~new_n3523_ | ~new_n3572_;
  assign new_n6420_ = ~pi0271 | ~new_n6394_;
  assign new_n6421_ = ~new_n6387_ | ~new_n3595_;
  assign new_n6422_ = ~new_n3663_ | ~new_n3582_;
  assign new_n6423_ = ~new_n6386_ | ~new_n3581_;
  assign new_n6424_ = ~new_n3523_ | ~new_n3571_;
  assign new_n6425_ = ~pi0272 | ~new_n6394_;
  assign new_n6426_ = ~new_n6387_ | ~new_n3594_;
  assign new_n6427_ = ~new_n3663_ | ~new_n3580_;
  assign new_n6428_ = ~new_n6386_ | ~new_n3579_;
  assign new_n6429_ = ~new_n3523_ | ~new_n3570_;
  assign new_n6430_ = ~pi0273 | ~new_n6394_;
  assign new_n6431_ = ~new_n6387_ | ~new_n3593_;
  assign new_n6432_ = ~new_n3663_ | ~new_n3578_;
  assign new_n6433_ = ~new_n6386_ | ~new_n3577_;
  assign new_n6434_ = ~new_n3523_ | ~new_n3569_;
  assign new_n6435_ = ~pi0274 | ~new_n6394_;
  assign new_n6436_ = ~new_n4353_;
  assign new_n6437_ = ~new_n4352_;
  assign new_n6438_ = ~new_n3616_ | ~new_n5809_;
  assign new_n6439_ = ~new_n4354_;
  assign new_n6440_ = ~new_n3665_ | ~new_n5813_;
  assign new_n6441_ = ~new_n4353_ | ~new_n6440_;
  assign new_n6442_ = ~new_n3645_ | ~new_n6441_;
  assign new_n6443_ = ~new_n6439_ | ~new_n6442_;
  assign new_n6444_ = ~pi0175 | ~new_n4352_;
  assign new_n6445_ = ~new_n4738_ | ~new_n6443_;
  assign new_n6446_ = ~new_n3645_ | ~new_n4292_;
  assign new_n6447_ = ~new_n6437_ | ~new_n3601_;
  assign new_n6448_ = ~new_n3666_ | ~new_n3592_;
  assign new_n6449_ = ~new_n6436_ | ~new_n3591_;
  assign new_n6450_ = ~new_n3522_ | ~new_n3576_;
  assign new_n6451_ = ~pi0275 | ~new_n6445_;
  assign new_n6452_ = ~new_n6437_ | ~new_n3599_;
  assign new_n6453_ = ~new_n3666_ | ~new_n3590_;
  assign new_n6454_ = ~new_n6436_ | ~new_n3589_;
  assign new_n6455_ = ~new_n3522_ | ~new_n3575_;
  assign new_n6456_ = ~pi0276 | ~new_n6445_;
  assign new_n6457_ = ~new_n6437_ | ~new_n3598_;
  assign new_n6458_ = ~new_n3666_ | ~new_n3588_;
  assign new_n6459_ = ~new_n6436_ | ~new_n3587_;
  assign new_n6460_ = ~new_n3522_ | ~new_n3574_;
  assign new_n6461_ = ~pi0277 | ~new_n6445_;
  assign new_n6462_ = ~new_n6437_ | ~new_n3597_;
  assign new_n6463_ = ~new_n3666_ | ~new_n3586_;
  assign new_n6464_ = ~new_n6436_ | ~new_n3585_;
  assign new_n6465_ = ~new_n3522_ | ~new_n3573_;
  assign new_n6466_ = ~pi0278 | ~new_n6445_;
  assign new_n6467_ = ~new_n6437_ | ~new_n3596_;
  assign new_n6468_ = ~new_n3666_ | ~new_n3584_;
  assign new_n6469_ = ~new_n6436_ | ~new_n3583_;
  assign new_n6470_ = ~new_n3522_ | ~new_n3572_;
  assign new_n6471_ = ~pi0279 | ~new_n6445_;
  assign new_n6472_ = ~new_n6437_ | ~new_n3595_;
  assign new_n6473_ = ~new_n3666_ | ~new_n3582_;
  assign new_n6474_ = ~new_n6436_ | ~new_n3581_;
  assign new_n6475_ = ~new_n3522_ | ~new_n3571_;
  assign new_n6476_ = ~pi0280 | ~new_n6445_;
  assign new_n6477_ = ~new_n6437_ | ~new_n3594_;
  assign new_n6478_ = ~new_n3666_ | ~new_n3580_;
  assign new_n6479_ = ~new_n6436_ | ~new_n3579_;
  assign new_n6480_ = ~new_n3522_ | ~new_n3570_;
  assign new_n6481_ = ~pi0281 | ~new_n6445_;
  assign new_n6482_ = ~new_n6437_ | ~new_n3593_;
  assign new_n6483_ = ~new_n3666_ | ~new_n3578_;
  assign new_n6484_ = ~new_n6436_ | ~new_n3577_;
  assign new_n6485_ = ~new_n3522_ | ~new_n3569_;
  assign new_n6486_ = ~pi0282 | ~new_n6445_;
  assign new_n6487_ = ~new_n4356_;
  assign new_n6488_ = ~new_n4355_;
  assign new_n6489_ = ~new_n3616_ | ~new_n5498_;
  assign new_n6490_ = ~new_n4357_;
  assign new_n6491_ = ~new_n3665_ | ~new_n5800_;
  assign new_n6492_ = ~new_n4356_ | ~new_n6491_;
  assign new_n6493_ = ~new_n3645_ | ~new_n6492_;
  assign new_n6494_ = ~new_n6490_ | ~new_n6493_;
  assign new_n6495_ = ~pi0175 | ~new_n4355_;
  assign new_n6496_ = ~new_n4755_ | ~new_n6494_;
  assign new_n6497_ = ~new_n3645_ | ~new_n4292_;
  assign new_n6498_ = ~new_n6488_ | ~new_n3601_;
  assign new_n6499_ = ~new_n3667_ | ~new_n3592_;
  assign new_n6500_ = ~new_n6487_ | ~new_n3591_;
  assign new_n6501_ = ~new_n3521_ | ~new_n3576_;
  assign new_n6502_ = ~pi0283 | ~new_n6496_;
  assign new_n6503_ = ~new_n6488_ | ~new_n3599_;
  assign new_n6504_ = ~new_n3667_ | ~new_n3590_;
  assign new_n6505_ = ~new_n6487_ | ~new_n3589_;
  assign new_n6506_ = ~new_n3521_ | ~new_n3575_;
  assign new_n6507_ = ~pi0284 | ~new_n6496_;
  assign new_n6508_ = ~new_n6488_ | ~new_n3598_;
  assign new_n6509_ = ~new_n3667_ | ~new_n3588_;
  assign new_n6510_ = ~new_n6487_ | ~new_n3587_;
  assign new_n6511_ = ~new_n3521_ | ~new_n3574_;
  assign new_n6512_ = ~pi0285 | ~new_n6496_;
  assign new_n6513_ = ~new_n6488_ | ~new_n3597_;
  assign new_n6514_ = ~new_n3667_ | ~new_n3586_;
  assign new_n6515_ = ~new_n6487_ | ~new_n3585_;
  assign new_n6516_ = ~new_n3521_ | ~new_n3573_;
  assign new_n6517_ = ~pi0286 | ~new_n6496_;
  assign new_n6518_ = ~new_n6488_ | ~new_n3596_;
  assign new_n6519_ = ~new_n3667_ | ~new_n3584_;
  assign new_n6520_ = ~new_n6487_ | ~new_n3583_;
  assign new_n6521_ = ~new_n3521_ | ~new_n3572_;
  assign new_n6522_ = ~pi0287 | ~new_n6496_;
  assign new_n6523_ = ~new_n6488_ | ~new_n3595_;
  assign new_n6524_ = ~new_n3667_ | ~new_n3582_;
  assign new_n6525_ = ~new_n6487_ | ~new_n3581_;
  assign new_n6526_ = ~new_n3521_ | ~new_n3571_;
  assign new_n6527_ = ~pi0288 | ~new_n6496_;
  assign new_n6528_ = ~new_n6488_ | ~new_n3594_;
  assign new_n6529_ = ~new_n3667_ | ~new_n3580_;
  assign new_n6530_ = ~new_n6487_ | ~new_n3579_;
  assign new_n6531_ = ~new_n3521_ | ~new_n3570_;
  assign new_n6532_ = ~pi0289 | ~new_n6496_;
  assign new_n6533_ = ~new_n6488_ | ~new_n3593_;
  assign new_n6534_ = ~new_n3667_ | ~new_n3578_;
  assign new_n6535_ = ~new_n6487_ | ~new_n3577_;
  assign new_n6536_ = ~new_n3521_ | ~new_n3569_;
  assign new_n6537_ = ~pi0290 | ~new_n6496_;
  assign new_n6538_ = ~new_n4359_;
  assign new_n6539_ = ~new_n4358_;
  assign new_n6540_ = ~new_n3616_ | ~new_n5499_;
  assign new_n6541_ = ~new_n4360_;
  assign new_n6542_ = ~new_n3665_ | ~new_n5801_;
  assign new_n6543_ = ~new_n4359_ | ~new_n6542_;
  assign new_n6544_ = ~new_n3645_ | ~new_n6543_;
  assign new_n6545_ = ~new_n6541_ | ~new_n6544_;
  assign new_n6546_ = ~pi0175 | ~new_n4358_;
  assign new_n6547_ = ~new_n4773_ | ~new_n6545_;
  assign new_n6548_ = ~new_n3645_ | ~new_n4292_;
  assign new_n6549_ = ~new_n6539_ | ~new_n3601_;
  assign new_n6550_ = ~new_n3668_ | ~new_n3592_;
  assign new_n6551_ = ~new_n6538_ | ~new_n3591_;
  assign new_n6552_ = ~new_n3520_ | ~new_n3576_;
  assign new_n6553_ = ~pi0291 | ~new_n6547_;
  assign new_n6554_ = ~new_n6539_ | ~new_n3599_;
  assign new_n6555_ = ~new_n3668_ | ~new_n3590_;
  assign new_n6556_ = ~new_n6538_ | ~new_n3589_;
  assign new_n6557_ = ~new_n3520_ | ~new_n3575_;
  assign new_n6558_ = ~pi0292 | ~new_n6547_;
  assign new_n6559_ = ~new_n6539_ | ~new_n3598_;
  assign new_n6560_ = ~new_n3668_ | ~new_n3588_;
  assign new_n6561_ = ~new_n6538_ | ~new_n3587_;
  assign new_n6562_ = ~new_n3520_ | ~new_n3574_;
  assign new_n6563_ = ~pi0293 | ~new_n6547_;
  assign new_n6564_ = ~new_n6539_ | ~new_n3597_;
  assign new_n6565_ = ~new_n3668_ | ~new_n3586_;
  assign new_n6566_ = ~new_n6538_ | ~new_n3585_;
  assign new_n6567_ = ~new_n3520_ | ~new_n3573_;
  assign new_n6568_ = ~pi0294 | ~new_n6547_;
  assign new_n6569_ = ~new_n6539_ | ~new_n3596_;
  assign new_n6570_ = ~new_n3668_ | ~new_n3584_;
  assign new_n6571_ = ~new_n6538_ | ~new_n3583_;
  assign new_n6572_ = ~new_n3520_ | ~new_n3572_;
  assign new_n6573_ = ~pi0295 | ~new_n6547_;
  assign new_n6574_ = ~new_n6539_ | ~new_n3595_;
  assign new_n6575_ = ~new_n3668_ | ~new_n3582_;
  assign new_n6576_ = ~new_n6538_ | ~new_n3581_;
  assign new_n6577_ = ~new_n3520_ | ~new_n3571_;
  assign new_n6578_ = ~pi0296 | ~new_n6547_;
  assign new_n6579_ = ~new_n6539_ | ~new_n3594_;
  assign new_n6580_ = ~new_n3668_ | ~new_n3580_;
  assign new_n6581_ = ~new_n6538_ | ~new_n3579_;
  assign new_n6582_ = ~new_n3520_ | ~new_n3570_;
  assign new_n6583_ = ~pi0297 | ~new_n6547_;
  assign new_n6584_ = ~new_n6539_ | ~new_n3593_;
  assign new_n6585_ = ~new_n3668_ | ~new_n3578_;
  assign new_n6586_ = ~new_n6538_ | ~new_n3577_;
  assign new_n6587_ = ~new_n3520_ | ~new_n3569_;
  assign new_n6588_ = ~pi0298 | ~new_n6547_;
  assign new_n6589_ = ~new_n4362_;
  assign new_n6590_ = ~new_n4361_;
  assign new_n6591_ = ~new_n4229_;
  assign new_n6592_ = ~new_n3665_ | ~new_n3652_;
  assign new_n6593_ = ~new_n4362_ | ~new_n6592_;
  assign new_n6594_ = ~new_n3645_ | ~new_n6593_;
  assign new_n6595_ = ~new_n6594_ | ~new_n4229_;
  assign new_n6596_ = ~pi0175 | ~new_n4361_;
  assign new_n6597_ = ~new_n4791_ | ~new_n6595_;
  assign new_n6598_ = ~new_n3645_ | ~new_n4292_;
  assign new_n6599_ = ~new_n6590_ | ~new_n3601_;
  assign new_n6600_ = ~new_n3669_ | ~new_n3592_;
  assign new_n6601_ = ~new_n6589_ | ~new_n3591_;
  assign new_n6602_ = ~new_n3519_ | ~new_n3576_;
  assign new_n6603_ = ~pi0299 | ~new_n6597_;
  assign new_n6604_ = ~new_n6590_ | ~new_n3599_;
  assign new_n6605_ = ~new_n3669_ | ~new_n3590_;
  assign new_n6606_ = ~new_n6589_ | ~new_n3589_;
  assign new_n6607_ = ~new_n3519_ | ~new_n3575_;
  assign new_n6608_ = ~pi0300 | ~new_n6597_;
  assign new_n6609_ = ~new_n6590_ | ~new_n3598_;
  assign new_n6610_ = ~new_n3669_ | ~new_n3588_;
  assign new_n6611_ = ~new_n6589_ | ~new_n3587_;
  assign new_n6612_ = ~new_n3519_ | ~new_n3574_;
  assign new_n6613_ = ~pi0301 | ~new_n6597_;
  assign new_n6614_ = ~new_n6590_ | ~new_n3597_;
  assign new_n6615_ = ~new_n3669_ | ~new_n3586_;
  assign new_n6616_ = ~new_n6589_ | ~new_n3585_;
  assign new_n6617_ = ~new_n3519_ | ~new_n3573_;
  assign new_n6618_ = ~pi0302 | ~new_n6597_;
  assign new_n6619_ = ~new_n6590_ | ~new_n3596_;
  assign new_n6620_ = ~new_n3669_ | ~new_n3584_;
  assign new_n6621_ = ~new_n6589_ | ~new_n3583_;
  assign new_n6622_ = ~new_n3519_ | ~new_n3572_;
  assign new_n6623_ = ~pi0303 | ~new_n6597_;
  assign new_n6624_ = ~new_n6590_ | ~new_n3595_;
  assign new_n6625_ = ~new_n3669_ | ~new_n3582_;
  assign new_n6626_ = ~new_n6589_ | ~new_n3581_;
  assign new_n6627_ = ~new_n3519_ | ~new_n3571_;
  assign new_n6628_ = ~pi0304 | ~new_n6597_;
  assign new_n6629_ = ~new_n6590_ | ~new_n3594_;
  assign new_n6630_ = ~new_n3669_ | ~new_n3580_;
  assign new_n6631_ = ~new_n6589_ | ~new_n3579_;
  assign new_n6632_ = ~new_n3519_ | ~new_n3570_;
  assign new_n6633_ = ~pi0305 | ~new_n6597_;
  assign new_n6634_ = ~new_n6590_ | ~new_n3593_;
  assign new_n6635_ = ~new_n3669_ | ~new_n3578_;
  assign new_n6636_ = ~new_n6589_ | ~new_n3577_;
  assign new_n6637_ = ~new_n3519_ | ~new_n3569_;
  assign new_n6638_ = ~pi0306 | ~new_n6597_;
  assign new_n6639_ = ~new_n3670_ | ~new_n5495_ | ~new_n4811_ | ~new_n9073_;
  assign new_n6640_ = ~new_n4365_;
  assign new_n6641_ = ~new_n5452_ | ~new_n4365_;
  assign new_n6642_ = ~new_n25105_ | ~new_n5459_;
  assign new_n6643_ = ~new_n27146_ | ~new_n5458_;
  assign new_n6644_ = ~new_n4411_;
  assign new_n6645_ = ~new_n27144_ | ~new_n5460_;
  assign new_n6646_ = ~new_n22221_ | ~new_n3512_;
  assign new_n6647_ = ~new_n4410_;
  assign new_n6648_ = ~new_n4410_ | ~new_n3786_;
  assign new_n6649_ = ~new_n21854_ | ~new_n3513_;
  assign new_n6650_ = ~new_n5450_ | ~new_n4411_;
  assign new_n6651_ = ~new_n21624_ | ~new_n5461_;
  assign new_n6652_ = ~new_n5446_;
  assign new_n6653_ = ~new_n3546_ | ~new_n5446_;
  assign new_n6654_ = ~pi0175 | ~new_n4277_;
  assign new_n6655_ = ~new_n5439_;
  assign new_n6656_ = ~new_n4251_ | ~new_n4253_;
  assign new_n6657_ = ~pi0308 | ~new_n6656_;
  assign new_n6658_ = ~new_n3637_ | ~new_n4251_;
  assign new_n6659_ = ~pi0309 | ~pi0310;
  assign new_n6660_ = ~new_n4379_;
  assign new_n6661_ = ~pi0309 | ~new_n5488_;
  assign new_n6662_ = ~new_n4380_;
  assign new_n6663_ = ~new_n6640_ | ~new_n4263_;
  assign new_n6664_ = ~new_n5644_ | ~new_n5678_ | ~new_n5763_;
  assign new_n6665_ = ~new_n5452_ | ~new_n6663_;
  assign new_n6666_ = ~new_n4260_ | ~new_n9130_ | ~new_n9129_;
  assign new_n6667_ = ~new_n5479_ | ~new_n5500_;
  assign new_n6668_ = ~new_n6665_ | ~new_n4821_;
  assign new_n6669_ = ~new_n5678_ | ~new_n5763_;
  assign new_n6670_ = ~new_n5763_ | ~new_n4374_;
  assign new_n6671_ = ~new_n5712_ | ~new_n6670_ | ~new_n4372_;
  assign new_n6672_ = ~new_n5729_ | ~new_n5661_;
  assign new_n6673_ = ~new_n5644_ | ~new_n6672_;
  assign new_n6674_ = ~new_n4268_ | ~new_n4259_ | ~new_n4374_;
  assign new_n6675_ = ~new_n5729_ | ~new_n5763_ | ~new_n4260_;
  assign new_n6676_ = ~new_n5480_ | ~new_n4259_;
  assign new_n6677_ = ~new_n6674_ | ~new_n4258_;
  assign new_n6678_ = ~new_n4376_;
  assign new_n6679_ = ~new_n4267_ | ~new_n4270_;
  assign new_n6680_ = ~new_n3608_ | ~new_n4264_;
  assign new_n6681_ = ~new_n4377_;
  assign new_n6682_ = ~new_n3618_ | ~new_n4260_;
  assign new_n6683_ = ~new_n4385_ | ~new_n4375_;
  assign new_n6684_ = ~new_n3612_ | ~new_n6683_;
  assign new_n6685_ = ~new_n3674_ | ~new_n4373_;
  assign new_n6686_ = ~pi0311 | ~new_n6685_;
  assign new_n6687_ = ~new_n6681_ | ~new_n6686_;
  assign new_n6688_ = ~new_n3606_ | ~new_n3617_ | ~new_n6679_;
  assign new_n6689_ = ~new_n4829_ | ~new_n9074_;
  assign new_n6690_ = ~new_n4382_;
  assign new_n6691_ = ~new_n4828_ | ~new_n6678_;
  assign new_n6692_ = ~new_n3607_ | ~new_n4815_ | ~new_n6679_;
  assign new_n6693_ = ~new_n4825_ | ~new_n6687_;
  assign new_n6694_ = ~new_n4826_ | ~new_n4376_;
  assign new_n6695_ = ~new_n6660_ | ~new_n6691_;
  assign new_n6696_ = ~new_n6662_ | ~new_n4382_;
  assign new_n6697_ = ~new_n27132_ | ~new_n3512_;
  assign new_n6698_ = ~new_n6693_ | ~new_n4832_;
  assign new_n6699_ = ~new_n4421_;
  assign new_n6700_ = ~new_n5501_ | ~new_n4421_;
  assign new_n6701_ = ~new_n5496_ | ~new_n6698_;
  assign new_n6702_ = ~new_n6701_ | ~new_n6700_;
  assign new_n6703_ = ~new_n4383_;
  assign new_n6704_ = ~new_n4381_;
  assign new_n6705_ = ~new_n6690_ | ~new_n6678_;
  assign new_n6706_ = ~new_n3607_ | ~new_n6704_ | ~new_n6679_;
  assign new_n6707_ = ~new_n6703_ | ~new_n6705_;
  assign new_n6708_ = ~new_n27133_ | ~new_n3512_;
  assign new_n6709_ = ~new_n4835_ | ~new_n9138_ | ~new_n9137_;
  assign new_n6710_ = ~new_n4443_ | ~pi0177 | ~new_n4442_;
  assign new_n6711_ = ~new_n5501_ | ~new_n4381_;
  assign new_n6712_ = ~new_n5496_ | ~new_n6709_;
  assign new_n6713_ = ~new_n4836_ | ~new_n6712_;
  assign new_n6714_ = ~new_n4384_;
  assign new_n6715_ = ~new_n5497_ | ~new_n5764_;
  assign new_n6716_ = ~new_n4387_;
  assign new_n6717_ = ~new_n4386_;
  assign new_n6718_ = ~new_n3622_ | ~new_n4386_;
  assign new_n6719_ = ~new_n6687_ | ~new_n4250_;
  assign new_n6720_ = ~new_n6714_ | ~new_n4387_;
  assign new_n6721_ = ~new_n27127_ | ~new_n3512_;
  assign new_n6722_ = ~new_n6719_ | ~new_n4837_;
  assign new_n6723_ = ~new_n9141_ | ~pi0177 | ~new_n4442_;
  assign new_n6724_ = ~new_n6714_ | ~new_n5501_;
  assign new_n6725_ = ~new_n5496_ | ~new_n6722_;
  assign new_n6726_ = ~new_n4839_ | ~new_n6725_;
  assign new_n6727_ = ~new_n6716_ | ~new_n6717_;
  assign new_n6728_ = ~pi0311 | ~new_n3512_;
  assign new_n6729_ = ~new_n6728_ | ~new_n9150_ | ~new_n9149_;
  assign new_n6730_ = ~new_n5501_ | ~new_n4249_;
  assign new_n6731_ = ~new_n5496_ | ~new_n6729_;
  assign new_n6732_ = ~new_n9144_ | ~pi0177;
  assign new_n6733_ = ~new_n4840_ | ~new_n6731_;
  assign new_n6734_ = ~new_n23877_ | ~new_n3609_ | ~pi0178;
  assign new_n6735_ = ~new_n4389_;
  assign new_n6736_ = ~pi0175 | ~new_n4288_;
  assign new_n6737_ = ~new_n4389_ | ~new_n6736_;
  assign new_n6738_ = ~new_n5471_ | ~new_n4279_;
  assign new_n6739_ = ~new_n5803_ | ~new_n4427_;
  assign new_n6740_ = ~new_n4338_ | ~new_n6739_;
  assign new_n6741_ = ~new_n4339_ | ~new_n6740_;
  assign new_n6742_ = ~new_n5478_ | ~new_n6741_;
  assign new_n6743_ = ~new_n6738_ | ~new_n4298_;
  assign new_n6744_ = ~new_n5806_ | ~pi0175;
  assign new_n6745_ = ~new_n4841_ | ~new_n6742_;
  assign new_n6746_ = ~new_n6745_ | ~new_n4389_;
  assign new_n6747_ = ~pi0313 | ~new_n6737_;
  assign new_n6748_ = ~new_n5804_ | ~pi0175 | ~new_n4287_;
  assign new_n6749_ = ~new_n5478_ | ~new_n9155_;
  assign new_n6750_ = ~new_n4426_ | ~new_n6738_;
  assign new_n6751_ = ~new_n4842_ | ~new_n6749_;
  assign new_n6752_ = ~pi0175 | ~new_n4286_;
  assign new_n6753_ = ~new_n4389_ | ~new_n6752_;
  assign new_n6754_ = ~pi0314 | ~new_n6753_;
  assign new_n6755_ = ~new_n6751_ | ~new_n4389_;
  assign new_n6756_ = ~new_n5478_ | ~new_n4312_;
  assign new_n6757_ = ~pi0175 | ~new_n4285_;
  assign new_n6758_ = ~new_n6757_ | ~new_n6756_;
  assign new_n6759_ = ~pi0316 | ~new_n6758_;
  assign new_n6760_ = ~new_n3649_ | ~new_n5478_;
  assign new_n6761_ = ~new_n6738_ | ~new_n4297_;
  assign new_n6762_ = ~new_n6760_ | ~new_n6761_ | ~new_n6759_;
  assign new_n6763_ = ~pi0175 | ~new_n4284_;
  assign new_n6764_ = ~new_n4389_ | ~new_n6763_;
  assign new_n6765_ = ~pi0315 | ~new_n6764_;
  assign new_n6766_ = ~new_n6762_ | ~new_n4389_;
  assign new_n6767_ = ~new_n4390_;
  assign new_n6768_ = ~new_n6767_ | ~new_n4389_;
  assign new_n6769_ = ~pi0175 | ~new_n4284_;
  assign new_n6770_ = ~new_n5493_ | ~new_n6769_;
  assign new_n6771_ = ~new_n6770_ | ~new_n4389_;
  assign new_n6772_ = ~pi0316 | ~new_n6768_;
  assign new_n6773_ = ~new_n25105_ | ~new_n3619_ | ~new_n5450_;
  assign new_n6774_ = ~new_n23443_ | ~new_n5500_;
  assign new_n6775_ = ~new_n6774_ | ~new_n6773_;
  assign new_n6776_ = ~new_n27144_ | ~new_n5746_ | ~new_n3786_;
  assign new_n6777_ = ~new_n22636_ | ~new_n4230_;
  assign new_n6778_ = ~new_n6777_ | ~new_n6776_;
  assign new_n6779_ = ~new_n21854_ | ~new_n5644_;
  assign new_n6780_ = ~new_n6779_ | ~new_n9157_ | ~new_n9156_;
  assign new_n6781_ = ~new_n21624_ | ~new_n4258_ | ~new_n4264_;
  assign new_n6782_ = ~new_n5505_ | ~new_n27146_;
  assign new_n6783_ = ~new_n5504_ | ~new_n22221_;
  assign new_n6784_ = ~new_n5695_ | ~new_n6780_;
  assign new_n6785_ = ~new_n6783_ | ~new_n6784_ | ~new_n4843_ | ~new_n3671_;
  assign new_n6786_ = ~new_n3546_ | ~new_n6785_;
  assign new_n6787_ = ~new_n4404_;
  assign new_n6788_ = ~new_n22720_ | ~new_n3551_;
  assign new_n6789_ = ~new_n24243_ | ~new_n3549_;
  assign new_n6790_ = ~new_n25993_ | ~new_n4376_;
  assign new_n6791_ = ~new_n5454_ | ~new_n25808_;
  assign new_n6792_ = ~new_n5455_ | ~new_n26393_;
  assign new_n6793_ = ~new_n5456_ | ~pi0317;
  assign new_n6794_ = ~new_n5457_ | ~pi0317;
  assign new_n6795_ = ~new_n3510_ | ~new_n21858_;
  assign new_n6796_ = ~new_n3511_ | ~new_n21030_;
  assign new_n6797_ = ~pi0317 | ~new_n5458_;
  assign new_n6798_ = ~pi0317 | ~new_n3512_;
  assign new_n6799_ = ~pi0317 | ~new_n5459_;
  assign new_n6800_ = ~pi0317 | ~new_n5460_;
  assign new_n6801_ = ~new_n25625_ | ~new_n5461_;
  assign new_n6802_ = ~new_n24922_ | ~new_n3513_;
  assign new_n6803_ = ~new_n3514_ | ~new_n26178_;
  assign new_n6804_ = ~new_n3515_ | ~new_n23258_;
  assign new_n6805_ = ~new_n5462_ | ~new_n25440_;
  assign new_n6806_ = ~new_n3518_ | ~new_n23447_;
  assign new_n6807_ = ~new_n26719_ | ~new_n3516_;
  assign new_n6808_ = ~new_n6790_ | ~new_n4854_ | ~new_n4849_ | ~new_n4848_;
  assign new_n6809_ = ~pi0508 | ~new_n3558_;
  assign new_n6810_ = ~new_n5474_ | ~new_n6808_;
  assign new_n6811_ = ~new_n6787_ | ~pi0317;
  assign new_n6812_ = ~new_n22654_ | ~new_n3551_;
  assign new_n6813_ = ~new_n24195_ | ~new_n3549_;
  assign new_n6814_ = ~new_n26073_ | ~new_n4376_;
  assign new_n6815_ = ~new_n25888_ | ~new_n5454_;
  assign new_n6816_ = ~new_n26473_ | ~new_n5455_;
  assign new_n6817_ = ~new_n23880_ | ~new_n5456_;
  assign new_n6818_ = ~new_n27327_ | ~new_n5457_;
  assign new_n6819_ = ~new_n21938_ | ~new_n3510_;
  assign new_n6820_ = ~new_n21096_ | ~new_n3511_;
  assign new_n6821_ = ~new_n24743_ | ~new_n5458_;
  assign new_n6822_ = ~new_n27148_ | ~new_n3512_;
  assign new_n6823_ = ~new_n21675_ | ~new_n5459_;
  assign new_n6824_ = ~new_n25261_ | ~new_n5460_;
  assign new_n6825_ = ~new_n25702_ | ~new_n5461_;
  assign new_n6826_ = ~new_n24999_ | ~new_n3513_;
  assign new_n6827_ = ~new_n26258_ | ~new_n3514_;
  assign new_n6828_ = ~new_n23338_ | ~new_n3515_;
  assign new_n6829_ = ~new_n25520_ | ~new_n5462_;
  assign new_n6830_ = ~new_n23527_ | ~new_n3518_;
  assign new_n6831_ = ~new_n26652_ | ~new_n3516_;
  assign new_n6832_ = ~new_n6814_ | ~new_n4856_ | ~new_n4861_ | ~new_n6812_ | ~new_n4855_;
  assign new_n6833_ = ~new_n3558_ | ~pi0509;
  assign new_n6834_ = ~new_n5474_ | ~new_n6832_;
  assign new_n6835_ = ~new_n6787_ | ~pi0318;
  assign new_n6836_ = ~new_n22726_ | ~new_n3551_;
  assign new_n6837_ = ~new_n24252_ | ~new_n3549_;
  assign new_n6838_ = ~new_n26062_ | ~new_n4376_;
  assign new_n6839_ = ~new_n25877_ | ~new_n5454_;
  assign new_n6840_ = ~new_n26462_ | ~new_n5455_;
  assign new_n6841_ = ~new_n23947_ | ~new_n5456_;
  assign new_n6842_ = ~new_n27394_ | ~new_n5457_;
  assign new_n6843_ = ~new_n21927_ | ~new_n3510_;
  assign new_n6844_ = ~new_n21085_ | ~new_n3511_;
  assign new_n6845_ = ~new_n24810_ | ~new_n5458_;
  assign new_n6846_ = ~new_n27215_ | ~new_n3512_;
  assign new_n6847_ = ~new_n21742_ | ~new_n5459_;
  assign new_n6848_ = ~new_n25328_ | ~new_n5460_;
  assign new_n6849_ = ~new_n25626_ | ~new_n5461_;
  assign new_n6850_ = ~new_n24923_ | ~new_n3513_;
  assign new_n6851_ = ~new_n26247_ | ~new_n3514_;
  assign new_n6852_ = ~new_n23327_ | ~new_n3515_;
  assign new_n6853_ = ~new_n25509_ | ~new_n5462_;
  assign new_n6854_ = ~new_n23516_ | ~new_n3518_;
  assign new_n6855_ = ~new_n26725_ | ~new_n3516_;
  assign new_n6856_ = ~new_n6838_ | ~new_n4869_ | ~new_n4862_ | ~new_n6836_ | ~new_n4866_;
  assign new_n6857_ = ~new_n3558_ | ~pi0510;
  assign new_n6858_ = ~new_n5474_ | ~new_n6856_;
  assign new_n6859_ = ~pi0319 | ~new_n6787_;
  assign new_n6860_ = ~new_n22652_ | ~new_n3551_;
  assign new_n6861_ = ~new_n24250_ | ~new_n3549_;
  assign new_n6862_ = ~new_n26059_ | ~new_n4376_;
  assign new_n6863_ = ~new_n25874_ | ~new_n5454_;
  assign new_n6864_ = ~new_n26459_ | ~new_n5455_;
  assign new_n6865_ = ~new_n23944_ | ~new_n5456_;
  assign new_n6866_ = ~new_n27391_ | ~new_n5457_;
  assign new_n6867_ = ~new_n21924_ | ~new_n3510_;
  assign new_n6868_ = ~new_n21082_ | ~new_n3511_;
  assign new_n6869_ = ~new_n24807_ | ~new_n5458_;
  assign new_n6870_ = ~new_n27212_ | ~new_n3512_;
  assign new_n6871_ = ~new_n21739_ | ~new_n5459_;
  assign new_n6872_ = ~new_n25325_ | ~new_n5460_;
  assign new_n6873_ = ~new_n25714_ | ~new_n5461_;
  assign new_n6874_ = ~new_n25011_ | ~new_n3513_;
  assign new_n6875_ = ~new_n26244_ | ~new_n3514_;
  assign new_n6876_ = ~new_n23324_ | ~new_n3515_;
  assign new_n6877_ = ~new_n25506_ | ~new_n5462_;
  assign new_n6878_ = ~new_n23513_ | ~new_n3518_;
  assign new_n6879_ = ~new_n26650_ | ~new_n3516_;
  assign new_n6880_ = ~new_n4871_ | ~new_n4877_ | ~new_n4870_ | ~new_n4874_ | ~new_n6862_;
  assign new_n6881_ = ~new_n3558_ | ~pi0511;
  assign new_n6882_ = ~new_n5474_ | ~new_n6880_;
  assign new_n6883_ = ~pi0320 | ~new_n6787_;
  assign new_n6884_ = ~new_n22653_ | ~new_n3551_;
  assign new_n6885_ = ~new_n24249_ | ~new_n3549_;
  assign new_n6886_ = ~new_n26058_ | ~new_n4376_;
  assign new_n6887_ = ~new_n25873_ | ~new_n5454_;
  assign new_n6888_ = ~new_n26458_ | ~new_n5455_;
  assign new_n6889_ = ~new_n23943_ | ~new_n5456_;
  assign new_n6890_ = ~new_n27390_ | ~new_n5457_;
  assign new_n6891_ = ~new_n21923_ | ~new_n3510_;
  assign new_n6892_ = ~new_n21081_ | ~new_n3511_;
  assign new_n6893_ = ~new_n24806_ | ~new_n5458_;
  assign new_n6894_ = ~new_n27211_ | ~new_n3512_;
  assign new_n6895_ = ~new_n21738_ | ~new_n5459_;
  assign new_n6896_ = ~new_n25324_ | ~new_n5460_;
  assign new_n6897_ = ~new_n25689_ | ~new_n5461_;
  assign new_n6898_ = ~new_n24986_ | ~new_n3513_;
  assign new_n6899_ = ~new_n26243_ | ~new_n3514_;
  assign new_n6900_ = ~new_n23323_ | ~new_n3515_;
  assign new_n6901_ = ~new_n25505_ | ~new_n5462_;
  assign new_n6902_ = ~new_n23512_ | ~new_n3518_;
  assign new_n6903_ = ~new_n26723_ | ~new_n3516_;
  assign new_n6904_ = ~new_n6886_ | ~new_n4885_ | ~new_n4878_ | ~new_n6884_ | ~new_n4882_;
  assign new_n6905_ = ~new_n3558_ | ~pi0512;
  assign new_n6906_ = ~new_n5474_ | ~new_n6904_;
  assign new_n6907_ = ~pi0321 | ~new_n6787_;
  assign new_n6908_ = ~new_n22724_ | ~new_n3551_;
  assign new_n6909_ = ~new_n24248_ | ~new_n3549_;
  assign new_n6910_ = ~new_n26057_ | ~new_n4376_;
  assign new_n6911_ = ~new_n25872_ | ~new_n5454_;
  assign new_n6912_ = ~new_n26457_ | ~new_n5455_;
  assign new_n6913_ = ~new_n23942_ | ~new_n5456_;
  assign new_n6914_ = ~new_n27389_ | ~new_n5457_;
  assign new_n6915_ = ~new_n21922_ | ~new_n3510_;
  assign new_n6916_ = ~new_n21080_ | ~new_n3511_;
  assign new_n6917_ = ~new_n24805_ | ~new_n5458_;
  assign new_n6918_ = ~new_n27210_ | ~new_n3512_;
  assign new_n6919_ = ~new_n21737_ | ~new_n5459_;
  assign new_n6920_ = ~new_n25323_ | ~new_n5460_;
  assign new_n6921_ = ~new_n25688_ | ~new_n5461_;
  assign new_n6922_ = ~new_n24985_ | ~new_n3513_;
  assign new_n6923_ = ~new_n26242_ | ~new_n3514_;
  assign new_n6924_ = ~new_n23322_ | ~new_n3515_;
  assign new_n6925_ = ~new_n25504_ | ~new_n5462_;
  assign new_n6926_ = ~new_n23511_ | ~new_n3518_;
  assign new_n6927_ = ~new_n26651_ | ~new_n3516_;
  assign new_n6928_ = ~new_n4890_ | ~new_n4893_ | ~new_n4886_ | ~new_n6909_ | ~new_n6910_;
  assign new_n6929_ = ~new_n3558_ | ~pi0513;
  assign new_n6930_ = ~new_n5474_ | ~new_n6928_;
  assign new_n6931_ = ~pi0322 | ~new_n6787_;
  assign new_n6932_ = ~new_n22723_ | ~new_n3551_;
  assign new_n6933_ = ~new_n24247_ | ~new_n3549_;
  assign new_n6934_ = ~new_n26056_ | ~new_n4376_;
  assign new_n6935_ = ~new_n25871_ | ~new_n5454_;
  assign new_n6936_ = ~new_n26456_ | ~new_n5455_;
  assign new_n6937_ = ~new_n23941_ | ~new_n5456_;
  assign new_n6938_ = ~new_n27388_ | ~new_n5457_;
  assign new_n6939_ = ~new_n21921_ | ~new_n3510_;
  assign new_n6940_ = ~new_n21079_ | ~new_n3511_;
  assign new_n6941_ = ~new_n24804_ | ~new_n5458_;
  assign new_n6942_ = ~new_n27209_ | ~new_n3512_;
  assign new_n6943_ = ~new_n21736_ | ~new_n5459_;
  assign new_n6944_ = ~new_n25322_ | ~new_n5460_;
  assign new_n6945_ = ~new_n25687_ | ~new_n5461_;
  assign new_n6946_ = ~new_n24984_ | ~new_n3513_;
  assign new_n6947_ = ~new_n26241_ | ~new_n3514_;
  assign new_n6948_ = ~new_n23321_ | ~new_n3515_;
  assign new_n6949_ = ~new_n25503_ | ~new_n5462_;
  assign new_n6950_ = ~new_n23510_ | ~new_n3518_;
  assign new_n6951_ = ~new_n26722_ | ~new_n3516_;
  assign new_n6952_ = ~new_n4898_ | ~new_n4901_ | ~new_n4894_ | ~new_n6933_ | ~new_n6934_;
  assign new_n6953_ = ~new_n3558_ | ~pi0514;
  assign new_n6954_ = ~new_n5474_ | ~new_n6952_;
  assign new_n6955_ = ~pi0323 | ~new_n6787_;
  assign new_n6956_ = ~new_n22722_ | ~new_n3551_;
  assign new_n6957_ = ~new_n24246_ | ~new_n3549_;
  assign new_n6958_ = ~new_n26055_ | ~new_n4376_;
  assign new_n6959_ = ~new_n25870_ | ~new_n5454_;
  assign new_n6960_ = ~new_n26455_ | ~new_n5455_;
  assign new_n6961_ = ~new_n23940_ | ~new_n5456_;
  assign new_n6962_ = ~new_n27387_ | ~new_n5457_;
  assign new_n6963_ = ~new_n21920_ | ~new_n3510_;
  assign new_n6964_ = ~new_n21078_ | ~new_n3511_;
  assign new_n6965_ = ~new_n24803_ | ~new_n5458_;
  assign new_n6966_ = ~new_n27208_ | ~new_n3512_;
  assign new_n6967_ = ~new_n21735_ | ~new_n5459_;
  assign new_n6968_ = ~new_n25321_ | ~new_n5460_;
  assign new_n6969_ = ~new_n25686_ | ~new_n5461_;
  assign new_n6970_ = ~new_n24983_ | ~new_n3513_;
  assign new_n6971_ = ~new_n26240_ | ~new_n3514_;
  assign new_n6972_ = ~new_n23320_ | ~new_n3515_;
  assign new_n6973_ = ~new_n25502_ | ~new_n5462_;
  assign new_n6974_ = ~new_n23509_ | ~new_n3518_;
  assign new_n6975_ = ~new_n26721_ | ~new_n3516_;
  assign new_n6976_ = ~new_n4906_ | ~new_n4909_ | ~new_n4902_ | ~new_n6957_ | ~new_n6958_;
  assign new_n6977_ = ~new_n3558_ | ~pi0515;
  assign new_n6978_ = ~new_n5474_ | ~new_n6976_;
  assign new_n6979_ = ~pi0324 | ~new_n6787_;
  assign new_n6980_ = ~new_n22721_ | ~new_n3551_;
  assign new_n6981_ = ~new_n24245_ | ~new_n3549_;
  assign new_n6982_ = ~new_n26054_ | ~new_n4376_;
  assign new_n6983_ = ~new_n25869_ | ~new_n5454_;
  assign new_n6984_ = ~new_n26454_ | ~new_n5455_;
  assign new_n6985_ = ~new_n23939_ | ~new_n5456_;
  assign new_n6986_ = ~new_n27386_ | ~new_n5457_;
  assign new_n6987_ = ~new_n21919_ | ~new_n3510_;
  assign new_n6988_ = ~new_n21077_ | ~new_n3511_;
  assign new_n6989_ = ~new_n24802_ | ~new_n5458_;
  assign new_n6990_ = ~new_n27207_ | ~new_n3512_;
  assign new_n6991_ = ~new_n21734_ | ~new_n5459_;
  assign new_n6992_ = ~new_n25320_ | ~new_n5460_;
  assign new_n6993_ = ~new_n25685_ | ~new_n5461_;
  assign new_n6994_ = ~new_n24982_ | ~new_n3513_;
  assign new_n6995_ = ~new_n26239_ | ~new_n3514_;
  assign new_n6996_ = ~new_n23319_ | ~new_n3515_;
  assign new_n6997_ = ~new_n25501_ | ~new_n5462_;
  assign new_n6998_ = ~new_n23508_ | ~new_n3518_;
  assign new_n6999_ = ~new_n26720_ | ~new_n3516_;
  assign new_n7000_ = ~new_n4913_ | ~new_n4916_ | ~new_n4910_ | ~new_n6981_ | ~new_n6982_;
  assign new_n7001_ = ~new_n3558_ | ~pi0516;
  assign new_n7002_ = ~new_n5474_ | ~new_n7000_;
  assign new_n7003_ = ~pi0325 | ~new_n6787_;
  assign new_n7004_ = ~new_n22741_ | ~new_n3551_;
  assign new_n7005_ = ~new_n24244_ | ~new_n3549_;
  assign new_n7006_ = ~new_n26053_ | ~new_n4376_;
  assign new_n7007_ = ~new_n25868_ | ~new_n5454_;
  assign new_n7008_ = ~new_n26453_ | ~new_n5455_;
  assign new_n7009_ = ~new_n23938_ | ~new_n5456_;
  assign new_n7010_ = ~new_n27385_ | ~new_n5457_;
  assign new_n7011_ = ~new_n21918_ | ~new_n3510_;
  assign new_n7012_ = ~new_n21076_ | ~new_n3511_;
  assign new_n7013_ = ~new_n24801_ | ~new_n5458_;
  assign new_n7014_ = ~new_n27206_ | ~new_n3512_;
  assign new_n7015_ = ~new_n21733_ | ~new_n5459_;
  assign new_n7016_ = ~new_n25319_ | ~new_n5460_;
  assign new_n7017_ = ~new_n25684_ | ~new_n5461_;
  assign new_n7018_ = ~new_n24981_ | ~new_n3513_;
  assign new_n7019_ = ~new_n26238_ | ~new_n3514_;
  assign new_n7020_ = ~new_n23318_ | ~new_n3515_;
  assign new_n7021_ = ~new_n25500_ | ~new_n5462_;
  assign new_n7022_ = ~new_n23507_ | ~new_n3518_;
  assign new_n7023_ = ~new_n26741_ | ~new_n3516_;
  assign new_n7024_ = ~new_n4920_ | ~new_n4923_ | ~new_n4917_ | ~new_n7005_ | ~new_n7006_;
  assign new_n7025_ = ~new_n3558_ | ~pi0517;
  assign new_n7026_ = ~new_n5474_ | ~new_n7024_;
  assign new_n7027_ = ~pi0326 | ~new_n6787_;
  assign new_n7028_ = ~new_n22639_ | ~new_n3551_;
  assign new_n7029_ = ~new_n24267_ | ~new_n3549_;
  assign new_n7030_ = ~new_n26083_ | ~new_n4376_;
  assign new_n7031_ = ~new_n25898_ | ~new_n5454_;
  assign new_n7032_ = ~new_n26483_ | ~new_n5455_;
  assign new_n7033_ = ~new_n23967_ | ~new_n5456_;
  assign new_n7034_ = ~new_n27414_ | ~new_n5457_;
  assign new_n7035_ = ~new_n21948_ | ~new_n3510_;
  assign new_n7036_ = ~new_n21106_ | ~new_n3511_;
  assign new_n7037_ = ~new_n24830_ | ~new_n5458_;
  assign new_n7038_ = ~new_n27235_ | ~new_n3512_;
  assign new_n7039_ = ~new_n21762_ | ~new_n5459_;
  assign new_n7040_ = ~new_n25348_ | ~new_n5460_;
  assign new_n7041_ = ~new_n25712_ | ~new_n5461_;
  assign new_n7042_ = ~new_n25009_ | ~new_n3513_;
  assign new_n7043_ = ~new_n26268_ | ~new_n3514_;
  assign new_n7044_ = ~new_n23348_ | ~new_n3515_;
  assign new_n7045_ = ~new_n25530_ | ~new_n5462_;
  assign new_n7046_ = ~new_n23537_ | ~new_n3518_;
  assign new_n7047_ = ~new_n26637_ | ~new_n3516_;
  assign new_n7048_ = ~new_n7030_ | ~new_n4924_ | ~new_n4930_ | ~new_n7028_ | ~new_n4927_;
  assign new_n7049_ = ~new_n3558_ | ~pi0518;
  assign new_n7050_ = ~new_n5474_ | ~new_n7048_;
  assign new_n7051_ = ~pi0327 | ~new_n6787_;
  assign new_n7052_ = ~new_n22719_ | ~new_n3551_;
  assign new_n7053_ = ~new_n24266_ | ~new_n3549_;
  assign new_n7054_ = ~new_n26082_ | ~new_n4376_;
  assign new_n7055_ = ~new_n25897_ | ~new_n5454_;
  assign new_n7056_ = ~new_n26482_ | ~new_n5455_;
  assign new_n7057_ = ~new_n23966_ | ~new_n5456_;
  assign new_n7058_ = ~new_n27413_ | ~new_n5457_;
  assign new_n7059_ = ~new_n21947_ | ~new_n3510_;
  assign new_n7060_ = ~new_n21105_ | ~new_n3511_;
  assign new_n7061_ = ~new_n24829_ | ~new_n5458_;
  assign new_n7062_ = ~new_n27234_ | ~new_n3512_;
  assign new_n7063_ = ~new_n21761_ | ~new_n5459_;
  assign new_n7064_ = ~new_n25347_ | ~new_n5460_;
  assign new_n7065_ = ~new_n25711_ | ~new_n5461_;
  assign new_n7066_ = ~new_n25008_ | ~new_n3513_;
  assign new_n7067_ = ~new_n26267_ | ~new_n3514_;
  assign new_n7068_ = ~new_n23347_ | ~new_n3515_;
  assign new_n7069_ = ~new_n25529_ | ~new_n5462_;
  assign new_n7070_ = ~new_n23536_ | ~new_n3518_;
  assign new_n7071_ = ~new_n26718_ | ~new_n3516_;
  assign new_n7072_ = ~new_n7054_ | ~new_n4937_ | ~new_n4931_ | ~new_n7052_ | ~new_n4934_;
  assign new_n7073_ = ~new_n3558_ | ~pi0519;
  assign new_n7074_ = ~new_n5474_ | ~new_n7072_;
  assign new_n7075_ = ~pi0328 | ~new_n6787_;
  assign new_n7076_ = ~new_n22640_ | ~new_n3551_;
  assign new_n7077_ = ~new_n24265_ | ~new_n3549_;
  assign new_n7078_ = ~new_n26081_ | ~new_n4376_;
  assign new_n7079_ = ~new_n25896_ | ~new_n5454_;
  assign new_n7080_ = ~new_n26481_ | ~new_n5455_;
  assign new_n7081_ = ~new_n23965_ | ~new_n5456_;
  assign new_n7082_ = ~new_n27412_ | ~new_n5457_;
  assign new_n7083_ = ~new_n21946_ | ~new_n3510_;
  assign new_n7084_ = ~new_n21104_ | ~new_n3511_;
  assign new_n7085_ = ~new_n24828_ | ~new_n5458_;
  assign new_n7086_ = ~new_n27233_ | ~new_n3512_;
  assign new_n7087_ = ~new_n21760_ | ~new_n5459_;
  assign new_n7088_ = ~new_n25346_ | ~new_n5460_;
  assign new_n7089_ = ~new_n25710_ | ~new_n5461_;
  assign new_n7090_ = ~new_n25007_ | ~new_n3513_;
  assign new_n7091_ = ~new_n26266_ | ~new_n3514_;
  assign new_n7092_ = ~new_n23346_ | ~new_n3515_;
  assign new_n7093_ = ~new_n25528_ | ~new_n5462_;
  assign new_n7094_ = ~new_n23535_ | ~new_n3518_;
  assign new_n7095_ = ~new_n26638_ | ~new_n3516_;
  assign new_n7096_ = ~new_n4941_ | ~new_n4944_ | ~new_n4938_ | ~new_n7077_ | ~new_n7078_;
  assign new_n7097_ = ~new_n3558_ | ~pi0520;
  assign new_n7098_ = ~new_n5474_ | ~new_n7096_;
  assign new_n7099_ = ~pi0329 | ~new_n6787_;
  assign new_n7100_ = ~new_n22641_ | ~new_n3551_;
  assign new_n7101_ = ~new_n24189_ | ~new_n3549_;
  assign new_n7102_ = ~new_n26080_ | ~new_n4376_;
  assign new_n7103_ = ~new_n25895_ | ~new_n5454_;
  assign new_n7104_ = ~new_n26480_ | ~new_n5455_;
  assign new_n7105_ = ~new_n23964_ | ~new_n5456_;
  assign new_n7106_ = ~new_n27411_ | ~new_n5457_;
  assign new_n7107_ = ~new_n21945_ | ~new_n3510_;
  assign new_n7108_ = ~new_n21103_ | ~new_n3511_;
  assign new_n7109_ = ~new_n24827_ | ~new_n5458_;
  assign new_n7110_ = ~new_n27232_ | ~new_n3512_;
  assign new_n7111_ = ~new_n21759_ | ~new_n5459_;
  assign new_n7112_ = ~new_n25345_ | ~new_n5460_;
  assign new_n7113_ = ~new_n25709_ | ~new_n5461_;
  assign new_n7114_ = ~new_n25006_ | ~new_n3513_;
  assign new_n7115_ = ~new_n26265_ | ~new_n3514_;
  assign new_n7116_ = ~new_n23345_ | ~new_n3515_;
  assign new_n7117_ = ~new_n25527_ | ~new_n5462_;
  assign new_n7118_ = ~new_n23534_ | ~new_n3518_;
  assign new_n7119_ = ~new_n26639_ | ~new_n3516_;
  assign new_n7120_ = ~new_n4948_ | ~new_n4951_ | ~new_n4945_ | ~new_n7101_ | ~new_n7102_;
  assign new_n7121_ = ~new_n3558_ | ~pi0521;
  assign new_n7122_ = ~new_n5474_ | ~new_n7120_;
  assign new_n7123_ = ~pi0330 | ~new_n6787_;
  assign new_n7124_ = ~new_n22718_ | ~new_n3551_;
  assign new_n7125_ = ~new_n24264_ | ~new_n3549_;
  assign new_n7126_ = ~new_n26079_ | ~new_n4376_;
  assign new_n7127_ = ~new_n25894_ | ~new_n5454_;
  assign new_n7128_ = ~new_n26479_ | ~new_n5455_;
  assign new_n7129_ = ~new_n23963_ | ~new_n5456_;
  assign new_n7130_ = ~new_n27410_ | ~new_n5457_;
  assign new_n7131_ = ~new_n21944_ | ~new_n3510_;
  assign new_n7132_ = ~new_n21102_ | ~new_n3511_;
  assign new_n7133_ = ~new_n24826_ | ~new_n5458_;
  assign new_n7134_ = ~new_n27231_ | ~new_n3512_;
  assign new_n7135_ = ~new_n21758_ | ~new_n5459_;
  assign new_n7136_ = ~new_n25344_ | ~new_n5460_;
  assign new_n7137_ = ~new_n25708_ | ~new_n5461_;
  assign new_n7138_ = ~new_n25005_ | ~new_n3513_;
  assign new_n7139_ = ~new_n26264_ | ~new_n3514_;
  assign new_n7140_ = ~new_n23344_ | ~new_n3515_;
  assign new_n7141_ = ~new_n25526_ | ~new_n5462_;
  assign new_n7142_ = ~new_n23533_ | ~new_n3518_;
  assign new_n7143_ = ~new_n26717_ | ~new_n3516_;
  assign new_n7144_ = ~new_n4958_ | ~new_n4955_;
  assign new_n7145_ = ~new_n3558_ | ~pi0522;
  assign new_n7146_ = ~new_n5474_ | ~new_n7144_;
  assign new_n7147_ = ~pi0331 | ~new_n6787_;
  assign new_n7148_ = ~new_n22642_ | ~new_n3551_;
  assign new_n7149_ = ~new_n24263_ | ~new_n3549_;
  assign new_n7150_ = ~new_n26078_ | ~new_n4376_;
  assign new_n7151_ = ~new_n25893_ | ~new_n5454_;
  assign new_n7152_ = ~new_n26478_ | ~new_n5455_;
  assign new_n7153_ = ~new_n23962_ | ~new_n5456_;
  assign new_n7154_ = ~new_n27409_ | ~new_n5457_;
  assign new_n7155_ = ~new_n21943_ | ~new_n3510_;
  assign new_n7156_ = ~new_n21101_ | ~new_n3511_;
  assign new_n7157_ = ~new_n24825_ | ~new_n5458_;
  assign new_n7158_ = ~new_n27230_ | ~new_n3512_;
  assign new_n7159_ = ~new_n21757_ | ~new_n5459_;
  assign new_n7160_ = ~new_n25343_ | ~new_n5460_;
  assign new_n7161_ = ~new_n25707_ | ~new_n5461_;
  assign new_n7162_ = ~new_n25004_ | ~new_n3513_;
  assign new_n7163_ = ~new_n26263_ | ~new_n3514_;
  assign new_n7164_ = ~new_n23343_ | ~new_n3515_;
  assign new_n7165_ = ~new_n25525_ | ~new_n5462_;
  assign new_n7166_ = ~new_n23532_ | ~new_n3518_;
  assign new_n7167_ = ~new_n26640_ | ~new_n3516_;
  assign new_n7168_ = ~new_n4966_ | ~new_n4963_;
  assign new_n7169_ = ~new_n3558_ | ~pi0523;
  assign new_n7170_ = ~new_n5474_ | ~new_n7168_;
  assign new_n7171_ = ~pi0332 | ~new_n6787_;
  assign new_n7172_ = ~new_n22717_ | ~new_n3551_;
  assign new_n7173_ = ~new_n24262_ | ~new_n3549_;
  assign new_n7174_ = ~new_n26077_ | ~new_n4376_;
  assign new_n7175_ = ~new_n25892_ | ~new_n5454_;
  assign new_n7176_ = ~new_n26477_ | ~new_n5455_;
  assign new_n7177_ = ~new_n23961_ | ~new_n5456_;
  assign new_n7178_ = ~new_n27408_ | ~new_n5457_;
  assign new_n7179_ = ~new_n21942_ | ~new_n3510_;
  assign new_n7180_ = ~new_n21100_ | ~new_n3511_;
  assign new_n7181_ = ~new_n24824_ | ~new_n5458_;
  assign new_n7182_ = ~new_n27229_ | ~new_n3512_;
  assign new_n7183_ = ~new_n21756_ | ~new_n5459_;
  assign new_n7184_ = ~new_n25342_ | ~new_n5460_;
  assign new_n7185_ = ~new_n25706_ | ~new_n5461_;
  assign new_n7186_ = ~new_n25003_ | ~new_n3513_;
  assign new_n7187_ = ~new_n26262_ | ~new_n3514_;
  assign new_n7188_ = ~new_n23342_ | ~new_n3515_;
  assign new_n7189_ = ~new_n25524_ | ~new_n5462_;
  assign new_n7190_ = ~new_n23531_ | ~new_n3518_;
  assign new_n7191_ = ~new_n26716_ | ~new_n3516_;
  assign new_n7192_ = ~new_n7174_ | ~new_n4974_ | ~new_n4968_ | ~new_n7172_ | ~new_n4971_;
  assign new_n7193_ = ~new_n3558_ | ~pi0524;
  assign new_n7194_ = ~new_n5474_ | ~new_n7192_;
  assign new_n7195_ = ~pi0333 | ~new_n6787_;
  assign new_n7196_ = ~new_n22643_ | ~new_n3551_;
  assign new_n7197_ = ~new_n24190_ | ~new_n3549_;
  assign new_n7198_ = ~new_n26076_ | ~new_n4376_;
  assign new_n7199_ = ~new_n25891_ | ~new_n5454_;
  assign new_n7200_ = ~new_n26476_ | ~new_n5455_;
  assign new_n7201_ = ~new_n23960_ | ~new_n5456_;
  assign new_n7202_ = ~new_n27407_ | ~new_n5457_;
  assign new_n7203_ = ~new_n21941_ | ~new_n3510_;
  assign new_n7204_ = ~new_n21099_ | ~new_n3511_;
  assign new_n7205_ = ~new_n24823_ | ~new_n5458_;
  assign new_n7206_ = ~new_n27228_ | ~new_n3512_;
  assign new_n7207_ = ~new_n21755_ | ~new_n5459_;
  assign new_n7208_ = ~new_n25341_ | ~new_n5460_;
  assign new_n7209_ = ~new_n25705_ | ~new_n5461_;
  assign new_n7210_ = ~new_n25002_ | ~new_n3513_;
  assign new_n7211_ = ~new_n26261_ | ~new_n3514_;
  assign new_n7212_ = ~new_n23341_ | ~new_n3515_;
  assign new_n7213_ = ~new_n25523_ | ~new_n5462_;
  assign new_n7214_ = ~new_n23530_ | ~new_n3518_;
  assign new_n7215_ = ~new_n26641_ | ~new_n3516_;
  assign new_n7216_ = ~new_n7198_ | ~new_n4976_ | ~new_n4980_ | ~new_n7196_ | ~new_n4975_;
  assign new_n7217_ = ~new_n3558_ | ~pi0525;
  assign new_n7218_ = ~new_n5474_ | ~new_n7216_;
  assign new_n7219_ = ~pi0334 | ~new_n6787_;
  assign new_n7220_ = ~new_n22716_ | ~new_n3551_;
  assign new_n7221_ = ~new_n24261_ | ~new_n3549_;
  assign new_n7222_ = ~new_n26075_ | ~new_n4376_;
  assign new_n7223_ = ~new_n25890_ | ~new_n5454_;
  assign new_n7224_ = ~new_n26475_ | ~new_n5455_;
  assign new_n7225_ = ~new_n23959_ | ~new_n5456_;
  assign new_n7226_ = ~new_n27406_ | ~new_n5457_;
  assign new_n7227_ = ~new_n21940_ | ~new_n3510_;
  assign new_n7228_ = ~new_n21098_ | ~new_n3511_;
  assign new_n7229_ = ~new_n24822_ | ~new_n5458_;
  assign new_n7230_ = ~new_n27227_ | ~new_n3512_;
  assign new_n7231_ = ~new_n21754_ | ~new_n5459_;
  assign new_n7232_ = ~new_n25340_ | ~new_n5460_;
  assign new_n7233_ = ~new_n25704_ | ~new_n5461_;
  assign new_n7234_ = ~new_n25001_ | ~new_n3513_;
  assign new_n7235_ = ~new_n26260_ | ~new_n3514_;
  assign new_n7236_ = ~new_n23340_ | ~new_n3515_;
  assign new_n7237_ = ~new_n25522_ | ~new_n5462_;
  assign new_n7238_ = ~new_n23529_ | ~new_n3518_;
  assign new_n7239_ = ~new_n26715_ | ~new_n3516_;
  assign new_n7240_ = ~new_n7222_ | ~new_n4987_ | ~new_n4981_ | ~new_n7220_ | ~new_n4984_;
  assign new_n7241_ = ~new_n3558_ | ~pi0526;
  assign new_n7242_ = ~new_n5474_ | ~new_n7240_;
  assign new_n7243_ = ~pi0335 | ~new_n6787_;
  assign new_n7244_ = ~new_n22644_ | ~new_n3551_;
  assign new_n7245_ = ~new_n24260_ | ~new_n3549_;
  assign new_n7246_ = ~new_n26074_ | ~new_n4376_;
  assign new_n7247_ = ~new_n25889_ | ~new_n5454_;
  assign new_n7248_ = ~new_n26474_ | ~new_n5455_;
  assign new_n7249_ = ~new_n23958_ | ~new_n5456_;
  assign new_n7250_ = ~new_n27405_ | ~new_n5457_;
  assign new_n7251_ = ~new_n21939_ | ~new_n3510_;
  assign new_n7252_ = ~new_n21097_ | ~new_n3511_;
  assign new_n7253_ = ~new_n24821_ | ~new_n5458_;
  assign new_n7254_ = ~new_n27226_ | ~new_n3512_;
  assign new_n7255_ = ~new_n21753_ | ~new_n5459_;
  assign new_n7256_ = ~new_n25339_ | ~new_n5460_;
  assign new_n7257_ = ~new_n25703_ | ~new_n5461_;
  assign new_n7258_ = ~new_n25000_ | ~new_n3513_;
  assign new_n7259_ = ~new_n26259_ | ~new_n3514_;
  assign new_n7260_ = ~new_n23339_ | ~new_n3515_;
  assign new_n7261_ = ~new_n25521_ | ~new_n5462_;
  assign new_n7262_ = ~new_n23528_ | ~new_n3518_;
  assign new_n7263_ = ~new_n26642_ | ~new_n3516_;
  assign new_n7264_ = ~new_n7246_ | ~new_n4989_ | ~new_n4993_ | ~new_n7244_ | ~new_n4988_;
  assign new_n7265_ = ~new_n3558_ | ~pi0527;
  assign new_n7266_ = ~new_n5474_ | ~new_n7264_;
  assign new_n7267_ = ~pi0336 | ~new_n6787_;
  assign new_n7268_ = ~new_n22645_ | ~new_n3551_;
  assign new_n7269_ = ~new_n24191_ | ~new_n3549_;
  assign new_n7270_ = ~new_n26072_ | ~new_n4376_;
  assign new_n7271_ = ~new_n25887_ | ~new_n5454_;
  assign new_n7272_ = ~new_n26472_ | ~new_n5455_;
  assign new_n7273_ = ~new_n23957_ | ~new_n5456_;
  assign new_n7274_ = ~new_n27404_ | ~new_n5457_;
  assign new_n7275_ = ~new_n21937_ | ~new_n3510_;
  assign new_n7276_ = ~new_n21095_ | ~new_n3511_;
  assign new_n7277_ = ~new_n24820_ | ~new_n5458_;
  assign new_n7278_ = ~new_n27225_ | ~new_n3512_;
  assign new_n7279_ = ~new_n21752_ | ~new_n5459_;
  assign new_n7280_ = ~new_n25338_ | ~new_n5460_;
  assign new_n7281_ = ~new_n25701_ | ~new_n5461_;
  assign new_n7282_ = ~new_n24998_ | ~new_n3513_;
  assign new_n7283_ = ~new_n26257_ | ~new_n3514_;
  assign new_n7284_ = ~new_n23337_ | ~new_n3515_;
  assign new_n7285_ = ~new_n25519_ | ~new_n5462_;
  assign new_n7286_ = ~new_n23526_ | ~new_n3518_;
  assign new_n7287_ = ~new_n26643_ | ~new_n3516_;
  assign new_n7288_ = ~new_n7269_ | ~new_n4997_;
  assign new_n7289_ = ~new_n3558_ | ~pi0528;
  assign new_n7290_ = ~new_n5474_ | ~new_n7288_;
  assign new_n7291_ = ~pi0337 | ~new_n6787_;
  assign new_n7292_ = ~new_n22646_ | ~new_n3551_;
  assign new_n7293_ = ~new_n24259_ | ~new_n3549_;
  assign new_n7294_ = ~new_n26071_ | ~new_n4376_;
  assign new_n7295_ = ~new_n25886_ | ~new_n5454_;
  assign new_n7296_ = ~new_n26471_ | ~new_n5455_;
  assign new_n7297_ = ~new_n23956_ | ~new_n5456_;
  assign new_n7298_ = ~new_n27403_ | ~new_n5457_;
  assign new_n7299_ = ~new_n21936_ | ~new_n3510_;
  assign new_n7300_ = ~new_n21094_ | ~new_n3511_;
  assign new_n7301_ = ~new_n24819_ | ~new_n5458_;
  assign new_n7302_ = ~new_n27224_ | ~new_n3512_;
  assign new_n7303_ = ~new_n21751_ | ~new_n5459_;
  assign new_n7304_ = ~new_n25337_ | ~new_n5460_;
  assign new_n7305_ = ~new_n25700_ | ~new_n5461_;
  assign new_n7306_ = ~new_n24997_ | ~new_n3513_;
  assign new_n7307_ = ~new_n26256_ | ~new_n3514_;
  assign new_n7308_ = ~new_n23336_ | ~new_n3515_;
  assign new_n7309_ = ~new_n25518_ | ~new_n5462_;
  assign new_n7310_ = ~new_n23525_ | ~new_n3518_;
  assign new_n7311_ = ~new_n26644_ | ~new_n3516_;
  assign new_n7312_ = ~new_n7293_ | ~new_n5005_;
  assign new_n7313_ = ~new_n3558_ | ~pi0529;
  assign new_n7314_ = ~new_n5474_ | ~new_n7312_;
  assign new_n7315_ = ~pi0338 | ~new_n6787_;
  assign new_n7316_ = ~new_n22715_ | ~new_n3551_;
  assign new_n7317_ = ~new_n24258_ | ~new_n3549_;
  assign new_n7318_ = ~new_n26070_ | ~new_n4376_;
  assign new_n7319_ = ~new_n25885_ | ~new_n5454_;
  assign new_n7320_ = ~new_n26470_ | ~new_n5455_;
  assign new_n7321_ = ~new_n23955_ | ~new_n5456_;
  assign new_n7322_ = ~new_n27402_ | ~new_n5457_;
  assign new_n7323_ = ~new_n21935_ | ~new_n3510_;
  assign new_n7324_ = ~new_n21093_ | ~new_n3511_;
  assign new_n7325_ = ~new_n24818_ | ~new_n5458_;
  assign new_n7326_ = ~new_n27223_ | ~new_n3512_;
  assign new_n7327_ = ~new_n21750_ | ~new_n5459_;
  assign new_n7328_ = ~new_n25336_ | ~new_n5460_;
  assign new_n7329_ = ~new_n25699_ | ~new_n5461_;
  assign new_n7330_ = ~new_n24996_ | ~new_n3513_;
  assign new_n7331_ = ~new_n26255_ | ~new_n3514_;
  assign new_n7332_ = ~new_n23335_ | ~new_n3515_;
  assign new_n7333_ = ~new_n25517_ | ~new_n5462_;
  assign new_n7334_ = ~new_n23524_ | ~new_n3518_;
  assign new_n7335_ = ~new_n26714_ | ~new_n3516_;
  assign new_n7336_ = ~new_n5018_ | ~new_n5013_;
  assign new_n7337_ = ~new_n3558_ | ~pi0530;
  assign new_n7338_ = ~new_n5474_ | ~new_n7336_;
  assign new_n7339_ = ~pi0339 | ~new_n6787_;
  assign new_n7340_ = ~new_n22647_ | ~new_n3551_;
  assign new_n7341_ = ~new_n24257_ | ~new_n3549_;
  assign new_n7342_ = ~new_n26069_ | ~new_n4376_;
  assign new_n7343_ = ~new_n25884_ | ~new_n5454_;
  assign new_n7344_ = ~new_n26469_ | ~new_n5455_;
  assign new_n7345_ = ~new_n23954_ | ~new_n5456_;
  assign new_n7346_ = ~new_n27401_ | ~new_n5457_;
  assign new_n7347_ = ~new_n21934_ | ~new_n3510_;
  assign new_n7348_ = ~new_n21092_ | ~new_n3511_;
  assign new_n7349_ = ~new_n24817_ | ~new_n5458_;
  assign new_n7350_ = ~new_n27222_ | ~new_n3512_;
  assign new_n7351_ = ~new_n21749_ | ~new_n5459_;
  assign new_n7352_ = ~new_n25335_ | ~new_n5460_;
  assign new_n7353_ = ~new_n25698_ | ~new_n5461_;
  assign new_n7354_ = ~new_n24995_ | ~new_n3513_;
  assign new_n7355_ = ~new_n26254_ | ~new_n3514_;
  assign new_n7356_ = ~new_n23334_ | ~new_n3515_;
  assign new_n7357_ = ~new_n25516_ | ~new_n5462_;
  assign new_n7358_ = ~new_n23523_ | ~new_n3518_;
  assign new_n7359_ = ~new_n26645_ | ~new_n3516_;
  assign new_n7360_ = ~new_n5028_ | ~new_n5023_;
  assign new_n7361_ = ~new_n3558_ | ~pi0531;
  assign new_n7362_ = ~new_n5474_ | ~new_n7360_;
  assign new_n7363_ = ~pi0340 | ~new_n6787_;
  assign new_n7364_ = ~new_n22714_ | ~new_n3551_;
  assign new_n7365_ = ~new_n24256_ | ~new_n3549_;
  assign new_n7366_ = ~new_n26068_ | ~new_n4376_;
  assign new_n7367_ = ~new_n25883_ | ~new_n5454_;
  assign new_n7368_ = ~new_n26468_ | ~new_n5455_;
  assign new_n7369_ = ~new_n23953_ | ~new_n5456_;
  assign new_n7370_ = ~new_n27400_ | ~new_n5457_;
  assign new_n7371_ = ~new_n21933_ | ~new_n3510_;
  assign new_n7372_ = ~new_n21091_ | ~new_n3511_;
  assign new_n7373_ = ~new_n24816_ | ~new_n5458_;
  assign new_n7374_ = ~new_n27221_ | ~new_n3512_;
  assign new_n7375_ = ~new_n21748_ | ~new_n5459_;
  assign new_n7376_ = ~new_n25334_ | ~new_n5460_;
  assign new_n7377_ = ~new_n25697_ | ~new_n5461_;
  assign new_n7378_ = ~new_n24994_ | ~new_n3513_;
  assign new_n7379_ = ~new_n26253_ | ~new_n3514_;
  assign new_n7380_ = ~new_n23333_ | ~new_n3515_;
  assign new_n7381_ = ~new_n25515_ | ~new_n5462_;
  assign new_n7382_ = ~new_n23522_ | ~new_n3518_;
  assign new_n7383_ = ~new_n26713_ | ~new_n3516_;
  assign new_n7384_ = ~new_n5038_ | ~new_n5033_;
  assign new_n7385_ = ~new_n3558_ | ~pi0532;
  assign new_n7386_ = ~new_n5474_ | ~new_n7384_;
  assign new_n7387_ = ~pi0341 | ~new_n6787_;
  assign new_n7388_ = ~new_n22648_ | ~new_n3551_;
  assign new_n7389_ = ~new_n24255_ | ~new_n3549_;
  assign new_n7390_ = ~new_n26067_ | ~new_n4376_;
  assign new_n7391_ = ~new_n25882_ | ~new_n5454_;
  assign new_n7392_ = ~new_n26467_ | ~new_n5455_;
  assign new_n7393_ = ~new_n23952_ | ~new_n5456_;
  assign new_n7394_ = ~new_n27399_ | ~new_n5457_;
  assign new_n7395_ = ~new_n21932_ | ~new_n3510_;
  assign new_n7396_ = ~new_n21090_ | ~new_n3511_;
  assign new_n7397_ = ~new_n24815_ | ~new_n5458_;
  assign new_n7398_ = ~new_n27220_ | ~new_n3512_;
  assign new_n7399_ = ~new_n21747_ | ~new_n5459_;
  assign new_n7400_ = ~new_n25333_ | ~new_n5460_;
  assign new_n7401_ = ~new_n25696_ | ~new_n5461_;
  assign new_n7402_ = ~new_n24993_ | ~new_n3513_;
  assign new_n7403_ = ~new_n26252_ | ~new_n3514_;
  assign new_n7404_ = ~new_n23332_ | ~new_n3515_;
  assign new_n7405_ = ~new_n25514_ | ~new_n5462_;
  assign new_n7406_ = ~new_n23521_ | ~new_n3518_;
  assign new_n7407_ = ~new_n26646_ | ~new_n3516_;
  assign new_n7408_ = ~new_n5048_ | ~new_n5043_;
  assign new_n7409_ = ~new_n3558_ | ~pi0533;
  assign new_n7410_ = ~new_n5474_ | ~new_n7408_;
  assign new_n7411_ = ~pi0342 | ~new_n6787_;
  assign new_n7412_ = ~new_n22649_ | ~new_n3551_;
  assign new_n7413_ = ~new_n24192_ | ~new_n3549_;
  assign new_n7414_ = ~new_n26066_ | ~new_n4376_;
  assign new_n7415_ = ~new_n25881_ | ~new_n5454_;
  assign new_n7416_ = ~new_n26466_ | ~new_n5455_;
  assign new_n7417_ = ~new_n23951_ | ~new_n5456_;
  assign new_n7418_ = ~new_n27398_ | ~new_n5457_;
  assign new_n7419_ = ~new_n21931_ | ~new_n3510_;
  assign new_n7420_ = ~new_n21089_ | ~new_n3511_;
  assign new_n7421_ = ~new_n24814_ | ~new_n5458_;
  assign new_n7422_ = ~new_n27219_ | ~new_n3512_;
  assign new_n7423_ = ~new_n21746_ | ~new_n5459_;
  assign new_n7424_ = ~new_n25332_ | ~new_n5460_;
  assign new_n7425_ = ~new_n25695_ | ~new_n5461_;
  assign new_n7426_ = ~new_n24992_ | ~new_n3513_;
  assign new_n7427_ = ~new_n26251_ | ~new_n3514_;
  assign new_n7428_ = ~new_n23331_ | ~new_n3515_;
  assign new_n7429_ = ~new_n25513_ | ~new_n5462_;
  assign new_n7430_ = ~new_n23520_ | ~new_n3518_;
  assign new_n7431_ = ~new_n26647_ | ~new_n3516_;
  assign new_n7432_ = ~new_n5050_ | ~new_n5058_ | ~new_n5053_ | ~new_n5051_ | ~new_n7414_;
  assign new_n7433_ = ~new_n3558_ | ~pi0534;
  assign new_n7434_ = ~new_n5474_ | ~new_n7432_;
  assign new_n7435_ = ~pi0343 | ~new_n6787_;
  assign new_n7436_ = ~new_n22713_ | ~new_n3551_;
  assign new_n7437_ = ~new_n24254_ | ~new_n3549_;
  assign new_n7438_ = ~new_n26065_ | ~new_n4376_;
  assign new_n7439_ = ~new_n25880_ | ~new_n5454_;
  assign new_n7440_ = ~new_n26465_ | ~new_n5455_;
  assign new_n7441_ = ~new_n23950_ | ~new_n5456_;
  assign new_n7442_ = ~new_n27397_ | ~new_n5457_;
  assign new_n7443_ = ~new_n21930_ | ~new_n3510_;
  assign new_n7444_ = ~new_n21088_ | ~new_n3511_;
  assign new_n7445_ = ~new_n24813_ | ~new_n5458_;
  assign new_n7446_ = ~new_n27218_ | ~new_n3512_;
  assign new_n7447_ = ~new_n21745_ | ~new_n5459_;
  assign new_n7448_ = ~new_n25331_ | ~new_n5460_;
  assign new_n7449_ = ~new_n25694_ | ~new_n5461_;
  assign new_n7450_ = ~new_n24991_ | ~new_n3513_;
  assign new_n7451_ = ~new_n26250_ | ~new_n3514_;
  assign new_n7452_ = ~new_n23330_ | ~new_n3515_;
  assign new_n7453_ = ~new_n25512_ | ~new_n5462_;
  assign new_n7454_ = ~new_n23519_ | ~new_n3518_;
  assign new_n7455_ = ~new_n26712_ | ~new_n3516_;
  assign new_n7456_ = ~new_n5059_ | ~new_n5067_ | ~new_n5062_ | ~new_n5060_ | ~new_n7438_;
  assign new_n7457_ = ~new_n3558_ | ~pi0535;
  assign new_n7458_ = ~new_n5474_ | ~new_n7456_;
  assign new_n7459_ = ~pi0344 | ~new_n6787_;
  assign new_n7460_ = ~new_n22650_ | ~new_n3551_;
  assign new_n7461_ = ~new_n24193_ | ~new_n3549_;
  assign new_n7462_ = ~new_n26064_ | ~new_n4376_;
  assign new_n7463_ = ~new_n25879_ | ~new_n5454_;
  assign new_n7464_ = ~new_n26464_ | ~new_n5455_;
  assign new_n7465_ = ~new_n23949_ | ~new_n5456_;
  assign new_n7466_ = ~new_n27396_ | ~new_n5457_;
  assign new_n7467_ = ~new_n21929_ | ~new_n3510_;
  assign new_n7468_ = ~new_n21087_ | ~new_n3511_;
  assign new_n7469_ = ~new_n24812_ | ~new_n5458_;
  assign new_n7470_ = ~new_n27217_ | ~new_n3512_;
  assign new_n7471_ = ~new_n21744_ | ~new_n5459_;
  assign new_n7472_ = ~new_n25330_ | ~new_n5460_;
  assign new_n7473_ = ~new_n25693_ | ~new_n5461_;
  assign new_n7474_ = ~new_n24990_ | ~new_n3513_;
  assign new_n7475_ = ~new_n26249_ | ~new_n3514_;
  assign new_n7476_ = ~new_n23329_ | ~new_n3515_;
  assign new_n7477_ = ~new_n25511_ | ~new_n5462_;
  assign new_n7478_ = ~new_n23518_ | ~new_n3518_;
  assign new_n7479_ = ~new_n26648_ | ~new_n3516_;
  assign new_n7480_ = ~new_n5068_ | ~new_n5076_ | ~new_n5071_ | ~new_n5069_ | ~new_n7462_;
  assign new_n7481_ = ~new_n3558_ | ~pi0536;
  assign new_n7482_ = ~new_n5474_ | ~new_n7480_;
  assign new_n7483_ = ~pi0345 | ~new_n6787_;
  assign new_n7484_ = ~new_n22651_ | ~new_n3551_;
  assign new_n7485_ = ~new_n24253_ | ~new_n3549_;
  assign new_n7486_ = ~new_n26063_ | ~new_n4376_;
  assign new_n7487_ = ~new_n25878_ | ~new_n5454_;
  assign new_n7488_ = ~new_n26463_ | ~new_n5455_;
  assign new_n7489_ = ~new_n23948_ | ~new_n5456_;
  assign new_n7490_ = ~new_n27395_ | ~new_n5457_;
  assign new_n7491_ = ~new_n21928_ | ~new_n3510_;
  assign new_n7492_ = ~new_n21086_ | ~new_n3511_;
  assign new_n7493_ = ~new_n24811_ | ~new_n5458_;
  assign new_n7494_ = ~new_n27216_ | ~new_n3512_;
  assign new_n7495_ = ~new_n21743_ | ~new_n5459_;
  assign new_n7496_ = ~new_n25329_ | ~new_n5460_;
  assign new_n7497_ = ~new_n25692_ | ~new_n5461_;
  assign new_n7498_ = ~new_n24989_ | ~new_n3513_;
  assign new_n7499_ = ~new_n26248_ | ~new_n3514_;
  assign new_n7500_ = ~new_n23328_ | ~new_n3515_;
  assign new_n7501_ = ~new_n25510_ | ~new_n5462_;
  assign new_n7502_ = ~new_n23517_ | ~new_n3518_;
  assign new_n7503_ = ~new_n26649_ | ~new_n3516_;
  assign new_n7504_ = ~new_n5077_ | ~new_n5085_ | ~new_n5080_ | ~new_n5078_ | ~new_n7486_;
  assign new_n7505_ = ~new_n3558_ | ~pi0537;
  assign new_n7506_ = ~new_n5474_ | ~new_n7504_;
  assign new_n7507_ = ~pi0346 | ~new_n6787_;
  assign new_n7508_ = ~new_n22712_ | ~new_n3551_;
  assign new_n7509_ = ~new_n24251_ | ~new_n3549_;
  assign new_n7510_ = ~new_n26061_ | ~new_n4376_;
  assign new_n7511_ = ~new_n25876_ | ~new_n5454_;
  assign new_n7512_ = ~new_n26461_ | ~new_n5455_;
  assign new_n7513_ = ~new_n23946_ | ~new_n5456_;
  assign new_n7514_ = ~new_n27393_ | ~new_n5457_;
  assign new_n7515_ = ~new_n21926_ | ~new_n3510_;
  assign new_n7516_ = ~new_n21084_ | ~new_n3511_;
  assign new_n7517_ = ~new_n24809_ | ~new_n5458_;
  assign new_n7518_ = ~new_n27214_ | ~new_n3512_;
  assign new_n7519_ = ~new_n21741_ | ~new_n5459_;
  assign new_n7520_ = ~new_n25327_ | ~new_n5460_;
  assign new_n7521_ = ~new_n25691_ | ~new_n5461_;
  assign new_n7522_ = ~new_n24988_ | ~new_n3513_;
  assign new_n7523_ = ~new_n26246_ | ~new_n3514_;
  assign new_n7524_ = ~new_n23326_ | ~new_n3515_;
  assign new_n7525_ = ~new_n25508_ | ~new_n5462_;
  assign new_n7526_ = ~new_n23515_ | ~new_n3518_;
  assign new_n7527_ = ~new_n26711_ | ~new_n3516_;
  assign new_n7528_ = ~new_n5086_ | ~new_n5094_ | ~new_n5089_ | ~new_n5087_ | ~new_n7510_;
  assign new_n7529_ = ~new_n3558_ | ~pi0538;
  assign new_n7530_ = ~new_n5474_ | ~new_n7528_;
  assign new_n7531_ = ~pi0347 | ~new_n6787_;
  assign new_n7532_ = ~new_n22725_ | ~new_n3551_;
  assign new_n7533_ = ~new_n24194_ | ~new_n3549_;
  assign new_n7534_ = ~new_n26060_ | ~new_n4376_;
  assign new_n7535_ = ~new_n25875_ | ~new_n5454_;
  assign new_n7536_ = ~new_n26460_ | ~new_n5455_;
  assign new_n7537_ = ~new_n23945_ | ~new_n5456_;
  assign new_n7538_ = ~new_n27392_ | ~new_n5457_;
  assign new_n7539_ = ~new_n21925_ | ~new_n3510_;
  assign new_n7540_ = ~new_n21083_ | ~new_n3511_;
  assign new_n7541_ = ~new_n24808_ | ~new_n5458_;
  assign new_n7542_ = ~new_n27213_ | ~new_n3512_;
  assign new_n7543_ = ~new_n21740_ | ~new_n5459_;
  assign new_n7544_ = ~new_n25326_ | ~new_n5460_;
  assign new_n7545_ = ~new_n25690_ | ~new_n5461_;
  assign new_n7546_ = ~new_n24987_ | ~new_n3513_;
  assign new_n7547_ = ~new_n26245_ | ~new_n3514_;
  assign new_n7548_ = ~new_n23325_ | ~new_n3515_;
  assign new_n7549_ = ~new_n25507_ | ~new_n5462_;
  assign new_n7550_ = ~new_n23514_ | ~new_n3518_;
  assign new_n7551_ = ~new_n26724_ | ~new_n3516_;
  assign new_n7552_ = ~new_n5106_ | ~new_n5101_;
  assign new_n7553_ = ~new_n3558_ | ~pi0539;
  assign new_n7554_ = ~pi0348 | ~new_n6787_;
  assign new_n7555_ = ~new_n22636_ | ~new_n3517_;
  assign new_n7556_ = ~new_n23443_ | ~new_n3516_;
  assign new_n7557_ = ~new_n7556_ | ~new_n7555_;
  assign new_n7558_ = ~new_n3546_ | ~new_n7557_;
  assign new_n7559_ = ~new_n4390_ | ~new_n4277_;
  assign new_n7560_ = ~new_n4405_;
  assign new_n7561_ = ~pi0349 | ~new_n3554_;
  assign new_n7562_ = ~pi0349 | ~new_n3553_;
  assign new_n7563_ = ~new_n3552_ | ~new_n22720_;
  assign new_n7564_ = ~new_n3550_ | ~new_n24243_;
  assign new_n7565_ = ~new_n3545_ | ~pi0508;
  assign new_n7566_ = ~pi0349 | ~new_n3544_;
  assign new_n7567_ = ~new_n3543_ | ~new_n26719_;
  assign new_n7568_ = ~pi0349 | ~new_n7560_;
  assign new_n7569_ = ~new_n22223_ | ~new_n3554_;
  assign new_n7570_ = ~pi0350 | ~new_n3553_;
  assign new_n7571_ = ~new_n3552_ | ~new_n22654_;
  assign new_n7572_ = ~new_n3550_ | ~new_n24195_;
  assign new_n7573_ = ~new_n3545_ | ~pi0509;
  assign new_n7574_ = ~new_n23655_ | ~new_n3544_;
  assign new_n7575_ = ~new_n3543_ | ~new_n26652_;
  assign new_n7576_ = ~pi0350 | ~new_n7560_;
  assign new_n7577_ = ~new_n22290_ | ~new_n3554_;
  assign new_n7578_ = ~new_n22463_ | ~new_n3553_;
  assign new_n7579_ = ~new_n3552_ | ~new_n22726_;
  assign new_n7580_ = ~new_n3550_ | ~new_n24252_;
  assign new_n7581_ = ~new_n3545_ | ~pi0510;
  assign new_n7582_ = ~new_n23722_ | ~new_n3544_;
  assign new_n7583_ = ~new_n3543_ | ~new_n26725_;
  assign new_n7584_ = ~pi0351 | ~new_n7560_;
  assign new_n7585_ = ~new_n22287_ | ~new_n3554_;
  assign new_n7586_ = ~new_n22525_ | ~new_n3553_;
  assign new_n7587_ = ~new_n3552_ | ~new_n22652_;
  assign new_n7588_ = ~new_n3550_ | ~new_n24250_;
  assign new_n7589_ = ~new_n3545_ | ~pi0511;
  assign new_n7590_ = ~new_n23719_ | ~new_n3544_;
  assign new_n7591_ = ~new_n3543_ | ~new_n26650_;
  assign new_n7592_ = ~pi0352 | ~new_n7560_;
  assign new_n7593_ = ~new_n22286_ | ~new_n3554_;
  assign new_n7594_ = ~new_n22524_ | ~new_n3553_;
  assign new_n7595_ = ~new_n3552_ | ~new_n22653_;
  assign new_n7596_ = ~new_n3550_ | ~new_n24249_;
  assign new_n7597_ = ~new_n3545_ | ~pi0512;
  assign new_n7598_ = ~new_n23718_ | ~new_n3544_;
  assign new_n7599_ = ~new_n3543_ | ~new_n26723_;
  assign new_n7600_ = ~pi0353 | ~new_n7560_;
  assign new_n7601_ = ~new_n22285_ | ~new_n3554_;
  assign new_n7602_ = ~new_n22523_ | ~new_n3553_;
  assign new_n7603_ = ~new_n3552_ | ~new_n22724_;
  assign new_n7604_ = ~new_n3550_ | ~new_n24248_;
  assign new_n7605_ = ~new_n3545_ | ~pi0513;
  assign new_n7606_ = ~new_n23717_ | ~new_n3544_;
  assign new_n7607_ = ~new_n3543_ | ~new_n26651_;
  assign new_n7608_ = ~pi0354 | ~new_n7560_;
  assign new_n7609_ = ~new_n22284_ | ~new_n3554_;
  assign new_n7610_ = ~new_n22522_ | ~new_n3553_;
  assign new_n7611_ = ~new_n3552_ | ~new_n22723_;
  assign new_n7612_ = ~new_n3550_ | ~new_n24247_;
  assign new_n7613_ = ~new_n3545_ | ~pi0514;
  assign new_n7614_ = ~new_n23716_ | ~new_n3544_;
  assign new_n7615_ = ~new_n3543_ | ~new_n26722_;
  assign new_n7616_ = ~pi0355 | ~new_n7560_;
  assign new_n7617_ = ~new_n22283_ | ~new_n3554_;
  assign new_n7618_ = ~new_n22521_ | ~new_n3553_;
  assign new_n7619_ = ~new_n3552_ | ~new_n22722_;
  assign new_n7620_ = ~new_n3550_ | ~new_n24246_;
  assign new_n7621_ = ~new_n3545_ | ~pi0515;
  assign new_n7622_ = ~new_n23715_ | ~new_n3544_;
  assign new_n7623_ = ~new_n3543_ | ~new_n26721_;
  assign new_n7624_ = ~pi0356 | ~new_n7560_;
  assign new_n7625_ = ~new_n22282_ | ~new_n3554_;
  assign new_n7626_ = ~new_n22520_ | ~new_n3553_;
  assign new_n7627_ = ~new_n3552_ | ~new_n22721_;
  assign new_n7628_ = ~new_n3550_ | ~new_n24245_;
  assign new_n7629_ = ~new_n3545_ | ~pi0516;
  assign new_n7630_ = ~new_n23714_ | ~new_n3544_;
  assign new_n7631_ = ~new_n3543_ | ~new_n26720_;
  assign new_n7632_ = ~pi0357 | ~new_n7560_;
  assign new_n7633_ = ~new_n22281_ | ~new_n3554_;
  assign new_n7634_ = ~new_n22519_ | ~new_n3553_;
  assign new_n7635_ = ~new_n3552_ | ~new_n22741_;
  assign new_n7636_ = ~new_n3550_ | ~new_n24244_;
  assign new_n7637_ = ~new_n3545_ | ~pi0517;
  assign new_n7638_ = ~new_n23713_ | ~new_n3544_;
  assign new_n7639_ = ~new_n3543_ | ~new_n26741_;
  assign new_n7640_ = ~pi0358 | ~new_n7560_;
  assign new_n7641_ = ~new_n22310_ | ~new_n3554_;
  assign new_n7642_ = ~new_n22547_ | ~new_n3553_;
  assign new_n7643_ = ~new_n3552_ | ~new_n22639_;
  assign new_n7644_ = ~new_n3550_ | ~new_n24267_;
  assign new_n7645_ = ~new_n3545_ | ~pi0518;
  assign new_n7646_ = ~new_n23742_ | ~new_n3544_;
  assign new_n7647_ = ~new_n3543_ | ~new_n26637_;
  assign new_n7648_ = ~pi0359 | ~new_n7560_;
  assign new_n7649_ = ~new_n22309_ | ~new_n3554_;
  assign new_n7650_ = ~new_n22546_ | ~new_n3553_;
  assign new_n7651_ = ~new_n3552_ | ~new_n22719_;
  assign new_n7652_ = ~new_n3550_ | ~new_n24266_;
  assign new_n7653_ = ~new_n3545_ | ~pi0519;
  assign new_n7654_ = ~new_n23741_ | ~new_n3544_;
  assign new_n7655_ = ~new_n3543_ | ~new_n26718_;
  assign new_n7656_ = ~pi0360 | ~new_n7560_;
  assign new_n7657_ = ~new_n22308_ | ~new_n3554_;
  assign new_n7658_ = ~new_n22545_ | ~new_n3553_;
  assign new_n7659_ = ~new_n3552_ | ~new_n22640_;
  assign new_n7660_ = ~new_n3550_ | ~new_n24265_;
  assign new_n7661_ = ~new_n3545_ | ~pi0520;
  assign new_n7662_ = ~new_n23740_ | ~new_n3544_;
  assign new_n7663_ = ~new_n3543_ | ~new_n26638_;
  assign new_n7664_ = ~pi0361 | ~new_n7560_;
  assign new_n7665_ = ~new_n22307_ | ~new_n3554_;
  assign new_n7666_ = ~new_n22544_ | ~new_n3553_;
  assign new_n7667_ = ~new_n3552_ | ~new_n22641_;
  assign new_n7668_ = ~new_n3550_ | ~new_n24189_;
  assign new_n7669_ = ~new_n3545_ | ~pi0521;
  assign new_n7670_ = ~new_n23739_ | ~new_n3544_;
  assign new_n7671_ = ~new_n3543_ | ~new_n26639_;
  assign new_n7672_ = ~pi0362 | ~new_n7560_;
  assign new_n7673_ = ~new_n22306_ | ~new_n3554_;
  assign new_n7674_ = ~new_n22543_ | ~new_n3553_;
  assign new_n7675_ = ~new_n3552_ | ~new_n22718_;
  assign new_n7676_ = ~new_n3550_ | ~new_n24264_;
  assign new_n7677_ = ~new_n3545_ | ~pi0522;
  assign new_n7678_ = ~new_n23738_ | ~new_n3544_;
  assign new_n7679_ = ~new_n3543_ | ~new_n26717_;
  assign new_n7680_ = ~pi0363 | ~new_n7560_;
  assign new_n7681_ = ~new_n22305_ | ~new_n3554_;
  assign new_n7682_ = ~new_n22542_ | ~new_n3553_;
  assign new_n7683_ = ~new_n3552_ | ~new_n22642_;
  assign new_n7684_ = ~new_n3550_ | ~new_n24263_;
  assign new_n7685_ = ~new_n3545_ | ~pi0523;
  assign new_n7686_ = ~new_n23737_ | ~new_n3544_;
  assign new_n7687_ = ~new_n3543_ | ~new_n26640_;
  assign new_n7688_ = ~pi0364 | ~new_n7560_;
  assign new_n7689_ = ~new_n22304_ | ~new_n3554_;
  assign new_n7690_ = ~new_n22541_ | ~new_n3553_;
  assign new_n7691_ = ~new_n3552_ | ~new_n22717_;
  assign new_n7692_ = ~new_n3550_ | ~new_n24262_;
  assign new_n7693_ = ~new_n3545_ | ~pi0524;
  assign new_n7694_ = ~new_n23736_ | ~new_n3544_;
  assign new_n7695_ = ~new_n3543_ | ~new_n26716_;
  assign new_n7696_ = ~pi0365 | ~new_n7560_;
  assign new_n7697_ = ~new_n22303_ | ~new_n3554_;
  assign new_n7698_ = ~new_n22540_ | ~new_n3553_;
  assign new_n7699_ = ~new_n3552_ | ~new_n22643_;
  assign new_n7700_ = ~new_n3550_ | ~new_n24190_;
  assign new_n7701_ = ~new_n3545_ | ~pi0525;
  assign new_n7702_ = ~new_n23735_ | ~new_n3544_;
  assign new_n7703_ = ~new_n3543_ | ~new_n26641_;
  assign new_n7704_ = ~pi0366 | ~new_n7560_;
  assign new_n7705_ = ~new_n22302_ | ~new_n3554_;
  assign new_n7706_ = ~new_n22539_ | ~new_n3553_;
  assign new_n7707_ = ~new_n3552_ | ~new_n22716_;
  assign new_n7708_ = ~new_n3550_ | ~new_n24261_;
  assign new_n7709_ = ~new_n3545_ | ~pi0526;
  assign new_n7710_ = ~new_n23734_ | ~new_n3544_;
  assign new_n7711_ = ~new_n3543_ | ~new_n26715_;
  assign new_n7712_ = ~pi0367 | ~new_n7560_;
  assign new_n7713_ = ~new_n22301_ | ~new_n3554_;
  assign new_n7714_ = ~new_n22538_ | ~new_n3553_;
  assign new_n7715_ = ~new_n3552_ | ~new_n22644_;
  assign new_n7716_ = ~new_n3550_ | ~new_n24260_;
  assign new_n7717_ = ~new_n3545_ | ~pi0527;
  assign new_n7718_ = ~new_n23733_ | ~new_n3544_;
  assign new_n7719_ = ~new_n3543_ | ~new_n26642_;
  assign new_n7720_ = ~pi0368 | ~new_n7560_;
  assign new_n7721_ = ~new_n22300_ | ~new_n3554_;
  assign new_n7722_ = ~new_n22537_ | ~new_n3553_;
  assign new_n7723_ = ~new_n3552_ | ~new_n22645_;
  assign new_n7724_ = ~new_n3550_ | ~new_n24191_;
  assign new_n7725_ = ~new_n3545_ | ~pi0528;
  assign new_n7726_ = ~new_n23732_ | ~new_n3544_;
  assign new_n7727_ = ~new_n3543_ | ~new_n26643_;
  assign new_n7728_ = ~pi0369 | ~new_n7560_;
  assign new_n7729_ = ~new_n22299_ | ~new_n3554_;
  assign new_n7730_ = ~new_n22536_ | ~new_n3553_;
  assign new_n7731_ = ~new_n3552_ | ~new_n22646_;
  assign new_n7732_ = ~new_n3550_ | ~new_n24259_;
  assign new_n7733_ = ~new_n3545_ | ~pi0529;
  assign new_n7734_ = ~new_n23731_ | ~new_n3544_;
  assign new_n7735_ = ~new_n3543_ | ~new_n26644_;
  assign new_n7736_ = ~pi0370 | ~new_n7560_;
  assign new_n7737_ = ~new_n22298_ | ~new_n3554_;
  assign new_n7738_ = ~new_n22535_ | ~new_n3553_;
  assign new_n7739_ = ~new_n3552_ | ~new_n22715_;
  assign new_n7740_ = ~new_n3550_ | ~new_n24258_;
  assign new_n7741_ = ~new_n3545_ | ~pi0530;
  assign new_n7742_ = ~new_n23730_ | ~new_n3544_;
  assign new_n7743_ = ~new_n3543_ | ~new_n26714_;
  assign new_n7744_ = ~pi0371 | ~new_n7560_;
  assign new_n7745_ = ~new_n22297_ | ~new_n3554_;
  assign new_n7746_ = ~new_n22534_ | ~new_n3553_;
  assign new_n7747_ = ~new_n3552_ | ~new_n22647_;
  assign new_n7748_ = ~new_n3550_ | ~new_n24257_;
  assign new_n7749_ = ~new_n3545_ | ~pi0531;
  assign new_n7750_ = ~new_n23729_ | ~new_n3544_;
  assign new_n7751_ = ~new_n3543_ | ~new_n26645_;
  assign new_n7752_ = ~pi0372 | ~new_n7560_;
  assign new_n7753_ = ~new_n22296_ | ~new_n3554_;
  assign new_n7754_ = ~new_n22533_ | ~new_n3553_;
  assign new_n7755_ = ~new_n3552_ | ~new_n22714_;
  assign new_n7756_ = ~new_n3550_ | ~new_n24256_;
  assign new_n7757_ = ~new_n3545_ | ~pi0532;
  assign new_n7758_ = ~new_n23728_ | ~new_n3544_;
  assign new_n7759_ = ~new_n3543_ | ~new_n26713_;
  assign new_n7760_ = ~pi0373 | ~new_n7560_;
  assign new_n7761_ = ~new_n22295_ | ~new_n3554_;
  assign new_n7762_ = ~new_n22532_ | ~new_n3553_;
  assign new_n7763_ = ~new_n3552_ | ~new_n22648_;
  assign new_n7764_ = ~new_n3550_ | ~new_n24255_;
  assign new_n7765_ = ~new_n3545_ | ~pi0533;
  assign new_n7766_ = ~new_n23727_ | ~new_n3544_;
  assign new_n7767_ = ~new_n3543_ | ~new_n26646_;
  assign new_n7768_ = ~pi0374 | ~new_n7560_;
  assign new_n7769_ = ~new_n22294_ | ~new_n3554_;
  assign new_n7770_ = ~new_n22531_ | ~new_n3553_;
  assign new_n7771_ = ~new_n3552_ | ~new_n22649_;
  assign new_n7772_ = ~new_n3550_ | ~new_n24192_;
  assign new_n7773_ = ~new_n3545_ | ~pi0534;
  assign new_n7774_ = ~new_n23726_ | ~new_n3544_;
  assign new_n7775_ = ~new_n3543_ | ~new_n26647_;
  assign new_n7776_ = ~pi0375 | ~new_n7560_;
  assign new_n7777_ = ~new_n22293_ | ~new_n3554_;
  assign new_n7778_ = ~new_n22530_ | ~new_n3553_;
  assign new_n7779_ = ~new_n3552_ | ~new_n22713_;
  assign new_n7780_ = ~new_n3550_ | ~new_n24254_;
  assign new_n7781_ = ~new_n3545_ | ~pi0535;
  assign new_n7782_ = ~new_n23725_ | ~new_n3544_;
  assign new_n7783_ = ~new_n3543_ | ~new_n26712_;
  assign new_n7784_ = ~pi0376 | ~new_n7560_;
  assign new_n7785_ = ~new_n22292_ | ~new_n3554_;
  assign new_n7786_ = ~new_n22529_ | ~new_n3553_;
  assign new_n7787_ = ~new_n3552_ | ~new_n22650_;
  assign new_n7788_ = ~new_n3550_ | ~new_n24193_;
  assign new_n7789_ = ~new_n3545_ | ~pi0536;
  assign new_n7790_ = ~new_n23724_ | ~new_n3544_;
  assign new_n7791_ = ~new_n3543_ | ~new_n26648_;
  assign new_n7792_ = ~pi0377 | ~new_n7560_;
  assign new_n7793_ = ~new_n22291_ | ~new_n3554_;
  assign new_n7794_ = ~new_n22528_ | ~new_n3553_;
  assign new_n7795_ = ~new_n3552_ | ~new_n22651_;
  assign new_n7796_ = ~new_n3550_ | ~new_n24253_;
  assign new_n7797_ = ~new_n3545_ | ~pi0537;
  assign new_n7798_ = ~new_n23723_ | ~new_n3544_;
  assign new_n7799_ = ~new_n3543_ | ~new_n26649_;
  assign new_n7800_ = ~pi0378 | ~new_n7560_;
  assign new_n7801_ = ~new_n22289_ | ~new_n3554_;
  assign new_n7802_ = ~new_n22527_ | ~new_n3553_;
  assign new_n7803_ = ~new_n3552_ | ~new_n22712_;
  assign new_n7804_ = ~new_n3550_ | ~new_n24251_;
  assign new_n7805_ = ~new_n3545_ | ~pi0538;
  assign new_n7806_ = ~new_n23721_ | ~new_n3544_;
  assign new_n7807_ = ~new_n3543_ | ~new_n26711_;
  assign new_n7808_ = ~pi0379 | ~new_n7560_;
  assign new_n7809_ = ~new_n22288_ | ~new_n3554_;
  assign new_n7810_ = ~new_n22526_ | ~new_n3553_;
  assign new_n7811_ = ~new_n3552_ | ~new_n22725_;
  assign new_n7812_ = ~new_n3550_ | ~new_n24194_;
  assign new_n7813_ = ~new_n3545_ | ~pi0539;
  assign new_n7814_ = ~new_n23720_ | ~new_n3544_;
  assign new_n7815_ = ~new_n3543_ | ~new_n26724_;
  assign new_n7816_ = ~pi0380 | ~new_n7560_;
  assign new_n7817_ = ~new_n27144_ | ~new_n5460_ | ~new_n3786_;
  assign new_n7818_ = ~new_n25105_ | ~new_n5459_;
  assign new_n7819_ = ~new_n7818_ | ~new_n7817_;
  assign new_n7820_ = ~pi0459 | ~new_n3563_;
  assign new_n7821_ = ~pi0085 | ~new_n3562_;
  assign new_n7822_ = ~pi0381 | ~new_n4406_;
  assign new_n7823_ = ~pi0458 | ~new_n3563_;
  assign new_n7824_ = ~pi0084 | ~new_n3562_;
  assign new_n7825_ = ~pi0382 | ~new_n4406_;
  assign new_n7826_ = ~pi0457 | ~new_n3563_;
  assign new_n7827_ = ~pi0083 | ~new_n3562_;
  assign new_n7828_ = ~pi0383 | ~new_n4406_;
  assign new_n7829_ = ~pi0456 | ~new_n3563_;
  assign new_n7830_ = ~pi0082 | ~new_n3562_;
  assign new_n7831_ = ~pi0384 | ~new_n4406_;
  assign new_n7832_ = ~pi0455 | ~new_n3563_;
  assign new_n7833_ = ~pi0081 | ~new_n3562_;
  assign new_n7834_ = ~pi0385 | ~new_n4406_;
  assign new_n7835_ = ~pi0454 | ~new_n3563_;
  assign new_n7836_ = ~pi0080 | ~new_n3562_;
  assign new_n7837_ = ~pi0386 | ~new_n4406_;
  assign new_n7838_ = ~pi0453 | ~new_n3563_;
  assign new_n7839_ = ~pi0079 | ~new_n3562_;
  assign new_n7840_ = ~pi0387 | ~new_n4406_;
  assign new_n7841_ = ~pi0452 | ~new_n3563_;
  assign new_n7842_ = ~pi0078 | ~new_n3562_;
  assign new_n7843_ = ~pi0388 | ~new_n4406_;
  assign new_n7844_ = ~pi0451 | ~new_n3563_;
  assign new_n7845_ = ~new_n3562_ | ~pi0077;
  assign new_n7846_ = ~pi0389 | ~new_n4406_;
  assign new_n7847_ = ~pi0450 | ~new_n3563_;
  assign new_n7848_ = ~new_n3562_ | ~pi0076;
  assign new_n7849_ = ~pi0390 | ~new_n4406_;
  assign new_n7850_ = ~pi0449 | ~new_n3563_;
  assign new_n7851_ = ~new_n3562_ | ~pi0075;
  assign new_n7852_ = ~pi0391 | ~new_n4406_;
  assign new_n7853_ = ~pi0448 | ~new_n3563_;
  assign new_n7854_ = ~new_n3562_ | ~pi0074;
  assign new_n7855_ = ~pi0392 | ~new_n4406_;
  assign new_n7856_ = ~pi0447 | ~new_n3563_;
  assign new_n7857_ = ~new_n3562_ | ~pi0073;
  assign new_n7858_ = ~pi0393 | ~new_n4406_;
  assign new_n7859_ = ~pi0446 | ~new_n3563_;
  assign new_n7860_ = ~new_n3562_ | ~pi0072;
  assign new_n7861_ = ~pi0394 | ~new_n4406_;
  assign new_n7862_ = ~pi0445 | ~new_n3563_;
  assign new_n7863_ = ~new_n3562_ | ~pi0071;
  assign new_n7864_ = ~pi0395 | ~new_n4406_;
  assign new_n7865_ = ~pi0444 | ~new_n3563_;
  assign new_n7866_ = ~new_n3562_ | ~pi0070;
  assign new_n7867_ = ~pi0396 | ~new_n4406_;
  assign new_n7868_ = ~pi0474 | ~new_n3563_;
  assign new_n7869_ = ~pi0084 | ~new_n3562_;
  assign new_n7870_ = ~pi0397 | ~new_n4406_;
  assign new_n7871_ = ~pi0473 | ~new_n3563_;
  assign new_n7872_ = ~pi0083 | ~new_n3562_;
  assign new_n7873_ = ~pi0398 | ~new_n4406_;
  assign new_n7874_ = ~pi0472 | ~new_n3563_;
  assign new_n7875_ = ~pi0082 | ~new_n3562_;
  assign new_n7876_ = ~pi0399 | ~new_n4406_;
  assign new_n7877_ = ~pi0471 | ~new_n3563_;
  assign new_n7878_ = ~pi0081 | ~new_n3562_;
  assign new_n7879_ = ~pi0400 | ~new_n4406_;
  assign new_n7880_ = ~pi0470 | ~new_n3563_;
  assign new_n7881_ = ~pi0080 | ~new_n3562_;
  assign new_n7882_ = ~pi0401 | ~new_n4406_;
  assign new_n7883_ = ~pi0469 | ~new_n3563_;
  assign new_n7884_ = ~pi0079 | ~new_n3562_;
  assign new_n7885_ = ~pi0402 | ~new_n4406_;
  assign new_n7886_ = ~pi0468 | ~new_n3563_;
  assign new_n7887_ = ~pi0078 | ~new_n3562_;
  assign new_n7888_ = ~pi0403 | ~new_n4406_;
  assign new_n7889_ = ~pi0467 | ~new_n3563_;
  assign new_n7890_ = ~new_n3562_ | ~pi0077;
  assign new_n7891_ = ~pi0404 | ~new_n4406_;
  assign new_n7892_ = ~pi0466 | ~new_n3563_;
  assign new_n7893_ = ~new_n3562_ | ~pi0076;
  assign new_n7894_ = ~pi0405 | ~new_n4406_;
  assign new_n7895_ = ~pi0465 | ~new_n3563_;
  assign new_n7896_ = ~new_n3562_ | ~pi0075;
  assign new_n7897_ = ~pi0406 | ~new_n4406_;
  assign new_n7898_ = ~pi0464 | ~new_n3563_;
  assign new_n7899_ = ~new_n3562_ | ~pi0074;
  assign new_n7900_ = ~pi0407 | ~new_n4406_;
  assign new_n7901_ = ~pi0463 | ~new_n3563_;
  assign new_n7902_ = ~new_n3562_ | ~pi0073;
  assign new_n7903_ = ~pi0408 | ~new_n4406_;
  assign new_n7904_ = ~pi0462 | ~new_n3563_;
  assign new_n7905_ = ~new_n3562_ | ~pi0072;
  assign new_n7906_ = ~pi0409 | ~new_n4406_;
  assign new_n7907_ = ~pi0461 | ~new_n3563_;
  assign new_n7908_ = ~new_n3562_ | ~pi0071;
  assign new_n7909_ = ~pi0410 | ~new_n4406_;
  assign new_n7910_ = ~pi0460 | ~new_n3563_;
  assign new_n7911_ = ~new_n3562_ | ~pi0070;
  assign new_n7912_ = ~pi0411 | ~new_n4406_;
  assign new_n7913_ = ~new_n5142_ | ~new_n4411_;
  assign new_n7914_ = ~new_n3609_ | ~new_n4277_;
  assign new_n7915_ = ~new_n4407_;
  assign new_n7916_ = ~new_n3566_ | ~pi0396;
  assign new_n7917_ = ~new_n3565_ | ~pi0444;
  assign new_n7918_ = ~pi0412 | ~new_n7915_;
  assign new_n7919_ = ~new_n3566_ | ~pi0395;
  assign new_n7920_ = ~new_n3565_ | ~pi0445;
  assign new_n7921_ = ~pi0413 | ~new_n7915_;
  assign new_n7922_ = ~new_n3566_ | ~pi0394;
  assign new_n7923_ = ~new_n3565_ | ~pi0446;
  assign new_n7924_ = ~pi0414 | ~new_n7915_;
  assign new_n7925_ = ~new_n3566_ | ~pi0393;
  assign new_n7926_ = ~new_n3565_ | ~pi0447;
  assign new_n7927_ = ~pi0415 | ~new_n7915_;
  assign new_n7928_ = ~new_n3566_ | ~pi0392;
  assign new_n7929_ = ~new_n3565_ | ~pi0448;
  assign new_n7930_ = ~pi0416 | ~new_n7915_;
  assign new_n7931_ = ~new_n3566_ | ~pi0391;
  assign new_n7932_ = ~new_n3565_ | ~pi0449;
  assign new_n7933_ = ~pi0417 | ~new_n7915_;
  assign new_n7934_ = ~new_n3566_ | ~pi0390;
  assign new_n7935_ = ~new_n3565_ | ~pi0450;
  assign new_n7936_ = ~pi0418 | ~new_n7915_;
  assign new_n7937_ = ~new_n3566_ | ~pi0389;
  assign new_n7938_ = ~new_n3565_ | ~pi0451;
  assign new_n7939_ = ~pi0419 | ~new_n7915_;
  assign new_n7940_ = ~new_n3566_ | ~pi0388;
  assign new_n7941_ = ~new_n3565_ | ~pi0452;
  assign new_n7942_ = ~pi0420 | ~new_n7915_;
  assign new_n7943_ = ~new_n3566_ | ~pi0387;
  assign new_n7944_ = ~new_n3565_ | ~pi0453;
  assign new_n7945_ = ~pi0421 | ~new_n7915_;
  assign new_n7946_ = ~new_n3566_ | ~pi0386;
  assign new_n7947_ = ~new_n3565_ | ~pi0454;
  assign new_n7948_ = ~pi0422 | ~new_n7915_;
  assign new_n7949_ = ~new_n3566_ | ~pi0385;
  assign new_n7950_ = ~new_n3565_ | ~pi0455;
  assign new_n7951_ = ~pi0423 | ~new_n7915_;
  assign new_n7952_ = ~new_n3566_ | ~pi0384;
  assign new_n7953_ = ~new_n3565_ | ~pi0456;
  assign new_n7954_ = ~pi0424 | ~new_n7915_;
  assign new_n7955_ = ~new_n3566_ | ~pi0383;
  assign new_n7956_ = ~new_n3565_ | ~pi0457;
  assign new_n7957_ = ~pi0425 | ~new_n7915_;
  assign new_n7958_ = ~new_n3566_ | ~pi0382;
  assign new_n7959_ = ~new_n3565_ | ~pi0458;
  assign new_n7960_ = ~pi0426 | ~new_n7915_;
  assign new_n7961_ = ~new_n3566_ | ~pi0381;
  assign new_n7962_ = ~new_n3565_ | ~pi0459;
  assign new_n7963_ = ~pi0427 | ~new_n7915_;
  assign new_n7964_ = ~new_n3603_ | ~pi0460;
  assign new_n7965_ = ~new_n3566_ | ~pi0411;
  assign new_n7966_ = ~pi0428 | ~new_n7915_;
  assign new_n7967_ = ~new_n3603_ | ~pi0461;
  assign new_n7968_ = ~new_n3566_ | ~pi0410;
  assign new_n7969_ = ~pi0429 | ~new_n7915_;
  assign new_n7970_ = ~new_n3603_ | ~pi0462;
  assign new_n7971_ = ~new_n3566_ | ~pi0409;
  assign new_n7972_ = ~pi0430 | ~new_n7915_;
  assign new_n7973_ = ~new_n3603_ | ~pi0463;
  assign new_n7974_ = ~new_n3566_ | ~pi0408;
  assign new_n7975_ = ~pi0431 | ~new_n7915_;
  assign new_n7976_ = ~new_n3603_ | ~pi0464;
  assign new_n7977_ = ~new_n3566_ | ~pi0407;
  assign new_n7978_ = ~pi0432 | ~new_n7915_;
  assign new_n7979_ = ~new_n3603_ | ~pi0465;
  assign new_n7980_ = ~new_n3566_ | ~pi0406;
  assign new_n7981_ = ~pi0433 | ~new_n7915_;
  assign new_n7982_ = ~new_n3603_ | ~pi0466;
  assign new_n7983_ = ~new_n3566_ | ~pi0405;
  assign new_n7984_ = ~pi0434 | ~new_n7915_;
  assign new_n7985_ = ~new_n3603_ | ~pi0467;
  assign new_n7986_ = ~new_n3566_ | ~pi0404;
  assign new_n7987_ = ~pi0435 | ~new_n7915_;
  assign new_n7988_ = ~new_n3603_ | ~pi0468;
  assign new_n7989_ = ~new_n3566_ | ~pi0403;
  assign new_n7990_ = ~pi0436 | ~new_n7915_;
  assign new_n7991_ = ~new_n3603_ | ~pi0469;
  assign new_n7992_ = ~new_n3566_ | ~pi0402;
  assign new_n7993_ = ~pi0437 | ~new_n7915_;
  assign new_n7994_ = ~new_n3603_ | ~pi0470;
  assign new_n7995_ = ~new_n3566_ | ~pi0401;
  assign new_n7996_ = ~pi0438 | ~new_n7915_;
  assign new_n7997_ = ~new_n3603_ | ~pi0471;
  assign new_n7998_ = ~new_n3566_ | ~pi0400;
  assign new_n7999_ = ~pi0439 | ~new_n7915_;
  assign new_n8000_ = ~new_n3603_ | ~pi0472;
  assign new_n8001_ = ~new_n3566_ | ~pi0399;
  assign new_n8002_ = ~pi0440 | ~new_n7915_;
  assign new_n8003_ = ~new_n3603_ | ~pi0473;
  assign new_n8004_ = ~new_n3566_ | ~pi0398;
  assign new_n8005_ = ~pi0441 | ~new_n7915_;
  assign new_n8006_ = ~new_n3603_ | ~pi0474;
  assign new_n8007_ = ~new_n3566_ | ~pi0397;
  assign new_n8008_ = ~pi0442 | ~new_n7915_;
  assign new_n8009_ = ~new_n3672_ | ~new_n4399_;
  assign new_n8010_ = ~new_n3602_ | ~pi0070;
  assign new_n8011_ = ~new_n3777_ | ~new_n3567_;
  assign new_n8012_ = ~new_n21426_ | ~new_n3556_;
  assign new_n8013_ = ~pi0444 | ~new_n4408_;
  assign new_n8014_ = ~new_n3602_ | ~pi0071;
  assign new_n8015_ = ~new_n3778_ | ~new_n3567_;
  assign new_n8016_ = ~new_n21492_ | ~new_n3556_;
  assign new_n8017_ = ~pi0445 | ~new_n4408_;
  assign new_n8018_ = ~new_n3602_ | ~pi0072;
  assign new_n8019_ = ~new_n3779_ | ~new_n3567_;
  assign new_n8020_ = ~new_n21481_ | ~new_n3556_;
  assign new_n8021_ = ~pi0446 | ~new_n4408_;
  assign new_n8022_ = ~new_n3602_ | ~pi0073;
  assign new_n8023_ = ~new_n3780_ | ~new_n3567_;
  assign new_n8024_ = ~new_n21478_ | ~new_n3556_;
  assign new_n8025_ = ~pi0447 | ~new_n4408_;
  assign new_n8026_ = ~new_n3602_ | ~pi0074;
  assign new_n8027_ = ~new_n3781_ | ~new_n3567_;
  assign new_n8028_ = ~new_n21477_ | ~new_n3556_;
  assign new_n8029_ = ~pi0448 | ~new_n4408_;
  assign new_n8030_ = ~new_n3602_ | ~pi0075;
  assign new_n8031_ = ~new_n3782_ | ~new_n3567_;
  assign new_n8032_ = ~new_n21476_ | ~new_n3556_;
  assign new_n8033_ = ~pi0449 | ~new_n4408_;
  assign new_n8034_ = ~new_n3602_ | ~pi0076;
  assign new_n8035_ = ~new_n3783_ | ~new_n3567_;
  assign new_n8036_ = ~new_n21475_ | ~new_n3556_;
  assign new_n8037_ = ~pi0450 | ~new_n4408_;
  assign new_n8038_ = ~new_n3602_ | ~pi0077;
  assign new_n8039_ = ~new_n3784_ | ~new_n3567_;
  assign new_n8040_ = ~new_n21474_ | ~new_n3556_;
  assign new_n8041_ = ~pi0451 | ~new_n4408_;
  assign new_n8042_ = ~new_n3602_ | ~pi0078;
  assign new_n8043_ = ~new_n3761_ | ~new_n3567_;
  assign new_n8044_ = ~new_n21473_ | ~new_n3556_;
  assign new_n8045_ = ~pi0452 | ~new_n4408_;
  assign new_n8046_ = ~new_n3602_ | ~pi0079;
  assign new_n8047_ = ~new_n3762_ | ~new_n3567_;
  assign new_n8048_ = ~new_n21472_ | ~new_n3556_;
  assign new_n8049_ = ~pi0453 | ~new_n4408_;
  assign new_n8050_ = ~new_n3602_ | ~pi0080;
  assign new_n8051_ = ~new_n3763_ | ~new_n3567_;
  assign new_n8052_ = ~new_n21502_ | ~new_n3556_;
  assign new_n8053_ = ~pi0454 | ~new_n4408_;
  assign new_n8054_ = ~new_n3602_ | ~pi0081;
  assign new_n8055_ = ~new_n3764_ | ~new_n3567_;
  assign new_n8056_ = ~new_n21501_ | ~new_n3556_;
  assign new_n8057_ = ~pi0455 | ~new_n4408_;
  assign new_n8058_ = ~new_n3602_ | ~pi0082;
  assign new_n8059_ = ~new_n3765_ | ~new_n3567_;
  assign new_n8060_ = ~new_n21500_ | ~new_n3556_;
  assign new_n8061_ = ~pi0456 | ~new_n4408_;
  assign new_n8062_ = ~new_n3602_ | ~pi0083;
  assign new_n8063_ = ~new_n3766_ | ~new_n3567_;
  assign new_n8064_ = ~new_n21499_ | ~new_n3556_;
  assign new_n8065_ = ~pi0457 | ~new_n4408_;
  assign new_n8066_ = ~new_n3602_ | ~pi0084;
  assign new_n8067_ = ~new_n3767_ | ~new_n3567_;
  assign new_n8068_ = ~new_n21498_ | ~new_n3556_;
  assign new_n8069_ = ~pi0458 | ~new_n4408_;
  assign new_n8070_ = ~new_n3602_ | ~pi0085;
  assign new_n8071_ = ~new_n3768_ | ~new_n3567_;
  assign new_n8072_ = ~new_n21497_ | ~new_n3556_;
  assign new_n8073_ = ~pi0459 | ~new_n4408_;
  assign new_n8074_ = ~new_n3604_ | ~pi0070;
  assign new_n8075_ = ~new_n3600_ | ~pi0086;
  assign new_n8076_ = ~new_n4218_ | ~new_n3567_;
  assign new_n8077_ = ~new_n21496_ | ~new_n3556_;
  assign new_n8078_ = ~pi0460 | ~new_n4408_;
  assign new_n8079_ = ~new_n3604_ | ~pi0071;
  assign new_n8080_ = ~new_n3600_ | ~pi0087;
  assign new_n8081_ = ~new_n4219_ | ~new_n3567_;
  assign new_n8082_ = ~new_n21495_ | ~new_n3556_;
  assign new_n8083_ = ~pi0461 | ~new_n4408_;
  assign new_n8084_ = ~new_n3604_ | ~pi0072;
  assign new_n8085_ = ~new_n3600_ | ~pi0088;
  assign new_n8086_ = ~new_n4220_ | ~new_n3567_;
  assign new_n8087_ = ~new_n21494_ | ~new_n3556_;
  assign new_n8088_ = ~pi0462 | ~new_n4408_;
  assign new_n8089_ = ~new_n3604_ | ~pi0073;
  assign new_n8090_ = ~new_n3600_ | ~pi0089;
  assign new_n8091_ = ~new_n4221_ | ~new_n3567_;
  assign new_n8092_ = ~new_n21493_ | ~new_n3556_;
  assign new_n8093_ = ~pi0463 | ~new_n4408_;
  assign new_n8094_ = ~new_n3604_ | ~pi0074;
  assign new_n8095_ = ~new_n3600_ | ~pi0090;
  assign new_n8096_ = ~new_n4222_ | ~new_n3567_;
  assign new_n8097_ = ~new_n21491_ | ~new_n3556_;
  assign new_n8098_ = ~pi0464 | ~new_n4408_;
  assign new_n8099_ = ~new_n3604_ | ~pi0075;
  assign new_n8100_ = ~new_n3600_ | ~pi0091;
  assign new_n8101_ = ~new_n4223_ | ~new_n3567_;
  assign new_n8102_ = ~new_n21490_ | ~new_n3556_;
  assign new_n8103_ = ~pi0465 | ~new_n4408_;
  assign new_n8104_ = ~new_n3604_ | ~pi0076;
  assign new_n8105_ = ~new_n3600_ | ~pi0092;
  assign new_n8106_ = ~new_n4224_ | ~new_n3567_;
  assign new_n8107_ = ~new_n21489_ | ~new_n3556_;
  assign new_n8108_ = ~pi0466 | ~new_n4408_;
  assign new_n8109_ = ~new_n3604_ | ~pi0077;
  assign new_n8110_ = ~new_n3600_ | ~pi0093;
  assign new_n8111_ = ~new_n21649_ | ~new_n3567_;
  assign new_n8112_ = ~new_n21488_ | ~new_n3556_;
  assign new_n8113_ = ~pi0467 | ~new_n4408_;
  assign new_n8114_ = ~new_n3604_ | ~pi0078;
  assign new_n8115_ = ~new_n3600_ | ~pi0094;
  assign new_n8116_ = ~new_n21648_ | ~new_n3567_;
  assign new_n8117_ = ~new_n21487_ | ~new_n3556_;
  assign new_n8118_ = ~pi0468 | ~new_n4408_;
  assign new_n8119_ = ~new_n3604_ | ~pi0079;
  assign new_n8120_ = ~new_n3600_ | ~pi0095;
  assign new_n8121_ = ~new_n21647_ | ~new_n3567_;
  assign new_n8122_ = ~new_n21486_ | ~new_n3556_;
  assign new_n8123_ = ~pi0469 | ~new_n4408_;
  assign new_n8124_ = ~new_n3604_ | ~pi0080;
  assign new_n8125_ = ~new_n3600_ | ~pi0096;
  assign new_n8126_ = ~new_n21646_ | ~new_n3567_;
  assign new_n8127_ = ~new_n21485_ | ~new_n3556_;
  assign new_n8128_ = ~pi0470 | ~new_n4408_;
  assign new_n8129_ = ~new_n3604_ | ~pi0081;
  assign new_n8130_ = ~new_n3600_ | ~pi0097;
  assign new_n8131_ = ~new_n21645_ | ~new_n3567_;
  assign new_n8132_ = ~new_n21484_ | ~new_n3556_;
  assign new_n8133_ = ~pi0471 | ~new_n4408_;
  assign new_n8134_ = ~new_n3604_ | ~pi0082;
  assign new_n8135_ = ~new_n3600_ | ~pi0098;
  assign new_n8136_ = ~new_n21644_ | ~new_n3567_;
  assign new_n8137_ = ~new_n21483_ | ~new_n3556_;
  assign new_n8138_ = ~pi0472 | ~new_n4408_;
  assign new_n8139_ = ~new_n3604_ | ~pi0083;
  assign new_n8140_ = ~new_n3600_ | ~pi0099;
  assign new_n8141_ = ~new_n21643_ | ~new_n3567_;
  assign new_n8142_ = ~new_n21482_ | ~new_n3556_;
  assign new_n8143_ = ~pi0473 | ~new_n4408_;
  assign new_n8144_ = ~new_n3604_ | ~pi0084;
  assign new_n8145_ = ~new_n3600_ | ~pi0100;
  assign new_n8146_ = ~new_n21642_ | ~new_n3567_;
  assign new_n8147_ = ~new_n21480_ | ~new_n3556_;
  assign new_n8148_ = ~pi0474 | ~new_n4408_;
  assign new_n8149_ = ~new_n3600_ | ~pi0101;
  assign new_n8150_ = ~new_n21479_ | ~new_n3556_;
  assign new_n8151_ = ~pi0475 | ~new_n4408_;
  assign new_n8152_ = ~new_n21624_ | ~new_n5461_;
  assign new_n8153_ = ~new_n4398_ | ~new_n8152_;
  assign new_n8154_ = ~pi0306 | ~new_n3564_;
  assign new_n8155_ = ~new_n21228_ | ~new_n3555_;
  assign new_n8156_ = ~pi0476 | ~new_n4409_;
  assign new_n8157_ = ~pi0305 | ~new_n3564_;
  assign new_n8158_ = ~new_n21294_ | ~new_n3555_;
  assign new_n8159_ = ~pi0477 | ~new_n4409_;
  assign new_n8160_ = ~pi0304 | ~new_n3564_;
  assign new_n8161_ = ~new_n21283_ | ~new_n3555_;
  assign new_n8162_ = ~pi0478 | ~new_n4409_;
  assign new_n8163_ = ~pi0303 | ~new_n3564_;
  assign new_n8164_ = ~new_n21280_ | ~new_n3555_;
  assign new_n8165_ = ~pi0479 | ~new_n4409_;
  assign new_n8166_ = ~pi0302 | ~new_n3564_;
  assign new_n8167_ = ~new_n21279_ | ~new_n3555_;
  assign new_n8168_ = ~pi0480 | ~new_n4409_;
  assign new_n8169_ = ~pi0301 | ~new_n3564_;
  assign new_n8170_ = ~new_n21278_ | ~new_n3555_;
  assign new_n8171_ = ~pi0481 | ~new_n4409_;
  assign new_n8172_ = ~pi0300 | ~new_n3564_;
  assign new_n8173_ = ~new_n21277_ | ~new_n3555_;
  assign new_n8174_ = ~pi0482 | ~new_n4409_;
  assign new_n8175_ = ~pi0299 | ~new_n3564_;
  assign new_n8176_ = ~new_n21276_ | ~new_n3555_;
  assign new_n8177_ = ~pi0483 | ~new_n4409_;
  assign new_n8178_ = ~new_n3761_ | ~new_n3564_;
  assign new_n8179_ = ~new_n21275_ | ~new_n3555_;
  assign new_n8180_ = ~pi0484 | ~new_n4409_;
  assign new_n8181_ = ~new_n3762_ | ~new_n3564_;
  assign new_n8182_ = ~new_n21274_ | ~new_n3555_;
  assign new_n8183_ = ~pi0485 | ~new_n4409_;
  assign new_n8184_ = ~new_n3763_ | ~new_n3564_;
  assign new_n8185_ = ~new_n21304_ | ~new_n3555_;
  assign new_n8186_ = ~pi0486 | ~new_n4409_;
  assign new_n8187_ = ~new_n3764_ | ~new_n3564_;
  assign new_n8188_ = ~new_n21303_ | ~new_n3555_;
  assign new_n8189_ = ~pi0487 | ~new_n4409_;
  assign new_n8190_ = ~new_n3765_ | ~new_n3564_;
  assign new_n8191_ = ~new_n21302_ | ~new_n3555_;
  assign new_n8192_ = ~pi0488 | ~new_n4409_;
  assign new_n8193_ = ~new_n3766_ | ~new_n3564_;
  assign new_n8194_ = ~new_n21301_ | ~new_n3555_;
  assign new_n8195_ = ~pi0489 | ~new_n4409_;
  assign new_n8196_ = ~new_n3767_ | ~new_n3564_;
  assign new_n8197_ = ~new_n21300_ | ~new_n3555_;
  assign new_n8198_ = ~pi0490 | ~new_n4409_;
  assign new_n8199_ = ~new_n3768_ | ~new_n3564_;
  assign new_n8200_ = ~new_n21299_ | ~new_n3555_;
  assign new_n8201_ = ~pi0491 | ~new_n4409_;
  assign new_n8202_ = ~new_n4218_ | ~new_n3564_;
  assign new_n8203_ = ~new_n21298_ | ~new_n3555_;
  assign new_n8204_ = ~pi0492 | ~new_n4409_;
  assign new_n8205_ = ~new_n4219_ | ~new_n3564_;
  assign new_n8206_ = ~new_n21297_ | ~new_n3555_;
  assign new_n8207_ = ~pi0493 | ~new_n4409_;
  assign new_n8208_ = ~new_n4220_ | ~new_n3564_;
  assign new_n8209_ = ~new_n21296_ | ~new_n3555_;
  assign new_n8210_ = ~pi0494 | ~new_n4409_;
  assign new_n8211_ = ~new_n4221_ | ~new_n3564_;
  assign new_n8212_ = ~new_n21295_ | ~new_n3555_;
  assign new_n8213_ = ~pi0495 | ~new_n4409_;
  assign new_n8214_ = ~new_n4222_ | ~new_n3564_;
  assign new_n8215_ = ~new_n21293_ | ~new_n3555_;
  assign new_n8216_ = ~pi0496 | ~new_n4409_;
  assign new_n8217_ = ~new_n4223_ | ~new_n3564_;
  assign new_n8218_ = ~new_n21292_ | ~new_n3555_;
  assign new_n8219_ = ~pi0497 | ~new_n4409_;
  assign new_n8220_ = ~new_n4224_ | ~new_n3564_;
  assign new_n8221_ = ~new_n21291_ | ~new_n3555_;
  assign new_n8222_ = ~pi0498 | ~new_n4409_;
  assign new_n8223_ = ~new_n27527_ | ~new_n3564_;
  assign new_n8224_ = ~new_n21290_ | ~new_n3555_;
  assign new_n8225_ = ~pi0499 | ~new_n4409_;
  assign new_n8226_ = ~new_n27526_ | ~new_n3564_;
  assign new_n8227_ = ~new_n21289_ | ~new_n3555_;
  assign new_n8228_ = ~pi0500 | ~new_n4409_;
  assign new_n8229_ = ~new_n27525_ | ~new_n3564_;
  assign new_n8230_ = ~new_n21288_ | ~new_n3555_;
  assign new_n8231_ = ~pi0501 | ~new_n4409_;
  assign new_n8232_ = ~new_n27524_ | ~new_n3564_;
  assign new_n8233_ = ~new_n21287_ | ~new_n3555_;
  assign new_n8234_ = ~pi0502 | ~new_n4409_;
  assign new_n8235_ = ~new_n27523_ | ~new_n3564_;
  assign new_n8236_ = ~new_n21286_ | ~new_n3555_;
  assign new_n8237_ = ~pi0503 | ~new_n4409_;
  assign new_n8238_ = ~new_n27522_ | ~new_n3564_;
  assign new_n8239_ = ~new_n21285_ | ~new_n3555_;
  assign new_n8240_ = ~pi0504 | ~new_n4409_;
  assign new_n8241_ = ~new_n27521_ | ~new_n3564_;
  assign new_n8242_ = ~new_n21284_ | ~new_n3555_;
  assign new_n8243_ = ~pi0505 | ~new_n4409_;
  assign new_n8244_ = ~new_n27520_ | ~new_n3564_;
  assign new_n8245_ = ~new_n21282_ | ~new_n3555_;
  assign new_n8246_ = ~pi0506 | ~new_n4409_;
  assign new_n8247_ = ~new_n21281_ | ~new_n3555_;
  assign new_n8248_ = ~pi0507 | ~new_n4409_;
  assign new_n8249_ = ~new_n6644_ | ~new_n6647_;
  assign new_n8250_ = ~new_n4416_;
  assign new_n8251_ = ~new_n4413_;
  assign new_n8252_ = pi0547 | new_n2971_;
  assign new_n8253_ = ~pi0476 | ~new_n3758_;
  assign new_n8254_ = ~pi0508 | ~new_n3757_;
  assign new_n8255_ = ~pi0476 | ~new_n9066_;
  assign new_n8256_ = ~new_n22197_ | ~new_n3611_;
  assign new_n8257_ = ~new_n24659_ | ~new_n3610_;
  assign new_n8258_ = ~pi0508 | ~new_n3561_;
  assign new_n8259_ = ~new_n3559_ | ~pi0349;
  assign new_n8260_ = ~pi0349 | ~new_n5475_;
  assign new_n8261_ = ~new_n3557_ | ~pi0349;
  assign new_n8262_ = ~new_n8250_ | ~pi0508;
  assign new_n8263_ = ~new_n25151_ | ~new_n3758_;
  assign new_n8264_ = ~new_n22900_ | ~new_n3757_;
  assign new_n8265_ = ~pi0477 | ~new_n9066_;
  assign new_n8266_ = ~new_n22209_ | ~new_n3611_;
  assign new_n8267_ = ~new_n24671_ | ~new_n3610_;
  assign new_n8268_ = ~new_n23079_ | ~new_n3561_;
  assign new_n8269_ = ~new_n3559_ | ~new_n22223_;
  assign new_n8270_ = ~new_n22087_ | ~new_n5475_;
  assign new_n8271_ = ~new_n3557_ | ~pi0350;
  assign new_n8272_ = ~new_n8250_ | ~pi0509;
  assign new_n8273_ = ~new_n25118_ | ~new_n3758_;
  assign new_n8274_ = ~new_n22967_ | ~new_n3757_;
  assign new_n8275_ = ~pi0478 | ~new_n9066_;
  assign new_n8276_ = ~new_n22208_ | ~new_n3611_;
  assign new_n8277_ = ~new_n24670_ | ~new_n3610_;
  assign new_n8278_ = ~new_n23146_ | ~new_n3561_;
  assign new_n8279_ = ~new_n3559_ | ~new_n22290_;
  assign new_n8280_ = ~new_n22054_ | ~new_n5475_;
  assign new_n8281_ = ~new_n3557_ | ~pi0351;
  assign new_n8282_ = ~new_n8250_ | ~pi0510;
  assign new_n8283_ = ~new_n25160_ | ~new_n3758_;
  assign new_n8284_ = ~new_n22964_ | ~new_n3757_;
  assign new_n8285_ = ~pi0479 | ~new_n9066_;
  assign new_n8286_ = ~new_n22207_ | ~new_n3611_;
  assign new_n8287_ = ~new_n24669_ | ~new_n3610_;
  assign new_n8288_ = ~new_n23143_ | ~new_n3561_;
  assign new_n8289_ = ~new_n3559_ | ~new_n22287_;
  assign new_n8290_ = ~new_n22096_ | ~new_n5475_;
  assign new_n8291_ = ~new_n3557_ | ~pi0352;
  assign new_n8292_ = ~new_n8250_ | ~pi0511;
  assign new_n8293_ = ~new_n25119_ | ~new_n3758_;
  assign new_n8294_ = ~new_n22963_ | ~new_n3757_;
  assign new_n8295_ = ~pi0480 | ~new_n9066_;
  assign new_n8296_ = ~new_n22206_ | ~new_n3611_;
  assign new_n8297_ = ~new_n24668_ | ~new_n3610_;
  assign new_n8298_ = ~new_n23142_ | ~new_n3561_;
  assign new_n8299_ = ~new_n3559_ | ~new_n22286_;
  assign new_n8300_ = ~new_n22055_ | ~new_n5475_;
  assign new_n8301_ = ~new_n3557_ | ~pi0353;
  assign new_n8302_ = ~new_n8250_ | ~pi0512;
  assign new_n8303_ = ~new_n25158_ | ~new_n3758_;
  assign new_n8304_ = ~new_n22962_ | ~new_n3757_;
  assign new_n8305_ = ~pi0481 | ~new_n9066_;
  assign new_n8306_ = ~new_n22198_ | ~new_n3611_;
  assign new_n8307_ = ~new_n24660_ | ~new_n3610_;
  assign new_n8308_ = ~new_n23141_ | ~new_n3561_;
  assign new_n8309_ = ~new_n3559_ | ~new_n22285_;
  assign new_n8310_ = ~new_n22094_ | ~new_n5475_;
  assign new_n8311_ = ~new_n3557_ | ~pi0354;
  assign new_n8312_ = ~new_n8250_ | ~pi0513;
  assign new_n8313_ = ~new_n25120_ | ~new_n3758_;
  assign new_n8314_ = ~new_n22961_ | ~new_n3757_;
  assign new_n8315_ = ~pi0482 | ~new_n9066_;
  assign new_n8316_ = ~new_n23140_ | ~new_n3561_;
  assign new_n8317_ = ~new_n3559_ | ~new_n22284_;
  assign new_n8318_ = ~new_n22056_ | ~new_n5475_;
  assign new_n8319_ = ~new_n3557_ | ~pi0355;
  assign new_n8320_ = ~new_n8250_ | ~pi0514;
  assign new_n8321_ = ~new_n25156_ | ~new_n3758_;
  assign new_n8322_ = ~new_n22960_ | ~new_n3757_;
  assign new_n8323_ = ~pi0483 | ~new_n9066_;
  assign new_n8324_ = ~new_n23139_ | ~new_n3561_;
  assign new_n8325_ = ~new_n3559_ | ~new_n22283_;
  assign new_n8326_ = ~new_n22092_ | ~new_n5475_;
  assign new_n8327_ = ~new_n3557_ | ~pi0356;
  assign new_n8328_ = ~new_n8250_ | ~pi0515;
  assign new_n8329_ = ~new_n25121_ | ~new_n3758_;
  assign new_n8330_ = ~new_n22959_ | ~new_n3757_;
  assign new_n8331_ = ~pi0484 | ~new_n9066_;
  assign new_n8332_ = ~new_n23138_ | ~new_n3561_;
  assign new_n8333_ = ~new_n3559_ | ~new_n22282_;
  assign new_n8334_ = ~new_n22057_ | ~new_n5475_;
  assign new_n8335_ = ~new_n3557_ | ~pi0357;
  assign new_n8336_ = ~new_n8250_ | ~pi0516;
  assign new_n8337_ = ~new_n25154_ | ~new_n3758_;
  assign new_n8338_ = ~new_n22958_ | ~new_n3757_;
  assign new_n8339_ = ~pi0485 | ~new_n9066_;
  assign new_n8340_ = ~new_n23137_ | ~new_n3561_;
  assign new_n8341_ = ~new_n3559_ | ~new_n22281_;
  assign new_n8342_ = ~new_n22090_ | ~new_n5475_;
  assign new_n8343_ = ~new_n3557_ | ~pi0358;
  assign new_n8344_ = ~new_n8250_ | ~pi0517;
  assign new_n8345_ = ~new_n25107_ | ~new_n3758_;
  assign new_n8346_ = ~new_n22987_ | ~new_n3757_;
  assign new_n8347_ = ~pi0486 | ~new_n9066_;
  assign new_n8348_ = ~new_n23166_ | ~new_n3561_;
  assign new_n8349_ = ~new_n3559_ | ~new_n22310_;
  assign new_n8350_ = ~new_n22043_ | ~new_n5475_;
  assign new_n8351_ = ~new_n3557_ | ~pi0359;
  assign new_n8352_ = ~new_n8250_ | ~pi0518;
  assign new_n8353_ = ~new_n25183_ | ~new_n3758_;
  assign new_n8354_ = ~new_n22986_ | ~new_n3757_;
  assign new_n8355_ = ~pi0487 | ~new_n9066_;
  assign new_n8356_ = ~new_n23165_ | ~new_n3561_;
  assign new_n8357_ = ~new_n3559_ | ~new_n22309_;
  assign new_n8358_ = ~new_n22119_ | ~new_n5475_;
  assign new_n8359_ = ~new_n3557_ | ~pi0360;
  assign new_n8360_ = ~new_n8250_ | ~pi0519;
  assign new_n8361_ = ~new_n25108_ | ~new_n3758_;
  assign new_n8362_ = ~new_n22985_ | ~new_n3757_;
  assign new_n8363_ = ~pi0488 | ~new_n9066_;
  assign new_n8364_ = ~new_n23164_ | ~new_n3561_;
  assign new_n8365_ = ~new_n3559_ | ~new_n22308_;
  assign new_n8366_ = ~new_n22044_ | ~new_n5475_;
  assign new_n8367_ = ~new_n3557_ | ~pi0361;
  assign new_n8368_ = ~new_n8250_ | ~pi0520;
  assign new_n8369_ = ~new_n25181_ | ~new_n3758_;
  assign new_n8370_ = ~new_n22984_ | ~new_n3757_;
  assign new_n8371_ = ~pi0489 | ~new_n9066_;
  assign new_n8372_ = ~new_n23163_ | ~new_n3561_;
  assign new_n8373_ = ~new_n3559_ | ~new_n22307_;
  assign new_n8374_ = ~new_n22117_ | ~new_n5475_;
  assign new_n8375_ = ~new_n3557_ | ~pi0362;
  assign new_n8376_ = ~new_n8250_ | ~pi0521;
  assign new_n8377_ = ~new_n25109_ | ~new_n3758_;
  assign new_n8378_ = ~new_n22983_ | ~new_n3757_;
  assign new_n8379_ = ~pi0490 | ~new_n9066_;
  assign new_n8380_ = ~new_n23162_ | ~new_n3561_;
  assign new_n8381_ = ~new_n3559_ | ~new_n22306_;
  assign new_n8382_ = ~new_n22045_ | ~new_n5475_;
  assign new_n8383_ = ~new_n3557_ | ~pi0363;
  assign new_n8384_ = ~new_n8250_ | ~pi0522;
  assign new_n8385_ = ~new_n25179_ | ~new_n3758_;
  assign new_n8386_ = ~new_n22982_ | ~new_n3757_;
  assign new_n8387_ = ~pi0491 | ~new_n9066_;
  assign new_n8388_ = ~new_n23161_ | ~new_n3561_;
  assign new_n8389_ = ~new_n3559_ | ~new_n22305_;
  assign new_n8390_ = ~new_n22115_ | ~new_n5475_;
  assign new_n8391_ = ~new_n3557_ | ~pi0364;
  assign new_n8392_ = ~new_n8250_ | ~pi0523;
  assign new_n8393_ = ~new_n25110_ | ~new_n3758_;
  assign new_n8394_ = ~new_n22981_ | ~new_n3757_;
  assign new_n8395_ = ~pi0492 | ~new_n9066_;
  assign new_n8396_ = ~new_n23160_ | ~new_n3561_;
  assign new_n8397_ = ~new_n3559_ | ~new_n22304_;
  assign new_n8398_ = ~new_n22046_ | ~new_n5475_;
  assign new_n8399_ = ~new_n3557_ | ~pi0365;
  assign new_n8400_ = ~new_n8250_ | ~pi0524;
  assign new_n8401_ = ~new_n25177_ | ~new_n3758_;
  assign new_n8402_ = ~new_n22980_ | ~new_n3757_;
  assign new_n8403_ = ~pi0493 | ~new_n9066_;
  assign new_n8404_ = ~new_n23159_ | ~new_n3561_;
  assign new_n8405_ = ~new_n3559_ | ~new_n22303_;
  assign new_n8406_ = ~new_n22113_ | ~new_n5475_;
  assign new_n8407_ = ~new_n3557_ | ~pi0366;
  assign new_n8408_ = ~new_n8250_ | ~pi0525;
  assign new_n8409_ = ~new_n25111_ | ~new_n3758_;
  assign new_n8410_ = ~new_n22979_ | ~new_n3757_;
  assign new_n8411_ = ~pi0494 | ~new_n9066_;
  assign new_n8412_ = ~new_n23158_ | ~new_n3561_;
  assign new_n8413_ = ~new_n3559_ | ~new_n22302_;
  assign new_n8414_ = ~new_n22047_ | ~new_n5475_;
  assign new_n8415_ = ~new_n3557_ | ~pi0367;
  assign new_n8416_ = ~new_n8250_ | ~pi0526;
  assign new_n8417_ = ~new_n25175_ | ~new_n3758_;
  assign new_n8418_ = ~new_n22978_ | ~new_n3757_;
  assign new_n8419_ = ~pi0495 | ~new_n9066_;
  assign new_n8420_ = ~new_n23157_ | ~new_n3561_;
  assign new_n8421_ = ~new_n3559_ | ~new_n22301_;
  assign new_n8422_ = ~new_n22111_ | ~new_n5475_;
  assign new_n8423_ = ~new_n3557_ | ~pi0368;
  assign new_n8424_ = ~new_n8250_ | ~pi0527;
  assign new_n8425_ = ~new_n25112_ | ~new_n3758_;
  assign new_n8426_ = ~new_n22977_ | ~new_n3757_;
  assign new_n8427_ = ~pi0496 | ~new_n9066_;
  assign new_n8428_ = ~new_n23156_ | ~new_n3561_;
  assign new_n8429_ = ~new_n3559_ | ~new_n22300_;
  assign new_n8430_ = ~new_n22048_ | ~new_n5475_;
  assign new_n8431_ = ~new_n3557_ | ~pi0369;
  assign new_n8432_ = ~new_n8250_ | ~pi0528;
  assign new_n8433_ = ~new_n25171_ | ~new_n3758_;
  assign new_n8434_ = ~new_n22976_ | ~new_n3757_;
  assign new_n8435_ = ~pi0497 | ~new_n9066_;
  assign new_n8436_ = ~new_n23155_ | ~new_n3561_;
  assign new_n8437_ = ~new_n3559_ | ~new_n22299_;
  assign new_n8438_ = ~new_n22107_ | ~new_n5475_;
  assign new_n8439_ = ~new_n3557_ | ~pi0370;
  assign new_n8440_ = ~new_n8250_ | ~pi0529;
  assign new_n8441_ = ~new_n25113_ | ~new_n3758_;
  assign new_n8442_ = ~new_n22975_ | ~new_n3757_;
  assign new_n8443_ = ~pi0498 | ~new_n9066_;
  assign new_n8444_ = ~new_n23154_ | ~new_n3561_;
  assign new_n8445_ = ~new_n3559_ | ~new_n22298_;
  assign new_n8446_ = ~new_n22049_ | ~new_n5475_;
  assign new_n8447_ = ~new_n3557_ | ~pi0371;
  assign new_n8448_ = ~new_n8250_ | ~pi0530;
  assign new_n8449_ = ~new_n25169_ | ~new_n3758_;
  assign new_n8450_ = ~new_n22974_ | ~new_n3757_;
  assign new_n8451_ = ~pi0499 | ~new_n9066_;
  assign new_n8452_ = ~new_n23153_ | ~new_n3561_;
  assign new_n8453_ = ~new_n3559_ | ~new_n22297_;
  assign new_n8454_ = ~new_n22105_ | ~new_n5475_;
  assign new_n8455_ = ~new_n3557_ | ~pi0372;
  assign new_n8456_ = ~new_n8250_ | ~pi0531;
  assign new_n8457_ = ~new_n25114_ | ~new_n3758_;
  assign new_n8458_ = ~new_n22973_ | ~new_n3757_;
  assign new_n8459_ = ~pi0500 | ~new_n9066_;
  assign new_n8460_ = ~new_n23152_ | ~new_n3561_;
  assign new_n8461_ = ~new_n3559_ | ~new_n22296_;
  assign new_n8462_ = ~new_n22050_ | ~new_n5475_;
  assign new_n8463_ = ~new_n3557_ | ~pi0373;
  assign new_n8464_ = ~new_n8250_ | ~pi0532;
  assign new_n8465_ = ~new_n25167_ | ~new_n3758_;
  assign new_n8466_ = ~new_n22972_ | ~new_n3757_;
  assign new_n8467_ = ~pi0501 | ~new_n9066_;
  assign new_n8468_ = ~new_n23151_ | ~new_n3561_;
  assign new_n8469_ = ~new_n3559_ | ~new_n22295_;
  assign new_n8470_ = ~new_n22103_ | ~new_n5475_;
  assign new_n8471_ = ~new_n3557_ | ~pi0374;
  assign new_n8472_ = ~new_n8250_ | ~pi0533;
  assign new_n8473_ = ~new_n25115_ | ~new_n3758_;
  assign new_n8474_ = ~new_n22971_ | ~new_n3757_;
  assign new_n8475_ = ~pi0502 | ~new_n9066_;
  assign new_n8476_ = ~new_n23150_ | ~new_n3561_;
  assign new_n8477_ = ~new_n3559_ | ~new_n22294_;
  assign new_n8478_ = ~new_n22051_ | ~new_n5475_;
  assign new_n8479_ = ~new_n3557_ | ~pi0375;
  assign new_n8480_ = ~new_n8250_ | ~pi0534;
  assign new_n8481_ = ~new_n25165_ | ~new_n3758_;
  assign new_n8482_ = ~new_n22970_ | ~new_n3757_;
  assign new_n8483_ = ~pi0503 | ~new_n9066_;
  assign new_n8484_ = ~new_n23149_ | ~new_n3561_;
  assign new_n8485_ = ~new_n3559_ | ~new_n22293_;
  assign new_n8486_ = ~new_n22101_ | ~new_n5475_;
  assign new_n8487_ = ~new_n3557_ | ~pi0376;
  assign new_n8488_ = ~new_n8250_ | ~pi0535;
  assign new_n8489_ = ~new_n25116_ | ~new_n3758_;
  assign new_n8490_ = ~new_n22969_ | ~new_n3757_;
  assign new_n8491_ = ~pi0504 | ~new_n9066_;
  assign new_n8492_ = ~new_n23148_ | ~new_n3561_;
  assign new_n8493_ = ~new_n3559_ | ~new_n22292_;
  assign new_n8494_ = ~new_n22052_ | ~new_n5475_;
  assign new_n8495_ = ~new_n3557_ | ~pi0377;
  assign new_n8496_ = ~new_n8250_ | ~pi0536;
  assign new_n8497_ = ~new_n25117_ | ~new_n3758_;
  assign new_n8498_ = ~new_n22968_ | ~new_n3757_;
  assign new_n8499_ = ~pi0505 | ~new_n9066_;
  assign new_n8500_ = ~new_n23147_ | ~new_n3561_;
  assign new_n8501_ = ~new_n3559_ | ~new_n22291_;
  assign new_n8502_ = ~new_n22053_ | ~new_n5475_;
  assign new_n8503_ = ~new_n3557_ | ~pi0378;
  assign new_n8504_ = ~new_n8250_ | ~pi0537;
  assign new_n8505_ = ~new_n25163_ | ~new_n3758_;
  assign new_n8506_ = ~new_n22966_ | ~new_n3757_;
  assign new_n8507_ = ~pi0506 | ~new_n9066_;
  assign new_n8508_ = ~new_n23145_ | ~new_n3561_;
  assign new_n8509_ = ~new_n3559_ | ~new_n22289_;
  assign new_n8510_ = ~new_n22099_ | ~new_n5475_;
  assign new_n8511_ = ~new_n3557_ | ~pi0379;
  assign new_n8512_ = ~new_n8250_ | ~pi0538;
  assign new_n8513_ = ~new_n5291_ | ~new_n3759_;
  assign new_n8514_ = ~new_n25152_ | ~new_n3758_;
  assign new_n8515_ = ~new_n22965_ | ~new_n3757_;
  assign new_n8516_ = ~pi0507 | ~new_n9066_;
  assign new_n8517_ = ~new_n23144_ | ~new_n3561_;
  assign new_n8518_ = ~new_n3559_ | ~new_n22288_;
  assign new_n8519_ = ~new_n8518_;
  assign new_n8520_ = ~new_n3557_ | ~pi0380;
  assign new_n8521_ = ~new_n8250_ | ~pi0539;
  assign new_n8522_ = ~pi0144 | ~pi0143;
  assign new_n8523_ = pi0509 | pi0508;
  assign new_n8524_ = ~new_n5441_;
  assign new_n8525_ = ~pi0545 | ~new_n5441_;
  assign new_n8526_ = ~new_n5779_ | ~new_n3546_;
  assign new_n8527_ = ~new_n3609_ | ~new_n3786_;
  assign new_n8528_ = ~new_n4279_ | ~new_n8527_;
  assign new_n8529_ = ~new_n8528_ | ~new_n4277_;
  assign new_n8530_ = ~new_n5443_;
  assign new_n8531_ = ~new_n5452_ | ~new_n3787_;
  assign new_n8532_ = ~new_n4268_ | ~new_n4274_;
  assign new_n8533_ = ~new_n5306_ | ~pi0176 | ~new_n9075_;
  assign new_n8534_ = ~pi0178 | ~new_n8533_;
  assign new_n8535_ = ~new_n4281_ | ~new_n8534_;
  assign new_n8536_ = ~new_n3546_ | ~new_n3760_;
  assign new_n8537_ = ~pi0551 | ~new_n8536_;
  assign new_n8538_ = ~new_n5503_ | ~pi0178;
  assign new_n8539_ = ~pi0552 | ~pi0142;
  assign new_n8540_ = ~new_n5444_;
  assign new_n8541_ = ~new_n4270_ | ~pi0176 | ~new_n4267_;
  assign new_n8542_ = ~new_n5644_ | ~pi0176;
  assign new_n8543_ = ~new_n3698_ | ~pi0179;
  assign new_n8544_ = ~new_n3697_ | ~pi0187;
  assign new_n8545_ = ~new_n3696_ | ~pi0195;
  assign new_n8546_ = ~new_n3695_ | ~pi0203;
  assign new_n8547_ = ~new_n3693_ | ~pi0211;
  assign new_n8548_ = ~new_n3692_ | ~pi0219;
  assign new_n8549_ = ~new_n3691_ | ~pi0227;
  assign new_n8550_ = ~new_n3690_ | ~pi0235;
  assign new_n8551_ = ~new_n3688_ | ~pi0243;
  assign new_n8552_ = ~new_n3687_ | ~pi0251;
  assign new_n8553_ = ~new_n3686_ | ~pi0259;
  assign new_n8554_ = ~new_n3685_ | ~pi0267;
  assign new_n8555_ = ~new_n3683_ | ~pi0275;
  assign new_n8556_ = ~new_n3681_ | ~pi0283;
  assign new_n8557_ = ~new_n3679_ | ~pi0291;
  assign new_n8558_ = ~new_n3677_ | ~pi0299;
  assign new_n8559_ = ~new_n3698_ | ~pi0180;
  assign new_n8560_ = ~new_n3697_ | ~pi0188;
  assign new_n8561_ = ~new_n3696_ | ~pi0196;
  assign new_n8562_ = ~new_n3695_ | ~pi0204;
  assign new_n8563_ = ~new_n3693_ | ~pi0212;
  assign new_n8564_ = ~new_n3692_ | ~pi0220;
  assign new_n8565_ = ~new_n3691_ | ~pi0228;
  assign new_n8566_ = ~new_n3690_ | ~pi0236;
  assign new_n8567_ = ~new_n3688_ | ~pi0244;
  assign new_n8568_ = ~new_n3687_ | ~pi0252;
  assign new_n8569_ = ~new_n3686_ | ~pi0260;
  assign new_n8570_ = ~new_n3685_ | ~pi0268;
  assign new_n8571_ = ~new_n3683_ | ~pi0276;
  assign new_n8572_ = ~new_n3681_ | ~pi0284;
  assign new_n8573_ = ~new_n3679_ | ~pi0292;
  assign new_n8574_ = ~new_n3677_ | ~pi0300;
  assign new_n8575_ = ~new_n3698_ | ~pi0181;
  assign new_n8576_ = ~new_n3697_ | ~pi0189;
  assign new_n8577_ = ~new_n3696_ | ~pi0197;
  assign new_n8578_ = ~new_n3695_ | ~pi0205;
  assign new_n8579_ = ~new_n3693_ | ~pi0213;
  assign new_n8580_ = ~new_n3692_ | ~pi0221;
  assign new_n8581_ = ~new_n3691_ | ~pi0229;
  assign new_n8582_ = ~new_n3690_ | ~pi0237;
  assign new_n8583_ = ~new_n3688_ | ~pi0245;
  assign new_n8584_ = ~new_n3687_ | ~pi0253;
  assign new_n8585_ = ~new_n3686_ | ~pi0261;
  assign new_n8586_ = ~new_n3685_ | ~pi0269;
  assign new_n8587_ = ~new_n3683_ | ~pi0277;
  assign new_n8588_ = ~new_n3681_ | ~pi0285;
  assign new_n8589_ = ~new_n3679_ | ~pi0293;
  assign new_n8590_ = ~new_n3677_ | ~pi0301;
  assign new_n8591_ = ~new_n3698_ | ~pi0182;
  assign new_n8592_ = ~new_n3697_ | ~pi0190;
  assign new_n8593_ = ~new_n3696_ | ~pi0198;
  assign new_n8594_ = ~new_n3695_ | ~pi0206;
  assign new_n8595_ = ~new_n3693_ | ~pi0214;
  assign new_n8596_ = ~new_n3692_ | ~pi0222;
  assign new_n8597_ = ~new_n3691_ | ~pi0230;
  assign new_n8598_ = ~new_n3690_ | ~pi0238;
  assign new_n8599_ = ~new_n3688_ | ~pi0246;
  assign new_n8600_ = ~new_n3687_ | ~pi0254;
  assign new_n8601_ = ~new_n3686_ | ~pi0262;
  assign new_n8602_ = ~new_n3685_ | ~pi0270;
  assign new_n8603_ = ~new_n3683_ | ~pi0278;
  assign new_n8604_ = ~new_n3681_ | ~pi0286;
  assign new_n8605_ = ~new_n3679_ | ~pi0294;
  assign new_n8606_ = ~new_n3677_ | ~pi0302;
  assign new_n8607_ = ~new_n3698_ | ~pi0183;
  assign new_n8608_ = ~new_n3697_ | ~pi0191;
  assign new_n8609_ = ~new_n3696_ | ~pi0199;
  assign new_n8610_ = ~new_n3695_ | ~pi0207;
  assign new_n8611_ = ~new_n3693_ | ~pi0215;
  assign new_n8612_ = ~new_n3692_ | ~pi0223;
  assign new_n8613_ = ~new_n3691_ | ~pi0231;
  assign new_n8614_ = ~new_n3690_ | ~pi0239;
  assign new_n8615_ = ~new_n3688_ | ~pi0247;
  assign new_n8616_ = ~new_n3687_ | ~pi0255;
  assign new_n8617_ = ~new_n3686_ | ~pi0263;
  assign new_n8618_ = ~new_n3685_ | ~pi0271;
  assign new_n8619_ = ~new_n3683_ | ~pi0279;
  assign new_n8620_ = ~new_n3681_ | ~pi0287;
  assign new_n8621_ = ~new_n3679_ | ~pi0295;
  assign new_n8622_ = ~new_n3677_ | ~pi0303;
  assign new_n8623_ = ~new_n3698_ | ~pi0184;
  assign new_n8624_ = ~new_n3697_ | ~pi0192;
  assign new_n8625_ = ~new_n3696_ | ~pi0200;
  assign new_n8626_ = ~new_n3695_ | ~pi0208;
  assign new_n8627_ = ~new_n3693_ | ~pi0216;
  assign new_n8628_ = ~new_n3692_ | ~pi0224;
  assign new_n8629_ = ~new_n3691_ | ~pi0232;
  assign new_n8630_ = ~new_n3690_ | ~pi0240;
  assign new_n8631_ = ~new_n3688_ | ~pi0248;
  assign new_n8632_ = ~new_n3687_ | ~pi0256;
  assign new_n8633_ = ~new_n3686_ | ~pi0264;
  assign new_n8634_ = ~new_n3685_ | ~pi0272;
  assign new_n8635_ = ~new_n3683_ | ~pi0280;
  assign new_n8636_ = ~new_n3681_ | ~pi0288;
  assign new_n8637_ = ~new_n3679_ | ~pi0296;
  assign new_n8638_ = ~new_n3677_ | ~pi0304;
  assign new_n8639_ = ~new_n3698_ | ~pi0185;
  assign new_n8640_ = ~new_n3697_ | ~pi0193;
  assign new_n8641_ = ~new_n3696_ | ~pi0201;
  assign new_n8642_ = ~new_n3695_ | ~pi0209;
  assign new_n8643_ = ~new_n3693_ | ~pi0217;
  assign new_n8644_ = ~new_n3692_ | ~pi0225;
  assign new_n8645_ = ~new_n3691_ | ~pi0233;
  assign new_n8646_ = ~new_n3690_ | ~pi0241;
  assign new_n8647_ = ~new_n3688_ | ~pi0249;
  assign new_n8648_ = ~new_n3687_ | ~pi0257;
  assign new_n8649_ = ~new_n3686_ | ~pi0265;
  assign new_n8650_ = ~new_n3685_ | ~pi0273;
  assign new_n8651_ = ~new_n3683_ | ~pi0281;
  assign new_n8652_ = ~new_n3681_ | ~pi0289;
  assign new_n8653_ = ~new_n3679_ | ~pi0297;
  assign new_n8654_ = ~new_n3677_ | ~pi0305;
  assign new_n8655_ = ~new_n3698_ | ~pi0186;
  assign new_n8656_ = ~new_n3697_ | ~pi0194;
  assign new_n8657_ = ~new_n3696_ | ~pi0202;
  assign new_n8658_ = ~new_n3695_ | ~pi0210;
  assign new_n8659_ = ~new_n3693_ | ~pi0218;
  assign new_n8660_ = ~new_n3692_ | ~pi0226;
  assign new_n8661_ = ~new_n3691_ | ~pi0234;
  assign new_n8662_ = ~new_n3690_ | ~pi0242;
  assign new_n8663_ = ~new_n3688_ | ~pi0250;
  assign new_n8664_ = ~new_n3687_ | ~pi0258;
  assign new_n8665_ = ~new_n3686_ | ~pi0266;
  assign new_n8666_ = ~new_n3685_ | ~pi0274;
  assign new_n8667_ = ~new_n3683_ | ~pi0282;
  assign new_n8668_ = ~new_n3681_ | ~pi0290;
  assign new_n8669_ = ~new_n3679_ | ~pi0298;
  assign new_n8670_ = ~new_n3677_ | ~pi0306;
  assign new_n8671_ = ~new_n5626_ | ~pi0310;
  assign new_n8672_ = ~new_n4422_;
  assign new_n8673_ = ~new_n3718_ | ~pi0299;
  assign new_n8674_ = ~new_n3717_ | ~pi0291;
  assign new_n8675_ = ~new_n3716_ | ~pi0283;
  assign new_n8676_ = ~new_n3715_ | ~pi0275;
  assign new_n8677_ = ~new_n3713_ | ~pi0267;
  assign new_n8678_ = ~new_n3712_ | ~pi0259;
  assign new_n8679_ = ~new_n3711_ | ~pi0251;
  assign new_n8680_ = ~new_n3710_ | ~pi0243;
  assign new_n8681_ = ~new_n3708_ | ~pi0235;
  assign new_n8682_ = ~new_n3707_ | ~pi0227;
  assign new_n8683_ = ~new_n3706_ | ~pi0219;
  assign new_n8684_ = ~new_n3705_ | ~pi0211;
  assign new_n8685_ = ~new_n3703_ | ~pi0203;
  assign new_n8686_ = ~new_n3702_ | ~pi0195;
  assign new_n8687_ = ~new_n3701_ | ~pi0187;
  assign new_n8688_ = ~new_n3700_ | ~pi0179;
  assign new_n8689_ = ~new_n3718_ | ~pi0300;
  assign new_n8690_ = ~new_n3717_ | ~pi0292;
  assign new_n8691_ = ~new_n3716_ | ~pi0284;
  assign new_n8692_ = ~new_n3715_ | ~pi0276;
  assign new_n8693_ = ~new_n3713_ | ~pi0268;
  assign new_n8694_ = ~new_n3712_ | ~pi0260;
  assign new_n8695_ = ~new_n3711_ | ~pi0252;
  assign new_n8696_ = ~new_n3710_ | ~pi0244;
  assign new_n8697_ = ~new_n3708_ | ~pi0236;
  assign new_n8698_ = ~new_n3707_ | ~pi0228;
  assign new_n8699_ = ~new_n3706_ | ~pi0220;
  assign new_n8700_ = ~new_n3705_ | ~pi0212;
  assign new_n8701_ = ~new_n3703_ | ~pi0204;
  assign new_n8702_ = ~new_n3702_ | ~pi0196;
  assign new_n8703_ = ~new_n3701_ | ~pi0188;
  assign new_n8704_ = ~new_n3700_ | ~pi0180;
  assign new_n8705_ = ~new_n3718_ | ~pi0301;
  assign new_n8706_ = ~new_n3717_ | ~pi0293;
  assign new_n8707_ = ~new_n3716_ | ~pi0285;
  assign new_n8708_ = ~new_n3715_ | ~pi0277;
  assign new_n8709_ = ~new_n3713_ | ~pi0269;
  assign new_n8710_ = ~new_n3712_ | ~pi0261;
  assign new_n8711_ = ~new_n3711_ | ~pi0253;
  assign new_n8712_ = ~new_n3710_ | ~pi0245;
  assign new_n8713_ = ~new_n3708_ | ~pi0237;
  assign new_n8714_ = ~new_n3707_ | ~pi0229;
  assign new_n8715_ = ~new_n3706_ | ~pi0221;
  assign new_n8716_ = ~new_n3705_ | ~pi0213;
  assign new_n8717_ = ~new_n3703_ | ~pi0205;
  assign new_n8718_ = ~new_n3702_ | ~pi0197;
  assign new_n8719_ = ~new_n3701_ | ~pi0189;
  assign new_n8720_ = ~new_n3700_ | ~pi0181;
  assign new_n8721_ = ~new_n3718_ | ~pi0302;
  assign new_n8722_ = ~new_n3717_ | ~pi0294;
  assign new_n8723_ = ~new_n3716_ | ~pi0286;
  assign new_n8724_ = ~new_n3715_ | ~pi0278;
  assign new_n8725_ = ~new_n3713_ | ~pi0270;
  assign new_n8726_ = ~new_n3712_ | ~pi0262;
  assign new_n8727_ = ~new_n3711_ | ~pi0254;
  assign new_n8728_ = ~new_n3710_ | ~pi0246;
  assign new_n8729_ = ~new_n3708_ | ~pi0238;
  assign new_n8730_ = ~new_n3707_ | ~pi0230;
  assign new_n8731_ = ~new_n3706_ | ~pi0222;
  assign new_n8732_ = ~new_n3705_ | ~pi0214;
  assign new_n8733_ = ~new_n3703_ | ~pi0206;
  assign new_n8734_ = ~new_n3702_ | ~pi0198;
  assign new_n8735_ = ~new_n3701_ | ~pi0190;
  assign new_n8736_ = ~new_n3700_ | ~pi0182;
  assign new_n8737_ = ~new_n3718_ | ~pi0303;
  assign new_n8738_ = ~new_n3717_ | ~pi0295;
  assign new_n8739_ = ~new_n3716_ | ~pi0287;
  assign new_n8740_ = ~new_n3715_ | ~pi0279;
  assign new_n8741_ = ~new_n3713_ | ~pi0271;
  assign new_n8742_ = ~new_n3712_ | ~pi0263;
  assign new_n8743_ = ~new_n3711_ | ~pi0255;
  assign new_n8744_ = ~new_n3710_ | ~pi0247;
  assign new_n8745_ = ~new_n3708_ | ~pi0239;
  assign new_n8746_ = ~new_n3707_ | ~pi0231;
  assign new_n8747_ = ~new_n3706_ | ~pi0223;
  assign new_n8748_ = ~new_n3705_ | ~pi0215;
  assign new_n8749_ = ~new_n3703_ | ~pi0207;
  assign new_n8750_ = ~new_n3702_ | ~pi0199;
  assign new_n8751_ = ~new_n3701_ | ~pi0191;
  assign new_n8752_ = ~new_n3700_ | ~pi0183;
  assign new_n8753_ = ~new_n3718_ | ~pi0304;
  assign new_n8754_ = ~new_n3717_ | ~pi0296;
  assign new_n8755_ = ~new_n3716_ | ~pi0288;
  assign new_n8756_ = ~new_n3715_ | ~pi0280;
  assign new_n8757_ = ~new_n3713_ | ~pi0272;
  assign new_n8758_ = ~new_n3712_ | ~pi0264;
  assign new_n8759_ = ~new_n3711_ | ~pi0256;
  assign new_n8760_ = ~new_n3710_ | ~pi0248;
  assign new_n8761_ = ~new_n3708_ | ~pi0240;
  assign new_n8762_ = ~new_n3707_ | ~pi0232;
  assign new_n8763_ = ~new_n3706_ | ~pi0224;
  assign new_n8764_ = ~new_n3705_ | ~pi0216;
  assign new_n8765_ = ~new_n3703_ | ~pi0208;
  assign new_n8766_ = ~new_n3702_ | ~pi0200;
  assign new_n8767_ = ~new_n3701_ | ~pi0192;
  assign new_n8768_ = ~new_n3700_ | ~pi0184;
  assign new_n8769_ = ~new_n3718_ | ~pi0305;
  assign new_n8770_ = ~new_n3717_ | ~pi0297;
  assign new_n8771_ = ~new_n3716_ | ~pi0289;
  assign new_n8772_ = ~new_n3715_ | ~pi0281;
  assign new_n8773_ = ~new_n3713_ | ~pi0273;
  assign new_n8774_ = ~new_n3712_ | ~pi0265;
  assign new_n8775_ = ~new_n3711_ | ~pi0257;
  assign new_n8776_ = ~new_n3710_ | ~pi0249;
  assign new_n8777_ = ~new_n3708_ | ~pi0241;
  assign new_n8778_ = ~new_n3707_ | ~pi0233;
  assign new_n8779_ = ~new_n3706_ | ~pi0225;
  assign new_n8780_ = ~new_n3705_ | ~pi0217;
  assign new_n8781_ = ~new_n3703_ | ~pi0209;
  assign new_n8782_ = ~new_n3702_ | ~pi0201;
  assign new_n8783_ = ~new_n3701_ | ~pi0193;
  assign new_n8784_ = ~new_n3700_ | ~pi0185;
  assign new_n8785_ = ~new_n3718_ | ~pi0306;
  assign new_n8786_ = ~new_n3717_ | ~pi0298;
  assign new_n8787_ = ~new_n3716_ | ~pi0290;
  assign new_n8788_ = ~new_n3715_ | ~pi0282;
  assign new_n8789_ = ~new_n3713_ | ~pi0274;
  assign new_n8790_ = ~new_n3712_ | ~pi0266;
  assign new_n8791_ = ~new_n3711_ | ~pi0258;
  assign new_n8792_ = ~new_n3710_ | ~pi0250;
  assign new_n8793_ = ~new_n3708_ | ~pi0242;
  assign new_n8794_ = ~new_n3707_ | ~pi0234;
  assign new_n8795_ = ~new_n3706_ | ~pi0226;
  assign new_n8796_ = ~new_n3705_ | ~pi0218;
  assign new_n8797_ = ~new_n3703_ | ~pi0210;
  assign new_n8798_ = ~new_n3702_ | ~pi0202;
  assign new_n8799_ = ~new_n3701_ | ~pi0194;
  assign new_n8800_ = ~new_n3700_ | ~pi0186;
  assign new_n8801_ = ~new_n5445_;
  assign new_n8802_ = ~new_n3738_ | ~pi0235;
  assign new_n8803_ = ~new_n3737_ | ~pi0227;
  assign new_n8804_ = ~new_n3736_ | ~pi0219;
  assign new_n8805_ = ~new_n3735_ | ~pi0211;
  assign new_n8806_ = ~new_n3733_ | ~pi0203;
  assign new_n8807_ = ~new_n3732_ | ~pi0195;
  assign new_n8808_ = ~new_n3731_ | ~pi0187;
  assign new_n8809_ = ~new_n3730_ | ~pi0179;
  assign new_n8810_ = ~new_n3728_ | ~pi0299;
  assign new_n8811_ = ~new_n3727_ | ~pi0291;
  assign new_n8812_ = ~new_n3726_ | ~pi0283;
  assign new_n8813_ = ~new_n3725_ | ~pi0275;
  assign new_n8814_ = ~new_n3723_ | ~pi0267;
  assign new_n8815_ = ~new_n3722_ | ~pi0259;
  assign new_n8816_ = ~new_n3721_ | ~pi0251;
  assign new_n8817_ = ~new_n3720_ | ~pi0243;
  assign new_n8818_ = ~new_n3738_ | ~pi0236;
  assign new_n8819_ = ~new_n3737_ | ~pi0228;
  assign new_n8820_ = ~new_n3736_ | ~pi0220;
  assign new_n8821_ = ~new_n3735_ | ~pi0212;
  assign new_n8822_ = ~new_n3733_ | ~pi0204;
  assign new_n8823_ = ~new_n3732_ | ~pi0196;
  assign new_n8824_ = ~new_n3731_ | ~pi0188;
  assign new_n8825_ = ~new_n3730_ | ~pi0180;
  assign new_n8826_ = ~new_n3728_ | ~pi0300;
  assign new_n8827_ = ~new_n3727_ | ~pi0292;
  assign new_n8828_ = ~new_n3726_ | ~pi0284;
  assign new_n8829_ = ~new_n3725_ | ~pi0276;
  assign new_n8830_ = ~new_n3723_ | ~pi0268;
  assign new_n8831_ = ~new_n3722_ | ~pi0260;
  assign new_n8832_ = ~new_n3721_ | ~pi0252;
  assign new_n8833_ = ~new_n3720_ | ~pi0244;
  assign new_n8834_ = ~new_n3738_ | ~pi0237;
  assign new_n8835_ = ~new_n3737_ | ~pi0229;
  assign new_n8836_ = ~new_n3736_ | ~pi0221;
  assign new_n8837_ = ~new_n3735_ | ~pi0213;
  assign new_n8838_ = ~new_n3733_ | ~pi0205;
  assign new_n8839_ = ~new_n3732_ | ~pi0197;
  assign new_n8840_ = ~new_n3731_ | ~pi0189;
  assign new_n8841_ = ~new_n3730_ | ~pi0181;
  assign new_n8842_ = ~new_n3728_ | ~pi0301;
  assign new_n8843_ = ~new_n3727_ | ~pi0293;
  assign new_n8844_ = ~new_n3726_ | ~pi0285;
  assign new_n8845_ = ~new_n3725_ | ~pi0277;
  assign new_n8846_ = ~new_n3723_ | ~pi0269;
  assign new_n8847_ = ~new_n3722_ | ~pi0261;
  assign new_n8848_ = ~new_n3721_ | ~pi0253;
  assign new_n8849_ = ~new_n3720_ | ~pi0245;
  assign new_n8850_ = ~new_n3738_ | ~pi0238;
  assign new_n8851_ = ~new_n3737_ | ~pi0230;
  assign new_n8852_ = ~new_n3736_ | ~pi0222;
  assign new_n8853_ = ~new_n3735_ | ~pi0214;
  assign new_n8854_ = ~new_n3733_ | ~pi0206;
  assign new_n8855_ = ~new_n3732_ | ~pi0198;
  assign new_n8856_ = ~new_n3731_ | ~pi0190;
  assign new_n8857_ = ~new_n3730_ | ~pi0182;
  assign new_n8858_ = ~new_n3728_ | ~pi0302;
  assign new_n8859_ = ~new_n3727_ | ~pi0294;
  assign new_n8860_ = ~new_n3726_ | ~pi0286;
  assign new_n8861_ = ~new_n3725_ | ~pi0278;
  assign new_n8862_ = ~new_n3723_ | ~pi0270;
  assign new_n8863_ = ~new_n3722_ | ~pi0262;
  assign new_n8864_ = ~new_n3721_ | ~pi0254;
  assign new_n8865_ = ~new_n3720_ | ~pi0246;
  assign new_n8866_ = ~new_n3738_ | ~pi0239;
  assign new_n8867_ = ~new_n3737_ | ~pi0231;
  assign new_n8868_ = ~new_n3736_ | ~pi0223;
  assign new_n8869_ = ~new_n3735_ | ~pi0215;
  assign new_n8870_ = ~new_n3733_ | ~pi0207;
  assign new_n8871_ = ~new_n3732_ | ~pi0199;
  assign new_n8872_ = ~new_n3731_ | ~pi0191;
  assign new_n8873_ = ~new_n3730_ | ~pi0183;
  assign new_n8874_ = ~new_n3728_ | ~pi0303;
  assign new_n8875_ = ~new_n3727_ | ~pi0295;
  assign new_n8876_ = ~new_n3726_ | ~pi0287;
  assign new_n8877_ = ~new_n3725_ | ~pi0279;
  assign new_n8878_ = ~new_n3723_ | ~pi0271;
  assign new_n8879_ = ~new_n3722_ | ~pi0263;
  assign new_n8880_ = ~new_n3721_ | ~pi0255;
  assign new_n8881_ = ~new_n3720_ | ~pi0247;
  assign new_n8882_ = ~new_n3738_ | ~pi0240;
  assign new_n8883_ = ~new_n3737_ | ~pi0232;
  assign new_n8884_ = ~new_n3736_ | ~pi0224;
  assign new_n8885_ = ~new_n3735_ | ~pi0216;
  assign new_n8886_ = ~new_n3733_ | ~pi0208;
  assign new_n8887_ = ~new_n3732_ | ~pi0200;
  assign new_n8888_ = ~new_n3731_ | ~pi0192;
  assign new_n8889_ = ~new_n3730_ | ~pi0184;
  assign new_n8890_ = ~new_n3728_ | ~pi0304;
  assign new_n8891_ = ~new_n3727_ | ~pi0296;
  assign new_n8892_ = ~new_n3726_ | ~pi0288;
  assign new_n8893_ = ~new_n3725_ | ~pi0280;
  assign new_n8894_ = ~new_n3723_ | ~pi0272;
  assign new_n8895_ = ~new_n3722_ | ~pi0264;
  assign new_n8896_ = ~new_n3721_ | ~pi0256;
  assign new_n8897_ = ~new_n3720_ | ~pi0248;
  assign new_n8898_ = ~new_n3738_ | ~pi0241;
  assign new_n8899_ = ~new_n3737_ | ~pi0233;
  assign new_n8900_ = ~new_n3736_ | ~pi0225;
  assign new_n8901_ = ~new_n3735_ | ~pi0217;
  assign new_n8902_ = ~new_n3733_ | ~pi0209;
  assign new_n8903_ = ~new_n3732_ | ~pi0201;
  assign new_n8904_ = ~new_n3731_ | ~pi0193;
  assign new_n8905_ = ~new_n3730_ | ~pi0185;
  assign new_n8906_ = ~new_n3728_ | ~pi0305;
  assign new_n8907_ = ~new_n3727_ | ~pi0297;
  assign new_n8908_ = ~new_n3726_ | ~pi0289;
  assign new_n8909_ = ~new_n3725_ | ~pi0281;
  assign new_n8910_ = ~new_n3723_ | ~pi0273;
  assign new_n8911_ = ~new_n3722_ | ~pi0265;
  assign new_n8912_ = ~new_n3721_ | ~pi0257;
  assign new_n8913_ = ~new_n3720_ | ~pi0249;
  assign new_n8914_ = ~new_n3738_ | ~pi0242;
  assign new_n8915_ = ~new_n3737_ | ~pi0234;
  assign new_n8916_ = ~new_n3736_ | ~pi0226;
  assign new_n8917_ = ~new_n3735_ | ~pi0218;
  assign new_n8918_ = ~new_n3733_ | ~pi0210;
  assign new_n8919_ = ~new_n3732_ | ~pi0202;
  assign new_n8920_ = ~new_n3731_ | ~pi0194;
  assign new_n8921_ = ~new_n3730_ | ~pi0186;
  assign new_n8922_ = ~new_n3728_ | ~pi0306;
  assign new_n8923_ = ~new_n3727_ | ~pi0298;
  assign new_n8924_ = ~new_n3726_ | ~pi0290;
  assign new_n8925_ = ~new_n3725_ | ~pi0282;
  assign new_n8926_ = ~new_n3723_ | ~pi0274;
  assign new_n8927_ = ~new_n3722_ | ~pi0266;
  assign new_n8928_ = ~new_n3721_ | ~pi0258;
  assign new_n8929_ = ~new_n3720_ | ~pi0250;
  assign new_n8930_ = ~pi0308 | ~new_n4253_;
  assign new_n8931_ = ~new_n4424_;
  assign new_n8932_ = ~new_n3756_ | ~pi0235;
  assign new_n8933_ = ~new_n3755_ | ~pi0227;
  assign new_n8934_ = ~new_n3754_ | ~pi0219;
  assign new_n8935_ = ~new_n3753_ | ~pi0211;
  assign new_n8936_ = ~new_n3751_ | ~pi0203;
  assign new_n8937_ = ~new_n3750_ | ~pi0195;
  assign new_n8938_ = ~new_n3749_ | ~pi0187;
  assign new_n8939_ = ~new_n3748_ | ~pi0179;
  assign new_n8940_ = ~new_n3747_ | ~pi0299;
  assign new_n8941_ = ~new_n3746_ | ~pi0291;
  assign new_n8942_ = ~new_n3745_ | ~pi0283;
  assign new_n8943_ = ~new_n3744_ | ~pi0275;
  assign new_n8944_ = ~new_n3742_ | ~pi0267;
  assign new_n8945_ = ~new_n3741_ | ~pi0259;
  assign new_n8946_ = ~new_n3740_ | ~pi0251;
  assign new_n8947_ = ~new_n3739_ | ~pi0243;
  assign new_n8948_ = ~new_n3756_ | ~pi0236;
  assign new_n8949_ = ~new_n3755_ | ~pi0228;
  assign new_n8950_ = ~new_n3754_ | ~pi0220;
  assign new_n8951_ = ~new_n3753_ | ~pi0212;
  assign new_n8952_ = ~new_n3751_ | ~pi0204;
  assign new_n8953_ = ~new_n3750_ | ~pi0196;
  assign new_n8954_ = ~new_n3749_ | ~pi0188;
  assign new_n8955_ = ~new_n3748_ | ~pi0180;
  assign new_n8956_ = ~new_n3747_ | ~pi0300;
  assign new_n8957_ = ~new_n3746_ | ~pi0292;
  assign new_n8958_ = ~new_n3745_ | ~pi0284;
  assign new_n8959_ = ~new_n3744_ | ~pi0276;
  assign new_n8960_ = ~new_n3742_ | ~pi0268;
  assign new_n8961_ = ~new_n3741_ | ~pi0260;
  assign new_n8962_ = ~new_n3740_ | ~pi0252;
  assign new_n8963_ = ~new_n3739_ | ~pi0244;
  assign new_n8964_ = ~new_n3756_ | ~pi0237;
  assign new_n8965_ = ~new_n3755_ | ~pi0229;
  assign new_n8966_ = ~new_n3754_ | ~pi0221;
  assign new_n8967_ = ~new_n3753_ | ~pi0213;
  assign new_n8968_ = ~new_n3751_ | ~pi0205;
  assign new_n8969_ = ~new_n3750_ | ~pi0197;
  assign new_n8970_ = ~new_n3749_ | ~pi0189;
  assign new_n8971_ = ~new_n3748_ | ~pi0181;
  assign new_n8972_ = ~new_n3747_ | ~pi0301;
  assign new_n8973_ = ~new_n3746_ | ~pi0293;
  assign new_n8974_ = ~new_n3745_ | ~pi0285;
  assign new_n8975_ = ~new_n3744_ | ~pi0277;
  assign new_n8976_ = ~new_n3742_ | ~pi0269;
  assign new_n8977_ = ~new_n3741_ | ~pi0261;
  assign new_n8978_ = ~new_n3740_ | ~pi0253;
  assign new_n8979_ = ~new_n3739_ | ~pi0245;
  assign new_n8980_ = ~new_n3756_ | ~pi0238;
  assign new_n8981_ = ~new_n3755_ | ~pi0230;
  assign new_n8982_ = ~new_n3754_ | ~pi0222;
  assign new_n8983_ = ~new_n3753_ | ~pi0214;
  assign new_n8984_ = ~new_n3751_ | ~pi0206;
  assign new_n8985_ = ~new_n3750_ | ~pi0198;
  assign new_n8986_ = ~new_n3749_ | ~pi0190;
  assign new_n8987_ = ~new_n3748_ | ~pi0182;
  assign new_n8988_ = ~new_n3747_ | ~pi0302;
  assign new_n8989_ = ~new_n3746_ | ~pi0294;
  assign new_n8990_ = ~new_n3745_ | ~pi0286;
  assign new_n8991_ = ~new_n3744_ | ~pi0278;
  assign new_n8992_ = ~new_n3742_ | ~pi0270;
  assign new_n8993_ = ~new_n3741_ | ~pi0262;
  assign new_n8994_ = ~new_n3740_ | ~pi0254;
  assign new_n8995_ = ~new_n3739_ | ~pi0246;
  assign new_n8996_ = ~new_n3756_ | ~pi0239;
  assign new_n8997_ = ~new_n3755_ | ~pi0231;
  assign new_n8998_ = ~new_n3754_ | ~pi0223;
  assign new_n8999_ = ~new_n3753_ | ~pi0215;
  assign new_n9000_ = ~new_n3751_ | ~pi0207;
  assign new_n9001_ = ~new_n3750_ | ~pi0199;
  assign new_n9002_ = ~new_n3749_ | ~pi0191;
  assign new_n9003_ = ~new_n3748_ | ~pi0183;
  assign new_n9004_ = ~new_n3747_ | ~pi0303;
  assign new_n9005_ = ~new_n3746_ | ~pi0295;
  assign new_n9006_ = ~new_n3745_ | ~pi0287;
  assign new_n9007_ = ~new_n3744_ | ~pi0279;
  assign new_n9008_ = ~new_n3742_ | ~pi0271;
  assign new_n9009_ = ~new_n3741_ | ~pi0263;
  assign new_n9010_ = ~new_n3740_ | ~pi0255;
  assign new_n9011_ = ~new_n3739_ | ~pi0247;
  assign new_n9012_ = ~new_n3756_ | ~pi0240;
  assign new_n9013_ = ~new_n3755_ | ~pi0232;
  assign new_n9014_ = ~new_n3754_ | ~pi0224;
  assign new_n9015_ = ~new_n3753_ | ~pi0216;
  assign new_n9016_ = ~new_n3751_ | ~pi0208;
  assign new_n9017_ = ~new_n3750_ | ~pi0200;
  assign new_n9018_ = ~new_n3749_ | ~pi0192;
  assign new_n9019_ = ~new_n3748_ | ~pi0184;
  assign new_n9020_ = ~new_n3747_ | ~pi0304;
  assign new_n9021_ = ~new_n3746_ | ~pi0296;
  assign new_n9022_ = ~new_n3745_ | ~pi0288;
  assign new_n9023_ = ~new_n3744_ | ~pi0280;
  assign new_n9024_ = ~new_n3742_ | ~pi0272;
  assign new_n9025_ = ~new_n3741_ | ~pi0264;
  assign new_n9026_ = ~new_n3740_ | ~pi0256;
  assign new_n9027_ = ~new_n3739_ | ~pi0248;
  assign new_n9028_ = ~new_n3756_ | ~pi0241;
  assign new_n9029_ = ~new_n3755_ | ~pi0233;
  assign new_n9030_ = ~new_n3754_ | ~pi0225;
  assign new_n9031_ = ~new_n3753_ | ~pi0217;
  assign new_n9032_ = ~new_n3751_ | ~pi0209;
  assign new_n9033_ = ~new_n3750_ | ~pi0201;
  assign new_n9034_ = ~new_n3749_ | ~pi0193;
  assign new_n9035_ = ~new_n3748_ | ~pi0185;
  assign new_n9036_ = ~new_n3747_ | ~pi0305;
  assign new_n9037_ = ~new_n3746_ | ~pi0297;
  assign new_n9038_ = ~new_n3745_ | ~pi0289;
  assign new_n9039_ = ~new_n3744_ | ~pi0281;
  assign new_n9040_ = ~new_n3742_ | ~pi0273;
  assign new_n9041_ = ~new_n3741_ | ~pi0265;
  assign new_n9042_ = ~new_n3740_ | ~pi0257;
  assign new_n9043_ = ~new_n3739_ | ~pi0249;
  assign new_n9044_ = ~new_n3756_ | ~pi0242;
  assign new_n9045_ = ~new_n3755_ | ~pi0234;
  assign new_n9046_ = ~new_n3754_ | ~pi0226;
  assign new_n9047_ = ~new_n3753_ | ~pi0218;
  assign new_n9048_ = ~new_n3751_ | ~pi0210;
  assign new_n9049_ = ~new_n3750_ | ~pi0202;
  assign new_n9050_ = ~new_n3749_ | ~pi0194;
  assign new_n9051_ = ~new_n3748_ | ~pi0186;
  assign new_n9052_ = ~new_n3747_ | ~pi0306;
  assign new_n9053_ = ~new_n3746_ | ~pi0298;
  assign new_n9054_ = ~new_n3745_ | ~pi0290;
  assign new_n9055_ = ~new_n3744_ | ~pi0282;
  assign new_n9056_ = ~new_n3742_ | ~pi0274;
  assign new_n9057_ = ~new_n3741_ | ~pi0266;
  assign new_n9058_ = ~new_n3740_ | ~pi0258;
  assign new_n9059_ = ~new_n3739_ | ~pi0250;
  assign new_n9060_ = ~pi0142 | ~new_n5448_;
  assign new_n9061_ = new_n2971_ | pi0176;
  assign new_n9062_ = ~new_n5095_ | ~new_n7553_;
  assign new_n9063_ = ~new_n5290_ | ~new_n3759_;
  assign new_n9064_ = ~new_n3560_ | ~new_n4412_;
  assign new_n9065_ = ~new_n3548_ | ~new_n8252_;
  assign new_n9066_ = ~new_n9065_ | ~new_n9064_ | ~new_n5473_;
  assign new_n9067_ = ~new_n4242_;
  assign new_n9068_ = ~new_n9067_ | ~new_n4244_;
  assign new_n9069_ = ~new_n5602_ | ~new_n5605_ | ~pi0141;
  assign new_n9070_ = ~pi0140 | ~new_n9060_;
  assign new_n9071_ = ~pi0141 | ~new_n5602_;
  assign new_n9072_ = ~new_n5661_ | ~new_n4262_;
  assign new_n9073_ = ~new_n5644_ | ~new_n5678_;
  assign new_n9074_ = ~new_n4364_ | ~new_n4375_;
  assign new_n9075_ = ~new_n8532_ | ~new_n4261_;
  assign new_n9076_ = ~pi0106 | ~new_n4233_;
  assign new_n9077_ = ~pi0540 | ~new_n5464_;
  assign new_n9078_ = ~pi0107 | ~new_n4233_;
  assign new_n9079_ = ~pi0541 | ~new_n5464_;
  assign new_n9080_ = ~pi0108 | ~new_n4233_;
  assign new_n9081_ = ~pi0542 | ~new_n5464_;
  assign new_n9082_ = ~pi0109 | ~new_n4233_;
  assign new_n9083_ = ~pi0543 | ~new_n5464_;
  assign new_n9084_ = ~new_n4235_ | ~pi0142 | ~pi0548;
  assign new_n9085_ = ~pi0140 | ~new_n4242_;
  assign new_n9086_ = ~new_n9085_ | ~new_n9084_;
  assign new_n9087_ = ~pi0141 | ~new_n9070_ | ~new_n5605_;
  assign new_n9088_ = ~new_n9086_ | ~new_n4232_;
  assign new_n9089_ = ~pi0140 | ~pi0142 | ~new_n4243_;
  assign new_n9090_ = ~new_n5615_ | ~new_n4235_;
  assign new_n9091_ = pi0142 | pi0141;
  assign new_n9092_ = ~pi0142 | ~new_n5502_;
  assign new_n9093_ = ~new_n4434_;
  assign new_n9094_ = ~new_n9093_ | ~pi0143;
  assign new_n9095_ = ~new_n4435_ | ~new_n4434_;
  assign new_n9096_ = ~new_n4434_ | ~new_n5620_;
  assign new_n9097_ = ~new_n9093_ | ~pi0144;
  assign new_n9098_ = ~new_n5661_ | ~new_n4367_;
  assign new_n9099_ = ~new_n4260_ | ~new_n4370_;
  assign new_n9100_ = ~new_n5661_ | ~new_n4369_;
  assign new_n9101_ = ~new_n4260_ | ~new_n4366_;
  assign new_n9102_ = ~new_n5695_ | ~new_n5774_;
  assign new_n9103_ = ~new_n5776_ | ~new_n4257_;
  assign new_n9104_ = ~new_n5437_ | ~new_n5773_;
  assign new_n9105_ = ~new_n5778_ | ~new_n5780_;
  assign new_n9106_ = ~new_n5661_ | ~new_n4393_;
  assign new_n9107_ = ~new_n4260_ | ~new_n4394_;
  assign new_n9108_ = ~pi0178 | ~new_n5783_;
  assign new_n9109_ = ~new_n5784_ | ~new_n4277_;
  assign new_n9110_ = ~pi0175 | ~new_n4278_;
  assign new_n9111_ = ~new_n3609_ | ~new_n5786_;
  assign new_n9112_ = pi0547 | pi0178;
  assign new_n9113_ = ~pi0178 | ~new_n9061_;
  assign new_n9114_ = ~pi0178 | ~new_n5794_;
  assign new_n9115_ = ~new_n4277_ | ~new_n5793_ | ~new_n5785_;
  assign new_n9116_ = ~pi0314 | ~new_n4286_;
  assign new_n9117_ = ~new_n5804_ | ~new_n4287_;
  assign new_n9118_ = ~new_n4425_;
  assign new_n9119_ = ~new_n9118_ | ~new_n5809_;
  assign new_n9120_ = ~new_n4425_ | ~new_n4294_;
  assign new_n9121_ = ~new_n4426_;
  assign new_n9122_ = ~new_n9121_ | ~new_n5813_;
  assign new_n9123_ = ~new_n4426_ | ~new_n4296_;
  assign new_n9124_ = ~new_n4427_;
  assign new_n9125_ = ~new_n4265_ | ~new_n4257_;
  assign new_n9126_ = ~new_n5695_ | ~new_n6639_;
  assign new_n9127_ = ~new_n4439_ | ~new_n5439_;
  assign new_n9128_ = ~new_n6655_ | ~pi0307;
  assign new_n9129_ = ~new_n4374_ | ~new_n4263_;
  assign new_n9130_ = ~new_n5729_ | ~new_n5746_;
  assign new_n9131_ = ~new_n5695_ | ~new_n6668_;
  assign new_n9132_ = ~new_n6671_ | ~new_n4257_;
  assign new_n9133_ = ~new_n4266_ | ~new_n5712_ | ~new_n6673_;
  assign new_n9134_ = ~new_n5746_ | ~new_n6669_ | ~new_n4263_;
  assign new_n9135_ = ~new_n6655_ | ~pi0308;
  assign new_n9136_ = ~new_n6702_ | ~new_n5439_;
  assign new_n9137_ = ~new_n4250_ | ~pi0309 | ~new_n4377_;
  assign new_n9138_ = ~pi0310 | ~new_n6687_ | ~new_n4253_;
  assign new_n9139_ = ~pi0318 | ~new_n5440_;
  assign new_n9140_ = ~new_n23872_ | ~pi0348;
  assign new_n9141_ = ~new_n4443_;
  assign new_n9142_ = ~pi0317 | ~new_n5440_;
  assign new_n9143_ = ~pi0317 | ~pi0348;
  assign new_n9144_ = ~new_n4442_;
  assign new_n9145_ = ~new_n6655_ | ~pi0309;
  assign new_n9146_ = ~new_n6713_ | ~new_n5439_;
  assign new_n9147_ = ~new_n6655_ | ~pi0310;
  assign new_n9148_ = ~new_n6726_ | ~new_n5439_;
  assign new_n9149_ = ~pi0311 | ~new_n4377_;
  assign new_n9150_ = ~new_n6727_ | ~new_n4249_;
  assign new_n9151_ = ~new_n6655_ | ~pi0311;
  assign new_n9152_ = ~new_n6733_ | ~new_n5439_;
  assign new_n9153_ = ~new_n9124_ | ~new_n5803_;
  assign new_n9154_ = ~new_n4427_ | ~new_n4299_;
  assign new_n9155_ = ~new_n9154_ | ~new_n9153_;
  assign new_n9156_ = ~new_n6778_ | ~new_n4260_;
  assign new_n9157_ = ~new_n5661_ | ~new_n6775_;
  assign new_n9158_ = ~pi0540 | ~new_n4417_;
  assign new_n9159_ = ~new_n4447_ | ~new_n5463_;
  assign new_n9160_ = pi0143 | pi0144;
  assign new_n9161_ = ~pi0143 | ~new_n4396_;
  assign new_n9162_ = ~new_n9161_ | ~new_n9160_;
  assign new_n9163_ = ~new_n9162_ | ~new_n4237_;
  assign new_n9164_ = ~pi0508 | ~pi0509;
  assign new_n9165_ = ~new_n9164_ | ~new_n9163_;
  assign new_n9166_ = ~pi0541 | ~new_n4417_;
  assign new_n9167_ = ~new_n9165_ | ~new_n5463_;
  assign new_n9168_ = ~pi0542 | ~new_n4417_;
  assign new_n9169_ = ~new_n5463_ | ~pi0509;
  assign new_n9170_ = ~pi0543 | ~new_n4417_;
  assign new_n9171_ = ~new_n5463_ | ~new_n8523_;
  assign new_n9172_ = ~new_n5464_ | ~new_n4420_;
  assign new_n9173_ = ~pi0544 | ~new_n4233_;
  assign new_n9174_ = ~new_n8524_ | ~new_n5773_;
  assign new_n9175_ = ~pi0546 | ~new_n5441_;
  assign new_n9176_ = ~new_n9093_ | ~pi0547;
  assign new_n9177_ = ~pi0035 | ~new_n4434_;
  assign new_n9178_ = ~new_n8530_ | ~pi0548;
  assign new_n9179_ = ~new_n8535_ | ~new_n5443_;
  assign new_n9180_ = ~new_n5464_ | ~new_n4419_;
  assign new_n9181_ = ~pi0549 | ~new_n4233_;
  assign new_n9182_ = ~pi0550 | ~new_n4233_;
  assign new_n9183_ = ~pi0554 | ~new_n5464_;
  assign new_n9184_ = ~new_n8540_ | ~pi0553;
  assign new_n9185_ = ~new_n8541_ | ~new_n5444_;
  assign new_n9186_ = ~new_n8540_ | ~pi0554;
  assign new_n9187_ = ~new_n8542_ | ~new_n5444_;
  assign new_n9188_ = ~pi0310 | ~new_n4253_;
  assign new_n9189_ = ~pi0309 | ~new_n4250_;
  assign new_n9190_ = ~new_n4428_;
  assign new_n9191_ = ~pi0308 | ~new_n5445_;
  assign new_n9192_ = ~new_n8801_ | ~new_n4256_;
  assign new_n9193_ = ~new_n4429_;
  assign new_n9194_ = ~pi0309 | ~new_n4363_;
  assign new_n9195_ = ~pi0545 | ~new_n4443_ | ~new_n4442_;
  assign new_n9196_ = ~pi0310 | ~new_n4363_;
  assign new_n9197_ = ~pi0545 | ~new_n4442_ | ~new_n9141_;
  assign new_n9198_ = ~pi0311 | ~new_n4363_;
  assign new_n9199_ = ~new_n9144_ | ~pi0545;
  assign new_n9200_ = ~new_n4459_ | ~new_n5446_;
  assign new_n9201_ = ~new_n6652_ | ~pi0307;
  assign new_n9202_ = ~new_n6652_ | ~pi0308;
  assign new_n9203_ = ~new_n6698_ | ~new_n5446_;
  assign new_n9204_ = ~new_n6652_ | ~pi0309;
  assign new_n9205_ = ~new_n6709_ | ~new_n5446_;
  assign new_n9206_ = ~new_n6652_ | ~pi0310;
  assign new_n9207_ = ~new_n6722_ | ~new_n5446_;
  assign new_n9208_ = ~new_n6652_ | ~pi0311;
  assign new_n9209_ = ~new_n6729_ | ~new_n5446_;
  assign new_n9210_ = ~new_n9286_ | ~new_n9373_;
  assign new_n9211_ = ~pi1218 | ~new_n9374_;
  assign new_n9212_ = ~new_n9258_ | ~new_n9288_;
  assign new_n9213_ = ~pi1246 | ~new_n9287_;
  assign new_n9214_ = ~new_n9279_ | ~new_n9359_;
  assign new_n9215_ = ~pi1225 | ~new_n9360_;
  assign new_n9216_ = ~new_n9270_ | ~new_n9341_;
  assign new_n9217_ = ~pi1234 | ~new_n9342_;
  assign new_n9218_ = ~new_n9266_ | ~new_n9333_;
  assign new_n9219_ = ~pi1238 | ~new_n9334_;
  assign new_n9220_ = ~new_n9281_ | ~new_n9363_;
  assign new_n9221_ = ~pi1223 | ~new_n9364_;
  assign new_n9222_ = ~new_n9284_ | ~new_n9369_;
  assign new_n9223_ = ~pi1220 | ~new_n9370_;
  assign new_n9224_ = ~new_n9275_ | ~new_n9351_;
  assign new_n9225_ = ~pi1229 | ~new_n9352_;
  assign new_n9226_ = ~new_n9262_ | ~new_n9325_;
  assign new_n9227_ = ~pi1242 | ~new_n9326_;
  assign new_n9228_ = ~new_n9285_ | ~new_n9371_;
  assign new_n9229_ = ~pi1219 | ~new_n9372_;
  assign new_n9230_ = ~new_n9274_ | ~new_n9349_;
  assign new_n9231_ = ~pi1230 | ~new_n9350_;
  assign new_n9232_ = ~new_n9263_ | ~new_n9327_;
  assign new_n9233_ = ~pi1241 | ~new_n9328_;
  assign new_n9234_ = ~new_n9278_ | ~new_n9357_;
  assign new_n9235_ = ~pi1226 | ~new_n9358_;
  assign new_n9236_ = ~new_n9271_ | ~new_n9343_;
  assign new_n9237_ = ~pi1233 | ~new_n9344_;
  assign new_n9238_ = ~new_n9267_ | ~new_n9335_;
  assign new_n9239_ = ~pi1237 | ~new_n9336_;
  assign new_n9240_ = ~new_n9280_ | ~new_n9361_;
  assign new_n9241_ = ~pi1224 | ~new_n9362_;
  assign new_n9242_ = ~new_n9276_ | ~new_n9353_;
  assign new_n9243_ = ~pi1228 | ~new_n9354_;
  assign new_n9244_ = ~new_n9269_ | ~new_n9339_;
  assign new_n9245_ = ~pi1235 | ~new_n9340_;
  assign new_n9246_ = ~pi1216 | ~new_n9375_;
  assign new_n9247_ = ~pi1217 | ~new_n9376_;
  assign new_n9248_ = ~new_n9272_ | ~new_n9345_;
  assign new_n9249_ = ~pi1232 | ~new_n9346_;
  assign new_n9250_ = ~new_n9265_ | ~new_n9331_;
  assign new_n9251_ = ~pi1239 | ~new_n9332_;
  assign new_n9252_ = ~new_n9260_ | ~new_n9321_;
  assign new_n9253_ = ~pi1244 | ~new_n9322_;
  assign new_n9254_ = ~new_n9259_ | ~new_n9320_;
  assign new_n9255_ = ~pi1245 | ~new_n9319_;
  assign new_n9256_ = ~new_n9283_ | ~new_n9368_;
  assign new_n9257_ = ~pi1221 | ~new_n9367_;
  assign new_n9258_ = ~new_n9287_;
  assign new_n9259_ = ~new_n9319_;
  assign new_n9260_ = ~new_n9322_;
  assign new_n9261_ = ~new_n9324_;
  assign new_n9262_ = ~new_n9326_;
  assign new_n9263_ = ~new_n9328_;
  assign new_n9264_ = ~new_n9330_;
  assign new_n9265_ = ~new_n9332_;
  assign new_n9266_ = ~new_n9334_;
  assign new_n9267_ = ~new_n9336_;
  assign new_n9268_ = ~new_n9338_;
  assign new_n9269_ = ~new_n9340_;
  assign new_n9270_ = ~new_n9342_;
  assign new_n9271_ = ~new_n9344_;
  assign new_n9272_ = ~new_n9346_;
  assign new_n9273_ = ~new_n9348_;
  assign new_n9274_ = ~new_n9350_;
  assign new_n9275_ = ~new_n9352_;
  assign new_n9276_ = ~new_n9354_;
  assign new_n9277_ = ~new_n9356_;
  assign new_n9278_ = ~new_n9358_;
  assign new_n9279_ = ~new_n9360_;
  assign new_n9280_ = ~new_n9362_;
  assign new_n9281_ = ~new_n9364_;
  assign new_n9282_ = ~new_n9366_;
  assign new_n9283_ = ~new_n9367_;
  assign new_n9284_ = ~new_n9370_;
  assign new_n9285_ = ~new_n9372_;
  assign new_n9286_ = ~new_n9374_;
  assign new_n9287_ = ~new_n9259_ | ~pi1245;
  assign new_n9288_ = ~pi1246;
  assign new_n9289_ = ~new_n2966_ | ~new_n2967_;
  assign new_n9290_ = ~new_n2968_ | ~new_n3499_;
  assign new_n9291_ = ~new_n3500_ | ~new_n3501_;
  assign new_n9292_ = ~new_n3502_ | ~new_n3503_;
  assign new_n9293_ = ~new_n3504_ | ~new_n3505_;
  assign new_n9294_ = ~new_n3506_ | ~new_n3507_;
  assign new_n9295_ = ~new_n9210_ | ~new_n9211_;
  assign new_n9296_ = ~new_n9212_ | ~new_n9213_;
  assign new_n9297_ = ~new_n9214_ | ~new_n9215_;
  assign new_n9298_ = ~new_n9216_ | ~new_n9217_;
  assign new_n9299_ = ~new_n9218_ | ~new_n9219_;
  assign new_n9300_ = ~new_n9220_ | ~new_n9221_;
  assign new_n9301_ = ~new_n9222_ | ~new_n9223_;
  assign new_n9302_ = ~new_n9224_ | ~new_n9225_;
  assign new_n9303_ = ~new_n9226_ | ~new_n9227_;
  assign new_n9304_ = ~new_n9228_ | ~new_n9229_;
  assign new_n9305_ = ~new_n9230_ | ~new_n9231_;
  assign new_n9306_ = ~new_n9232_ | ~new_n9233_;
  assign new_n9307_ = ~new_n9234_ | ~new_n9235_;
  assign new_n9308_ = ~new_n9236_ | ~new_n9237_;
  assign new_n9309_ = ~new_n9238_ | ~new_n9239_;
  assign new_n9310_ = ~new_n9240_ | ~new_n9241_;
  assign new_n9311_ = ~new_n9242_ | ~new_n9243_;
  assign new_n9312_ = ~new_n9244_ | ~new_n9245_;
  assign new_n9313_ = ~new_n9246_ | ~new_n9247_;
  assign new_n9314_ = ~new_n9248_ | ~new_n9249_;
  assign new_n9315_ = ~new_n9250_ | ~new_n9251_;
  assign new_n9316_ = ~new_n9252_ | ~new_n9253_;
  assign new_n9317_ = ~new_n9254_ | ~new_n9255_;
  assign new_n9318_ = ~new_n9256_ | ~new_n9257_;
  assign new_n9319_ = ~pi1244 | ~new_n9260_;
  assign new_n9320_ = ~pi1245;
  assign new_n9321_ = ~pi1244;
  assign new_n9322_ = ~pi1243 | ~new_n9261_;
  assign new_n9323_ = ~pi1243;
  assign new_n9324_ = ~pi1242 | ~new_n9262_;
  assign new_n9325_ = ~pi1242;
  assign new_n9326_ = ~pi1241 | ~new_n9263_;
  assign new_n9327_ = ~pi1241;
  assign new_n9328_ = ~pi1240 | ~new_n9264_;
  assign new_n9329_ = ~pi1240;
  assign new_n9330_ = ~pi1239 | ~new_n9265_;
  assign new_n9331_ = ~pi1239;
  assign new_n9332_ = ~pi1238 | ~new_n9266_;
  assign new_n9333_ = ~pi1238;
  assign new_n9334_ = ~pi1237 | ~new_n9267_;
  assign new_n9335_ = ~pi1237;
  assign new_n9336_ = ~pi1236 | ~new_n9268_;
  assign new_n9337_ = ~pi1236;
  assign new_n9338_ = ~pi1235 | ~new_n9269_;
  assign new_n9339_ = ~pi1235;
  assign new_n9340_ = ~pi1234 | ~new_n9270_;
  assign new_n9341_ = ~pi1234;
  assign new_n9342_ = ~pi1233 | ~new_n9271_;
  assign new_n9343_ = ~pi1233;
  assign new_n9344_ = ~pi1232 | ~new_n9272_;
  assign new_n9345_ = ~pi1232;
  assign new_n9346_ = ~pi1231 | ~new_n9273_;
  assign new_n9347_ = ~pi1231;
  assign new_n9348_ = ~pi1230 | ~new_n9274_;
  assign new_n9349_ = ~pi1230;
  assign new_n9350_ = ~pi1229 | ~new_n9275_;
  assign new_n9351_ = ~pi1229;
  assign new_n9352_ = ~pi1228 | ~new_n9276_;
  assign new_n9353_ = ~pi1228;
  assign new_n9354_ = ~pi1227 | ~new_n9277_;
  assign new_n9355_ = ~pi1227;
  assign new_n9356_ = ~pi1226 | ~new_n9278_;
  assign new_n9357_ = ~pi1226;
  assign new_n9358_ = ~pi1225 | ~new_n9279_;
  assign new_n9359_ = ~pi1225;
  assign new_n9360_ = ~pi1224 | ~new_n9280_;
  assign new_n9361_ = ~pi1224;
  assign new_n9362_ = ~pi1223 | ~new_n9281_;
  assign new_n9363_ = ~pi1223;
  assign new_n9364_ = ~pi1222 | ~new_n9282_;
  assign new_n9365_ = ~pi1222;
  assign new_n9366_ = ~new_n9283_ | ~pi1221;
  assign new_n9367_ = ~pi1220 | ~new_n9284_;
  assign new_n9368_ = ~pi1221;
  assign new_n9369_ = ~pi1220;
  assign new_n9370_ = ~pi1219 | ~new_n9285_;
  assign new_n9371_ = ~pi1219;
  assign new_n9372_ = ~pi1218 | ~new_n9286_;
  assign new_n9373_ = ~pi1218;
  assign new_n9374_ = ~pi1217 | ~pi1216;
  assign new_n9375_ = ~pi1217;
  assign new_n9376_ = ~pi1216;
  assign new_n9377_ = ~new_n33511_ & ~new_n33510_ & ~new_n33512_ & ~new_n33513_;
  assign new_n9378_ = ~new_n33497_ & ~new_n9377_;
  assign new_n9379_ = ~new_n20979_ | ~new_n33689_;
  assign new_n9380_ = ~pi1231 | ~new_n33688_;
  assign new_n9381_ = ~new_n15528_ | ~new_n33707_;
  assign new_n9382_ = ~pi1240 | ~new_n33706_;
  assign new_n9383_ = ~new_n20988_ | ~new_n33671_;
  assign new_n9384_ = ~pi1222 | ~new_n33670_;
  assign new_n9385_ = ~new_n20983_ | ~new_n33681_;
  assign new_n9386_ = ~pi1227 | ~new_n33680_;
  assign new_n9387_ = ~new_n15532_ | ~new_n33699_;
  assign new_n9388_ = ~pi1236 | ~new_n33698_;
  assign new_n9389_ = ~new_n15525_ | ~new_n33713_;
  assign new_n9390_ = ~pi1243 | ~new_n33712_;
  assign new_n9391_ = ~pi1215 | ~new_n33662_;
  assign new_n9392_ = ~pi1216 | ~new_n33660_;
  assign new_n9393_ = new_n14914_ & new_n9658_ & new_n10341_;
  assign new_n9394_ = new_n11384_ & new_n9480_;
  assign new_n9395_ = pi0627 & new_n14902_ & new_n14914_;
  assign new_n9396_ = new_n9488_ & new_n14902_;
  assign new_n9397_ = pi0627 & new_n10294_;
  assign new_n9398_ = new_n10753_ & new_n9499_;
  assign new_n9399_ = new_n11472_ & pi0627;
  assign new_n9400_ = new_n11452_ & new_n10306_;
  assign new_n9401_ = ~new_n2973_ & ~pi0996;
  assign new_n9402_ = new_n29495_ & new_n9397_;
  assign new_n9403_ = new_n9439_ & new_n11484_;
  assign new_n9404_ = pi0625 & new_n10576_;
  assign new_n9405_ = pi0625 & new_n10587_;
  assign new_n9406_ = new_n11484_ & pi0624;
  assign new_n9407_ = pi0626 & new_n10587_;
  assign new_n9408_ = new_n9405_ & new_n11458_;
  assign new_n9409_ = new_n9404_ & new_n11461_;
  assign new_n9410_ = new_n9405_ & new_n11469_;
  assign new_n9411_ = new_n9488_ & new_n10578_;
  assign new_n9412_ = new_n11031_ & new_n10578_;
  assign new_n9413_ = new_n11030_ & new_n10578_;
  assign new_n9414_ = new_n11460_ & new_n10578_;
  assign new_n9415_ = new_n11509_ & pi0627;
  assign new_n9416_ = new_n11482_ & new_n10562_;
  assign new_n9417_ = new_n10914_ & new_n9477_;
  assign new_n9418_ = new_n9408_ & new_n11452_;
  assign new_n9419_ = pi0624 & new_n10587_;
  assign new_n9420_ = new_n11481_ & new_n14906_;
  assign new_n9421_ = new_n11482_ & new_n14906_;
  assign new_n9422_ = new_n10576_ & new_n10311_;
  assign new_n9423_ = new_n9407_ & new_n10688_;
  assign new_n9424_ = new_n9407_ & new_n10569_;
  assign new_n9425_ = new_n9409_ & new_n11458_;
  assign new_n9426_ = new_n9409_ & new_n11469_;
  assign new_n9427_ = new_n9404_ & new_n11477_;
  assign new_n9428_ = new_n12981_ & new_n10578_;
  assign new_n9429_ = new_n9404_ & new_n12716_;
  assign new_n9430_ = new_n9404_ & new_n12718_;
  assign new_n9431_ = new_n9404_ & new_n12720_;
  assign new_n9432_ = new_n9410_ & new_n10586_;
  assign new_n9433_ = new_n13612_ & new_n9410_;
  assign new_n9434_ = new_n11481_ & new_n10562_;
  assign new_n9435_ = new_n11483_ & new_n9657_;
  assign new_n9436_ = new_n11483_ & new_n14914_;
  assign new_n9437_ = new_n10582_ & new_n10325_;
  assign new_n9438_ = new_n11482_ & new_n11642_;
  assign new_n9439_ = new_n11471_ & pi0996;
  assign new_n9440_ = new_n3076_ & new_n11484_;
  assign new_n9441_ = new_n3065_ & new_n11484_;
  assign new_n9442_ = new_n3054_ & new_n11484_;
  assign new_n9443_ = new_n3051_ & new_n11484_;
  assign new_n9444_ = new_n3050_ & new_n11484_;
  assign new_n9445_ = new_n3049_ & new_n11484_;
  assign new_n9446_ = new_n3048_ & new_n11484_;
  assign new_n9447_ = new_n3047_ & new_n11484_;
  assign new_n9448_ = new_n3060_ & new_n9403_;
  assign new_n9449_ = new_n3069_ & new_n9403_;
  assign new_n9450_ = new_n3059_ & new_n9403_;
  assign new_n9451_ = new_n3068_ & new_n9403_;
  assign new_n9452_ = new_n3058_ & new_n9403_;
  assign new_n9453_ = new_n3067_ & new_n9403_;
  assign new_n9454_ = new_n3057_ & new_n9403_;
  assign new_n9455_ = new_n3066_ & new_n9403_;
  assign new_n9456_ = new_n3056_ & new_n9403_;
  assign new_n9457_ = new_n3064_ & new_n9403_;
  assign new_n9458_ = new_n3055_ & new_n9403_;
  assign new_n9459_ = new_n3063_ & new_n9403_;
  assign new_n9460_ = new_n3053_ & new_n9403_;
  assign new_n9461_ = new_n3062_ & new_n9403_;
  assign new_n9462_ = new_n3052_ & new_n9403_;
  assign new_n9463_ = new_n3061_ & new_n9403_;
  assign new_n9464_ = new_n9406_ & new_n10296_;
  assign new_n9465_ = new_n9406_ & new_n10319_;
  assign new_n9466_ = new_n9406_ & new_n10562_;
  assign new_n9467_ = new_n9406_ & new_n10320_;
  assign new_n9468_ = new_n9416_ & new_n10320_;
  assign new_n9469_ = new_n9406_ & new_n9657_;
  assign new_n9470_ = new_n9406_ & new_n9658_;
  assign new_n9471_ = pi0627 & new_n10582_;
  assign new_n9472_ = new_n9406_ & new_n10294_;
  assign new_n9473_ = new_n9406_ & new_n10321_;
  assign new_n9474_ = new_n9416_ & new_n10336_;
  assign new_n9475_ = new_n9416_ & new_n14910_;
  assign new_n9476_ = new_n9397_ & new_n10582_;
  assign new_n9477_ = new_n14900_ & new_n14908_;
  assign new_n9478_ = new_n9405_ & new_n14912_;
  assign new_n9479_ = new_n14900_ & new_n10319_;
  assign new_n9480_ = new_n11380_ & new_n10562_;
  assign new_n9481_ = new_n10621_ & new_n10469_;
  assign new_n9482_ = new_n11688_ & new_n10621_;
  assign new_n9483_ = new_n15108_ & new_n10469_;
  assign new_n9484_ = new_n11688_ & new_n15108_;
  assign new_n9485_ = new_n10284_ & new_n10348_;
  assign new_n9486_ = new_n11691_ & new_n10348_;
  assign new_n9487_ = new_n30327_ & new_n11465_;
  assign new_n9488_ = pi0627 & new_n9657_;
  assign new_n9489_ = pi0625 & pi0626;
  assign new_n9490_ = new_n10319_ & new_n10562_;
  assign new_n9491_ = new_n9395_ & new_n14912_;
  assign new_n9492_ = new_n9479_ & new_n11642_ & new_n9498_;
  assign new_n9493_ = pi0758 & pi0759 & new_n10313_;
  assign new_n9494_ = pi0758 & pi0760 & new_n10312_;
  assign new_n9495_ = pi0758 & new_n10312_ & new_n10313_;
  assign new_n9496_ = pi0759 & new_n10317_ & new_n10313_;
  assign new_n9497_ = pi0760 & new_n10317_ & new_n10312_;
  assign new_n9498_ = new_n10562_ & new_n10296_;
  assign new_n9499_ = new_n14904_ & new_n9658_ & new_n10320_;
  assign new_n9500_ = new_n11434_ & new_n15094_ & new_n15093_;
  assign new_n9501_ = new_n28333_ & new_n10358_;
  assign new_n9502_ = new_n10620_ & new_n10467_;
  assign new_n9503_ = new_n28369_ & new_n28333_;
  assign new_n9504_ = new_n11678_ & new_n9503_;
  assign new_n9505_ = pi0763 & pi0762;
  assign new_n9506_ = pi0763 & new_n10350_;
  assign new_n9507_ = new_n27644_ & new_n27643_;
  assign new_n9508_ = new_n27553_ & new_n27642_;
  assign new_n9509_ = new_n10361_ & new_n11698_;
  assign new_n9510_ = new_n11674_ & new_n9503_;
  assign new_n9511_ = new_n27553_ & new_n10364_;
  assign new_n9512_ = new_n10380_ & new_n11756_;
  assign new_n9513_ = new_n11675_ & new_n9503_;
  assign new_n9514_ = new_n27642_ & new_n10365_;
  assign new_n9515_ = new_n10395_ & new_n11815_;
  assign new_n9516_ = new_n11676_ & new_n28362_;
  assign new_n9517_ = ~new_n28362_ & ~new_n28361_;
  assign new_n9518_ = new_n9517_ & new_n9503_;
  assign new_n9519_ = ~pi0765 & ~pi0764;
  assign new_n9520_ = ~new_n27642_ & ~new_n27553_;
  assign new_n9521_ = new_n10407_ & new_n11872_;
  assign new_n9522_ = new_n15105_ & new_n10467_;
  assign new_n9523_ = new_n11679_ & new_n11678_;
  assign new_n9524_ = new_n27643_ & new_n10363_;
  assign new_n9525_ = new_n10420_ & new_n11930_;
  assign new_n9526_ = new_n11679_ & new_n11674_;
  assign new_n9527_ = new_n10432_ & new_n11987_;
  assign new_n9528_ = new_n11679_ & new_n11675_;
  assign new_n9529_ = new_n10443_ & new_n12045_;
  assign new_n9530_ = new_n11679_ & new_n9517_;
  assign new_n9531_ = new_n10455_ & new_n12102_;
  assign new_n9532_ = new_n11681_ & new_n10620_;
  assign new_n9533_ = new_n27644_ & new_n10362_;
  assign new_n9534_ = new_n10468_ & new_n10466_;
  assign new_n9535_ = new_n11674_ & new_n9501_;
  assign new_n9536_ = new_n10481_ & new_n12215_;
  assign new_n9537_ = new_n11675_ & new_n9501_;
  assign new_n9538_ = new_n10492_ & new_n12273_;
  assign new_n9539_ = new_n9517_ & new_n9501_;
  assign new_n9540_ = new_n10504_ & new_n12330_;
  assign new_n9541_ = new_n11681_ & new_n15105_;
  assign new_n9542_ = ~new_n28333_ & ~new_n28369_;
  assign new_n9543_ = new_n9542_ & new_n11678_;
  assign new_n9544_ = ~pi0762 & ~pi0763;
  assign new_n9545_ = ~new_n27643_ & ~new_n27644_;
  assign new_n9546_ = new_n10515_ & new_n12388_;
  assign new_n9547_ = new_n9542_ & new_n11674_;
  assign new_n9548_ = new_n10527_ & new_n12445_;
  assign new_n9549_ = new_n9542_ & new_n11675_;
  assign new_n9550_ = new_n10538_ & new_n12503_;
  assign new_n9551_ = new_n9542_ & new_n9517_;
  assign new_n9552_ = new_n10550_ & new_n12560_;
  assign new_n9553_ = new_n10910_ & new_n15110_ & new_n15109_;
  assign new_n9554_ = new_n12621_ & new_n12620_;
  assign new_n9555_ = new_n10923_ & new_n10922_ & new_n14937_;
  assign new_n9556_ = new_n15123_ & new_n15141_;
  assign new_n9557_ = new_n12657_ & pi0760;
  assign new_n9558_ = new_n9556_ & new_n9557_;
  assign new_n9559_ = new_n12657_ & new_n10313_;
  assign new_n9560_ = new_n9556_ & new_n9559_;
  assign new_n9561_ = new_n15123_ & new_n10623_;
  assign new_n9562_ = new_n9561_ & new_n9557_;
  assign new_n9563_ = new_n9561_ & new_n9559_;
  assign new_n9564_ = pi0760 & new_n10571_;
  assign new_n9565_ = new_n9556_ & new_n9564_;
  assign new_n9566_ = new_n10313_ & new_n10571_;
  assign new_n9567_ = new_n9556_ & new_n9566_;
  assign new_n9568_ = new_n9561_ & new_n9564_;
  assign new_n9569_ = new_n9561_ & new_n9566_;
  assign new_n9570_ = new_n10623_ & new_n10622_;
  assign new_n9571_ = new_n9566_ & new_n9570_;
  assign new_n9572_ = new_n9564_ & new_n9570_;
  assign new_n9573_ = new_n15141_ & new_n10622_;
  assign new_n9574_ = new_n9566_ & new_n9573_;
  assign new_n9575_ = new_n9564_ & new_n9573_;
  assign new_n9576_ = new_n9570_ & new_n9559_;
  assign new_n9577_ = new_n9570_ & new_n9557_;
  assign new_n9578_ = new_n9559_ & new_n9573_;
  assign new_n9579_ = new_n9557_ & new_n9573_;
  assign new_n9580_ = ~new_n29006_ & ~new_n29002_;
  assign new_n9581_ = ~pi0760 & ~new_n29007_;
  assign new_n9582_ = new_n9580_ & new_n9581_;
  assign new_n9583_ = pi0760 & new_n10570_;
  assign new_n9584_ = new_n9580_ & new_n9583_;
  assign new_n9585_ = new_n29002_ & new_n10567_;
  assign new_n9586_ = new_n9585_ & new_n9581_;
  assign new_n9587_ = new_n9585_ & new_n9583_;
  assign new_n9588_ = new_n29007_ & new_n10573_;
  assign new_n9589_ = new_n9580_ & new_n9588_;
  assign new_n9590_ = pi0760 & new_n29007_;
  assign new_n9591_ = new_n9580_ & new_n9590_;
  assign new_n9592_ = new_n9585_ & new_n9588_;
  assign new_n9593_ = new_n9585_ & new_n9590_;
  assign new_n9594_ = new_n29006_ & new_n10572_;
  assign new_n9595_ = new_n9581_ & new_n9594_;
  assign new_n9596_ = new_n9583_ & new_n9594_;
  assign new_n9597_ = new_n29002_ & new_n29006_;
  assign new_n9598_ = new_n9581_ & new_n9597_;
  assign new_n9599_ = new_n9583_ & new_n9597_;
  assign new_n9600_ = new_n9594_ & new_n9588_;
  assign new_n9601_ = new_n9594_ & new_n9590_;
  assign new_n9602_ = new_n9588_ & new_n9597_;
  assign new_n9603_ = new_n9590_ & new_n9597_;
  assign new_n9604_ = new_n15141_ & new_n10313_;
  assign new_n9605_ = new_n11450_ & new_n10624_;
  assign new_n9606_ = new_n9605_ & new_n9604_;
  assign new_n9607_ = new_n15141_ & pi0760;
  assign new_n9608_ = new_n9605_ & new_n9607_;
  assign new_n9609_ = new_n10623_ & new_n10313_;
  assign new_n9610_ = new_n9605_ & new_n9609_;
  assign new_n9611_ = pi0760 & new_n10623_;
  assign new_n9612_ = new_n9605_ & new_n9611_;
  assign new_n9613_ = new_n10624_ & new_n10594_;
  assign new_n9614_ = new_n9613_ & new_n9604_;
  assign new_n9615_ = new_n9613_ & new_n9607_;
  assign new_n9616_ = new_n9613_ & new_n9609_;
  assign new_n9617_ = new_n9613_ & new_n9611_;
  assign new_n9618_ = new_n11450_ & new_n15190_;
  assign new_n9619_ = new_n9618_ & new_n9604_;
  assign new_n9620_ = new_n9618_ & new_n9607_;
  assign new_n9621_ = new_n9618_ & new_n9609_;
  assign new_n9622_ = new_n9618_ & new_n9611_;
  assign new_n9623_ = new_n15190_ & new_n10594_;
  assign new_n9624_ = new_n9604_ & new_n9623_;
  assign new_n9625_ = new_n9607_ & new_n9623_;
  assign new_n9626_ = new_n9609_ & new_n9623_;
  assign new_n9627_ = new_n9611_ & new_n9623_;
  assign new_n9628_ = pi0956 & new_n9432_;
  assign new_n9629_ = new_n9418_ & new_n9401_;
  assign new_n9630_ = new_n10591_ & new_n10590_ & new_n11498_ & new_n14622_;
  assign new_n9631_ = new_n12631_ & new_n9477_;
  assign new_n9632_ = ~new_n11315_ | ~new_n11314_;
  assign new_n9633_ = ~new_n11313_ | ~new_n11312_;
  assign new_n9634_ = ~new_n11311_ | ~new_n11310_;
  assign new_n9635_ = ~new_n11309_ | ~new_n11308_;
  assign new_n9636_ = ~new_n11307_ | ~new_n11306_;
  assign new_n9637_ = ~new_n11305_ | ~new_n11304_;
  assign new_n9638_ = ~new_n11303_ | ~new_n11302_;
  assign new_n9639_ = ~new_n11301_ | ~new_n11300_;
  assign new_n9640_ = ~new_n11298_ | ~new_n11296_ | ~new_n11297_ | ~new_n11299_;
  assign new_n9641_ = ~new_n11294_ | ~new_n11292_ | ~new_n11293_ | ~new_n11295_;
  assign new_n9642_ = ~new_n11290_ | ~new_n11288_ | ~new_n11289_ | ~new_n11291_;
  assign new_n9643_ = ~new_n11286_ | ~new_n11284_ | ~new_n11285_ | ~new_n11287_;
  assign new_n9644_ = ~new_n11282_ | ~new_n11280_ | ~new_n11281_ | ~new_n11283_;
  assign new_n9645_ = ~new_n11278_ | ~new_n11276_ | ~new_n11277_ | ~new_n11279_;
  assign new_n9646_ = ~new_n11274_ | ~new_n11272_ | ~new_n11273_ | ~new_n11275_;
  assign new_n9647_ = ~new_n11270_ | ~new_n11268_ | ~new_n11269_ | ~new_n11271_;
  assign new_n9648_ = ~new_n11266_ | ~new_n11264_ | ~new_n11265_ | ~new_n11267_;
  assign new_n9649_ = ~new_n11262_ | ~new_n11260_ | ~new_n11261_ | ~new_n11263_;
  assign new_n9650_ = ~new_n11258_ | ~new_n11256_ | ~new_n11257_ | ~new_n11259_;
  assign new_n9651_ = ~new_n11254_ | ~new_n11252_ | ~new_n11253_ | ~new_n11255_;
  assign new_n9652_ = ~new_n11250_ | ~new_n11248_ | ~new_n11249_ | ~new_n11251_;
  assign new_n9653_ = ~new_n11246_ | ~new_n11244_ | ~new_n11245_ | ~new_n11247_;
  assign new_n9654_ = ~new_n11242_ | ~new_n11240_ | ~new_n11241_ | ~new_n11243_;
  assign new_n9655_ = ~new_n11238_ | ~new_n11236_ | ~new_n11237_ | ~new_n11239_;
  assign new_n9656_ = pi0756 & new_n10560_;
  assign new_n9657_ = ~new_n10747_ | ~new_n10746_;
  assign new_n9658_ = ~new_n10735_ | ~new_n10734_;
  assign new_n9659_ = ~new_n11391_ | ~new_n14494_;
  assign new_n9660_ = ~new_n11392_ | ~new_n14497_;
  assign new_n9661_ = ~new_n11394_ | ~new_n14503_;
  assign new_n9662_ = ~new_n11395_ | ~new_n14506_;
  assign new_n9663_ = ~new_n11396_ | ~new_n14509_;
  assign new_n9664_ = ~new_n11397_ | ~new_n14512_;
  assign new_n9665_ = ~new_n11398_ | ~new_n14515_;
  assign new_n9666_ = ~new_n11399_ | ~new_n14518_;
  assign new_n9667_ = ~new_n11400_ | ~new_n14521_;
  assign new_n9668_ = ~new_n11401_ | ~new_n14524_;
  assign new_n9669_ = ~new_n11402_ | ~new_n14527_;
  assign new_n9670_ = ~new_n11403_ | ~new_n14530_;
  assign new_n9671_ = ~new_n11405_ | ~new_n14536_;
  assign new_n9672_ = ~new_n11406_ | ~new_n14539_;
  assign new_n9673_ = ~new_n11407_ | ~new_n14542_;
  assign new_n9674_ = ~new_n11408_ | ~new_n14545_;
  assign new_n9675_ = ~new_n11409_ | ~new_n14549_ | ~new_n14548_;
  assign new_n9676_ = ~new_n11410_ | ~new_n14553_ | ~new_n14552_;
  assign new_n9677_ = ~new_n11411_ | ~new_n14557_ | ~new_n14556_;
  assign new_n9678_ = ~new_n11412_ | ~new_n14561_ | ~new_n14560_;
  assign new_n9679_ = ~new_n11413_ | ~new_n14565_ | ~new_n14564_;
  assign new_n9680_ = ~new_n11414_ | ~new_n14569_ | ~new_n14568_;
  assign new_n9681_ = ~new_n11385_ | ~new_n14475_ | ~new_n14474_;
  assign new_n9682_ = ~new_n11386_ | ~new_n14479_ | ~new_n14478_;
  assign new_n9683_ = ~new_n11387_ | ~new_n14482_;
  assign new_n9684_ = ~new_n11388_ | ~new_n14485_;
  assign new_n9685_ = ~new_n11389_ | ~new_n14488_;
  assign new_n9686_ = ~new_n11390_ | ~new_n14491_;
  assign new_n9687_ = ~new_n11393_ | ~new_n14500_;
  assign new_n9688_ = ~new_n11404_ | ~new_n14533_;
  assign new_n9689_ = ~new_n11415_ | ~new_n14572_;
  assign new_n9690_ = ~new_n11416_ | ~new_n14575_ | ~new_n10341_;
  assign new_n9691_ = new_n9393_ & new_n10283_;
  assign new_n9692_ = new_n9393_ & new_n14258_;
  assign new_n9693_ = new_n9393_ & new_n14292_;
  assign new_n9694_ = new_n9393_ & new_n14326_;
  assign new_n9695_ = ~new_n14464_ | ~new_n14463_;
  assign new_n9696_ = ~new_n11379_ | ~new_n14465_;
  assign new_n9697_ = ~new_n11381_ | ~new_n14468_;
  assign new_n9698_ = ~new_n11383_ | ~new_n14470_;
  assign new_n9699_ = new_n9395_ & new_n9639_;
  assign new_n9700_ = new_n9395_ & new_n9638_;
  assign new_n9701_ = new_n9395_ & new_n9637_;
  assign new_n9702_ = new_n9395_ & new_n9636_;
  assign new_n9703_ = new_n9395_ & new_n9635_;
  assign new_n9704_ = new_n9395_ & new_n9634_;
  assign new_n9705_ = new_n9395_ & new_n9633_;
  assign new_n9706_ = new_n9395_ & new_n9632_;
  assign new_n9707_ = new_n9655_ & new_n9396_;
  assign new_n9708_ = new_n9654_ & new_n9396_;
  assign new_n9709_ = new_n9653_ & new_n9396_;
  assign new_n9710_ = new_n9652_ & new_n9396_;
  assign new_n9711_ = new_n9651_ & new_n9396_;
  assign new_n9712_ = new_n9650_ & new_n9396_;
  assign new_n9713_ = new_n9649_ & new_n9396_;
  assign new_n9714_ = new_n9648_ & new_n9396_;
  assign new_n9715_ = pi0748 & new_n9396_;
  assign new_n9716_ = pi0749 & new_n9396_;
  assign new_n9717_ = pi0750 & new_n9396_;
  assign new_n9718_ = pi0751 & new_n9396_;
  assign new_n9719_ = pi0752 & new_n9396_;
  assign new_n9720_ = pi0753 & new_n9396_;
  assign new_n9721_ = pi0754 & new_n9396_;
  assign new_n9722_ = ~new_n14207_ | ~new_n11316_;
  assign new_n9723_ = new_n9396_ & new_n28262_;
  assign new_n9724_ = new_n28263_ & new_n9396_;
  assign new_n9725_ = new_n28268_ & new_n9396_;
  assign new_n9726_ = new_n28266_ & new_n9396_;
  assign new_n9727_ = new_n28265_ & new_n9396_;
  assign new_n9728_ = new_n28269_ & new_n9396_;
  assign new_n9729_ = new_n28264_ & new_n9396_;
  assign new_n9730_ = ~new_n14183_ | ~new_n14182_;
  assign new_n9731_ = ~new_n14185_ | ~new_n14184_;
  assign new_n9732_ = ~new_n14187_ | ~new_n14186_;
  assign new_n9733_ = ~new_n14189_ | ~new_n14188_;
  assign new_n9734_ = ~new_n14194_ | ~new_n14193_;
  assign new_n9735_ = ~new_n14196_ | ~new_n14195_;
  assign new_n9736_ = ~new_n14198_ | ~new_n14197_;
  assign new_n9737_ = ~new_n14200_ | ~new_n14199_;
  assign new_n9738_ = ~new_n20992_ | ~new_n33663_;
  assign new_n9739_ = pi0756 & new_n10595_;
  assign new_n9740_ = ~new_n14179_ | ~new_n14180_ | ~new_n14181_;
  assign new_n9741_ = ~new_n14190_ | ~new_n14191_ | ~new_n14192_;
  assign new_n9742_ = ~new_n14201_ | ~new_n14202_ | ~new_n14203_;
  assign new_n9743_ = ~new_n14204_ | ~new_n14205_ | ~new_n14206_;
  assign new_n9744_ = ~new_n14768_ | ~new_n14767_;
  assign new_n9745_ = ~new_n14770_ | ~new_n14769_;
  assign new_n9746_ = ~new_n11431_ | ~new_n14771_;
  assign new_n9747_ = ~new_n10591_ | ~new_n14773_ | ~new_n14774_;
  assign new_n9748_ = ~new_n11432_ | ~new_n14775_;
  assign new_n9749_ = new_n29038_ & new_n14764_;
  assign new_n9750_ = new_n29039_ & new_n14764_;
  assign new_n9751_ = new_n29040_ & new_n14764_;
  assign new_n9752_ = ~pi0627 | ~new_n14765_;
  assign new_n9753_ = ~new_n11448_ | ~new_n14912_ | ~pi0627;
  assign new_n9754_ = ~pi0627 | ~new_n14766_;
  assign new_n9755_ = ~new_n11449_ | ~new_n14912_ | ~pi0627;
  assign new_n9756_ = ~new_n9397_ | ~new_n9657_;
  assign new_n9757_ = ~new_n14660_ | ~new_n14658_ | ~new_n14659_ | ~new_n14661_;
  assign new_n9758_ = ~new_n14664_ | ~new_n14662_ | ~new_n14663_ | ~new_n14665_;
  assign new_n9759_ = ~new_n14672_ | ~new_n14670_ | ~new_n14671_ | ~new_n14673_;
  assign new_n9760_ = ~new_n14676_ | ~new_n14674_ | ~new_n14675_ | ~new_n14677_;
  assign new_n9761_ = ~new_n14680_ | ~new_n14678_ | ~new_n14679_ | ~new_n14681_;
  assign new_n9762_ = ~new_n14684_ | ~new_n14682_ | ~new_n14683_ | ~new_n14685_;
  assign new_n9763_ = ~new_n14688_ | ~new_n14686_ | ~new_n14687_ | ~new_n14689_;
  assign new_n9764_ = ~new_n14692_ | ~new_n14690_ | ~new_n14691_ | ~new_n14693_;
  assign new_n9765_ = ~new_n14696_ | ~new_n14694_ | ~new_n14695_ | ~new_n14697_;
  assign new_n9766_ = ~new_n14700_ | ~new_n14698_ | ~new_n14699_ | ~new_n14701_;
  assign new_n9767_ = ~new_n14704_ | ~new_n14702_ | ~new_n14703_ | ~new_n14705_;
  assign new_n9768_ = ~new_n14708_ | ~new_n14706_ | ~new_n14707_ | ~new_n14709_;
  assign new_n9769_ = ~new_n14716_ | ~new_n14714_ | ~new_n14715_ | ~new_n14717_;
  assign new_n9770_ = ~new_n14720_ | ~new_n14718_ | ~new_n14719_ | ~new_n14721_;
  assign new_n9771_ = ~new_n14724_ | ~new_n14722_ | ~new_n14723_ | ~new_n14725_;
  assign new_n9772_ = ~new_n14728_ | ~new_n14726_ | ~new_n14727_ | ~new_n14729_;
  assign new_n9773_ = ~new_n14732_ | ~new_n14730_ | ~new_n14731_ | ~new_n14733_;
  assign new_n9774_ = ~new_n14736_ | ~new_n14734_ | ~new_n14735_ | ~new_n14737_;
  assign new_n9775_ = ~new_n14740_ | ~new_n14738_ | ~new_n14739_ | ~new_n14741_;
  assign new_n9776_ = ~new_n14744_ | ~new_n14742_ | ~new_n14743_ | ~new_n14745_;
  assign new_n9777_ = ~new_n14748_ | ~new_n14746_ | ~new_n14747_ | ~new_n14749_;
  assign new_n9778_ = ~new_n14752_ | ~new_n14750_ | ~new_n14751_ | ~new_n14753_;
  assign new_n9779_ = ~new_n14636_ | ~new_n14634_ | ~new_n14635_ | ~new_n14637_;
  assign new_n9780_ = ~new_n14640_ | ~new_n14638_ | ~new_n14639_ | ~new_n14641_;
  assign new_n9781_ = ~new_n14644_ | ~new_n14642_ | ~new_n14643_ | ~new_n14645_;
  assign new_n9782_ = ~new_n14648_ | ~new_n14646_ | ~new_n14647_ | ~new_n14649_;
  assign new_n9783_ = ~new_n14652_ | ~new_n14650_ | ~new_n14651_ | ~new_n14653_;
  assign new_n9784_ = ~new_n14656_ | ~new_n14654_ | ~new_n14655_ | ~new_n14657_;
  assign new_n9785_ = ~new_n14668_ | ~new_n14666_ | ~new_n14667_ | ~new_n14669_;
  assign new_n9786_ = ~new_n14712_ | ~new_n14710_ | ~new_n14711_ | ~new_n14713_;
  assign new_n9787_ = ~new_n14756_ | ~new_n14754_ | ~new_n14755_ | ~new_n14757_;
  assign new_n9788_ = ~new_n14927_ | ~new_n14758_ | ~new_n11429_ | ~new_n11430_ | ~new_n14762_;
  assign new_n9789_ = ~new_n14624_ | ~new_n14623_;
  assign new_n9790_ = ~new_n11421_ | ~new_n14625_;
  assign new_n9791_ = ~new_n11423_ | ~new_n14629_;
  assign new_n9792_ = new_n14929_ & new_n14778_;
  assign new_n9793_ = new_n14914_ & new_n10321_ & pi0756;
  assign new_n9794_ = ~new_n10327_ | ~new_n14613_;
  assign new_n9795_ = ~new_n10327_ | ~new_n14614_;
  assign new_n9796_ = ~new_n10327_ | ~new_n14615_;
  assign new_n9797_ = ~new_n10327_ | ~new_n14616_;
  assign new_n9798_ = ~new_n10327_ | ~new_n14617_;
  assign new_n9799_ = new_n11469_ & new_n10283_;
  assign new_n9800_ = new_n11469_ & new_n14258_;
  assign new_n9801_ = new_n11469_ & new_n14292_;
  assign new_n9802_ = ~new_n14604_ | ~new_n14603_;
  assign new_n9803_ = ~new_n14606_ | ~new_n14605_;
  assign new_n9804_ = ~new_n14608_ | ~new_n14607_;
  assign new_n9805_ = ~new_n14610_ | ~new_n14609_;
  assign new_n9806_ = ~new_n14612_ | ~new_n14611_;
  assign new_n9807_ = ~new_n11488_ | ~new_n14580_;
  assign new_n9808_ = ~new_n11488_ | ~new_n14581_;
  assign new_n9809_ = ~new_n11488_ | ~new_n14582_;
  assign new_n9810_ = ~new_n11488_ | ~new_n14583_;
  assign new_n9811_ = ~new_n11488_ | ~new_n14584_;
  assign new_n9812_ = ~new_n11488_ | ~new_n14585_;
  assign new_n9813_ = ~new_n11488_ | ~new_n14586_;
  assign new_n9814_ = ~new_n11488_ | ~new_n14587_;
  assign new_n9815_ = ~new_n11488_ | ~new_n14588_;
  assign new_n9816_ = ~new_n11488_ | ~new_n14589_;
  assign new_n9817_ = ~new_n11488_ | ~new_n14590_;
  assign new_n9818_ = ~new_n11488_ | ~new_n14591_;
  assign new_n9819_ = ~new_n11488_ | ~new_n14592_;
  assign new_n9820_ = ~new_n11488_ | ~new_n14593_;
  assign new_n9821_ = ~new_n11488_ | ~new_n14594_;
  assign new_n9822_ = ~new_n11488_ | ~new_n14595_;
  assign new_n9823_ = ~new_n11488_ | ~new_n14596_;
  assign new_n9824_ = ~new_n11488_ | ~new_n14597_;
  assign new_n9825_ = ~new_n11488_ | ~new_n14598_;
  assign new_n9826_ = ~new_n11488_ | ~new_n14599_;
  assign new_n9827_ = ~new_n11488_ | ~new_n14600_;
  assign new_n9828_ = ~new_n11488_ | ~new_n14601_;
  assign new_n9829_ = ~new_n11488_ | ~new_n14578_;
  assign new_n9830_ = ~new_n11488_ | ~new_n14579_;
  assign new_n9831_ = new_n10283_ & new_n30569_;
  assign new_n9832_ = new_n10283_ & new_n30522_;
  assign new_n9833_ = new_n10283_ & new_n30521_;
  assign new_n9834_ = new_n10283_ & new_n30573_;
  assign new_n9835_ = new_n10283_ & new_n30520_;
  assign new_n9836_ = new_n10283_ & new_n30575_;
  assign new_n9837_ = new_n10283_ & new_n30519_;
  assign new_n9838_ = new_n10283_ & new_n30577_;
  assign new_n9839_ = new_n10283_ & new_n30518_;
  assign new_n9840_ = new_n10283_ & new_n30579_;
  assign new_n9841_ = new_n10283_ & new_n30517_;
  assign new_n9842_ = new_n10283_ & new_n30581_;
  assign new_n9843_ = new_n10283_ & new_n30516_;
  assign new_n9844_ = new_n10283_ & new_n30585_;
  assign new_n9845_ = new_n10283_ & new_n30515_;
  assign new_n9846_ = new_n10283_ & new_n30587_;
  assign new_n9847_ = new_n10283_ & new_n30514_;
  assign new_n9848_ = new_n10283_ & new_n30589_;
  assign new_n9849_ = new_n10283_ & new_n30513_;
  assign new_n9850_ = new_n10283_ & new_n30591_;
  assign new_n9851_ = new_n10283_ & new_n30512_;
  assign new_n9852_ = new_n10283_ & new_n30593_;
  assign new_n9853_ = new_n10283_ & new_n30526_;
  assign new_n9854_ = pi0757 & new_n10560_;
  assign po1062 = ~new_n11231_ | ~new_n13902_;
  assign po1060 = ~new_n14958_ | ~new_n13897_;
  assign po1059 = ~new_n13896_ | ~new_n13895_;
  assign po1057 = ~new_n11504_ | ~new_n15181_ | ~new_n15180_;
  assign po1055 = ~new_n11504_ | ~new_n15177_ | ~new_n15176_;
  assign po1053 = ~new_n13881_ | ~new_n13880_;
  assign po1051 = ~new_n10589_ | ~new_n15169_ | ~new_n15168_;
  assign po1050 = ~new_n13878_ | ~new_n10589_ | ~new_n11493_;
  assign po1049 = ~new_n11439_ | ~new_n13877_;
  assign po1048 = ~new_n11493_ | ~new_n15165_ | ~new_n15164_;
  assign po1047 = ~new_n13868_ | ~new_n13869_ | ~new_n13871_ | ~new_n11209_ | ~new_n13870_;
  assign po1046 = ~new_n13860_ | ~new_n13861_ | ~new_n13863_ | ~new_n11207_ | ~new_n13862_;
  assign po1045 = ~new_n13852_ | ~new_n13853_ | ~new_n13855_ | ~new_n11205_ | ~new_n13854_;
  assign po1044 = ~new_n13844_ | ~new_n13845_ | ~new_n13847_ | ~new_n11203_ | ~new_n13846_;
  assign po1043 = ~new_n13836_ | ~new_n13837_ | ~new_n13839_ | ~new_n11201_ | ~new_n13838_;
  assign po1042 = ~new_n13828_ | ~new_n13829_ | ~new_n13831_ | ~new_n11199_ | ~new_n13830_;
  assign po1041 = ~new_n13820_ | ~new_n13821_ | ~new_n11197_ | ~new_n13823_ | ~new_n13822_;
  assign po1040 = ~new_n13813_ | ~new_n11193_;
  assign po1039 = ~new_n13805_ | ~new_n11190_;
  assign po1038 = ~new_n13796_ | ~new_n11189_ | ~new_n13797_ | ~new_n13799_ | ~new_n13798_;
  assign po1037 = ~new_n11187_ | ~new_n11185_;
  assign po1036 = ~new_n11184_ | ~new_n11182_;
  assign po1035 = ~new_n11181_ | ~new_n11179_;
  assign po1034 = ~new_n11177_ | ~new_n11175_;
  assign po1033 = ~new_n11173_ | ~new_n11171_;
  assign po1032 = ~new_n11169_ | ~new_n11167_;
  assign po1031 = ~new_n11165_ | ~new_n11163_;
  assign po1030 = ~new_n13734_ | ~new_n11160_ | ~new_n13737_ | ~new_n13733_ | ~new_n11159_;
  assign po1029 = ~new_n13726_ | ~new_n11157_ | ~new_n13729_ | ~new_n13725_ | ~new_n11156_;
  assign po1028 = ~new_n13718_ | ~new_n11154_ | ~new_n13721_ | ~new_n13717_ | ~new_n11153_;
  assign po1027 = ~new_n13711_ | ~new_n11151_ | ~new_n13713_ | ~new_n11150_ | ~new_n13710_;
  assign po1026 = ~new_n13703_ | ~new_n11148_ | ~new_n13705_ | ~new_n11147_ | ~new_n13702_;
  assign po1025 = ~new_n13695_ | ~new_n11145_ | ~new_n13697_ | ~new_n11144_ | ~new_n13694_;
  assign po1024 = ~new_n13687_ | ~new_n11142_ | ~new_n13689_ | ~new_n11141_ | ~new_n13686_;
  assign po1023 = ~new_n13679_ | ~new_n11139_ | ~new_n13681_ | ~new_n11138_ | ~new_n13678_;
  assign po1022 = ~new_n13671_ | ~new_n11136_ | ~new_n13673_ | ~new_n11135_ | ~new_n13670_;
  assign po1021 = ~new_n11134_ | ~new_n11132_;
  assign po1020 = ~new_n11130_ | ~new_n11128_;
  assign po1019 = ~new_n11123_ | ~new_n11125_ | ~new_n13647_ | ~new_n13643_;
  assign po1018 = ~new_n11119_ | ~new_n11121_ | ~new_n13638_ | ~new_n13634_;
  assign po1017 = ~new_n11115_ | ~new_n11117_ | ~new_n13629_ | ~new_n13625_;
  assign po1016 = ~new_n11111_ | ~new_n11113_ | ~new_n13620_ | ~new_n13616_;
  assign po1015 = ~new_n13606_ | ~new_n13605_;
  assign po1014 = ~new_n13602_ | ~new_n13603_ | ~new_n13604_;
  assign po1013 = ~new_n13599_ | ~new_n13600_ | ~new_n13601_;
  assign po1012 = ~new_n13596_ | ~new_n13597_ | ~new_n13598_;
  assign po1011 = ~new_n13593_ | ~new_n13594_ | ~new_n13595_;
  assign po1010 = ~new_n13590_ | ~new_n13591_ | ~new_n13592_;
  assign po1009 = ~new_n13587_ | ~new_n13588_ | ~new_n13589_;
  assign po1008 = ~new_n13584_ | ~new_n13585_ | ~new_n13586_;
  assign po1007 = ~new_n13581_ | ~new_n13582_ | ~new_n13583_;
  assign po1006 = ~new_n13578_ | ~new_n13579_ | ~new_n13580_;
  assign po1005 = ~new_n13575_ | ~new_n13576_ | ~new_n13577_;
  assign po1004 = ~new_n13572_ | ~new_n13573_ | ~new_n13574_;
  assign po1003 = ~new_n13569_ | ~new_n13570_ | ~new_n13571_;
  assign po1002 = ~new_n13566_ | ~new_n13567_ | ~new_n13568_;
  assign po1001 = ~new_n13563_ | ~new_n13564_ | ~new_n13565_;
  assign po1000 = ~new_n13560_ | ~new_n13561_ | ~new_n13562_;
  assign po0999 = ~new_n13557_ | ~new_n13558_ | ~new_n13559_;
  assign po0998 = ~new_n13554_ | ~new_n13555_ | ~new_n13556_;
  assign po0997 = ~new_n13551_ | ~new_n13552_ | ~new_n13553_;
  assign po0996 = ~new_n13548_ | ~new_n13549_ | ~new_n13550_;
  assign po0995 = ~new_n13545_ | ~new_n13546_ | ~new_n13547_;
  assign po0994 = ~new_n13542_ | ~new_n13543_ | ~new_n13544_;
  assign po0993 = ~new_n13539_ | ~new_n13540_ | ~new_n13541_;
  assign po0992 = ~new_n13536_ | ~new_n13537_ | ~new_n13538_;
  assign po0991 = ~new_n13535_ | ~new_n13534_ | ~new_n13533_;
  assign po0990 = ~new_n13532_ | ~new_n13531_ | ~new_n13530_;
  assign po0989 = ~new_n13529_ | ~new_n13528_ | ~new_n13527_;
  assign po0988 = ~new_n13526_ | ~new_n13525_ | ~new_n13524_;
  assign po0987 = ~new_n13523_ | ~new_n13522_ | ~new_n13521_;
  assign po0986 = ~new_n13520_ | ~new_n13519_ | ~new_n13518_;
  assign po0985 = ~new_n13517_ | ~new_n13516_ | ~new_n13515_;
  assign po0984 = ~new_n13514_ | ~new_n13513_ | ~new_n13512_;
  assign po0983 = ~new_n13508_ | ~new_n13509_ | ~new_n13507_;
  assign po0982 = ~new_n13503_ | ~new_n13504_ | ~new_n13505_ | ~new_n13506_ | ~new_n13502_;
  assign po0981 = ~new_n13498_ | ~new_n13499_ | ~new_n13500_ | ~new_n13501_ | ~new_n13497_;
  assign po0980 = ~new_n13493_ | ~new_n13494_ | ~new_n13495_ | ~new_n13496_ | ~new_n13492_;
  assign po0979 = ~new_n13488_ | ~new_n13489_ | ~new_n13490_ | ~new_n13491_ | ~new_n13487_;
  assign po0978 = ~new_n13483_ | ~new_n13484_ | ~new_n13485_ | ~new_n13486_ | ~new_n13482_;
  assign po0977 = ~new_n13478_ | ~new_n13479_ | ~new_n13480_ | ~new_n13481_ | ~new_n13477_;
  assign po0976 = ~new_n13473_ | ~new_n13474_ | ~new_n13475_ | ~new_n13476_ | ~new_n13472_;
  assign po0975 = ~new_n13468_ | ~new_n13469_ | ~new_n13470_ | ~new_n13471_ | ~new_n13467_;
  assign po0974 = ~new_n13463_ | ~new_n13464_ | ~new_n13465_ | ~new_n13466_ | ~new_n13462_;
  assign po0973 = ~new_n13458_ | ~new_n13459_ | ~new_n13460_ | ~new_n13461_ | ~new_n13457_;
  assign po0972 = ~new_n13453_ | ~new_n13454_ | ~new_n13455_ | ~new_n13456_ | ~new_n13452_;
  assign po0971 = ~new_n13448_ | ~new_n13449_ | ~new_n13450_ | ~new_n13451_ | ~new_n13447_;
  assign po0970 = ~new_n13443_ | ~new_n13444_ | ~new_n13445_ | ~new_n13446_ | ~new_n13442_;
  assign po0969 = ~new_n13438_ | ~new_n13439_ | ~new_n13440_ | ~new_n13441_ | ~new_n13437_;
  assign po0968 = ~new_n13433_ | ~new_n13434_ | ~new_n13435_ | ~new_n13436_ | ~new_n13432_;
  assign po0967 = ~new_n13428_ | ~new_n13429_ | ~new_n13430_ | ~new_n13431_;
  assign po0966 = ~new_n13424_ | ~new_n13425_ | ~new_n13426_ | ~new_n13427_;
  assign po0965 = ~new_n13420_ | ~new_n13421_ | ~new_n13422_ | ~new_n13423_;
  assign po0964 = ~new_n13416_ | ~new_n13417_ | ~new_n13418_ | ~new_n13419_;
  assign po0963 = ~new_n13412_ | ~new_n13413_ | ~new_n13414_ | ~new_n13415_;
  assign po0962 = ~new_n13408_ | ~new_n13409_ | ~new_n13410_ | ~new_n13411_;
  assign po0961 = ~new_n13405_ | ~new_n11109_ | ~new_n13404_;
  assign po0960 = ~new_n13401_ | ~new_n11108_ | ~new_n13400_;
  assign po0959 = ~new_n13397_ | ~new_n11107_ | ~new_n13396_;
  assign po0958 = ~new_n11106_ | ~new_n13393_ | ~new_n13392_;
  assign po0957 = ~new_n11105_ | ~new_n13389_ | ~new_n13388_;
  assign po0956 = ~new_n11104_ | ~new_n13385_ | ~new_n13384_;
  assign po0955 = ~new_n11103_ | ~new_n13381_ | ~new_n13380_;
  assign po0954 = ~new_n11102_ | ~new_n13377_ | ~new_n13376_;
  assign po0953 = ~new_n11101_ | ~new_n13373_ | ~new_n13372_;
  assign po0952 = ~new_n11100_ | ~new_n13369_ | ~new_n13368_;
  assign po0951 = pi0892 & new_n13273_;
  assign po0950 = ~new_n13366_ | ~new_n13365_ | ~new_n13364_;
  assign po0949 = ~new_n13363_ | ~new_n13362_ | ~new_n13361_;
  assign po0948 = ~new_n13360_ | ~new_n13359_ | ~new_n13358_;
  assign po0947 = ~new_n13357_ | ~new_n13356_ | ~new_n13355_;
  assign po0946 = ~new_n13354_ | ~new_n13353_ | ~new_n13352_;
  assign po0945 = ~new_n13351_ | ~new_n13350_ | ~new_n13349_;
  assign po0944 = ~new_n13348_ | ~new_n13347_ | ~new_n13346_;
  assign po0943 = ~new_n13345_ | ~new_n13344_ | ~new_n13343_;
  assign po0942 = ~new_n13342_ | ~new_n13341_ | ~new_n13340_;
  assign po0941 = ~new_n13339_ | ~new_n13338_ | ~new_n13337_;
  assign po0940 = ~new_n13336_ | ~new_n13335_ | ~new_n13334_;
  assign po0939 = ~new_n13333_ | ~new_n13332_ | ~new_n13331_;
  assign po0938 = ~new_n13330_ | ~new_n13329_ | ~new_n13328_;
  assign po0937 = ~new_n13327_ | ~new_n13326_ | ~new_n13325_;
  assign po0936 = ~new_n13324_ | ~new_n13323_ | ~new_n13322_;
  assign po0935 = ~new_n13321_ | ~new_n13320_ | ~new_n13319_;
  assign po0934 = ~new_n13318_ | ~new_n13317_ | ~new_n13316_;
  assign po0933 = ~new_n13315_ | ~new_n13314_ | ~new_n13313_;
  assign po0932 = ~new_n13312_ | ~new_n13311_ | ~new_n13310_;
  assign po0931 = ~new_n13309_ | ~new_n13308_ | ~new_n13307_;
  assign po0930 = ~new_n13306_ | ~new_n13305_ | ~new_n13304_;
  assign po0929 = ~new_n13303_ | ~new_n13302_ | ~new_n13301_;
  assign po0928 = ~new_n13300_ | ~new_n13299_ | ~new_n13298_;
  assign po0927 = ~new_n13297_ | ~new_n13296_ | ~new_n13295_;
  assign po0926 = ~new_n13294_ | ~new_n13293_ | ~new_n13292_;
  assign po0925 = ~new_n13291_ | ~new_n13290_ | ~new_n13289_;
  assign po0924 = ~new_n13288_ | ~new_n13287_ | ~new_n13286_;
  assign po0923 = ~new_n13285_ | ~new_n13284_ | ~new_n13283_;
  assign po0922 = ~new_n13282_ | ~new_n13281_ | ~new_n13280_;
  assign po0921 = ~new_n13279_ | ~new_n13278_ | ~new_n13277_;
  assign po0920 = ~new_n13276_ | ~new_n13275_ | ~new_n13274_;
  assign po0919 = ~new_n13267_ | ~new_n13266_ | ~new_n13265_;
  assign po0918 = ~new_n13264_ | ~new_n13263_ | ~new_n13262_;
  assign po0917 = ~new_n13261_ | ~new_n13260_ | ~new_n13259_;
  assign po0916 = ~new_n13258_ | ~new_n13257_ | ~new_n13256_;
  assign po0915 = ~new_n13255_ | ~new_n13254_ | ~new_n13253_;
  assign po0914 = ~new_n13252_ | ~new_n13251_ | ~new_n13250_;
  assign po0913 = ~new_n13249_ | ~new_n13248_ | ~new_n13247_;
  assign po0912 = ~new_n13246_ | ~new_n13245_ | ~new_n13244_;
  assign po0911 = ~new_n13243_ | ~new_n13242_ | ~new_n13241_;
  assign po0910 = ~new_n13240_ | ~new_n13239_ | ~new_n13238_;
  assign po0909 = ~new_n13237_ | ~new_n13236_ | ~new_n13235_;
  assign po0908 = ~new_n13234_ | ~new_n13233_ | ~new_n13232_;
  assign po0907 = ~new_n13231_ | ~new_n13230_ | ~new_n13229_;
  assign po0906 = ~new_n13228_ | ~new_n13227_ | ~new_n13226_;
  assign po0905 = ~new_n13225_ | ~new_n13224_ | ~new_n13223_;
  assign po0904 = ~new_n13222_ | ~new_n13221_ | ~new_n13220_;
  assign po0903 = ~new_n13219_ | ~new_n13218_ | ~new_n13217_;
  assign po0902 = ~new_n13216_ | ~new_n13215_ | ~new_n13214_;
  assign po0901 = ~new_n13213_ | ~new_n13212_ | ~new_n13211_;
  assign po0900 = ~new_n13210_ | ~new_n13209_ | ~new_n13208_;
  assign po0899 = ~new_n13207_ | ~new_n13206_ | ~new_n13205_;
  assign po0898 = ~new_n13204_ | ~new_n13203_ | ~new_n13202_;
  assign po0897 = ~new_n13201_ | ~new_n13200_ | ~new_n13199_;
  assign po0896 = ~new_n13198_ | ~new_n13197_ | ~new_n13196_;
  assign po0895 = ~new_n13195_ | ~new_n13194_ | ~new_n13193_;
  assign po0894 = ~new_n13192_ | ~new_n13191_ | ~new_n13190_;
  assign po0893 = ~new_n13189_ | ~new_n13188_ | ~new_n13187_;
  assign po0892 = ~new_n13186_ | ~new_n13185_ | ~new_n13184_;
  assign po0891 = ~new_n13183_ | ~new_n13182_ | ~new_n13181_;
  assign po0890 = ~new_n13180_ | ~new_n13179_ | ~new_n13178_;
  assign po0889 = ~new_n13177_ | ~new_n13176_ | ~new_n13175_;
  assign po0888 = ~new_n11095_ | ~new_n11094_;
  assign po0887 = ~new_n11093_ | ~new_n11092_;
  assign po0886 = ~new_n11091_ | ~new_n11090_;
  assign po0885 = ~new_n11089_ | ~new_n11088_;
  assign po0884 = ~new_n11087_ | ~new_n11086_;
  assign po0883 = ~new_n11085_ | ~new_n11084_;
  assign po0882 = ~new_n11083_ | ~new_n11082_;
  assign po0881 = ~new_n11081_ | ~new_n11080_;
  assign po0880 = ~new_n11079_ | ~new_n11078_;
  assign po0879 = ~new_n11077_ | ~new_n11076_;
  assign po0878 = ~new_n11075_ | ~new_n11074_;
  assign po0877 = ~new_n11073_ | ~new_n11072_;
  assign po0876 = ~new_n11071_ | ~new_n11070_;
  assign po0875 = ~new_n11069_ | ~new_n11068_;
  assign po0874 = ~new_n11067_ | ~new_n11066_;
  assign po0873 = ~new_n11065_ | ~new_n11064_;
  assign po0872 = ~new_n11063_ | ~new_n11062_;
  assign po0871 = ~new_n11061_ | ~new_n11060_;
  assign po0870 = ~new_n11059_ | ~new_n11058_;
  assign po0869 = ~new_n11057_ | ~new_n11056_;
  assign po0868 = ~new_n11055_ | ~new_n11054_;
  assign po0867 = ~new_n11053_ | ~new_n11052_;
  assign po0866 = ~new_n11051_ | ~new_n11050_;
  assign po0865 = ~new_n11049_ | ~new_n11048_;
  assign po0864 = ~new_n11047_ | ~new_n11046_;
  assign po0863 = ~new_n11045_ | ~new_n11044_;
  assign po0862 = ~new_n11043_ | ~new_n11042_;
  assign po0861 = ~new_n11041_ | ~new_n11040_;
  assign po0860 = ~new_n11039_ | ~new_n11038_;
  assign po0859 = ~new_n11037_ | ~new_n11036_;
  assign po0858 = ~new_n11035_ | ~new_n11034_;
  assign po0857 = ~new_n11033_ | ~new_n11032_;
  assign po0856 = ~new_n12974_ | ~new_n12969_ | ~new_n11028_ | ~new_n11029_ | ~new_n12973_;
  assign po0855 = ~new_n12966_ | ~new_n12961_ | ~new_n11026_ | ~new_n11027_ | ~new_n12965_;
  assign po0854 = ~new_n12957_ | ~new_n11024_ | ~new_n11025_ | ~new_n12958_;
  assign po0853 = ~new_n12950_ | ~new_n11021_ | ~new_n11022_ | ~new_n11023_ | ~new_n12949_;
  assign po0852 = ~new_n12942_ | ~new_n11018_ | ~new_n11019_ | ~new_n11020_ | ~new_n12941_;
  assign po0851 = ~new_n12934_ | ~new_n11015_ | ~new_n11016_ | ~new_n11017_ | ~new_n12933_;
  assign po0850 = ~new_n12926_ | ~new_n11012_ | ~new_n11013_ | ~new_n11014_ | ~new_n12925_;
  assign po0849 = ~new_n12918_ | ~new_n11009_ | ~new_n11010_ | ~new_n11011_ | ~new_n12917_;
  assign po0848 = ~new_n12910_ | ~new_n11006_ | ~new_n11007_ | ~new_n11008_ | ~new_n12909_;
  assign po0847 = ~new_n12902_ | ~new_n11003_ | ~new_n11004_ | ~new_n11005_ | ~new_n12901_;
  assign po0846 = ~new_n12894_ | ~new_n11000_ | ~new_n11001_ | ~new_n11002_ | ~new_n12893_;
  assign po0845 = ~new_n12886_ | ~new_n10997_ | ~new_n10998_ | ~new_n10999_ | ~new_n12885_;
  assign po0844 = ~new_n12878_ | ~new_n10994_ | ~new_n10995_ | ~new_n10996_ | ~new_n12877_;
  assign po0843 = ~new_n12870_ | ~new_n10991_ | ~new_n10992_ | ~new_n10993_ | ~new_n12869_;
  assign po0842 = ~new_n12862_ | ~new_n10988_ | ~new_n10989_ | ~new_n10990_ | ~new_n12861_;
  assign po0841 = ~new_n12854_ | ~new_n10985_ | ~new_n10986_ | ~new_n10987_ | ~new_n12853_;
  assign po0840 = ~new_n12846_ | ~new_n10982_ | ~new_n10983_ | ~new_n10984_ | ~new_n12845_;
  assign po0839 = ~new_n12838_ | ~new_n10979_ | ~new_n10980_ | ~new_n10981_ | ~new_n12837_;
  assign po0838 = ~new_n12830_ | ~new_n10976_ | ~new_n10977_ | ~new_n10978_ | ~new_n12829_;
  assign po0837 = ~new_n12822_ | ~new_n10973_ | ~new_n10974_ | ~new_n10975_ | ~new_n12821_;
  assign po0836 = ~new_n12814_ | ~new_n10970_ | ~new_n10971_ | ~new_n10972_ | ~new_n12813_;
  assign po0835 = ~new_n12806_ | ~new_n10967_ | ~new_n10968_ | ~new_n10969_ | ~new_n12805_;
  assign po0834 = ~new_n12798_ | ~new_n10964_ | ~new_n10965_ | ~new_n10966_ | ~new_n12797_;
  assign po0833 = ~new_n12790_ | ~new_n10961_ | ~new_n10962_ | ~new_n10963_ | ~new_n12789_;
  assign po0832 = ~new_n12782_ | ~new_n10958_ | ~new_n10959_ | ~new_n10960_ | ~new_n12781_;
  assign po0831 = ~new_n12774_ | ~new_n10955_ | ~new_n10956_ | ~new_n10957_ | ~new_n12773_;
  assign po0830 = ~new_n12766_ | ~new_n10952_ | ~new_n10953_ | ~new_n10954_ | ~new_n12765_;
  assign po0829 = ~new_n12758_ | ~new_n10949_ | ~new_n10950_ | ~new_n10951_ | ~new_n12757_;
  assign po0828 = ~new_n12750_ | ~new_n10946_ | ~new_n10947_ | ~new_n10948_ | ~new_n12749_;
  assign po0827 = ~new_n12742_ | ~new_n10943_ | ~new_n10944_ | ~new_n10945_ | ~new_n12741_;
  assign po0826 = ~new_n12734_ | ~new_n10940_ | ~new_n10941_ | ~new_n10942_ | ~new_n12733_;
  assign po0825 = ~new_n12726_ | ~new_n10937_ | ~new_n10938_ | ~new_n10939_ | ~new_n12725_;
  assign po0820 = pi0761 & new_n12684_;
  assign po0814 = ~new_n10906_ | ~new_n12611_ | ~new_n12610_;
  assign po0813 = ~new_n10905_ | ~new_n12606_ | ~new_n12605_;
  assign po0812 = ~new_n10904_ | ~new_n12601_ | ~new_n12600_;
  assign po0811 = ~new_n10903_ | ~new_n12596_ | ~new_n12595_;
  assign po0810 = ~new_n10902_ | ~new_n12591_ | ~new_n12590_;
  assign po0809 = ~new_n10901_ | ~new_n12586_ | ~new_n12585_;
  assign po0808 = ~new_n10900_ | ~new_n12581_ | ~new_n12580_;
  assign po0807 = ~new_n10899_ | ~new_n12576_ | ~new_n12575_;
  assign po0806 = ~new_n10897_ | ~new_n12554_ | ~new_n12553_;
  assign po0805 = ~new_n10896_ | ~new_n12549_ | ~new_n12548_;
  assign po0804 = ~new_n10895_ | ~new_n12544_ | ~new_n12543_;
  assign po0803 = ~new_n10894_ | ~new_n12539_ | ~new_n12538_;
  assign po0802 = ~new_n10893_ | ~new_n12534_ | ~new_n12533_;
  assign po0801 = ~new_n10892_ | ~new_n12529_ | ~new_n12528_;
  assign po0800 = ~new_n10891_ | ~new_n12524_ | ~new_n12523_;
  assign po0799 = ~new_n10890_ | ~new_n12519_ | ~new_n12518_;
  assign po0798 = ~new_n10888_ | ~new_n12496_ | ~new_n12495_;
  assign po0797 = ~new_n10887_ | ~new_n12491_ | ~new_n12490_;
  assign po0796 = ~new_n10886_ | ~new_n12486_ | ~new_n12485_;
  assign po0795 = ~new_n10885_ | ~new_n12481_ | ~new_n12480_;
  assign po0794 = ~new_n10884_ | ~new_n12476_ | ~new_n12475_;
  assign po0793 = ~new_n10883_ | ~new_n12471_ | ~new_n12470_;
  assign po0792 = ~new_n10882_ | ~new_n12466_ | ~new_n12465_;
  assign po0791 = ~new_n10881_ | ~new_n12461_ | ~new_n12460_;
  assign po0790 = ~new_n10879_ | ~new_n12439_ | ~new_n12438_;
  assign po0789 = ~new_n10878_ | ~new_n12434_ | ~new_n12433_;
  assign po0788 = ~new_n10877_ | ~new_n12429_ | ~new_n12428_;
  assign po0787 = ~new_n10876_ | ~new_n12424_ | ~new_n12423_;
  assign po0786 = ~new_n10875_ | ~new_n12419_ | ~new_n12418_;
  assign po0785 = ~new_n10874_ | ~new_n12414_ | ~new_n12413_;
  assign po0784 = ~new_n10873_ | ~new_n12409_ | ~new_n12408_;
  assign po0783 = ~new_n10872_ | ~new_n12404_ | ~new_n12403_;
  assign po0782 = ~new_n10870_ | ~new_n12381_ | ~new_n12380_;
  assign po0781 = ~new_n10869_ | ~new_n12376_ | ~new_n12375_;
  assign po0780 = ~new_n10868_ | ~new_n12371_ | ~new_n12370_;
  assign po0779 = ~new_n10867_ | ~new_n12366_ | ~new_n12365_;
  assign po0778 = ~new_n10866_ | ~new_n12361_ | ~new_n12360_;
  assign po0777 = ~new_n10865_ | ~new_n12356_ | ~new_n12355_;
  assign po0776 = ~new_n10864_ | ~new_n12351_ | ~new_n12350_;
  assign po0775 = ~new_n10863_ | ~new_n12346_ | ~new_n12345_;
  assign po0774 = ~new_n10861_ | ~new_n12324_ | ~new_n12323_;
  assign po0773 = ~new_n10860_ | ~new_n12319_ | ~new_n12318_;
  assign po0772 = ~new_n10859_ | ~new_n12314_ | ~new_n12313_;
  assign po0771 = ~new_n10858_ | ~new_n12309_ | ~new_n12308_;
  assign po0770 = ~new_n10857_ | ~new_n12304_ | ~new_n12303_;
  assign po0769 = ~new_n10856_ | ~new_n12299_ | ~new_n12298_;
  assign po0768 = ~new_n10855_ | ~new_n12294_ | ~new_n12293_;
  assign po0767 = ~new_n10854_ | ~new_n12289_ | ~new_n12288_;
  assign po0766 = ~new_n10852_ | ~new_n12266_ | ~new_n12265_;
  assign po0765 = ~new_n10851_ | ~new_n12261_ | ~new_n12260_;
  assign po0764 = ~new_n10850_ | ~new_n12256_ | ~new_n12255_;
  assign po0763 = ~new_n10849_ | ~new_n12251_ | ~new_n12250_;
  assign po0762 = ~new_n10848_ | ~new_n12246_ | ~new_n12245_;
  assign po0761 = ~new_n10847_ | ~new_n12241_ | ~new_n12240_;
  assign po0760 = ~new_n10846_ | ~new_n12236_ | ~new_n12235_;
  assign po0759 = ~new_n10845_ | ~new_n12231_ | ~new_n12230_;
  assign po0758 = ~new_n10843_ | ~new_n12209_ | ~new_n12208_;
  assign po0757 = ~new_n10842_ | ~new_n12204_ | ~new_n12203_;
  assign po0756 = ~new_n10841_ | ~new_n12199_ | ~new_n12198_;
  assign po0755 = ~new_n10840_ | ~new_n12194_ | ~new_n12193_;
  assign po0754 = ~new_n10839_ | ~new_n12189_ | ~new_n12188_;
  assign po0753 = ~new_n10838_ | ~new_n12184_ | ~new_n12183_;
  assign po0752 = ~new_n10837_ | ~new_n12179_ | ~new_n12178_;
  assign po0751 = ~new_n10836_ | ~new_n12174_ | ~new_n12173_;
  assign po0750 = ~new_n10834_ | ~new_n12153_ | ~new_n12152_;
  assign po0749 = ~new_n10833_ | ~new_n12148_ | ~new_n12147_;
  assign po0748 = ~new_n10832_ | ~new_n12143_ | ~new_n12142_;
  assign po0747 = ~new_n10831_ | ~new_n12138_ | ~new_n12137_;
  assign po0746 = ~new_n10830_ | ~new_n12133_ | ~new_n12132_;
  assign po0745 = ~new_n10829_ | ~new_n12128_ | ~new_n12127_;
  assign po0744 = ~new_n10828_ | ~new_n12123_ | ~new_n12122_;
  assign po0743 = ~new_n10827_ | ~new_n12118_ | ~new_n12117_;
  assign po0742 = ~new_n10825_ | ~new_n12096_ | ~new_n12095_;
  assign po0741 = ~new_n10824_ | ~new_n12091_ | ~new_n12090_;
  assign po0740 = ~new_n10823_ | ~new_n12086_ | ~new_n12085_;
  assign po0739 = ~new_n10822_ | ~new_n12081_ | ~new_n12080_;
  assign po0738 = ~new_n10821_ | ~new_n12076_ | ~new_n12075_;
  assign po0737 = ~new_n10820_ | ~new_n12071_ | ~new_n12070_;
  assign po0736 = ~new_n10819_ | ~new_n12066_ | ~new_n12065_;
  assign po0735 = ~new_n10818_ | ~new_n12061_ | ~new_n12060_;
  assign po0734 = ~new_n10816_ | ~new_n12038_ | ~new_n12037_;
  assign po0733 = ~new_n10815_ | ~new_n12033_ | ~new_n12032_;
  assign po0732 = ~new_n10814_ | ~new_n12028_ | ~new_n12027_;
  assign po0731 = ~new_n10813_ | ~new_n12023_ | ~new_n12022_;
  assign po0730 = ~new_n10812_ | ~new_n12018_ | ~new_n12017_;
  assign po0729 = ~new_n10811_ | ~new_n12013_ | ~new_n12012_;
  assign po0728 = ~new_n10810_ | ~new_n12008_ | ~new_n12007_;
  assign po0727 = ~new_n10809_ | ~new_n12003_ | ~new_n12002_;
  assign po0726 = ~new_n10807_ | ~new_n11981_ | ~new_n11980_;
  assign po0725 = ~new_n10806_ | ~new_n11976_ | ~new_n11975_;
  assign po0724 = ~new_n10805_ | ~new_n11971_ | ~new_n11970_;
  assign po0723 = ~new_n10804_ | ~new_n11966_ | ~new_n11965_;
  assign po0722 = ~new_n10803_ | ~new_n11961_ | ~new_n11960_;
  assign po0721 = ~new_n10802_ | ~new_n11956_ | ~new_n11955_;
  assign po0720 = ~new_n10801_ | ~new_n11951_ | ~new_n11950_;
  assign po0719 = ~new_n10800_ | ~new_n11946_ | ~new_n11945_;
  assign po0718 = ~new_n10798_ | ~new_n11923_ | ~new_n11922_;
  assign po0717 = ~new_n10797_ | ~new_n11918_ | ~new_n11917_;
  assign po0716 = ~new_n10796_ | ~new_n11913_ | ~new_n11912_;
  assign po0715 = ~new_n10795_ | ~new_n11908_ | ~new_n11907_;
  assign po0714 = ~new_n10794_ | ~new_n11903_ | ~new_n11902_;
  assign po0713 = ~new_n10793_ | ~new_n11898_ | ~new_n11897_;
  assign po0712 = ~new_n10792_ | ~new_n11893_ | ~new_n11892_;
  assign po0711 = ~new_n10791_ | ~new_n11888_ | ~new_n11887_;
  assign po0710 = ~new_n10789_ | ~new_n11866_ | ~new_n11865_;
  assign po0709 = ~new_n10788_ | ~new_n11861_ | ~new_n11860_;
  assign po0708 = ~new_n10787_ | ~new_n11856_ | ~new_n11855_;
  assign po0707 = ~new_n10786_ | ~new_n11851_ | ~new_n11850_;
  assign po0706 = ~new_n10785_ | ~new_n11846_ | ~new_n11845_;
  assign po0705 = ~new_n10784_ | ~new_n11841_ | ~new_n11840_;
  assign po0704 = ~new_n10783_ | ~new_n11836_ | ~new_n11835_;
  assign po0703 = ~new_n10782_ | ~new_n11831_ | ~new_n11830_;
  assign po0702 = ~new_n10780_ | ~new_n11807_ | ~new_n11806_;
  assign po0701 = ~new_n10779_ | ~new_n11802_ | ~new_n11801_;
  assign po0700 = ~new_n10778_ | ~new_n11797_ | ~new_n11796_;
  assign po0699 = ~new_n10777_ | ~new_n11792_ | ~new_n11791_;
  assign po0698 = ~new_n10776_ | ~new_n11787_ | ~new_n11786_;
  assign po0697 = ~new_n10775_ | ~new_n11782_ | ~new_n11781_;
  assign po0696 = ~new_n10774_ | ~new_n11777_ | ~new_n11776_;
  assign po0695 = ~new_n10773_ | ~new_n11772_ | ~new_n11771_;
  assign po0694 = ~new_n10771_ | ~new_n11749_ | ~new_n11748_;
  assign po0693 = ~new_n10770_ | ~new_n11744_ | ~new_n11743_;
  assign po0692 = ~new_n10769_ | ~new_n11739_ | ~new_n11738_;
  assign po0691 = ~new_n10768_ | ~new_n11734_ | ~new_n11733_;
  assign po0690 = ~new_n10767_ | ~new_n11729_ | ~new_n11728_;
  assign po0689 = ~new_n10766_ | ~new_n11724_ | ~new_n11723_;
  assign po0688 = ~new_n10765_ | ~new_n11719_ | ~new_n11718_;
  assign po0687 = ~new_n10764_ | ~new_n11714_ | ~new_n11713_;
  assign po0686 = ~new_n10762_ | ~new_n15102_ | ~new_n15101_;
  assign po0685 = ~new_n11669_ | ~new_n11495_ | ~new_n11668_ | ~new_n11670_;
  assign po0684 = ~new_n10757_ | ~new_n11666_;
  assign po0682 = pi0623 & new_n14958_;
  assign po0681 = pi0622 & new_n14958_;
  assign po0680 = pi0621 & new_n14958_;
  assign po0679 = pi0620 & new_n14958_;
  assign po0678 = pi0619 & new_n14958_;
  assign po0677 = pi0618 & new_n14958_;
  assign po0676 = pi0617 & new_n14958_;
  assign po0675 = pi0616 & new_n14958_;
  assign po0674 = pi0615 & new_n14958_;
  assign po0673 = pi0614 & new_n14958_;
  assign po0672 = pi0613 & new_n14958_;
  assign po0671 = pi0612 & new_n14958_;
  assign po0670 = pi0611 & new_n14958_;
  assign po0669 = pi0610 & new_n14958_;
  assign po0668 = pi0609 & new_n14958_;
  assign po0667 = pi0608 & new_n14958_;
  assign po0666 = pi0607 & new_n14958_;
  assign po0665 = pi0606 & new_n14958_;
  assign po0664 = pi0605 & new_n14958_;
  assign po0663 = pi0604 & new_n14958_;
  assign po0662 = pi0603 & new_n14958_;
  assign po0661 = pi0602 & new_n14958_;
  assign po0660 = pi0601 & new_n14958_;
  assign po0659 = pi0600 & new_n14958_;
  assign po0658 = pi0599 & new_n14958_;
  assign po0657 = pi0598 & new_n14958_;
  assign po0656 = pi0597 & new_n14958_;
  assign po0655 = pi0596 & new_n14958_;
  assign po0654 = pi0595 & new_n14958_;
  assign po0653 = pi0594 & new_n14958_;
  assign po0650 = ~new_n11629_ | ~new_n14955_ | ~new_n14954_;
  assign po0649 = ~new_n10732_ | ~new_n14953_ | ~new_n14952_;
  assign po0648 = ~new_n10731_ | ~new_n11620_;
  assign po0647 = ~new_n11608_ | ~new_n11607_ | ~new_n11606_;
  assign po0646 = ~new_n11605_ | ~new_n11604_ | ~new_n11603_;
  assign po0645 = ~new_n11602_ | ~new_n11601_ | ~new_n11600_;
  assign po0644 = ~new_n11599_ | ~new_n11598_ | ~new_n11597_;
  assign po0643 = ~new_n11596_ | ~new_n11595_ | ~new_n11594_;
  assign po0642 = ~new_n11593_ | ~new_n11592_ | ~new_n11591_;
  assign po0641 = ~new_n11590_ | ~new_n11589_ | ~new_n11588_;
  assign po0640 = ~new_n11587_ | ~new_n11586_ | ~new_n11585_;
  assign po0639 = ~new_n11584_ | ~new_n11583_ | ~new_n11582_;
  assign po0638 = ~new_n11581_ | ~new_n11580_ | ~new_n11579_;
  assign po0637 = ~new_n11578_ | ~new_n11577_ | ~new_n11576_;
  assign po0636 = ~new_n11575_ | ~new_n11574_ | ~new_n11573_;
  assign po0635 = ~new_n11572_ | ~new_n11571_ | ~new_n11570_;
  assign po0634 = ~new_n11569_ | ~new_n11568_ | ~new_n11567_;
  assign po0633 = ~new_n11566_ | ~new_n11565_ | ~new_n11564_;
  assign po0632 = ~new_n11563_ | ~new_n11562_ | ~new_n11561_;
  assign po0631 = ~new_n11560_ | ~new_n11559_ | ~new_n11558_;
  assign po0630 = ~new_n11557_ | ~new_n11556_ | ~new_n11555_;
  assign po0629 = ~new_n11554_ | ~new_n11553_ | ~new_n11552_;
  assign po0628 = ~new_n11551_ | ~new_n11550_ | ~new_n11549_;
  assign po0627 = ~new_n11548_ | ~new_n11547_ | ~new_n11546_;
  assign po0626 = ~new_n11545_ | ~new_n11544_ | ~new_n11543_;
  assign po0625 = ~new_n11542_ | ~new_n11541_ | ~new_n11540_;
  assign po0624 = ~new_n11539_ | ~new_n11538_ | ~new_n11537_;
  assign po0623 = ~new_n11536_ | ~new_n11535_ | ~new_n11534_;
  assign po0622 = ~new_n11533_ | ~new_n11532_ | ~new_n11531_;
  assign po0621 = ~new_n11530_ | ~new_n11529_ | ~new_n11528_;
  assign po0620 = ~new_n11527_ | ~new_n11526_ | ~new_n11525_;
  assign po0619 = ~new_n11524_ | ~new_n11523_ | ~new_n11522_;
  assign po0618 = ~new_n11521_ | ~new_n11520_ | ~new_n11519_;
  assign new_n10283_ = ~new_n11234_ | ~new_n11232_ | ~new_n11233_ | ~new_n11235_;
  assign new_n10284_ = ~new_n10390_ | ~new_n10376_;
  assign new_n10285_ = ~pi0589;
  assign new_n10286_ = ~new_n9481_ | ~new_n10284_;
  assign new_n10287_ = ~new_n9481_ | ~new_n11691_;
  assign new_n10288_ = ~new_n9483_ | ~new_n10284_;
  assign new_n10289_ = ~new_n9483_ | ~new_n11691_;
  assign new_n10290_ = ~new_n9482_ | ~new_n10284_;
  assign new_n10291_ = ~new_n9482_ | ~new_n11691_;
  assign new_n10292_ = ~new_n9484_ | ~new_n10284_;
  assign new_n10293_ = ~new_n9484_ | ~new_n11691_;
  assign new_n10294_ = ~new_n10749_ | ~new_n10748_;
  assign new_n10295_ = ~new_n9631_ | ~new_n11470_;
  assign new_n10296_ = ~new_n10737_ | ~new_n10736_;
  assign new_n10297_ = ~pi0997;
  assign new_n10298_ = ~new_n15091_ | ~new_n11649_ | ~new_n11650_ | ~new_n15092_;
  assign new_n10299_ = ~pi0590;
  assign new_n10300_ = ~pi0590 | ~new_n10307_;
  assign new_n10301_ = ~new_n11480_ | ~new_n10285_;
  assign new_n10302_ = ~new_n11480_ | ~pi0589;
  assign new_n10303_ = ~pi0590 | ~new_n10285_;
  assign new_n10304_ = pi0589 | pi0590;
  assign new_n10305_ = ~pi0033;
  assign new_n10306_ = ~new_n2973_;
  assign new_n10307_ = ~pi0591;
  assign new_n10308_ = ~pi0997 | ~new_n10305_;
  assign new_n10309_ = pi0033 | pi0997;
  assign new_n10310_ = ~pi0626;
  assign new_n10311_ = ~pi0625;
  assign new_n10312_ = ~pi0759;
  assign new_n10313_ = ~pi0760;
  assign new_n10314_ = ~pi0757;
  assign new_n10315_ = ~pi0760 | ~pi0759 | ~new_n10317_;
  assign new_n10316_ = pi0759 | pi0758 | pi0760;
  assign new_n10317_ = ~pi0758;
  assign new_n10318_ = ~pi0758 | ~pi0760 | ~pi0759;
  assign new_n10319_ = ~new_n10741_ | ~new_n10740_;
  assign new_n10320_ = ~new_n10743_ | ~new_n10742_;
  assign new_n10321_ = ~new_n10745_ | ~new_n10744_;
  assign new_n10322_ = ~new_n14900_ | ~new_n14902_ | ~new_n14904_;
  assign new_n10323_ = ~new_n11517_ | ~new_n9498_ | ~new_n14910_;
  assign new_n10324_ = ~new_n10294_ | ~new_n14914_;
  assign new_n10325_ = ~pi0627;
  assign new_n10326_ = ~new_n11465_ | ~new_n10750_;
  assign new_n10327_ = ~new_n10294_ | ~new_n9657_;
  assign new_n10328_ = ~new_n29402_;
  assign new_n10329_ = ~new_n9499_ | ~new_n9498_ | ~new_n14900_;
  assign new_n10330_ = ~new_n9657_ | ~new_n14912_;
  assign new_n10331_ = ~new_n11636_ | ~new_n10307_;
  assign new_n10332_ = ~new_n10754_ | ~new_n9500_;
  assign new_n10333_ = ~new_n29132_;
  assign new_n10334_ = ~new_n9398_ | ~new_n10321_;
  assign new_n10335_ = ~new_n14912_ | ~new_n14914_;
  assign new_n10336_ = ~new_n14902_ | ~new_n9658_;
  assign new_n10337_ = ~new_n9492_ | ~new_n11469_;
  assign new_n10338_ = ~new_n28599_;
  assign new_n10339_ = ~new_n14935_ | ~new_n11651_ | ~new_n11655_ | ~new_n29406_ | ~new_n11485_;
  assign new_n10340_ = ~pi0627 | ~new_n11660_;
  assign new_n10341_ = ~pi0624;
  assign new_n10342_ = ~pi0627 | ~new_n10311_;
  assign new_n10343_ = ~pi0996;
  assign new_n10344_ = pi0624 | pi0626;
  assign new_n10345_ = ~pi0625 | ~new_n10310_;
  assign new_n10346_ = ~pi0624 | ~new_n28599_;
  assign new_n10347_ = ~new_n11697_ | ~new_n10325_;
  assign new_n10348_ = ~pi0765;
  assign new_n10349_ = ~pi0764;
  assign new_n10350_ = ~pi0762;
  assign new_n10351_ = ~pi0763;
  assign new_n10352_ = ~pi0764 | ~pi0765;
  assign new_n10353_ = ~new_n11683_ | ~new_n9505_;
  assign new_n10354_ = pi0624 | pi0625;
  assign new_n10355_ = ~new_n28362_;
  assign new_n10356_ = ~new_n28361_;
  assign new_n10357_ = ~new_n28333_;
  assign new_n10358_ = ~new_n28369_;
  assign new_n10359_ = ~new_n28361_ | ~new_n28362_;
  assign new_n10360_ = ~new_n10393_ | ~new_n10355_;
  assign new_n10361_ = ~new_n11677_ | ~new_n9502_;
  assign new_n10362_ = ~new_n27643_;
  assign new_n10363_ = ~new_n27644_;
  assign new_n10364_ = ~new_n27642_;
  assign new_n10365_ = ~new_n27553_;
  assign new_n10366_ = ~new_n10353_ | ~new_n11692_;
  assign new_n10367_ = ~new_n10611_ | ~new_n10353_;
  assign new_n10368_ = ~pi0628;
  assign new_n10369_ = ~pi0629;
  assign new_n10370_ = ~pi0630;
  assign new_n10371_ = ~pi0631;
  assign new_n10372_ = ~pi0632;
  assign new_n10373_ = ~pi0633;
  assign new_n10374_ = ~pi0634;
  assign new_n10375_ = ~pi0635;
  assign new_n10376_ = ~pi0764 | ~new_n10348_;
  assign new_n10377_ = ~new_n11690_ | ~new_n9505_;
  assign new_n10378_ = ~new_n28361_ | ~new_n10355_;
  assign new_n10379_ = ~new_n28362_ | ~new_n10393_;
  assign new_n10380_ = ~new_n11750_ | ~new_n9502_;
  assign new_n10381_ = ~new_n10610_ | ~new_n10377_;
  assign new_n10382_ = ~pi0636;
  assign new_n10383_ = ~pi0637;
  assign new_n10384_ = ~pi0638;
  assign new_n10385_ = ~pi0639;
  assign new_n10386_ = ~pi0640;
  assign new_n10387_ = ~pi0641;
  assign new_n10388_ = ~pi0642;
  assign new_n10389_ = ~pi0643;
  assign new_n10390_ = ~pi0765 | ~new_n10349_;
  assign new_n10391_ = ~new_n11689_ | ~new_n9505_;
  assign new_n10392_ = ~new_n28362_ | ~new_n10356_;
  assign new_n10393_ = ~new_n10378_ | ~new_n10392_;
  assign new_n10394_ = ~new_n11676_ | ~new_n10355_;
  assign new_n10395_ = ~new_n11808_ | ~new_n9502_;
  assign new_n10396_ = ~new_n10391_ | ~new_n11811_;
  assign new_n10397_ = ~new_n10609_ | ~new_n10391_;
  assign new_n10398_ = ~pi0644;
  assign new_n10399_ = ~pi0645;
  assign new_n10400_ = ~pi0646;
  assign new_n10401_ = ~pi0647;
  assign new_n10402_ = ~pi0648;
  assign new_n10403_ = ~pi0649;
  assign new_n10404_ = ~pi0650;
  assign new_n10405_ = ~pi0651;
  assign new_n10406_ = ~new_n9519_ | ~new_n9505_;
  assign new_n10407_ = ~new_n9516_ | ~new_n9502_;
  assign new_n10408_ = ~new_n10608_ | ~new_n10406_;
  assign new_n10409_ = ~pi0652;
  assign new_n10410_ = ~pi0653;
  assign new_n10411_ = ~pi0654;
  assign new_n10412_ = ~pi0655;
  assign new_n10413_ = ~pi0656;
  assign new_n10414_ = ~pi0657;
  assign new_n10415_ = ~pi0658;
  assign new_n10416_ = ~pi0659;
  assign new_n10417_ = ~pi0762 | ~new_n10351_;
  assign new_n10418_ = ~new_n11686_ | ~new_n11683_;
  assign new_n10419_ = ~new_n28369_ | ~new_n10357_;
  assign new_n10420_ = ~new_n9522_ | ~new_n11677_;
  assign new_n10421_ = ~new_n10418_ | ~new_n11926_;
  assign new_n10422_ = ~new_n10607_ | ~new_n10418_;
  assign new_n10423_ = ~pi0660;
  assign new_n10424_ = ~pi0661;
  assign new_n10425_ = ~pi0662;
  assign new_n10426_ = ~pi0663;
  assign new_n10427_ = ~pi0664;
  assign new_n10428_ = ~pi0665;
  assign new_n10429_ = ~pi0666;
  assign new_n10430_ = ~pi0667;
  assign new_n10431_ = ~new_n11686_ | ~new_n11690_;
  assign new_n10432_ = ~new_n9522_ | ~new_n11750_;
  assign new_n10433_ = ~new_n10606_ | ~new_n10431_;
  assign new_n10434_ = ~pi0668;
  assign new_n10435_ = ~pi0669;
  assign new_n10436_ = ~pi0670;
  assign new_n10437_ = ~pi0671;
  assign new_n10438_ = ~pi0672;
  assign new_n10439_ = ~pi0673;
  assign new_n10440_ = ~pi0674;
  assign new_n10441_ = ~pi0675;
  assign new_n10442_ = ~new_n11686_ | ~new_n11689_;
  assign new_n10443_ = ~new_n9522_ | ~new_n11808_;
  assign new_n10444_ = ~new_n10442_ | ~new_n12041_;
  assign new_n10445_ = ~new_n10605_ | ~new_n10442_;
  assign new_n10446_ = ~pi0676;
  assign new_n10447_ = ~pi0677;
  assign new_n10448_ = ~pi0678;
  assign new_n10449_ = ~pi0679;
  assign new_n10450_ = ~pi0680;
  assign new_n10451_ = ~pi0681;
  assign new_n10452_ = ~pi0682;
  assign new_n10453_ = ~pi0683;
  assign new_n10454_ = ~new_n11686_ | ~new_n9519_;
  assign new_n10455_ = ~new_n9522_ | ~new_n9516_;
  assign new_n10456_ = ~new_n10604_ | ~new_n10454_;
  assign new_n10457_ = ~pi0684;
  assign new_n10458_ = ~pi0685;
  assign new_n10459_ = ~pi0686;
  assign new_n10460_ = ~pi0687;
  assign new_n10461_ = ~pi0688;
  assign new_n10462_ = ~pi0689;
  assign new_n10463_ = ~pi0690;
  assign new_n10464_ = ~pi0691;
  assign new_n10465_ = ~new_n9506_ | ~new_n11683_;
  assign new_n10466_ = ~new_n9501_ | ~new_n11678_;
  assign new_n10467_ = ~new_n10466_ | ~new_n10419_ | ~new_n11680_;
  assign new_n10468_ = ~new_n9532_ | ~new_n11677_;
  assign new_n10469_ = ~new_n10465_ | ~new_n10417_ | ~new_n11687_;
  assign new_n10470_ = ~new_n10465_ | ~new_n12155_;
  assign new_n10471_ = ~new_n10603_ | ~new_n10465_;
  assign new_n10472_ = ~pi0692;
  assign new_n10473_ = ~pi0693;
  assign new_n10474_ = ~pi0694;
  assign new_n10475_ = ~pi0695;
  assign new_n10476_ = ~pi0696;
  assign new_n10477_ = ~pi0697;
  assign new_n10478_ = ~pi0698;
  assign new_n10479_ = ~pi0699;
  assign new_n10480_ = ~new_n11690_ | ~new_n9506_;
  assign new_n10481_ = ~new_n9532_ | ~new_n11750_;
  assign new_n10482_ = ~new_n10602_ | ~new_n10480_;
  assign new_n10483_ = ~pi0700;
  assign new_n10484_ = ~pi0701;
  assign new_n10485_ = ~pi0702;
  assign new_n10486_ = ~pi0703;
  assign new_n10487_ = ~pi0704;
  assign new_n10488_ = ~pi0705;
  assign new_n10489_ = ~pi0706;
  assign new_n10490_ = ~pi0707;
  assign new_n10491_ = ~new_n11689_ | ~new_n9506_;
  assign new_n10492_ = ~new_n9532_ | ~new_n11808_;
  assign new_n10493_ = ~new_n10491_ | ~new_n12269_;
  assign new_n10494_ = ~new_n10601_ | ~new_n10491_;
  assign new_n10495_ = ~pi0708;
  assign new_n10496_ = ~pi0709;
  assign new_n10497_ = ~pi0710;
  assign new_n10498_ = ~pi0711;
  assign new_n10499_ = ~pi0712;
  assign new_n10500_ = ~pi0713;
  assign new_n10501_ = ~pi0714;
  assign new_n10502_ = ~pi0715;
  assign new_n10503_ = ~new_n9519_ | ~new_n9506_;
  assign new_n10504_ = ~new_n9532_ | ~new_n9516_;
  assign new_n10505_ = ~new_n10600_ | ~new_n10503_;
  assign new_n10506_ = ~pi0716;
  assign new_n10507_ = ~pi0717;
  assign new_n10508_ = ~pi0718;
  assign new_n10509_ = ~pi0719;
  assign new_n10510_ = ~pi0720;
  assign new_n10511_ = ~pi0721;
  assign new_n10512_ = ~pi0722;
  assign new_n10513_ = ~pi0723;
  assign new_n10514_ = ~new_n9544_ | ~new_n11683_;
  assign new_n10515_ = ~new_n9541_ | ~new_n11677_;
  assign new_n10516_ = ~new_n10514_ | ~new_n12384_;
  assign new_n10517_ = ~new_n10599_ | ~new_n10514_;
  assign new_n10518_ = ~pi0724;
  assign new_n10519_ = ~pi0725;
  assign new_n10520_ = ~pi0726;
  assign new_n10521_ = ~pi0727;
  assign new_n10522_ = ~pi0728;
  assign new_n10523_ = ~pi0729;
  assign new_n10524_ = ~pi0730;
  assign new_n10525_ = ~pi0731;
  assign new_n10526_ = ~new_n9544_ | ~new_n11690_;
  assign new_n10527_ = ~new_n9541_ | ~new_n11750_;
  assign new_n10528_ = ~new_n10598_ | ~new_n10526_;
  assign new_n10529_ = ~pi0732;
  assign new_n10530_ = ~pi0733;
  assign new_n10531_ = ~pi0734;
  assign new_n10532_ = ~pi0735;
  assign new_n10533_ = ~pi0736;
  assign new_n10534_ = ~pi0737;
  assign new_n10535_ = ~pi0738;
  assign new_n10536_ = ~pi0739;
  assign new_n10537_ = ~new_n9544_ | ~new_n11689_;
  assign new_n10538_ = ~new_n9541_ | ~new_n11808_;
  assign new_n10539_ = ~new_n10537_ | ~new_n12499_;
  assign new_n10540_ = ~new_n10597_ | ~new_n10537_;
  assign new_n10541_ = ~pi0740;
  assign new_n10542_ = ~pi0741;
  assign new_n10543_ = ~pi0742;
  assign new_n10544_ = ~pi0743;
  assign new_n10545_ = ~pi0744;
  assign new_n10546_ = ~pi0745;
  assign new_n10547_ = ~pi0746;
  assign new_n10548_ = ~pi0747;
  assign new_n10549_ = ~new_n9544_ | ~new_n9519_;
  assign new_n10550_ = ~new_n9541_ | ~new_n9516_;
  assign new_n10551_ = ~new_n10596_ | ~new_n10549_;
  assign new_n10552_ = ~pi0748;
  assign new_n10553_ = ~pi0749;
  assign new_n10554_ = ~pi0750;
  assign new_n10555_ = ~pi0751;
  assign new_n10556_ = ~pi0752;
  assign new_n10557_ = ~pi0753;
  assign new_n10558_ = ~pi0754;
  assign new_n10559_ = ~pi0755;
  assign new_n10560_ = ~pi0994;
  assign new_n10561_ = ~new_n30327_;
  assign new_n10562_ = ~new_n10739_ | ~new_n10738_;
  assign new_n10563_ = ~new_n9492_ | ~new_n11470_;
  assign new_n10564_ = ~new_n11516_ | ~new_n11468_;
  assign new_n10565_ = ~new_n11470_ | ~new_n11516_;
  assign new_n10566_ = ~new_n14904_ | ~new_n14910_ | ~new_n10320_ | ~new_n14906_;
  assign new_n10567_ = ~new_n29006_;
  assign new_n10568_ = ~new_n10324_ | ~new_n10330_;
  assign new_n10569_ = ~new_n10688_;
  assign new_n10570_ = ~new_n29007_;
  assign new_n10571_ = ~new_n10315_ | ~new_n12656_;
  assign new_n10572_ = ~new_n29002_;
  assign new_n10573_ = ~pi0760;
  assign new_n10574_ = ~new_n12683_ | ~new_n11496_ | ~new_n10347_;
  assign new_n10575_ = ~new_n11471_ | ~new_n10310_;
  assign new_n10576_ = ~new_n12713_ | ~new_n12712_;
  assign new_n10577_ = ~pi0627 | ~new_n14914_;
  assign new_n10578_ = ~new_n12978_ | ~new_n12977_;
  assign new_n10579_ = ~new_n11096_ | ~new_n9487_;
  assign new_n10580_ = ~new_n11097_ | ~new_n9398_;
  assign new_n10581_ = ~pi0625 | ~new_n10325_;
  assign new_n10582_ = ~new_n13272_ | ~new_n13271_;
  assign new_n10583_ = ~new_n9415_ | ~new_n13367_;
  assign new_n10584_ = ~new_n9415_ | ~new_n13511_;
  assign new_n10585_ = ~pi0956;
  assign new_n10586_ = pi0996 | new_n2973_;
  assign new_n10587_ = ~new_n11110_ | ~new_n11503_;
  assign new_n10588_ = ~new_n11218_ | ~new_n11212_ | ~new_n11215_ | ~new_n11222_;
  assign new_n10589_ = ~new_n11479_ | ~pi0958;
  assign new_n10590_ = ~new_n9397_ | ~new_n11461_;
  assign new_n10591_ = ~new_n11468_ | ~pi0627;
  assign new_n10592_ = ~pi1000;
  assign new_n10593_ = ~pi1002;
  assign new_n10594_ = ~new_n11446_ | ~new_n10316_;
  assign new_n10595_ = ~new_n11456_ | ~new_n10617_;
  assign new_n10596_ = ~new_n9545_ | ~new_n9520_;
  assign new_n10597_ = ~new_n9545_ | ~new_n9514_;
  assign new_n10598_ = ~new_n9545_ | ~new_n9511_;
  assign new_n10599_ = ~new_n9545_ | ~new_n9508_;
  assign new_n10600_ = ~new_n9533_ | ~new_n9520_;
  assign new_n10601_ = ~new_n9533_ | ~new_n9514_;
  assign new_n10602_ = ~new_n9533_ | ~new_n9511_;
  assign new_n10603_ = ~new_n9533_ | ~new_n9508_;
  assign new_n10604_ = ~new_n9524_ | ~new_n9520_;
  assign new_n10605_ = ~new_n9524_ | ~new_n9514_;
  assign new_n10606_ = ~new_n9524_ | ~new_n9511_;
  assign new_n10607_ = ~new_n9524_ | ~new_n9508_;
  assign new_n10608_ = ~new_n9520_ | ~new_n9507_;
  assign new_n10609_ = ~new_n9514_ | ~new_n9507_;
  assign new_n10610_ = ~new_n9511_ | ~new_n9507_;
  assign new_n10611_ = ~new_n9507_ | ~new_n9508_;
  assign new_n10612_ = ~new_n14906_ | ~new_n10341_;
  assign new_n10613_ = ~new_n10283_;
  assign new_n10614_ = pi0627 | pi0626;
  assign new_n10615_ = ~new_n10562_ | ~new_n12612_ | ~new_n10336_;
  assign new_n10616_ = ~new_n11460_ | ~new_n14912_;
  assign new_n10617_ = ~new_n11460_ | ~new_n10320_;
  assign new_n10618_ = ~new_n11465_ | ~new_n13886_;
  assign new_n10619_ = ~new_n9631_ | ~new_n11469_;
  assign new_n10620_ = ~new_n15104_ | ~new_n15103_;
  assign new_n10621_ = ~new_n15107_ | ~new_n15106_;
  assign new_n10622_ = ~new_n15122_ | ~new_n15121_;
  assign new_n10623_ = ~new_n15140_ | ~new_n15139_;
  assign new_n10624_ = ~new_n15189_ | ~new_n15188_;
  assign new_n10625_ = ~new_n15192_ | ~new_n15191_;
  assign po0614 = ~new_n14941_ | ~new_n14940_;
  assign po0615 = ~new_n14943_ | ~new_n14942_;
  assign po0616 = ~new_n14945_ | ~new_n14944_;
  assign po0617 = ~new_n14947_ | ~new_n14946_;
  assign new_n10630_ = ~new_n14957_ | ~new_n14956_;
  assign new_n10631_ = new_n10304_ & new_n11442_;
  assign po0651 = ~new_n14960_ | ~new_n14959_;
  assign po0652 = ~new_n14962_ | ~new_n14961_;
  assign po0683 = ~new_n15100_ | ~new_n15099_;
  assign new_n10635_ = new_n10907_ & new_n11475_;
  assign po0815 = ~new_n15114_ | ~new_n15113_;
  assign po0816 = ~new_n15125_ | ~new_n15124_;
  assign new_n10638_ = ~new_n15127_ | ~new_n15126_;
  assign new_n10639_ = ~new_n15130_ | ~new_n15129_;
  assign po0817 = ~new_n15135_ | ~new_n15134_;
  assign po0818 = ~new_n15143_ | ~new_n15142_;
  assign po0819 = ~new_n15145_ | ~new_n15144_;
  assign po0821 = ~new_n15147_ | ~new_n15146_;
  assign po0822 = ~new_n15152_ | ~new_n15151_;
  assign po0823 = ~new_n15154_ | ~new_n15153_;
  assign po0824 = ~new_n15156_ | ~new_n15155_;
  assign new_n10647_ = ~pi0958 & ~pi0593;
  assign new_n10648_ = new_n11224_ & new_n14939_;
  assign po1052 = ~new_n15171_ | ~new_n15170_;
  assign po1054 = ~new_n15175_ | ~new_n15174_;
  assign po1056 = ~new_n15179_ | ~new_n15178_;
  assign po1058 = ~new_n15183_ | ~new_n15182_;
  assign po1061 = ~new_n15185_ | ~new_n15184_;
  assign new_n10654_ = ~new_n15323_ | ~new_n15322_;
  assign new_n10655_ = ~new_n15325_ | ~new_n15324_;
  assign new_n10656_ = ~new_n15327_ | ~new_n15326_;
  assign new_n10657_ = new_n11475_ & new_n29005_;
  assign new_n10658_ = ~new_n15329_ | ~new_n15328_;
  assign new_n10659_ = ~new_n15331_ | ~new_n15330_;
  assign new_n10660_ = ~new_n15333_ | ~new_n15332_;
  assign new_n10661_ = ~new_n15335_ | ~new_n15334_;
  assign new_n10662_ = ~new_n15337_ | ~new_n15336_;
  assign new_n10663_ = ~new_n15339_ | ~new_n15338_;
  assign new_n10664_ = ~new_n15341_ | ~new_n15340_;
  assign new_n10665_ = ~new_n15343_ | ~new_n15342_;
  assign new_n10666_ = ~new_n15345_ | ~new_n15344_;
  assign new_n10667_ = ~new_n15347_ | ~new_n15346_;
  assign new_n10668_ = ~new_n15349_ | ~new_n15348_;
  assign new_n10669_ = ~new_n15351_ | ~new_n15350_;
  assign new_n10670_ = ~new_n15353_ | ~new_n15352_;
  assign new_n10671_ = ~new_n15355_ | ~new_n15354_;
  assign new_n10672_ = ~new_n15357_ | ~new_n15356_;
  assign new_n10673_ = ~new_n15359_ | ~new_n15358_;
  assign new_n10674_ = ~new_n15361_ | ~new_n15360_;
  assign new_n10675_ = ~new_n15363_ | ~new_n15362_;
  assign new_n10676_ = ~new_n15365_ | ~new_n15364_;
  assign new_n10677_ = ~new_n15367_ | ~new_n15366_;
  assign new_n10678_ = ~new_n15369_ | ~new_n15368_;
  assign new_n10679_ = ~new_n15371_ | ~new_n15370_;
  assign new_n10680_ = ~new_n15373_ | ~new_n15372_;
  assign new_n10681_ = ~new_n15375_ | ~new_n15374_;
  assign new_n10682_ = ~new_n15377_ | ~new_n15376_;
  assign new_n10683_ = ~new_n15379_ | ~new_n15378_;
  assign new_n10684_ = ~new_n15381_ | ~new_n15380_;
  assign new_n10685_ = ~new_n15383_ | ~new_n15382_;
  assign new_n10686_ = ~new_n15385_ | ~new_n15384_;
  assign new_n10687_ = ~new_n15387_ | ~new_n15386_;
  assign new_n10688_ = ~new_n15391_ | ~new_n15390_;
  assign new_n10689_ = ~new_n15393_ | ~new_n15392_;
  assign new_n10690_ = ~new_n15395_ | ~new_n15394_;
  assign new_n10691_ = ~new_n15397_ | ~new_n15396_;
  assign new_n10692_ = ~new_n15399_ | ~new_n15398_;
  assign new_n10693_ = ~new_n15401_ | ~new_n15400_;
  assign new_n10694_ = ~new_n15403_ | ~new_n15402_;
  assign new_n10695_ = ~new_n15405_ | ~new_n15404_;
  assign new_n10696_ = ~new_n15407_ | ~new_n15406_;
  assign new_n10697_ = ~new_n15409_ | ~new_n15408_;
  assign new_n10698_ = ~new_n15411_ | ~new_n15410_;
  assign new_n10699_ = ~new_n15413_ | ~new_n15412_;
  assign new_n10700_ = ~new_n15415_ | ~new_n15414_;
  assign new_n10701_ = ~new_n15417_ | ~new_n15416_;
  assign new_n10702_ = ~new_n15419_ | ~new_n15418_;
  assign new_n10703_ = ~new_n15421_ | ~new_n15420_;
  assign new_n10704_ = ~new_n15423_ | ~new_n15422_;
  assign new_n10705_ = ~new_n15425_ | ~new_n15424_;
  assign new_n10706_ = ~new_n15427_ | ~new_n15426_;
  assign new_n10707_ = ~new_n15429_ | ~new_n15428_;
  assign new_n10708_ = ~new_n15431_ | ~new_n15430_;
  assign new_n10709_ = ~new_n15433_ | ~new_n15432_;
  assign new_n10710_ = ~new_n15435_ | ~new_n15434_;
  assign new_n10711_ = ~new_n15437_ | ~new_n15436_;
  assign new_n10712_ = ~new_n15439_ | ~new_n15438_;
  assign new_n10713_ = ~new_n15441_ | ~new_n15440_;
  assign new_n10714_ = ~new_n15443_ | ~new_n15442_;
  assign new_n10715_ = ~new_n15445_ | ~new_n15444_;
  assign new_n10716_ = ~new_n15447_ | ~new_n15446_;
  assign new_n10717_ = ~new_n15449_ | ~new_n15448_;
  assign new_n10718_ = ~new_n15451_ | ~new_n15450_;
  assign new_n10719_ = ~new_n15453_ | ~new_n15452_;
  assign new_n10720_ = ~new_n15455_ | ~new_n15454_;
  assign new_n10721_ = ~new_n15457_ | ~new_n15456_;
  assign new_n10722_ = ~new_n15459_ | ~new_n15458_;
  assign new_n10723_ = ~new_n15461_ | ~new_n15460_;
  assign new_n10724_ = ~new_n15463_ | ~new_n15462_;
  assign new_n10725_ = ~new_n15465_ | ~new_n15464_;
  assign new_n10726_ = ~new_n15467_ | ~new_n15466_;
  assign new_n10727_ = ~new_n15469_ | ~new_n15468_;
  assign new_n10728_ = ~new_n15471_ | ~new_n15470_;
  assign new_n10729_ = ~new_n15473_ | ~new_n15472_;
  assign new_n10730_ = ~new_n15475_ | ~new_n15474_;
  assign new_n10731_ = new_n11619_ & new_n10302_;
  assign new_n10732_ = new_n11624_ & new_n10301_;
  assign new_n10733_ = pi0997 & pi0591;
  assign new_n10734_ = new_n14824_ & new_n14792_ & new_n14808_ & new_n14840_;
  assign new_n10735_ = new_n14888_ & new_n14856_ & new_n14872_ & new_n14909_;
  assign new_n10736_ = new_n14823_ & new_n14791_ & new_n14807_ & new_n14839_;
  assign new_n10737_ = new_n14887_ & new_n14855_ & new_n14871_ & new_n14907_;
  assign new_n10738_ = new_n14822_ & new_n14790_ & new_n14806_ & new_n14838_;
  assign new_n10739_ = new_n14886_ & new_n14854_ & new_n14870_ & new_n14905_;
  assign new_n10740_ = new_n14821_ & new_n14789_ & new_n14805_ & new_n14837_;
  assign new_n10741_ = new_n14885_ & new_n14853_ & new_n14869_ & new_n14903_;
  assign new_n10742_ = new_n14820_ & new_n14788_ & new_n14804_ & new_n14836_;
  assign new_n10743_ = new_n14884_ & new_n14852_ & new_n14868_ & new_n14901_;
  assign new_n10744_ = new_n14819_ & new_n14787_ & new_n14803_ & new_n14835_;
  assign new_n10745_ = new_n14883_ & new_n14851_ & new_n14867_ & new_n14899_;
  assign new_n10746_ = new_n14826_ & new_n14794_ & new_n14810_ & new_n14842_;
  assign new_n10747_ = new_n14890_ & new_n14858_ & new_n14874_ & new_n14913_;
  assign new_n10748_ = new_n14825_ & new_n14793_ & new_n14809_ & new_n14841_;
  assign new_n10749_ = new_n14889_ & new_n14857_ & new_n14873_ & new_n14911_;
  assign new_n10750_ = new_n10751_ & new_n11458_;
  assign new_n10751_ = pi0627 & new_n11636_;
  assign new_n10752_ = new_n9401_ & new_n10307_;
  assign new_n10753_ = new_n10562_ & new_n14908_;
  assign new_n10754_ = new_n11640_ & new_n11639_;
  assign new_n10755_ = pi0625 & new_n10614_;
  assign new_n10756_ = new_n10755_ & new_n11659_;
  assign new_n10757_ = new_n11665_ & new_n10345_;
  assign new_n10758_ = new_n11507_ & new_n10306_;
  assign new_n10759_ = pi0624 & new_n10310_;
  assign new_n10760_ = ~pi0625 & ~pi0626;
  assign new_n10761_ = new_n11506_ & new_n11494_;
  assign new_n10762_ = new_n10761_ & new_n11673_;
  assign new_n10763_ = new_n11484_ & new_n11702_ & new_n11703_;
  assign new_n10764_ = new_n11712_ & new_n11711_ & new_n11710_;
  assign new_n10765_ = new_n11717_ & new_n11716_ & new_n11715_;
  assign new_n10766_ = new_n11722_ & new_n11721_ & new_n11720_;
  assign new_n10767_ = new_n11727_ & new_n11726_ & new_n11725_;
  assign new_n10768_ = new_n11732_ & new_n11731_ & new_n11730_;
  assign new_n10769_ = new_n11737_ & new_n11736_ & new_n11735_;
  assign new_n10770_ = new_n11742_ & new_n11741_ & new_n11740_;
  assign new_n10771_ = new_n11747_ & new_n11746_ & new_n11745_;
  assign new_n10772_ = new_n11484_ & new_n11760_ & new_n11761_;
  assign new_n10773_ = new_n11770_ & new_n11769_ & new_n11768_;
  assign new_n10774_ = new_n11775_ & new_n11774_ & new_n11773_;
  assign new_n10775_ = new_n11780_ & new_n11779_ & new_n11778_;
  assign new_n10776_ = new_n11785_ & new_n11784_ & new_n11783_;
  assign new_n10777_ = new_n11790_ & new_n11789_ & new_n11788_;
  assign new_n10778_ = new_n11795_ & new_n11794_ & new_n11793_;
  assign new_n10779_ = new_n11800_ & new_n11799_ & new_n11798_;
  assign new_n10780_ = new_n11805_ & new_n11804_ & new_n11803_;
  assign new_n10781_ = new_n11484_ & new_n11819_ & new_n11820_;
  assign new_n10782_ = new_n11829_ & new_n11828_ & new_n11827_;
  assign new_n10783_ = new_n11834_ & new_n11833_ & new_n11832_;
  assign new_n10784_ = new_n11839_ & new_n11838_ & new_n11837_;
  assign new_n10785_ = new_n11844_ & new_n11843_ & new_n11842_;
  assign new_n10786_ = new_n11849_ & new_n11848_ & new_n11847_;
  assign new_n10787_ = new_n11854_ & new_n11853_ & new_n11852_;
  assign new_n10788_ = new_n11859_ & new_n11858_ & new_n11857_;
  assign new_n10789_ = new_n11864_ & new_n11863_ & new_n11862_;
  assign new_n10790_ = new_n11484_ & new_n11876_ & new_n11877_;
  assign new_n10791_ = new_n11886_ & new_n11885_ & new_n11884_;
  assign new_n10792_ = new_n11891_ & new_n11890_ & new_n11889_;
  assign new_n10793_ = new_n11896_ & new_n11895_ & new_n11894_;
  assign new_n10794_ = new_n11901_ & new_n11900_ & new_n11899_;
  assign new_n10795_ = new_n11906_ & new_n11905_ & new_n11904_;
  assign new_n10796_ = new_n11911_ & new_n11910_ & new_n11909_;
  assign new_n10797_ = new_n11916_ & new_n11915_ & new_n11914_;
  assign new_n10798_ = new_n11921_ & new_n11920_ & new_n11919_;
  assign new_n10799_ = new_n11484_ & new_n11934_ & new_n11935_;
  assign new_n10800_ = new_n11944_ & new_n11943_ & new_n11942_;
  assign new_n10801_ = new_n11949_ & new_n11948_ & new_n11947_;
  assign new_n10802_ = new_n11954_ & new_n11953_ & new_n11952_;
  assign new_n10803_ = new_n11959_ & new_n11958_ & new_n11957_;
  assign new_n10804_ = new_n11964_ & new_n11963_ & new_n11962_;
  assign new_n10805_ = new_n11969_ & new_n11968_ & new_n11967_;
  assign new_n10806_ = new_n11974_ & new_n11973_ & new_n11972_;
  assign new_n10807_ = new_n11979_ & new_n11978_ & new_n11977_;
  assign new_n10808_ = new_n11484_ & new_n11991_ & new_n11992_;
  assign new_n10809_ = new_n12001_ & new_n12000_ & new_n11999_;
  assign new_n10810_ = new_n12006_ & new_n12005_ & new_n12004_;
  assign new_n10811_ = new_n12011_ & new_n12010_ & new_n12009_;
  assign new_n10812_ = new_n12016_ & new_n12015_ & new_n12014_;
  assign new_n10813_ = new_n12021_ & new_n12020_ & new_n12019_;
  assign new_n10814_ = new_n12026_ & new_n12025_ & new_n12024_;
  assign new_n10815_ = new_n12031_ & new_n12030_ & new_n12029_;
  assign new_n10816_ = new_n12036_ & new_n12035_ & new_n12034_;
  assign new_n10817_ = new_n11484_ & new_n12049_ & new_n12050_;
  assign new_n10818_ = new_n12059_ & new_n12058_ & new_n12057_;
  assign new_n10819_ = new_n12064_ & new_n12063_ & new_n12062_;
  assign new_n10820_ = new_n12069_ & new_n12068_ & new_n12067_;
  assign new_n10821_ = new_n12074_ & new_n12073_ & new_n12072_;
  assign new_n10822_ = new_n12079_ & new_n12078_ & new_n12077_;
  assign new_n10823_ = new_n12084_ & new_n12083_ & new_n12082_;
  assign new_n10824_ = new_n12089_ & new_n12088_ & new_n12087_;
  assign new_n10825_ = new_n12094_ & new_n12093_ & new_n12092_;
  assign new_n10826_ = new_n11484_ & new_n12106_ & new_n12107_;
  assign new_n10827_ = new_n12116_ & new_n12115_ & new_n12114_;
  assign new_n10828_ = new_n12121_ & new_n12120_ & new_n12119_;
  assign new_n10829_ = new_n12126_ & new_n12125_ & new_n12124_;
  assign new_n10830_ = new_n12131_ & new_n12130_ & new_n12129_;
  assign new_n10831_ = new_n12136_ & new_n12135_ & new_n12134_;
  assign new_n10832_ = new_n12141_ & new_n12140_ & new_n12139_;
  assign new_n10833_ = new_n12146_ & new_n12145_ & new_n12144_;
  assign new_n10834_ = new_n12151_ & new_n12150_ & new_n12149_;
  assign new_n10835_ = new_n11484_ & new_n12162_ & new_n12163_;
  assign new_n10836_ = new_n12172_ & new_n12171_ & new_n12170_;
  assign new_n10837_ = new_n12177_ & new_n12176_ & new_n12175_;
  assign new_n10838_ = new_n12182_ & new_n12181_ & new_n12180_;
  assign new_n10839_ = new_n12187_ & new_n12186_ & new_n12185_;
  assign new_n10840_ = new_n12192_ & new_n12191_ & new_n12190_;
  assign new_n10841_ = new_n12197_ & new_n12196_ & new_n12195_;
  assign new_n10842_ = new_n12202_ & new_n12201_ & new_n12200_;
  assign new_n10843_ = new_n12207_ & new_n12206_ & new_n12205_;
  assign new_n10844_ = new_n11484_ & new_n12219_ & new_n12220_;
  assign new_n10845_ = new_n12229_ & new_n12228_ & new_n12227_;
  assign new_n10846_ = new_n12234_ & new_n12233_ & new_n12232_;
  assign new_n10847_ = new_n12239_ & new_n12238_ & new_n12237_;
  assign new_n10848_ = new_n12244_ & new_n12243_ & new_n12242_;
  assign new_n10849_ = new_n12249_ & new_n12248_ & new_n12247_;
  assign new_n10850_ = new_n12254_ & new_n12253_ & new_n12252_;
  assign new_n10851_ = new_n12259_ & new_n12258_ & new_n12257_;
  assign new_n10852_ = new_n12264_ & new_n12263_ & new_n12262_;
  assign new_n10853_ = new_n11484_ & new_n12277_ & new_n12278_;
  assign new_n10854_ = new_n12287_ & new_n12286_ & new_n12285_;
  assign new_n10855_ = new_n12292_ & new_n12291_ & new_n12290_;
  assign new_n10856_ = new_n12297_ & new_n12296_ & new_n12295_;
  assign new_n10857_ = new_n12302_ & new_n12301_ & new_n12300_;
  assign new_n10858_ = new_n12307_ & new_n12306_ & new_n12305_;
  assign new_n10859_ = new_n12312_ & new_n12311_ & new_n12310_;
  assign new_n10860_ = new_n12317_ & new_n12316_ & new_n12315_;
  assign new_n10861_ = new_n12322_ & new_n12321_ & new_n12320_;
  assign new_n10862_ = new_n11484_ & new_n12334_ & new_n12335_;
  assign new_n10863_ = new_n12344_ & new_n12343_ & new_n12342_;
  assign new_n10864_ = new_n12349_ & new_n12348_ & new_n12347_;
  assign new_n10865_ = new_n12354_ & new_n12353_ & new_n12352_;
  assign new_n10866_ = new_n12359_ & new_n12358_ & new_n12357_;
  assign new_n10867_ = new_n12364_ & new_n12363_ & new_n12362_;
  assign new_n10868_ = new_n12369_ & new_n12368_ & new_n12367_;
  assign new_n10869_ = new_n12374_ & new_n12373_ & new_n12372_;
  assign new_n10870_ = new_n12379_ & new_n12378_ & new_n12377_;
  assign new_n10871_ = new_n11484_ & new_n12392_ & new_n12393_;
  assign new_n10872_ = new_n12402_ & new_n12401_ & new_n12400_;
  assign new_n10873_ = new_n12407_ & new_n12406_ & new_n12405_;
  assign new_n10874_ = new_n12412_ & new_n12411_ & new_n12410_;
  assign new_n10875_ = new_n12417_ & new_n12416_ & new_n12415_;
  assign new_n10876_ = new_n12422_ & new_n12421_ & new_n12420_;
  assign new_n10877_ = new_n12427_ & new_n12426_ & new_n12425_;
  assign new_n10878_ = new_n12432_ & new_n12431_ & new_n12430_;
  assign new_n10879_ = new_n12437_ & new_n12436_ & new_n12435_;
  assign new_n10880_ = new_n11484_ & new_n12449_ & new_n12450_;
  assign new_n10881_ = new_n12459_ & new_n12458_ & new_n12457_;
  assign new_n10882_ = new_n12464_ & new_n12463_ & new_n12462_;
  assign new_n10883_ = new_n12469_ & new_n12468_ & new_n12467_;
  assign new_n10884_ = new_n12474_ & new_n12473_ & new_n12472_;
  assign new_n10885_ = new_n12479_ & new_n12478_ & new_n12477_;
  assign new_n10886_ = new_n12484_ & new_n12483_ & new_n12482_;
  assign new_n10887_ = new_n12489_ & new_n12488_ & new_n12487_;
  assign new_n10888_ = new_n12494_ & new_n12493_ & new_n12492_;
  assign new_n10889_ = new_n11484_ & new_n12507_ & new_n12508_;
  assign new_n10890_ = new_n12517_ & new_n12516_ & new_n12515_;
  assign new_n10891_ = new_n12522_ & new_n12521_ & new_n12520_;
  assign new_n10892_ = new_n12527_ & new_n12526_ & new_n12525_;
  assign new_n10893_ = new_n12532_ & new_n12531_ & new_n12530_;
  assign new_n10894_ = new_n12537_ & new_n12536_ & new_n12535_;
  assign new_n10895_ = new_n12542_ & new_n12541_ & new_n12540_;
  assign new_n10896_ = new_n12547_ & new_n12546_ & new_n12545_;
  assign new_n10897_ = new_n12552_ & new_n12551_ & new_n12550_;
  assign new_n10898_ = new_n11484_ & new_n12564_ & new_n12565_;
  assign new_n10899_ = new_n12574_ & new_n12573_ & new_n12572_;
  assign new_n10900_ = new_n12579_ & new_n12578_ & new_n12577_;
  assign new_n10901_ = new_n12584_ & new_n12583_ & new_n12582_;
  assign new_n10902_ = new_n12589_ & new_n12588_ & new_n12587_;
  assign new_n10903_ = new_n12594_ & new_n12593_ & new_n12592_;
  assign new_n10904_ = new_n12599_ & new_n12598_ & new_n12597_;
  assign new_n10905_ = new_n12604_ & new_n12603_ & new_n12602_;
  assign new_n10906_ = new_n12609_ & new_n12608_ & new_n12607_;
  assign new_n10907_ = new_n29005_ & new_n11507_;
  assign new_n10908_ = pi0994 & pi0627;
  assign new_n10909_ = new_n12614_ & new_n12612_;
  assign new_n10910_ = new_n10909_ & new_n12617_;
  assign new_n10911_ = new_n11501_ & new_n11497_;
  assign new_n10912_ = new_n15111_ & new_n9553_ & new_n10911_ & new_n15112_;
  assign new_n10913_ = new_n12624_ & new_n11496_;
  assign new_n10914_ = new_n10562_ & new_n14910_;
  assign new_n10915_ = new_n14902_ & new_n10319_;
  assign new_n10916_ = new_n10915_ & new_n11470_;
  assign new_n10917_ = new_n11470_ & new_n10320_;
  assign new_n10918_ = new_n14900_ & new_n12634_;
  assign new_n10919_ = new_n14904_ & new_n10562_;
  assign new_n10920_ = new_n10322_ & new_n12628_ & new_n12629_;
  assign new_n10921_ = new_n12640_ & new_n10295_;
  assign new_n10922_ = new_n10921_ & new_n12642_ & new_n12641_;
  assign new_n10923_ = new_n14938_ & new_n12643_;
  assign new_n10924_ = new_n12649_ & new_n12648_;
  assign new_n10925_ = new_n10924_ & new_n12650_;
  assign new_n10926_ = new_n11437_ & new_n12658_;
  assign new_n10927_ = new_n11642_ & new_n9490_;
  assign new_n10928_ = new_n10623_ & new_n14900_;
  assign new_n10929_ = new_n12668_ & new_n12667_;
  assign new_n10930_ = new_n14900_ & new_n10313_;
  assign new_n10931_ = new_n12676_ & new_n12675_;
  assign new_n10932_ = new_n12690_ & new_n12691_;
  assign new_n10933_ = new_n12694_ & new_n12695_;
  assign new_n10934_ = new_n12699_ & new_n12700_;
  assign new_n10935_ = new_n11497_ & new_n11501_ & new_n12709_;
  assign new_n10936_ = new_n12715_ & new_n10619_;
  assign new_n10937_ = new_n12722_ & new_n12721_;
  assign new_n10938_ = new_n12724_ & new_n12723_;
  assign new_n10939_ = new_n12728_ & new_n12727_;
  assign new_n10940_ = new_n12730_ & new_n12729_;
  assign new_n10941_ = new_n12732_ & new_n12731_;
  assign new_n10942_ = new_n12736_ & new_n12735_;
  assign new_n10943_ = new_n12738_ & new_n12737_;
  assign new_n10944_ = new_n12740_ & new_n12739_;
  assign new_n10945_ = new_n12744_ & new_n12743_;
  assign new_n10946_ = new_n12746_ & new_n12745_;
  assign new_n10947_ = new_n12748_ & new_n12747_;
  assign new_n10948_ = new_n12752_ & new_n12751_;
  assign new_n10949_ = new_n12754_ & new_n12753_;
  assign new_n10950_ = new_n12756_ & new_n12755_;
  assign new_n10951_ = new_n12760_ & new_n12759_;
  assign new_n10952_ = new_n12762_ & new_n12761_;
  assign new_n10953_ = new_n12764_ & new_n12763_;
  assign new_n10954_ = new_n12768_ & new_n12767_;
  assign new_n10955_ = new_n12770_ & new_n12769_;
  assign new_n10956_ = new_n12772_ & new_n12771_;
  assign new_n10957_ = new_n12776_ & new_n12775_;
  assign new_n10958_ = new_n12778_ & new_n12777_;
  assign new_n10959_ = new_n12780_ & new_n12779_;
  assign new_n10960_ = new_n12784_ & new_n12783_;
  assign new_n10961_ = new_n12786_ & new_n12785_;
  assign new_n10962_ = new_n12788_ & new_n12787_;
  assign new_n10963_ = new_n12792_ & new_n12791_;
  assign new_n10964_ = new_n12794_ & new_n12793_;
  assign new_n10965_ = new_n12796_ & new_n12795_;
  assign new_n10966_ = new_n12800_ & new_n12799_;
  assign new_n10967_ = new_n12802_ & new_n12801_;
  assign new_n10968_ = new_n12804_ & new_n12803_;
  assign new_n10969_ = new_n12808_ & new_n12807_;
  assign new_n10970_ = new_n12810_ & new_n12809_;
  assign new_n10971_ = new_n12812_ & new_n12811_;
  assign new_n10972_ = new_n12816_ & new_n12815_;
  assign new_n10973_ = new_n12818_ & new_n12817_;
  assign new_n10974_ = new_n12820_ & new_n12819_;
  assign new_n10975_ = new_n12824_ & new_n12823_;
  assign new_n10976_ = new_n12826_ & new_n12825_;
  assign new_n10977_ = new_n12828_ & new_n12827_;
  assign new_n10978_ = new_n12832_ & new_n12831_;
  assign new_n10979_ = new_n12834_ & new_n12833_;
  assign new_n10980_ = new_n12836_ & new_n12835_;
  assign new_n10981_ = new_n12840_ & new_n12839_;
  assign new_n10982_ = new_n12842_ & new_n12841_;
  assign new_n10983_ = new_n12844_ & new_n12843_;
  assign new_n10984_ = new_n12848_ & new_n12847_;
  assign new_n10985_ = new_n12850_ & new_n12849_;
  assign new_n10986_ = new_n12852_ & new_n12851_;
  assign new_n10987_ = new_n12856_ & new_n12855_;
  assign new_n10988_ = new_n12858_ & new_n12857_;
  assign new_n10989_ = new_n12860_ & new_n12859_;
  assign new_n10990_ = new_n12864_ & new_n12863_;
  assign new_n10991_ = new_n12866_ & new_n12865_;
  assign new_n10992_ = new_n12868_ & new_n12867_;
  assign new_n10993_ = new_n12872_ & new_n12871_;
  assign new_n10994_ = new_n12874_ & new_n12873_;
  assign new_n10995_ = new_n12876_ & new_n12875_;
  assign new_n10996_ = new_n12880_ & new_n12879_;
  assign new_n10997_ = new_n12882_ & new_n12881_;
  assign new_n10998_ = new_n12884_ & new_n12883_;
  assign new_n10999_ = new_n12888_ & new_n12887_;
  assign new_n11000_ = new_n12890_ & new_n12889_;
  assign new_n11001_ = new_n12892_ & new_n12891_;
  assign new_n11002_ = new_n12896_ & new_n12895_;
  assign new_n11003_ = new_n12898_ & new_n12897_;
  assign new_n11004_ = new_n12900_ & new_n12899_;
  assign new_n11005_ = new_n12904_ & new_n12903_;
  assign new_n11006_ = new_n12906_ & new_n12905_;
  assign new_n11007_ = new_n12908_ & new_n12907_;
  assign new_n11008_ = new_n12912_ & new_n12911_;
  assign new_n11009_ = new_n12914_ & new_n12913_;
  assign new_n11010_ = new_n12916_ & new_n12915_;
  assign new_n11011_ = new_n12920_ & new_n12919_;
  assign new_n11012_ = new_n12922_ & new_n12921_;
  assign new_n11013_ = new_n12924_ & new_n12923_;
  assign new_n11014_ = new_n12928_ & new_n12927_;
  assign new_n11015_ = new_n12930_ & new_n12929_;
  assign new_n11016_ = new_n12932_ & new_n12931_;
  assign new_n11017_ = new_n12936_ & new_n12935_;
  assign new_n11018_ = new_n12938_ & new_n12937_;
  assign new_n11019_ = new_n12940_ & new_n12939_;
  assign new_n11020_ = new_n12944_ & new_n12943_;
  assign new_n11021_ = new_n12946_ & new_n12945_;
  assign new_n11022_ = new_n12948_ & new_n12947_;
  assign new_n11023_ = new_n12952_ & new_n12951_;
  assign new_n11024_ = new_n12955_ & new_n12953_ & new_n12954_ & new_n12956_;
  assign new_n11025_ = new_n12960_ & new_n12959_;
  assign new_n11026_ = new_n12962_ & new_n12964_ & new_n12963_;
  assign new_n11027_ = new_n12968_ & new_n12967_;
  assign new_n11028_ = new_n12970_ & new_n12972_ & new_n12971_;
  assign new_n11029_ = new_n12976_ & new_n12975_;
  assign new_n11030_ = pi0626 & pi0996;
  assign new_n11031_ = ~pi0625 & ~pi0626;
  assign new_n11032_ = new_n12984_ & new_n12983_ & new_n12982_;
  assign new_n11033_ = new_n12987_ & new_n12986_ & new_n12985_;
  assign new_n11034_ = new_n12990_ & new_n12989_ & new_n12988_;
  assign new_n11035_ = new_n12993_ & new_n12992_ & new_n12991_;
  assign new_n11036_ = new_n12996_ & new_n12995_ & new_n12994_;
  assign new_n11037_ = new_n12999_ & new_n12998_ & new_n12997_;
  assign new_n11038_ = new_n13002_ & new_n13001_ & new_n13000_;
  assign new_n11039_ = new_n13005_ & new_n13004_ & new_n13003_;
  assign new_n11040_ = new_n13008_ & new_n13007_ & new_n13006_;
  assign new_n11041_ = new_n13011_ & new_n13010_ & new_n13009_;
  assign new_n11042_ = new_n13014_ & new_n13013_ & new_n13012_;
  assign new_n11043_ = new_n13017_ & new_n13016_ & new_n13015_;
  assign new_n11044_ = new_n13020_ & new_n13019_ & new_n13018_;
  assign new_n11045_ = new_n13023_ & new_n13022_ & new_n13021_;
  assign new_n11046_ = new_n13026_ & new_n13025_ & new_n13024_;
  assign new_n11047_ = new_n13029_ & new_n13028_ & new_n13027_;
  assign new_n11048_ = new_n13032_ & new_n13031_ & new_n13030_;
  assign new_n11049_ = new_n13035_ & new_n13034_ & new_n13033_;
  assign new_n11050_ = new_n13038_ & new_n13037_ & new_n13036_;
  assign new_n11051_ = new_n13041_ & new_n13040_ & new_n13039_;
  assign new_n11052_ = new_n13044_ & new_n13043_ & new_n13042_;
  assign new_n11053_ = new_n13047_ & new_n13046_ & new_n13045_;
  assign new_n11054_ = new_n13050_ & new_n13049_ & new_n13048_;
  assign new_n11055_ = new_n13053_ & new_n13052_ & new_n13051_;
  assign new_n11056_ = new_n13056_ & new_n13055_ & new_n13054_;
  assign new_n11057_ = new_n13059_ & new_n13058_ & new_n13057_;
  assign new_n11058_ = new_n13062_ & new_n13061_ & new_n13060_;
  assign new_n11059_ = new_n13065_ & new_n13064_ & new_n13063_;
  assign new_n11060_ = new_n13068_ & new_n13067_ & new_n13066_;
  assign new_n11061_ = new_n13071_ & new_n13070_ & new_n13069_;
  assign new_n11062_ = new_n13074_ & new_n13073_ & new_n13072_;
  assign new_n11063_ = new_n13077_ & new_n13076_ & new_n13075_;
  assign new_n11064_ = new_n13080_ & new_n13079_ & new_n13078_;
  assign new_n11065_ = new_n13083_ & new_n13082_ & new_n13081_;
  assign new_n11066_ = new_n13086_ & new_n13085_ & new_n13084_;
  assign new_n11067_ = new_n13089_ & new_n13088_ & new_n13087_;
  assign new_n11068_ = new_n13092_ & new_n13091_ & new_n13090_;
  assign new_n11069_ = new_n13095_ & new_n13094_ & new_n13093_;
  assign new_n11070_ = new_n13098_ & new_n13097_ & new_n13096_;
  assign new_n11071_ = new_n13101_ & new_n13100_ & new_n13099_;
  assign new_n11072_ = new_n13104_ & new_n13103_ & new_n13102_;
  assign new_n11073_ = new_n13107_ & new_n13106_ & new_n13105_;
  assign new_n11074_ = new_n13110_ & new_n13109_ & new_n13108_;
  assign new_n11075_ = new_n13113_ & new_n13112_ & new_n13111_;
  assign new_n11076_ = new_n13116_ & new_n13115_ & new_n13114_;
  assign new_n11077_ = new_n13119_ & new_n13118_ & new_n13117_;
  assign new_n11078_ = new_n13122_ & new_n13121_ & new_n13120_;
  assign new_n11079_ = new_n13125_ & new_n13124_ & new_n13123_;
  assign new_n11080_ = new_n13128_ & new_n13127_ & new_n13126_;
  assign new_n11081_ = new_n13131_ & new_n13130_ & new_n13129_;
  assign new_n11082_ = new_n13134_ & new_n13133_ & new_n13132_;
  assign new_n11083_ = new_n13137_ & new_n13136_ & new_n13135_;
  assign new_n11084_ = new_n13140_ & new_n13139_ & new_n13138_;
  assign new_n11085_ = new_n13143_ & new_n13142_ & new_n13141_;
  assign new_n11086_ = new_n13146_ & new_n13145_ & new_n13144_;
  assign new_n11087_ = new_n13149_ & new_n13148_ & new_n13147_;
  assign new_n11088_ = new_n13152_ & new_n13151_ & new_n13150_;
  assign new_n11089_ = new_n13155_ & new_n13154_ & new_n13153_;
  assign new_n11090_ = new_n13158_ & new_n13157_ & new_n13156_;
  assign new_n11091_ = new_n13161_ & new_n13160_ & new_n13159_;
  assign new_n11092_ = new_n13164_ & new_n13163_ & new_n13162_;
  assign new_n11093_ = new_n13166_ & new_n13167_ & new_n13165_;
  assign new_n11094_ = new_n13170_ & new_n13169_ & new_n13168_;
  assign new_n11095_ = new_n13173_ & new_n13172_ & new_n13171_;
  assign new_n11096_ = new_n9397_ & new_n11509_ & new_n13174_;
  assign new_n11097_ = new_n14912_ & new_n10321_ & pi0627;
  assign new_n11098_ = new_n9657_ & new_n11509_;
  assign new_n11099_ = new_n9415_ & new_n11458_;
  assign new_n11100_ = new_n13371_ & new_n13370_;
  assign new_n11101_ = new_n13375_ & new_n13374_;
  assign new_n11102_ = new_n13379_ & new_n13378_;
  assign new_n11103_ = new_n13383_ & new_n13382_;
  assign new_n11104_ = new_n13387_ & new_n13386_;
  assign new_n11105_ = new_n13391_ & new_n13390_;
  assign new_n11106_ = new_n13395_ & new_n13394_;
  assign new_n11107_ = new_n13399_ & new_n13398_;
  assign new_n11108_ = new_n13403_ & new_n13402_;
  assign new_n11109_ = new_n13407_ & new_n13406_;
  assign new_n11110_ = new_n13610_ & new_n11495_ & new_n11494_;
  assign new_n11111_ = new_n11112_ & new_n13615_ & new_n13614_;
  assign new_n11112_ = new_n13618_ & new_n13617_;
  assign new_n11113_ = new_n11114_ & new_n13619_;
  assign new_n11114_ = new_n13622_ & new_n13621_;
  assign new_n11115_ = new_n11116_ & new_n13624_ & new_n13623_;
  assign new_n11116_ = new_n13627_ & new_n13626_;
  assign new_n11117_ = new_n11118_ & new_n13628_;
  assign new_n11118_ = new_n13631_ & new_n13630_;
  assign new_n11119_ = new_n11120_ & new_n13633_ & new_n13632_;
  assign new_n11120_ = new_n13636_ & new_n13635_;
  assign new_n11121_ = new_n11122_ & new_n13637_;
  assign new_n11122_ = new_n13640_ & new_n13639_;
  assign new_n11123_ = new_n11124_ & new_n13642_ & new_n13641_;
  assign new_n11124_ = new_n13645_ & new_n13644_;
  assign new_n11125_ = new_n11126_ & new_n13646_;
  assign new_n11126_ = new_n13649_ & new_n13648_;
  assign new_n11127_ = new_n13651_ & new_n13650_ & new_n11487_;
  assign new_n11128_ = new_n11129_ & new_n13656_;
  assign new_n11129_ = new_n13658_ & new_n13657_;
  assign new_n11130_ = new_n13653_ & new_n13655_ & new_n13654_ & new_n11127_ & new_n13652_;
  assign new_n11131_ = new_n13660_ & new_n13659_ & new_n11487_;
  assign new_n11132_ = new_n11133_ & new_n13665_;
  assign new_n11133_ = new_n13667_ & new_n13666_;
  assign new_n11134_ = new_n13662_ & new_n13664_ & new_n13663_ & new_n11131_ & new_n13661_;
  assign new_n11135_ = new_n13669_ & new_n13668_ & new_n11487_;
  assign new_n11136_ = new_n11137_ & new_n13672_;
  assign new_n11137_ = new_n13675_ & new_n13674_;
  assign new_n11138_ = new_n13677_ & new_n13676_ & new_n11487_;
  assign new_n11139_ = new_n11140_ & new_n13680_;
  assign new_n11140_ = new_n13683_ & new_n13682_;
  assign new_n11141_ = new_n13685_ & new_n13684_ & new_n11487_;
  assign new_n11142_ = new_n11143_ & new_n13688_;
  assign new_n11143_ = new_n13691_ & new_n13690_;
  assign new_n11144_ = new_n13693_ & new_n13692_ & new_n11487_;
  assign new_n11145_ = new_n11146_ & new_n13696_;
  assign new_n11146_ = new_n13699_ & new_n13698_;
  assign new_n11147_ = new_n13701_ & new_n13700_ & new_n11487_;
  assign new_n11148_ = new_n11149_ & new_n13704_;
  assign new_n11149_ = new_n13707_ & new_n13706_;
  assign new_n11150_ = new_n13709_ & new_n13708_ & new_n11487_;
  assign new_n11151_ = new_n11152_ & new_n13712_;
  assign new_n11152_ = new_n13715_ & new_n13714_;
  assign new_n11153_ = new_n13719_ & new_n13716_ & new_n11487_;
  assign new_n11154_ = new_n11155_ & new_n13720_;
  assign new_n11155_ = new_n13723_ & new_n13722_;
  assign new_n11156_ = new_n13727_ & new_n13724_ & new_n11487_;
  assign new_n11157_ = new_n11158_ & new_n13728_;
  assign new_n11158_ = new_n13731_ & new_n13730_;
  assign new_n11159_ = new_n13735_ & new_n13732_ & new_n11487_;
  assign new_n11160_ = new_n11161_ & new_n13736_;
  assign new_n11161_ = new_n13739_ & new_n13738_;
  assign new_n11162_ = new_n13740_ & new_n11487_;
  assign new_n11163_ = new_n11164_ & new_n13744_;
  assign new_n11164_ = new_n13747_ & new_n13746_;
  assign new_n11165_ = new_n11162_ & new_n13745_ & new_n13741_ & new_n13743_ & new_n13742_;
  assign new_n11166_ = new_n13748_ & new_n11487_;
  assign new_n11167_ = new_n11168_ & new_n13752_;
  assign new_n11168_ = new_n13755_ & new_n13754_;
  assign new_n11169_ = new_n11166_ & new_n13753_ & new_n13749_ & new_n13751_ & new_n13750_;
  assign new_n11170_ = new_n13756_ & new_n11487_;
  assign new_n11171_ = new_n11172_ & new_n13760_;
  assign new_n11172_ = new_n13763_ & new_n13762_;
  assign new_n11173_ = new_n11170_ & new_n13761_ & new_n13757_ & new_n13759_ & new_n13758_;
  assign new_n11174_ = new_n13764_ & new_n11487_;
  assign new_n11175_ = new_n11176_ & new_n13768_;
  assign new_n11176_ = new_n13771_ & new_n13770_;
  assign new_n11177_ = new_n11174_ & new_n13769_ & new_n13765_ & new_n13767_ & new_n13766_;
  assign new_n11178_ = new_n13772_ & new_n11487_;
  assign new_n11179_ = new_n11180_ & new_n13776_;
  assign new_n11180_ = new_n13779_ & new_n13778_;
  assign new_n11181_ = new_n11178_ & new_n13777_ & new_n13773_ & new_n13775_ & new_n13774_;
  assign new_n11182_ = new_n11183_ & new_n13784_;
  assign new_n11183_ = new_n13787_ & new_n13786_;
  assign new_n11184_ = new_n13780_ & new_n13785_ & new_n13781_ & new_n13783_ & new_n13782_;
  assign new_n11185_ = new_n11186_ & new_n13792_;
  assign new_n11186_ = new_n13795_ & new_n13794_;
  assign new_n11187_ = new_n13788_ & new_n13793_ & new_n13789_ & new_n13791_ & new_n13790_;
  assign new_n11188_ = new_n13803_ & new_n13802_;
  assign new_n11189_ = new_n13801_ & new_n11188_ & new_n13800_;
  assign new_n11190_ = new_n13804_ & new_n11191_ & new_n13809_ & new_n13807_ & new_n13806_;
  assign new_n11191_ = new_n11192_ & new_n13808_;
  assign new_n11192_ = new_n13811_ & new_n13810_;
  assign new_n11193_ = new_n13812_ & new_n11194_ & new_n13817_ & new_n13815_ & new_n13814_;
  assign new_n11194_ = new_n11195_ & new_n13816_;
  assign new_n11195_ = new_n13819_ & new_n13818_;
  assign new_n11196_ = new_n13827_ & new_n13826_;
  assign new_n11197_ = new_n13825_ & new_n11196_ & new_n13824_;
  assign new_n11198_ = new_n13835_ & new_n13834_;
  assign new_n11199_ = new_n13833_ & new_n11198_ & new_n13832_;
  assign new_n11200_ = new_n13843_ & new_n13842_;
  assign new_n11201_ = new_n13841_ & new_n11200_ & new_n13840_;
  assign new_n11202_ = new_n13851_ & new_n13850_;
  assign new_n11203_ = new_n13849_ & new_n11202_ & new_n13848_;
  assign new_n11204_ = new_n13859_ & new_n13858_;
  assign new_n11205_ = new_n13857_ & new_n11204_ & new_n13856_;
  assign new_n11206_ = new_n13867_ & new_n13866_;
  assign new_n11207_ = new_n13865_ & new_n11206_ & new_n13864_;
  assign new_n11208_ = new_n13875_ & new_n13874_;
  assign new_n11209_ = new_n13873_ & new_n11208_ & new_n13872_;
  assign new_n11210_ = ~pi0595 & ~pi0594 & ~pi0597 & ~pi0596;
  assign new_n11211_ = ~pi0599 & ~pi0598 & ~pi0601 & ~pi0600;
  assign new_n11212_ = new_n11211_ & new_n11210_;
  assign new_n11213_ = ~pi0603 & ~pi0602 & ~pi0605 & ~pi0604;
  assign new_n11214_ = ~pi0607 & ~pi0606 & ~pi0609 & ~pi0608;
  assign new_n11215_ = new_n11214_ & new_n11213_;
  assign new_n11216_ = ~pi0611 & ~pi0610 & ~pi0613 & ~pi0612;
  assign new_n11217_ = ~pi0615 & ~pi0614 & ~pi0617 & ~pi0616;
  assign new_n11218_ = new_n11217_ & new_n11216_;
  assign new_n11219_ = ~pi0618 & ~pi0619;
  assign new_n11220_ = ~pi0620 & ~pi0621;
  assign new_n11221_ = ~pi0622 & ~pi0623;
  assign new_n11222_ = new_n13876_ & new_n11219_ & new_n11220_ & new_n11221_;
  assign new_n11223_ = ~pi0957 & ~pi0592 & ~pi0593;
  assign new_n11224_ = ~pi0958 & ~pi0593;
  assign new_n11225_ = new_n13885_ & new_n14914_;
  assign new_n11226_ = new_n13889_ & new_n10342_;
  assign new_n11227_ = new_n11226_ & new_n13890_;
  assign new_n11228_ = pi0626 & new_n10306_;
  assign new_n11229_ = new_n13882_ & new_n13883_ & new_n10354_;
  assign new_n11230_ = new_n9415_ & new_n10294_;
  assign new_n11231_ = new_n13901_ & new_n10575_;
  assign new_n11232_ = new_n13905_ & new_n13903_ & new_n13904_ & new_n13906_;
  assign new_n11233_ = new_n13909_ & new_n13907_ & new_n13908_ & new_n13910_;
  assign new_n11234_ = new_n13913_ & new_n13911_ & new_n13912_ & new_n13914_;
  assign new_n11235_ = new_n13917_ & new_n13915_ & new_n13916_ & new_n13918_;
  assign new_n11236_ = new_n13921_ & new_n13919_ & new_n13920_ & new_n13922_;
  assign new_n11237_ = new_n13925_ & new_n13923_ & new_n13924_ & new_n13926_;
  assign new_n11238_ = new_n13929_ & new_n13927_ & new_n13928_ & new_n13930_;
  assign new_n11239_ = new_n13933_ & new_n13931_ & new_n13932_ & new_n13934_;
  assign new_n11240_ = new_n13937_ & new_n13935_ & new_n13936_ & new_n13938_;
  assign new_n11241_ = new_n13941_ & new_n13939_ & new_n13940_ & new_n13942_;
  assign new_n11242_ = new_n13945_ & new_n13943_ & new_n13944_ & new_n13946_;
  assign new_n11243_ = new_n13949_ & new_n13947_ & new_n13948_ & new_n13950_;
  assign new_n11244_ = new_n13953_ & new_n13951_ & new_n13952_ & new_n13954_;
  assign new_n11245_ = new_n13957_ & new_n13955_ & new_n13956_ & new_n13958_;
  assign new_n11246_ = new_n13961_ & new_n13959_ & new_n13960_ & new_n13962_;
  assign new_n11247_ = new_n13965_ & new_n13963_ & new_n13964_ & new_n13966_;
  assign new_n11248_ = new_n13969_ & new_n13967_ & new_n13968_ & new_n13970_;
  assign new_n11249_ = new_n13973_ & new_n13971_ & new_n13972_ & new_n13974_;
  assign new_n11250_ = new_n13977_ & new_n13975_ & new_n13976_ & new_n13978_;
  assign new_n11251_ = new_n13981_ & new_n13979_ & new_n13980_ & new_n13982_;
  assign new_n11252_ = new_n13985_ & new_n13983_ & new_n13984_ & new_n13986_;
  assign new_n11253_ = new_n13989_ & new_n13987_ & new_n13988_ & new_n13990_;
  assign new_n11254_ = new_n13993_ & new_n13991_ & new_n13992_ & new_n13994_;
  assign new_n11255_ = new_n13997_ & new_n13995_ & new_n13996_ & new_n13998_;
  assign new_n11256_ = new_n14001_ & new_n13999_ & new_n14000_ & new_n14002_;
  assign new_n11257_ = new_n14005_ & new_n14003_ & new_n14004_ & new_n14006_;
  assign new_n11258_ = new_n14009_ & new_n14007_ & new_n14008_ & new_n14010_;
  assign new_n11259_ = new_n14013_ & new_n14011_ & new_n14012_ & new_n14014_;
  assign new_n11260_ = new_n14017_ & new_n14015_ & new_n14016_ & new_n14018_;
  assign new_n11261_ = new_n14021_ & new_n14019_ & new_n14020_ & new_n14022_;
  assign new_n11262_ = new_n14025_ & new_n14023_ & new_n14024_ & new_n14026_;
  assign new_n11263_ = new_n14029_ & new_n14027_ & new_n14028_ & new_n14030_;
  assign new_n11264_ = new_n14033_ & new_n14031_ & new_n14032_ & new_n14034_;
  assign new_n11265_ = new_n14037_ & new_n14035_ & new_n14036_ & new_n14038_;
  assign new_n11266_ = new_n14041_ & new_n14039_ & new_n14040_ & new_n14042_;
  assign new_n11267_ = new_n14045_ & new_n14043_ & new_n14044_ & new_n14046_;
  assign new_n11268_ = new_n14051_ & new_n14049_ & new_n14050_ & new_n14052_;
  assign new_n11269_ = new_n14055_ & new_n14053_ & new_n14054_ & new_n14056_;
  assign new_n11270_ = new_n14059_ & new_n14057_ & new_n14058_ & new_n14060_;
  assign new_n11271_ = new_n14063_ & new_n14061_ & new_n14062_ & new_n14064_;
  assign new_n11272_ = new_n14067_ & new_n14065_ & new_n14066_ & new_n14068_;
  assign new_n11273_ = new_n14071_ & new_n14069_ & new_n14070_ & new_n14072_;
  assign new_n11274_ = new_n14075_ & new_n14073_ & new_n14074_ & new_n14076_;
  assign new_n11275_ = new_n14079_ & new_n14077_ & new_n14078_ & new_n14080_;
  assign new_n11276_ = new_n14083_ & new_n14081_ & new_n14082_ & new_n14084_;
  assign new_n11277_ = new_n14087_ & new_n14085_ & new_n14086_ & new_n14088_;
  assign new_n11278_ = new_n14091_ & new_n14089_ & new_n14090_ & new_n14092_;
  assign new_n11279_ = new_n14095_ & new_n14093_ & new_n14094_ & new_n14096_;
  assign new_n11280_ = new_n14099_ & new_n14097_ & new_n14098_ & new_n14100_;
  assign new_n11281_ = new_n14103_ & new_n14101_ & new_n14102_ & new_n14104_;
  assign new_n11282_ = new_n14107_ & new_n14105_ & new_n14106_ & new_n14108_;
  assign new_n11283_ = new_n14111_ & new_n14109_ & new_n14110_ & new_n14112_;
  assign new_n11284_ = new_n14115_ & new_n14113_ & new_n14114_ & new_n14116_;
  assign new_n11285_ = new_n14119_ & new_n14117_ & new_n14118_ & new_n14120_;
  assign new_n11286_ = new_n14123_ & new_n14121_ & new_n14122_ & new_n14124_;
  assign new_n11287_ = new_n14127_ & new_n14125_ & new_n14126_ & new_n14128_;
  assign new_n11288_ = new_n14131_ & new_n14129_ & new_n14130_ & new_n14132_;
  assign new_n11289_ = new_n14135_ & new_n14133_ & new_n14134_ & new_n14136_;
  assign new_n11290_ = new_n14139_ & new_n14137_ & new_n14138_ & new_n14140_;
  assign new_n11291_ = new_n14143_ & new_n14141_ & new_n14142_ & new_n14144_;
  assign new_n11292_ = new_n14147_ & new_n14145_ & new_n14146_ & new_n14148_;
  assign new_n11293_ = new_n14151_ & new_n14149_ & new_n14150_ & new_n14152_;
  assign new_n11294_ = new_n14155_ & new_n14153_ & new_n14154_ & new_n14156_;
  assign new_n11295_ = new_n14159_ & new_n14157_ & new_n14158_ & new_n14160_;
  assign new_n11296_ = new_n14163_ & new_n14161_ & new_n14162_ & new_n14164_;
  assign new_n11297_ = new_n14167_ & new_n14165_ & new_n14166_ & new_n14168_;
  assign new_n11298_ = new_n14171_ & new_n14169_ & new_n14170_ & new_n14172_;
  assign new_n11299_ = new_n14175_ & new_n14173_ & new_n14174_ & new_n14176_;
  assign new_n11300_ = new_n14827_ & new_n14795_ & new_n14811_ & new_n14843_;
  assign new_n11301_ = new_n14891_ & new_n14859_ & new_n14875_ & new_n14915_;
  assign new_n11302_ = new_n14828_ & new_n14796_ & new_n14812_ & new_n14844_;
  assign new_n11303_ = new_n14892_ & new_n14860_ & new_n14876_ & new_n14916_;
  assign new_n11304_ = new_n14829_ & new_n14797_ & new_n14813_ & new_n14845_;
  assign new_n11305_ = new_n14893_ & new_n14861_ & new_n14877_ & new_n14917_;
  assign new_n11306_ = new_n14830_ & new_n14798_ & new_n14814_ & new_n14846_;
  assign new_n11307_ = new_n14894_ & new_n14862_ & new_n14878_ & new_n14918_;
  assign new_n11308_ = new_n14831_ & new_n14799_ & new_n14815_ & new_n14847_;
  assign new_n11309_ = new_n14895_ & new_n14863_ & new_n14879_ & new_n14919_;
  assign new_n11310_ = new_n14832_ & new_n14800_ & new_n14816_ & new_n14848_;
  assign new_n11311_ = new_n14896_ & new_n14864_ & new_n14880_ & new_n14920_;
  assign new_n11312_ = new_n14833_ & new_n14801_ & new_n14817_ & new_n14849_;
  assign new_n11313_ = new_n14897_ & new_n14865_ & new_n14881_ & new_n14921_;
  assign new_n11314_ = new_n14834_ & new_n14802_ & new_n14818_ & new_n14850_;
  assign new_n11315_ = new_n14898_ & new_n14866_ & new_n14882_ & new_n14922_;
  assign new_n11316_ = new_n14902_ & new_n11317_;
  assign new_n11317_ = pi0627 & pi0625 & new_n10341_;
  assign new_n11318_ = new_n14210_ & new_n14208_ & new_n14209_ & new_n14211_;
  assign new_n11319_ = new_n14214_ & new_n14212_ & new_n14213_ & new_n14215_;
  assign new_n11320_ = new_n14218_ & new_n14216_ & new_n14217_ & new_n14219_;
  assign new_n11321_ = new_n14222_ & new_n14220_ & new_n14221_ & new_n14223_;
  assign new_n11322_ = new_n14227_ & new_n14225_ & new_n14226_ & new_n14228_;
  assign new_n11323_ = new_n14231_ & new_n14229_ & new_n14230_ & new_n14232_;
  assign new_n11324_ = new_n14235_ & new_n14233_ & new_n14234_ & new_n14236_;
  assign new_n11325_ = new_n14239_ & new_n14237_ & new_n14238_ & new_n14240_;
  assign new_n11326_ = new_n14244_ & new_n14242_ & new_n14243_ & new_n14245_;
  assign new_n11327_ = new_n14248_ & new_n14246_ & new_n14247_ & new_n14249_;
  assign new_n11328_ = new_n14252_ & new_n14250_ & new_n14251_ & new_n14253_;
  assign new_n11329_ = new_n14256_ & new_n14254_ & new_n14255_ & new_n14257_;
  assign new_n11330_ = new_n14261_ & new_n14259_ & new_n14260_ & new_n14262_;
  assign new_n11331_ = new_n14265_ & new_n14263_ & new_n14264_ & new_n14266_;
  assign new_n11332_ = new_n14269_ & new_n14267_ & new_n14268_ & new_n14270_;
  assign new_n11333_ = new_n14273_ & new_n14271_ & new_n14272_ & new_n14274_;
  assign new_n11334_ = new_n14278_ & new_n14276_ & new_n14277_ & new_n14279_;
  assign new_n11335_ = new_n14282_ & new_n14280_ & new_n14281_ & new_n14283_;
  assign new_n11336_ = new_n14286_ & new_n14284_ & new_n14285_ & new_n14287_;
  assign new_n11337_ = new_n14290_ & new_n14288_ & new_n14289_ & new_n14291_;
  assign new_n11338_ = new_n14295_ & new_n14293_ & new_n14294_ & new_n14296_;
  assign new_n11339_ = new_n14299_ & new_n14297_ & new_n14298_ & new_n14300_;
  assign new_n11340_ = new_n14303_ & new_n14301_ & new_n14302_ & new_n14304_;
  assign new_n11341_ = new_n14307_ & new_n14305_ & new_n14306_ & new_n14308_;
  assign new_n11342_ = new_n14312_ & new_n14310_ & new_n14311_ & new_n14313_;
  assign new_n11343_ = new_n14316_ & new_n14314_ & new_n14315_ & new_n14317_;
  assign new_n11344_ = new_n14320_ & new_n14318_ & new_n14319_ & new_n14321_;
  assign new_n11345_ = new_n14324_ & new_n14322_ & new_n14323_ & new_n14325_;
  assign new_n11346_ = new_n14329_ & new_n14327_ & new_n14328_ & new_n14330_;
  assign new_n11347_ = new_n14333_ & new_n14331_ & new_n14332_ & new_n14334_;
  assign new_n11348_ = new_n14337_ & new_n14335_ & new_n14336_ & new_n14338_;
  assign new_n11349_ = new_n14341_ & new_n14339_ & new_n14340_ & new_n14342_;
  assign new_n11350_ = new_n14346_ & new_n14344_ & new_n14345_ & new_n14347_;
  assign new_n11351_ = new_n14350_ & new_n14348_ & new_n14349_ & new_n14351_;
  assign new_n11352_ = new_n14354_ & new_n14352_ & new_n14353_ & new_n14355_;
  assign new_n11353_ = new_n14358_ & new_n14356_ & new_n14357_ & new_n14359_;
  assign new_n11354_ = new_n14363_ & new_n14361_ & new_n14362_ & new_n14364_;
  assign new_n11355_ = new_n14367_ & new_n14365_ & new_n14366_ & new_n14368_;
  assign new_n11356_ = new_n14371_ & new_n14369_ & new_n14370_ & new_n14372_;
  assign new_n11357_ = new_n14375_ & new_n14373_ & new_n14374_ & new_n14376_;
  assign new_n11358_ = new_n14380_ & new_n14378_ & new_n14379_ & new_n14381_;
  assign new_n11359_ = new_n14384_ & new_n14382_ & new_n14383_ & new_n14385_;
  assign new_n11360_ = new_n14388_ & new_n14386_ & new_n14387_ & new_n14389_;
  assign new_n11361_ = new_n14392_ & new_n14390_ & new_n14391_ & new_n14393_;
  assign new_n11362_ = new_n14397_ & new_n14395_ & new_n14396_ & new_n14398_;
  assign new_n11363_ = new_n14401_ & new_n14399_ & new_n14400_ & new_n14402_;
  assign new_n11364_ = new_n14405_ & new_n14403_ & new_n14404_ & new_n14406_;
  assign new_n11365_ = new_n14409_ & new_n14407_ & new_n14408_ & new_n14410_;
  assign new_n11366_ = new_n14414_ & new_n14412_ & new_n14413_ & new_n14415_;
  assign new_n11367_ = new_n14418_ & new_n14416_ & new_n14417_ & new_n14419_;
  assign new_n11368_ = new_n14422_ & new_n14420_ & new_n14421_ & new_n14423_;
  assign new_n11369_ = new_n14426_ & new_n14424_ & new_n14425_ & new_n14427_;
  assign new_n11370_ = new_n14431_ & new_n14429_ & new_n14430_ & new_n14432_;
  assign new_n11371_ = new_n14435_ & new_n14433_ & new_n14434_ & new_n14436_;
  assign new_n11372_ = new_n14439_ & new_n14437_ & new_n14438_ & new_n14440_;
  assign new_n11373_ = new_n14443_ & new_n14441_ & new_n14442_ & new_n14444_;
  assign new_n11374_ = new_n14448_ & new_n14446_ & new_n14447_ & new_n14449_;
  assign new_n11375_ = new_n14452_ & new_n14450_ & new_n14451_ & new_n14453_;
  assign new_n11376_ = new_n14456_ & new_n14454_ & new_n14455_ & new_n14457_;
  assign new_n11377_ = new_n14460_ & new_n14458_ & new_n14459_ & new_n14461_;
  assign new_n11378_ = new_n9657_ & new_n10341_;
  assign new_n11379_ = new_n14466_ & new_n11454_;
  assign new_n11380_ = new_n11636_ & new_n10341_;
  assign new_n11381_ = new_n14469_ & new_n14467_ & new_n11455_;
  assign new_n11382_ = new_n14471_ & new_n10612_;
  assign new_n11383_ = new_n11454_ & new_n11382_;
  assign new_n11384_ = new_n14910_ & new_n14914_;
  assign new_n11385_ = new_n14477_ & new_n14476_;
  assign new_n11386_ = new_n14481_ & new_n14480_;
  assign new_n11387_ = new_n14483_ & new_n14484_;
  assign new_n11388_ = new_n14486_ & new_n14487_;
  assign new_n11389_ = new_n14489_ & new_n14490_;
  assign new_n11390_ = new_n14492_ & new_n14493_;
  assign new_n11391_ = new_n14495_ & new_n14496_;
  assign new_n11392_ = new_n14498_ & new_n14499_;
  assign new_n11393_ = new_n14501_ & new_n14502_;
  assign new_n11394_ = new_n14504_ & new_n14505_;
  assign new_n11395_ = new_n14507_ & new_n14508_;
  assign new_n11396_ = new_n14510_ & new_n14511_;
  assign new_n11397_ = new_n14513_ & new_n14514_;
  assign new_n11398_ = new_n14516_ & new_n14517_;
  assign new_n11399_ = new_n14519_ & new_n14520_;
  assign new_n11400_ = new_n14522_ & new_n14523_;
  assign new_n11401_ = new_n14525_ & new_n14526_;
  assign new_n11402_ = new_n14528_ & new_n14529_;
  assign new_n11403_ = new_n14531_ & new_n14532_;
  assign new_n11404_ = new_n14534_ & new_n14535_;
  assign new_n11405_ = new_n14537_ & new_n14538_;
  assign new_n11406_ = new_n14540_ & new_n14541_;
  assign new_n11407_ = new_n14543_ & new_n14544_;
  assign new_n11408_ = new_n14546_ & new_n14547_;
  assign new_n11409_ = new_n14551_ & new_n14550_;
  assign new_n11410_ = new_n14555_ & new_n14554_;
  assign new_n11411_ = new_n14559_ & new_n14558_;
  assign new_n11412_ = new_n14563_ & new_n14562_;
  assign new_n11413_ = new_n14567_ & new_n14566_;
  assign new_n11414_ = new_n14571_ & new_n14570_;
  assign new_n11415_ = new_n14573_ & new_n14574_;
  assign new_n11416_ = new_n14577_ & new_n14576_;
  assign new_n11417_ = new_n10296_ & new_n13886_;
  assign new_n11418_ = new_n14904_ & new_n10296_;
  assign new_n11419_ = new_n9397_ & new_n14914_;
  assign new_n11420_ = new_n14619_ & new_n14620_ & new_n14621_;
  assign new_n11421_ = new_n14626_ & new_n10310_;
  assign new_n11422_ = new_n9397_ & new_n11636_;
  assign new_n11423_ = new_n10618_ & new_n14627_ & new_n14628_ & new_n11513_ & new_n10580_;
  assign new_n11424_ = new_n14620_ & new_n11463_;
  assign new_n11425_ = new_n11424_ & new_n14619_;
  assign new_n11426_ = new_n14621_ & new_n11499_;
  assign new_n11427_ = new_n14631_ & new_n14630_;
  assign new_n11428_ = pi0627 & new_n14777_;
  assign new_n11429_ = new_n11499_ & new_n10590_ & new_n11498_ & new_n10614_;
  assign new_n11430_ = new_n14760_ & new_n14759_;
  assign new_n11431_ = new_n14772_ & new_n10577_;
  assign new_n11432_ = new_n14776_ & new_n10577_;
  assign new_n11433_ = new_n14949_ & new_n14948_;
  assign new_n11434_ = new_n15096_ & new_n15095_;
  assign new_n11435_ = ~new_n10913_ | ~new_n12623_;
  assign new_n11436_ = new_n15120_ & new_n15119_;
  assign new_n11437_ = new_n15133_ & new_n15132_;
  assign new_n11438_ = new_n15161_ & new_n15160_;
  assign new_n11439_ = new_n15167_ & new_n15166_;
  assign new_n11440_ = new_n15173_ & new_n15172_;
  assign new_n11441_ = ~new_n9415_ | ~new_n10332_;
  assign new_n11442_ = ~pi0035;
  assign new_n11443_ = ~new_n11503_ | ~new_n11229_;
  assign new_n11444_ = ~new_n10575_ | ~new_n11503_;
  assign new_n11445_ = new_n15187_ & new_n15186_;
  assign new_n11446_ = ~pi0758 | ~new_n14047_;
  assign new_n11447_ = ~new_n9554_ | ~new_n10912_;
  assign new_n11448_ = ~new_n29042_;
  assign new_n11449_ = ~new_n29021_;
  assign new_n11450_ = ~new_n10594_;
  assign new_n11451_ = ~pi0033 | ~new_n10306_;
  assign new_n11452_ = ~new_n10331_;
  assign new_n11453_ = ~new_n10612_;
  assign new_n11454_ = ~new_n11378_ | ~new_n11642_;
  assign new_n11455_ = ~new_n14910_ | ~new_n9657_ | ~new_n10341_;
  assign new_n11456_ = ~new_n9488_ | ~new_n10320_;
  assign new_n11457_ = ~new_n10617_;
  assign new_n11458_ = ~new_n10324_;
  assign new_n11459_ = ~new_n10591_;
  assign new_n11460_ = ~new_n10577_;
  assign new_n11461_ = ~new_n10329_;
  assign new_n11462_ = ~new_n10580_;
  assign new_n11463_ = ~new_n9491_ | ~new_n9417_ | ~new_n10319_;
  assign new_n11464_ = ~new_n10618_;
  assign new_n11465_ = ~new_n10323_;
  assign new_n11466_ = ~new_n10326_;
  assign new_n11467_ = ~new_n10590_;
  assign new_n11468_ = ~new_n10330_;
  assign new_n11469_ = ~new_n10327_;
  assign new_n11470_ = ~new_n10335_;
  assign new_n11471_ = ~new_n10354_;
  assign new_n11472_ = ~new_n10619_;
  assign new_n11473_ = ~new_n10295_;
  assign new_n11474_ = ~new_n10564_;
  assign new_n11475_ = ~new_n10565_;
  assign new_n11476_ = ~new_n10337_;
  assign new_n11477_ = ~new_n10563_;
  assign new_n11478_ = ~new_n10916_ | ~new_n9417_;
  assign new_n11479_ = ~new_n10588_;
  assign new_n11480_ = ~new_n10300_;
  assign new_n11481_ = ~new_n10584_;
  assign new_n11482_ = ~new_n10583_;
  assign new_n11483_ = ~new_n10579_;
  assign new_n11484_ = ~new_n10347_;
  assign new_n11485_ = ~new_n28821_;
  assign new_n11486_ = ~new_n11471_ | ~new_n10343_;
  assign new_n11487_ = ~new_n11502_ | ~new_n10587_;
  assign new_n11488_ = ~new_n29020_ | ~new_n9658_;
  assign new_n11489_ = ~new_n9408_ | ~new_n10331_;
  assign new_n11490_ = ~new_n10302_;
  assign new_n11491_ = ~new_n10301_;
  assign new_n11492_ = ~new_n10466_;
  assign new_n11493_ = ~new_n11223_ | ~new_n11479_;
  assign new_n11494_ = ~new_n10759_ | ~new_n11515_;
  assign new_n11495_ = ~new_n10343_ | ~new_n10325_ | ~new_n10311_ | ~pi0626;
  assign new_n11496_ = ~new_n10908_ | ~new_n9489_;
  assign new_n11497_ = ~new_n9487_ | ~new_n9400_;
  assign new_n11498_ = ~new_n9397_ | ~new_n10321_;
  assign new_n11499_ = ~new_n11419_ | ~new_n14618_;
  assign new_n11500_ = ~new_n10616_;
  assign new_n11501_ = ~new_n9479_ | ~new_n10336_;
  assign new_n11502_ = ~new_n10575_;
  assign new_n11503_ = ~new_n9415_ | ~new_n13609_;
  assign new_n11504_ = ~new_n11615_ | ~new_n10307_;
  assign new_n11505_ = ~new_n9489_ | ~new_n10333_;
  assign new_n11506_ = ~new_n11515_ | ~new_n2973_;
  assign new_n11507_ = ~new_n10344_;
  assign new_n11508_ = ~new_n10581_;
  assign new_n11509_ = ~new_n10345_;
  assign new_n11510_ = ~new_n10346_;
  assign new_n11511_ = ~new_n10917_ | ~new_n9417_;
  assign new_n11512_ = ~new_n10614_;
  assign new_n11513_ = ~new_n11457_ | ~new_n9417_ | ~new_n14912_;
  assign new_n11514_ = ~new_n10303_;
  assign new_n11515_ = ~new_n10342_;
  assign new_n11516_ = ~new_n10334_;
  assign new_n11517_ = ~new_n10322_;
  assign new_n11518_ = ~new_n10589_;
  assign new_n11519_ = ~pi0988 | ~new_n11491_;
  assign new_n11520_ = ~pi0987 | ~new_n11490_;
  assign new_n11521_ = ~pi0559 | ~new_n10300_;
  assign new_n11522_ = ~pi0987 | ~new_n11491_;
  assign new_n11523_ = ~pi0986 | ~new_n11490_;
  assign new_n11524_ = ~pi0560 | ~new_n10300_;
  assign new_n11525_ = ~pi0986 | ~new_n11491_;
  assign new_n11526_ = ~pi0985 | ~new_n11490_;
  assign new_n11527_ = ~pi0561 | ~new_n10300_;
  assign new_n11528_ = ~pi0985 | ~new_n11491_;
  assign new_n11529_ = ~pi0984 | ~new_n11490_;
  assign new_n11530_ = ~pi0562 | ~new_n10300_;
  assign new_n11531_ = ~pi0984 | ~new_n11491_;
  assign new_n11532_ = ~pi0983 | ~new_n11490_;
  assign new_n11533_ = ~pi0563 | ~new_n10300_;
  assign new_n11534_ = ~pi0983 | ~new_n11491_;
  assign new_n11535_ = ~pi0982 | ~new_n11490_;
  assign new_n11536_ = ~pi0564 | ~new_n10300_;
  assign new_n11537_ = ~pi0982 | ~new_n11491_;
  assign new_n11538_ = ~pi0981 | ~new_n11490_;
  assign new_n11539_ = ~pi0565 | ~new_n10300_;
  assign new_n11540_ = ~pi0981 | ~new_n11491_;
  assign new_n11541_ = ~pi0980 | ~new_n11490_;
  assign new_n11542_ = ~pi0566 | ~new_n10300_;
  assign new_n11543_ = ~pi0980 | ~new_n11491_;
  assign new_n11544_ = ~pi0979 | ~new_n11490_;
  assign new_n11545_ = ~pi0567 | ~new_n10300_;
  assign new_n11546_ = ~pi0979 | ~new_n11491_;
  assign new_n11547_ = ~pi0978 | ~new_n11490_;
  assign new_n11548_ = ~pi0568 | ~new_n10300_;
  assign new_n11549_ = ~pi0978 | ~new_n11491_;
  assign new_n11550_ = ~pi0977 | ~new_n11490_;
  assign new_n11551_ = ~pi0569 | ~new_n10300_;
  assign new_n11552_ = ~pi0977 | ~new_n11491_;
  assign new_n11553_ = ~pi0976 | ~new_n11490_;
  assign new_n11554_ = ~pi0570 | ~new_n10300_;
  assign new_n11555_ = ~pi0976 | ~new_n11491_;
  assign new_n11556_ = ~pi0975 | ~new_n11490_;
  assign new_n11557_ = ~pi0571 | ~new_n10300_;
  assign new_n11558_ = ~pi0975 | ~new_n11491_;
  assign new_n11559_ = ~pi0974 | ~new_n11490_;
  assign new_n11560_ = ~pi0572 | ~new_n10300_;
  assign new_n11561_ = ~pi0974 | ~new_n11491_;
  assign new_n11562_ = ~pi0973 | ~new_n11490_;
  assign new_n11563_ = ~pi0573 | ~new_n10300_;
  assign new_n11564_ = ~pi0973 | ~new_n11491_;
  assign new_n11565_ = ~pi0972 | ~new_n11490_;
  assign new_n11566_ = ~pi0574 | ~new_n10300_;
  assign new_n11567_ = ~pi0972 | ~new_n11491_;
  assign new_n11568_ = ~pi0971 | ~new_n11490_;
  assign new_n11569_ = ~pi0575 | ~new_n10300_;
  assign new_n11570_ = ~pi0971 | ~new_n11491_;
  assign new_n11571_ = ~pi0970 | ~new_n11490_;
  assign new_n11572_ = ~pi0576 | ~new_n10300_;
  assign new_n11573_ = ~pi0970 | ~new_n11491_;
  assign new_n11574_ = ~pi0969 | ~new_n11490_;
  assign new_n11575_ = ~pi0577 | ~new_n10300_;
  assign new_n11576_ = ~pi0969 | ~new_n11491_;
  assign new_n11577_ = ~pi0968 | ~new_n11490_;
  assign new_n11578_ = ~pi0578 | ~new_n10300_;
  assign new_n11579_ = ~pi0968 | ~new_n11491_;
  assign new_n11580_ = ~pi0967 | ~new_n11490_;
  assign new_n11581_ = ~pi0579 | ~new_n10300_;
  assign new_n11582_ = ~pi0967 | ~new_n11491_;
  assign new_n11583_ = ~pi0966 | ~new_n11490_;
  assign new_n11584_ = ~pi0580 | ~new_n10300_;
  assign new_n11585_ = ~pi0966 | ~new_n11491_;
  assign new_n11586_ = ~pi0965 | ~new_n11490_;
  assign new_n11587_ = ~pi0581 | ~new_n10300_;
  assign new_n11588_ = ~pi0965 | ~new_n11491_;
  assign new_n11589_ = ~pi0964 | ~new_n11490_;
  assign new_n11590_ = ~pi0582 | ~new_n10300_;
  assign new_n11591_ = ~pi0964 | ~new_n11491_;
  assign new_n11592_ = ~pi0963 | ~new_n11490_;
  assign new_n11593_ = ~pi0583 | ~new_n10300_;
  assign new_n11594_ = ~pi0963 | ~new_n11491_;
  assign new_n11595_ = ~pi0962 | ~new_n11490_;
  assign new_n11596_ = ~pi0584 | ~new_n10300_;
  assign new_n11597_ = ~pi0962 | ~new_n11491_;
  assign new_n11598_ = ~pi0961 | ~new_n11490_;
  assign new_n11599_ = ~pi0585 | ~new_n10300_;
  assign new_n11600_ = ~pi0961 | ~new_n11491_;
  assign new_n11601_ = ~pi0960 | ~new_n11490_;
  assign new_n11602_ = ~pi0586 | ~new_n10300_;
  assign new_n11603_ = ~pi0960 | ~new_n11491_;
  assign new_n11604_ = ~pi0959 | ~new_n11490_;
  assign new_n11605_ = ~pi0587 | ~new_n10300_;
  assign new_n11606_ = ~pi0959 | ~new_n11491_;
  assign new_n11607_ = ~pi0958 | ~new_n11490_;
  assign new_n11608_ = ~pi0588 | ~new_n10300_;
  assign new_n11609_ = ~new_n10308_;
  assign new_n11610_ = ~new_n11609_ | ~new_n10306_;
  assign new_n11611_ = ~pi0034 | ~new_n11514_;
  assign new_n11612_ = ~new_n10309_;
  assign new_n11613_ = ~new_n11612_ | ~new_n10306_;
  assign new_n11614_ = ~new_n11433_ | ~new_n14932_;
  assign new_n11615_ = ~new_n10304_;
  assign new_n11616_ = ~new_n11615_ | ~pi0033 | ~new_n10297_;
  assign new_n11617_ = ~new_n2973_ | ~pi0590 | ~new_n10309_;
  assign new_n11618_ = ~new_n11617_ | ~new_n11616_;
  assign new_n11619_ = ~new_n11618_ | ~pi0591 | ~new_n11611_;
  assign new_n11620_ = ~pi0589 | ~new_n11614_;
  assign new_n11621_ = ~pi0591 | ~new_n11451_;
  assign new_n11622_ = ~new_n11621_ | ~pi0589;
  assign new_n11623_ = ~new_n14933_ | ~new_n14951_ | ~new_n14950_;
  assign new_n11624_ = ~new_n2973_ | ~new_n11480_;
  assign new_n11625_ = ~new_n10733_ | ~new_n14934_;
  assign new_n11626_ = ~pi0589 | ~new_n10308_;
  assign new_n11627_ = ~pi0034 | ~new_n10307_;
  assign new_n11628_ = ~new_n11627_ | ~new_n11626_;
  assign new_n11629_ = ~new_n11628_ | ~new_n10299_;
  assign new_n11630_ = ~new_n11442_ | ~new_n10304_;
  assign new_n11631_ = ~new_n10318_;
  assign new_n11632_ = ~pi0760 | ~pi0759;
  assign new_n11633_ = ~new_n10315_;
  assign new_n11634_ = ~new_n10316_;
  assign new_n11635_ = ~pi0589 | ~new_n10299_;
  assign new_n11636_ = ~new_n10303_ | ~new_n11635_;
  assign new_n11637_ = ~new_n10568_;
  assign new_n11638_ = ~new_n10335_ | ~new_n10327_;
  assign new_n11639_ = ~new_n11638_ | ~new_n10306_;
  assign new_n11640_ = ~new_n9400_ | ~new_n10568_;
  assign new_n11641_ = ~new_n10332_;
  assign new_n11642_ = ~new_n10336_;
  assign new_n11643_ = ~new_n11465_ | ~new_n10294_;
  assign new_n11644_ = ~new_n10565_ | ~new_n11643_;
  assign new_n11645_ = ~new_n10564_ | ~new_n10563_;
  assign new_n11646_ = ~new_n29132_ | ~new_n11469_;
  assign new_n11647_ = ~new_n11458_ | ~new_n10328_;
  assign new_n11648_ = ~new_n11647_ | ~new_n11646_;
  assign new_n11649_ = ~new_n11461_ | ~new_n11648_;
  assign new_n11650_ = ~new_n11644_ | ~new_n10561_;
  assign new_n11651_ = ~new_n10298_;
  assign new_n11652_ = ~new_n11469_ | ~new_n10333_;
  assign new_n11653_ = ~new_n29402_ | ~new_n11458_;
  assign new_n11654_ = ~new_n11653_ | ~new_n11652_;
  assign new_n11655_ = ~new_n11461_ | ~new_n11654_;
  assign new_n11656_ = pi0995 | pi0994;
  assign new_n11657_ = ~new_n10339_;
  assign new_n11658_ = ~new_n11657_ | ~new_n10310_;
  assign new_n11659_ = ~new_n10752_ | ~new_n11466_;
  assign new_n11660_ = ~new_n10756_ | ~new_n15098_ | ~new_n15097_;
  assign new_n11661_ = ~new_n10340_;
  assign new_n11662_ = ~new_n11515_ | ~new_n10306_;
  assign new_n11663_ = ~pi0996 | ~new_n10325_;
  assign new_n11664_ = ~new_n11663_ | ~new_n11662_;
  assign new_n11665_ = ~pi0626 | ~new_n11664_;
  assign new_n11666_ = ~pi0625 | ~new_n10340_;
  assign new_n11667_ = ~new_n11660_ | ~new_n11506_;
  assign new_n11668_ = ~new_n10758_ | ~new_n11661_;
  assign new_n11669_ = ~pi0626 | ~new_n11667_;
  assign new_n11670_ = ~new_n9415_ | ~new_n11660_;
  assign new_n11671_ = ~new_n10760_ | ~new_n11510_;
  assign new_n11672_ = ~new_n11660_ | ~new_n11505_;
  assign new_n11673_ = ~new_n9415_ | ~new_n10339_;
  assign new_n11674_ = ~new_n10378_;
  assign new_n11675_ = ~new_n10392_;
  assign new_n11676_ = ~new_n10393_;
  assign new_n11677_ = ~new_n10360_;
  assign new_n11678_ = ~new_n10359_;
  assign new_n11679_ = ~new_n10419_;
  assign new_n11680_ = ~new_n28369_ | ~new_n10359_;
  assign new_n11681_ = ~new_n10467_;
  assign new_n11682_ = ~new_n10361_;
  assign new_n11683_ = ~new_n10352_;
  assign new_n11684_ = ~new_n10353_;
  assign new_n11685_ = ~new_n10465_;
  assign new_n11686_ = ~new_n10417_;
  assign new_n11687_ = ~pi0762 | ~new_n10352_;
  assign new_n11688_ = ~new_n10469_;
  assign new_n11689_ = ~new_n10390_;
  assign new_n11690_ = ~new_n10376_;
  assign new_n11691_ = ~new_n10284_;
  assign new_n11692_ = ~new_n9481_ | ~new_n9485_;
  assign new_n11693_ = ~new_n10366_;
  assign new_n11694_ = ~new_n10611_;
  assign new_n11695_ = ~new_n10367_;
  assign new_n11696_ = ~pi0626 | ~new_n10311_;
  assign new_n11697_ = ~new_n10346_ | ~new_n11696_ | ~new_n10345_;
  assign new_n11698_ = ~new_n11678_ | ~new_n9503_;
  assign new_n11699_ = ~new_n9509_ | ~new_n9403_;
  assign new_n11700_ = ~new_n11486_ | ~new_n11699_;
  assign new_n11701_ = ~new_n11693_ | ~new_n11700_;
  assign new_n11702_ = ~new_n11695_ | ~pi0625;
  assign new_n11703_ = ~pi0624 | ~new_n10353_;
  assign new_n11704_ = ~new_n11701_ | ~new_n10763_;
  assign new_n11705_ = ~new_n9509_ | ~new_n9439_;
  assign new_n11706_ = ~new_n11486_ | ~new_n11705_;
  assign new_n11707_ = ~new_n11706_ | ~new_n10366_;
  assign new_n11708_ = ~pi0625 | ~new_n10367_;
  assign new_n11709_ = ~new_n11708_ | ~new_n11707_;
  assign new_n11710_ = ~new_n9466_ | ~new_n11684_;
  assign new_n11711_ = ~new_n9463_ | ~new_n9504_;
  assign new_n11712_ = ~new_n9462_ | ~new_n11682_;
  assign new_n11713_ = ~new_n9447_ | ~new_n11709_;
  assign new_n11714_ = ~pi0628 | ~new_n11704_;
  assign new_n11715_ = ~new_n9467_ | ~new_n11684_;
  assign new_n11716_ = ~new_n9461_ | ~new_n9504_;
  assign new_n11717_ = ~new_n9460_ | ~new_n11682_;
  assign new_n11718_ = ~new_n9446_ | ~new_n11709_;
  assign new_n11719_ = ~pi0629 | ~new_n11704_;
  assign new_n11720_ = ~new_n9470_ | ~new_n11684_;
  assign new_n11721_ = ~new_n9459_ | ~new_n9504_;
  assign new_n11722_ = ~new_n9458_ | ~new_n11682_;
  assign new_n11723_ = ~new_n9445_ | ~new_n11709_;
  assign new_n11724_ = ~pi0630 | ~new_n11704_;
  assign new_n11725_ = ~new_n9465_ | ~new_n11684_;
  assign new_n11726_ = ~new_n9457_ | ~new_n9504_;
  assign new_n11727_ = ~new_n9456_ | ~new_n11682_;
  assign new_n11728_ = ~new_n9444_ | ~new_n11709_;
  assign new_n11729_ = ~pi0631 | ~new_n11704_;
  assign new_n11730_ = ~new_n9464_ | ~new_n11684_;
  assign new_n11731_ = ~new_n9455_ | ~new_n9504_;
  assign new_n11732_ = ~new_n9454_ | ~new_n11682_;
  assign new_n11733_ = ~new_n9443_ | ~new_n11709_;
  assign new_n11734_ = ~pi0632 | ~new_n11704_;
  assign new_n11735_ = ~new_n9473_ | ~new_n11684_;
  assign new_n11736_ = ~new_n9453_ | ~new_n9504_;
  assign new_n11737_ = ~new_n9452_ | ~new_n11682_;
  assign new_n11738_ = ~new_n9442_ | ~new_n11709_;
  assign new_n11739_ = ~pi0633 | ~new_n11704_;
  assign new_n11740_ = ~new_n9469_ | ~new_n11684_;
  assign new_n11741_ = ~new_n9451_ | ~new_n9504_;
  assign new_n11742_ = ~new_n9450_ | ~new_n11682_;
  assign new_n11743_ = ~new_n9441_ | ~new_n11709_;
  assign new_n11744_ = ~pi0634 | ~new_n11704_;
  assign new_n11745_ = ~new_n9472_ | ~new_n11684_;
  assign new_n11746_ = ~new_n9449_ | ~new_n9504_;
  assign new_n11747_ = ~new_n9448_ | ~new_n11682_;
  assign new_n11748_ = ~new_n9440_ | ~new_n11709_;
  assign new_n11749_ = ~pi0635 | ~new_n11704_;
  assign new_n11750_ = ~new_n10379_;
  assign new_n11751_ = ~new_n10380_;
  assign new_n11752_ = ~new_n10377_;
  assign new_n11753_ = ~new_n10286_;
  assign new_n11754_ = ~new_n10610_;
  assign new_n11755_ = ~new_n10381_;
  assign new_n11756_ = ~new_n11674_ | ~new_n9503_;
  assign new_n11757_ = ~new_n9512_ | ~new_n9403_;
  assign new_n11758_ = ~new_n11486_ | ~new_n11757_;
  assign new_n11759_ = ~new_n11758_ | ~new_n10286_;
  assign new_n11760_ = ~new_n11755_ | ~pi0625;
  assign new_n11761_ = ~pi0624 | ~new_n10377_;
  assign new_n11762_ = ~new_n11759_ | ~new_n10772_;
  assign new_n11763_ = ~new_n9512_ | ~new_n9439_;
  assign new_n11764_ = ~new_n11486_ | ~new_n11763_;
  assign new_n11765_ = ~new_n11764_ | ~new_n11753_;
  assign new_n11766_ = ~pi0625 | ~new_n10381_;
  assign new_n11767_ = ~new_n11766_ | ~new_n11765_;
  assign new_n11768_ = ~new_n11752_ | ~new_n9466_;
  assign new_n11769_ = ~new_n9510_ | ~new_n9463_;
  assign new_n11770_ = ~new_n11751_ | ~new_n9462_;
  assign new_n11771_ = ~new_n9447_ | ~new_n11767_;
  assign new_n11772_ = ~pi0636 | ~new_n11762_;
  assign new_n11773_ = ~new_n11752_ | ~new_n9467_;
  assign new_n11774_ = ~new_n9510_ | ~new_n9461_;
  assign new_n11775_ = ~new_n11751_ | ~new_n9460_;
  assign new_n11776_ = ~new_n9446_ | ~new_n11767_;
  assign new_n11777_ = ~pi0637 | ~new_n11762_;
  assign new_n11778_ = ~new_n11752_ | ~new_n9470_;
  assign new_n11779_ = ~new_n9510_ | ~new_n9459_;
  assign new_n11780_ = ~new_n11751_ | ~new_n9458_;
  assign new_n11781_ = ~new_n9445_ | ~new_n11767_;
  assign new_n11782_ = ~pi0638 | ~new_n11762_;
  assign new_n11783_ = ~new_n11752_ | ~new_n9465_;
  assign new_n11784_ = ~new_n9510_ | ~new_n9457_;
  assign new_n11785_ = ~new_n11751_ | ~new_n9456_;
  assign new_n11786_ = ~new_n9444_ | ~new_n11767_;
  assign new_n11787_ = ~pi0639 | ~new_n11762_;
  assign new_n11788_ = ~new_n11752_ | ~new_n9464_;
  assign new_n11789_ = ~new_n9510_ | ~new_n9455_;
  assign new_n11790_ = ~new_n11751_ | ~new_n9454_;
  assign new_n11791_ = ~new_n9443_ | ~new_n11767_;
  assign new_n11792_ = ~pi0640 | ~new_n11762_;
  assign new_n11793_ = ~new_n11752_ | ~new_n9473_;
  assign new_n11794_ = ~new_n9510_ | ~new_n9453_;
  assign new_n11795_ = ~new_n11751_ | ~new_n9452_;
  assign new_n11796_ = ~new_n9442_ | ~new_n11767_;
  assign new_n11797_ = ~pi0641 | ~new_n11762_;
  assign new_n11798_ = ~new_n11752_ | ~new_n9469_;
  assign new_n11799_ = ~new_n9510_ | ~new_n9451_;
  assign new_n11800_ = ~new_n11751_ | ~new_n9450_;
  assign new_n11801_ = ~new_n9441_ | ~new_n11767_;
  assign new_n11802_ = ~pi0642 | ~new_n11762_;
  assign new_n11803_ = ~new_n11752_ | ~new_n9472_;
  assign new_n11804_ = ~new_n9510_ | ~new_n9449_;
  assign new_n11805_ = ~new_n11751_ | ~new_n9448_;
  assign new_n11806_ = ~new_n9440_ | ~new_n11767_;
  assign new_n11807_ = ~pi0643 | ~new_n11762_;
  assign new_n11808_ = ~new_n10394_;
  assign new_n11809_ = ~new_n10395_;
  assign new_n11810_ = ~new_n10391_;
  assign new_n11811_ = ~new_n9486_ | ~new_n9481_;
  assign new_n11812_ = ~new_n10396_;
  assign new_n11813_ = ~new_n10609_;
  assign new_n11814_ = ~new_n10397_;
  assign new_n11815_ = ~new_n11675_ | ~new_n9503_;
  assign new_n11816_ = ~new_n9515_ | ~new_n9403_;
  assign new_n11817_ = ~new_n11486_ | ~new_n11816_;
  assign new_n11818_ = ~new_n11812_ | ~new_n11817_;
  assign new_n11819_ = ~new_n11814_ | ~pi0625;
  assign new_n11820_ = ~pi0624 | ~new_n10391_;
  assign new_n11821_ = ~new_n11818_ | ~new_n10781_;
  assign new_n11822_ = ~new_n9515_ | ~new_n9439_;
  assign new_n11823_ = ~new_n11486_ | ~new_n11822_;
  assign new_n11824_ = ~new_n11823_ | ~new_n10396_;
  assign new_n11825_ = ~pi0625 | ~new_n10397_;
  assign new_n11826_ = ~new_n11825_ | ~new_n11824_;
  assign new_n11827_ = ~new_n11810_ | ~new_n9466_;
  assign new_n11828_ = ~new_n9513_ | ~new_n9463_;
  assign new_n11829_ = ~new_n11809_ | ~new_n9462_;
  assign new_n11830_ = ~new_n9447_ | ~new_n11826_;
  assign new_n11831_ = ~pi0644 | ~new_n11821_;
  assign new_n11832_ = ~new_n11810_ | ~new_n9467_;
  assign new_n11833_ = ~new_n9513_ | ~new_n9461_;
  assign new_n11834_ = ~new_n11809_ | ~new_n9460_;
  assign new_n11835_ = ~new_n9446_ | ~new_n11826_;
  assign new_n11836_ = ~pi0645 | ~new_n11821_;
  assign new_n11837_ = ~new_n11810_ | ~new_n9470_;
  assign new_n11838_ = ~new_n9513_ | ~new_n9459_;
  assign new_n11839_ = ~new_n11809_ | ~new_n9458_;
  assign new_n11840_ = ~new_n9445_ | ~new_n11826_;
  assign new_n11841_ = ~pi0646 | ~new_n11821_;
  assign new_n11842_ = ~new_n11810_ | ~new_n9465_;
  assign new_n11843_ = ~new_n9513_ | ~new_n9457_;
  assign new_n11844_ = ~new_n11809_ | ~new_n9456_;
  assign new_n11845_ = ~new_n9444_ | ~new_n11826_;
  assign new_n11846_ = ~pi0647 | ~new_n11821_;
  assign new_n11847_ = ~new_n11810_ | ~new_n9464_;
  assign new_n11848_ = ~new_n9513_ | ~new_n9455_;
  assign new_n11849_ = ~new_n11809_ | ~new_n9454_;
  assign new_n11850_ = ~new_n9443_ | ~new_n11826_;
  assign new_n11851_ = ~pi0648 | ~new_n11821_;
  assign new_n11852_ = ~new_n11810_ | ~new_n9473_;
  assign new_n11853_ = ~new_n9513_ | ~new_n9453_;
  assign new_n11854_ = ~new_n11809_ | ~new_n9452_;
  assign new_n11855_ = ~new_n9442_ | ~new_n11826_;
  assign new_n11856_ = ~pi0649 | ~new_n11821_;
  assign new_n11857_ = ~new_n11810_ | ~new_n9469_;
  assign new_n11858_ = ~new_n9513_ | ~new_n9451_;
  assign new_n11859_ = ~new_n11809_ | ~new_n9450_;
  assign new_n11860_ = ~new_n9441_ | ~new_n11826_;
  assign new_n11861_ = ~pi0650 | ~new_n11821_;
  assign new_n11862_ = ~new_n11810_ | ~new_n9472_;
  assign new_n11863_ = ~new_n9513_ | ~new_n9449_;
  assign new_n11864_ = ~new_n11809_ | ~new_n9448_;
  assign new_n11865_ = ~new_n9440_ | ~new_n11826_;
  assign new_n11866_ = ~pi0651 | ~new_n11821_;
  assign new_n11867_ = ~new_n10407_;
  assign new_n11868_ = ~new_n10406_;
  assign new_n11869_ = ~new_n10287_;
  assign new_n11870_ = ~new_n10608_;
  assign new_n11871_ = ~new_n10408_;
  assign new_n11872_ = ~new_n9517_ | ~new_n9503_;
  assign new_n11873_ = ~new_n9521_ | ~new_n9403_;
  assign new_n11874_ = ~new_n11486_ | ~new_n11873_;
  assign new_n11875_ = ~new_n11874_ | ~new_n10287_;
  assign new_n11876_ = ~new_n11871_ | ~pi0625;
  assign new_n11877_ = ~pi0624 | ~new_n10406_;
  assign new_n11878_ = ~new_n11875_ | ~new_n10790_;
  assign new_n11879_ = ~new_n9521_ | ~new_n9439_;
  assign new_n11880_ = ~new_n11486_ | ~new_n11879_;
  assign new_n11881_ = ~new_n11880_ | ~new_n11869_;
  assign new_n11882_ = ~pi0625 | ~new_n10408_;
  assign new_n11883_ = ~new_n11882_ | ~new_n11881_;
  assign new_n11884_ = ~new_n11868_ | ~new_n9466_;
  assign new_n11885_ = ~new_n9518_ | ~new_n9463_;
  assign new_n11886_ = ~new_n11867_ | ~new_n9462_;
  assign new_n11887_ = ~new_n9447_ | ~new_n11883_;
  assign new_n11888_ = ~pi0652 | ~new_n11878_;
  assign new_n11889_ = ~new_n11868_ | ~new_n9467_;
  assign new_n11890_ = ~new_n9518_ | ~new_n9461_;
  assign new_n11891_ = ~new_n11867_ | ~new_n9460_;
  assign new_n11892_ = ~new_n9446_ | ~new_n11883_;
  assign new_n11893_ = ~pi0653 | ~new_n11878_;
  assign new_n11894_ = ~new_n11868_ | ~new_n9470_;
  assign new_n11895_ = ~new_n9518_ | ~new_n9459_;
  assign new_n11896_ = ~new_n11867_ | ~new_n9458_;
  assign new_n11897_ = ~new_n9445_ | ~new_n11883_;
  assign new_n11898_ = ~pi0654 | ~new_n11878_;
  assign new_n11899_ = ~new_n11868_ | ~new_n9465_;
  assign new_n11900_ = ~new_n9518_ | ~new_n9457_;
  assign new_n11901_ = ~new_n11867_ | ~new_n9456_;
  assign new_n11902_ = ~new_n9444_ | ~new_n11883_;
  assign new_n11903_ = ~pi0655 | ~new_n11878_;
  assign new_n11904_ = ~new_n11868_ | ~new_n9464_;
  assign new_n11905_ = ~new_n9518_ | ~new_n9455_;
  assign new_n11906_ = ~new_n11867_ | ~new_n9454_;
  assign new_n11907_ = ~new_n9443_ | ~new_n11883_;
  assign new_n11908_ = ~pi0656 | ~new_n11878_;
  assign new_n11909_ = ~new_n11868_ | ~new_n9473_;
  assign new_n11910_ = ~new_n9518_ | ~new_n9453_;
  assign new_n11911_ = ~new_n11867_ | ~new_n9452_;
  assign new_n11912_ = ~new_n9442_ | ~new_n11883_;
  assign new_n11913_ = ~pi0657 | ~new_n11878_;
  assign new_n11914_ = ~new_n11868_ | ~new_n9469_;
  assign new_n11915_ = ~new_n9518_ | ~new_n9451_;
  assign new_n11916_ = ~new_n11867_ | ~new_n9450_;
  assign new_n11917_ = ~new_n9441_ | ~new_n11883_;
  assign new_n11918_ = ~pi0658 | ~new_n11878_;
  assign new_n11919_ = ~new_n11868_ | ~new_n9472_;
  assign new_n11920_ = ~new_n9518_ | ~new_n9449_;
  assign new_n11921_ = ~new_n11867_ | ~new_n9448_;
  assign new_n11922_ = ~new_n9440_ | ~new_n11883_;
  assign new_n11923_ = ~pi0659 | ~new_n11878_;
  assign new_n11924_ = ~new_n10420_;
  assign new_n11925_ = ~new_n10418_;
  assign new_n11926_ = ~new_n9483_ | ~new_n9485_;
  assign new_n11927_ = ~new_n10421_;
  assign new_n11928_ = ~new_n10607_;
  assign new_n11929_ = ~new_n10422_;
  assign new_n11930_ = ~new_n11679_ | ~new_n11678_;
  assign new_n11931_ = ~new_n9525_ | ~new_n9403_;
  assign new_n11932_ = ~new_n11486_ | ~new_n11931_;
  assign new_n11933_ = ~new_n11927_ | ~new_n11932_;
  assign new_n11934_ = ~new_n11929_ | ~pi0625;
  assign new_n11935_ = ~pi0624 | ~new_n10418_;
  assign new_n11936_ = ~new_n11933_ | ~new_n10799_;
  assign new_n11937_ = ~new_n9525_ | ~new_n9439_;
  assign new_n11938_ = ~new_n11486_ | ~new_n11937_;
  assign new_n11939_ = ~new_n11938_ | ~new_n10421_;
  assign new_n11940_ = ~pi0625 | ~new_n10422_;
  assign new_n11941_ = ~new_n11940_ | ~new_n11939_;
  assign new_n11942_ = ~new_n11925_ | ~new_n9466_;
  assign new_n11943_ = ~new_n9523_ | ~new_n9463_;
  assign new_n11944_ = ~new_n11924_ | ~new_n9462_;
  assign new_n11945_ = ~new_n9447_ | ~new_n11941_;
  assign new_n11946_ = ~pi0660 | ~new_n11936_;
  assign new_n11947_ = ~new_n11925_ | ~new_n9467_;
  assign new_n11948_ = ~new_n9523_ | ~new_n9461_;
  assign new_n11949_ = ~new_n11924_ | ~new_n9460_;
  assign new_n11950_ = ~new_n9446_ | ~new_n11941_;
  assign new_n11951_ = ~pi0661 | ~new_n11936_;
  assign new_n11952_ = ~new_n11925_ | ~new_n9470_;
  assign new_n11953_ = ~new_n9523_ | ~new_n9459_;
  assign new_n11954_ = ~new_n11924_ | ~new_n9458_;
  assign new_n11955_ = ~new_n9445_ | ~new_n11941_;
  assign new_n11956_ = ~pi0662 | ~new_n11936_;
  assign new_n11957_ = ~new_n11925_ | ~new_n9465_;
  assign new_n11958_ = ~new_n9523_ | ~new_n9457_;
  assign new_n11959_ = ~new_n11924_ | ~new_n9456_;
  assign new_n11960_ = ~new_n9444_ | ~new_n11941_;
  assign new_n11961_ = ~pi0663 | ~new_n11936_;
  assign new_n11962_ = ~new_n11925_ | ~new_n9464_;
  assign new_n11963_ = ~new_n9523_ | ~new_n9455_;
  assign new_n11964_ = ~new_n11924_ | ~new_n9454_;
  assign new_n11965_ = ~new_n9443_ | ~new_n11941_;
  assign new_n11966_ = ~pi0664 | ~new_n11936_;
  assign new_n11967_ = ~new_n11925_ | ~new_n9473_;
  assign new_n11968_ = ~new_n9523_ | ~new_n9453_;
  assign new_n11969_ = ~new_n11924_ | ~new_n9452_;
  assign new_n11970_ = ~new_n9442_ | ~new_n11941_;
  assign new_n11971_ = ~pi0665 | ~new_n11936_;
  assign new_n11972_ = ~new_n11925_ | ~new_n9469_;
  assign new_n11973_ = ~new_n9523_ | ~new_n9451_;
  assign new_n11974_ = ~new_n11924_ | ~new_n9450_;
  assign new_n11975_ = ~new_n9441_ | ~new_n11941_;
  assign new_n11976_ = ~pi0666 | ~new_n11936_;
  assign new_n11977_ = ~new_n11925_ | ~new_n9472_;
  assign new_n11978_ = ~new_n9523_ | ~new_n9449_;
  assign new_n11979_ = ~new_n11924_ | ~new_n9448_;
  assign new_n11980_ = ~new_n9440_ | ~new_n11941_;
  assign new_n11981_ = ~pi0667 | ~new_n11936_;
  assign new_n11982_ = ~new_n10432_;
  assign new_n11983_ = ~new_n10431_;
  assign new_n11984_ = ~new_n10288_;
  assign new_n11985_ = ~new_n10606_;
  assign new_n11986_ = ~new_n10433_;
  assign new_n11987_ = ~new_n11679_ | ~new_n11674_;
  assign new_n11988_ = ~new_n9527_ | ~new_n9403_;
  assign new_n11989_ = ~new_n11486_ | ~new_n11988_;
  assign new_n11990_ = ~new_n11989_ | ~new_n10288_;
  assign new_n11991_ = ~new_n11986_ | ~pi0625;
  assign new_n11992_ = ~pi0624 | ~new_n10431_;
  assign new_n11993_ = ~new_n11990_ | ~new_n10808_;
  assign new_n11994_ = ~new_n9527_ | ~new_n9439_;
  assign new_n11995_ = ~new_n11486_ | ~new_n11994_;
  assign new_n11996_ = ~new_n11995_ | ~new_n11984_;
  assign new_n11997_ = ~pi0625 | ~new_n10433_;
  assign new_n11998_ = ~new_n11997_ | ~new_n11996_;
  assign new_n11999_ = ~new_n11983_ | ~new_n9466_;
  assign new_n12000_ = ~new_n9526_ | ~new_n9463_;
  assign new_n12001_ = ~new_n11982_ | ~new_n9462_;
  assign new_n12002_ = ~new_n9447_ | ~new_n11998_;
  assign new_n12003_ = ~pi0668 | ~new_n11993_;
  assign new_n12004_ = ~new_n11983_ | ~new_n9467_;
  assign new_n12005_ = ~new_n9526_ | ~new_n9461_;
  assign new_n12006_ = ~new_n11982_ | ~new_n9460_;
  assign new_n12007_ = ~new_n9446_ | ~new_n11998_;
  assign new_n12008_ = ~pi0669 | ~new_n11993_;
  assign new_n12009_ = ~new_n11983_ | ~new_n9470_;
  assign new_n12010_ = ~new_n9526_ | ~new_n9459_;
  assign new_n12011_ = ~new_n11982_ | ~new_n9458_;
  assign new_n12012_ = ~new_n9445_ | ~new_n11998_;
  assign new_n12013_ = ~pi0670 | ~new_n11993_;
  assign new_n12014_ = ~new_n11983_ | ~new_n9465_;
  assign new_n12015_ = ~new_n9526_ | ~new_n9457_;
  assign new_n12016_ = ~new_n11982_ | ~new_n9456_;
  assign new_n12017_ = ~new_n9444_ | ~new_n11998_;
  assign new_n12018_ = ~pi0671 | ~new_n11993_;
  assign new_n12019_ = ~new_n11983_ | ~new_n9464_;
  assign new_n12020_ = ~new_n9526_ | ~new_n9455_;
  assign new_n12021_ = ~new_n11982_ | ~new_n9454_;
  assign new_n12022_ = ~new_n9443_ | ~new_n11998_;
  assign new_n12023_ = ~pi0672 | ~new_n11993_;
  assign new_n12024_ = ~new_n11983_ | ~new_n9473_;
  assign new_n12025_ = ~new_n9526_ | ~new_n9453_;
  assign new_n12026_ = ~new_n11982_ | ~new_n9452_;
  assign new_n12027_ = ~new_n9442_ | ~new_n11998_;
  assign new_n12028_ = ~pi0673 | ~new_n11993_;
  assign new_n12029_ = ~new_n11983_ | ~new_n9469_;
  assign new_n12030_ = ~new_n9526_ | ~new_n9451_;
  assign new_n12031_ = ~new_n11982_ | ~new_n9450_;
  assign new_n12032_ = ~new_n9441_ | ~new_n11998_;
  assign new_n12033_ = ~pi0674 | ~new_n11993_;
  assign new_n12034_ = ~new_n11983_ | ~new_n9472_;
  assign new_n12035_ = ~new_n9526_ | ~new_n9449_;
  assign new_n12036_ = ~new_n11982_ | ~new_n9448_;
  assign new_n12037_ = ~new_n9440_ | ~new_n11998_;
  assign new_n12038_ = ~pi0675 | ~new_n11993_;
  assign new_n12039_ = ~new_n10443_;
  assign new_n12040_ = ~new_n10442_;
  assign new_n12041_ = ~new_n9483_ | ~new_n9486_;
  assign new_n12042_ = ~new_n10444_;
  assign new_n12043_ = ~new_n10605_;
  assign new_n12044_ = ~new_n10445_;
  assign new_n12045_ = ~new_n11679_ | ~new_n11675_;
  assign new_n12046_ = ~new_n9529_ | ~new_n9403_;
  assign new_n12047_ = ~new_n11486_ | ~new_n12046_;
  assign new_n12048_ = ~new_n12042_ | ~new_n12047_;
  assign new_n12049_ = ~new_n12044_ | ~pi0625;
  assign new_n12050_ = ~pi0624 | ~new_n10442_;
  assign new_n12051_ = ~new_n12048_ | ~new_n10817_;
  assign new_n12052_ = ~new_n9529_ | ~new_n9439_;
  assign new_n12053_ = ~new_n11486_ | ~new_n12052_;
  assign new_n12054_ = ~new_n12053_ | ~new_n10444_;
  assign new_n12055_ = ~pi0625 | ~new_n10445_;
  assign new_n12056_ = ~new_n12055_ | ~new_n12054_;
  assign new_n12057_ = ~new_n12040_ | ~new_n9466_;
  assign new_n12058_ = ~new_n9528_ | ~new_n9463_;
  assign new_n12059_ = ~new_n12039_ | ~new_n9462_;
  assign new_n12060_ = ~new_n9447_ | ~new_n12056_;
  assign new_n12061_ = ~pi0676 | ~new_n12051_;
  assign new_n12062_ = ~new_n12040_ | ~new_n9467_;
  assign new_n12063_ = ~new_n9528_ | ~new_n9461_;
  assign new_n12064_ = ~new_n12039_ | ~new_n9460_;
  assign new_n12065_ = ~new_n9446_ | ~new_n12056_;
  assign new_n12066_ = ~pi0677 | ~new_n12051_;
  assign new_n12067_ = ~new_n12040_ | ~new_n9470_;
  assign new_n12068_ = ~new_n9528_ | ~new_n9459_;
  assign new_n12069_ = ~new_n12039_ | ~new_n9458_;
  assign new_n12070_ = ~new_n9445_ | ~new_n12056_;
  assign new_n12071_ = ~pi0678 | ~new_n12051_;
  assign new_n12072_ = ~new_n12040_ | ~new_n9465_;
  assign new_n12073_ = ~new_n9528_ | ~new_n9457_;
  assign new_n12074_ = ~new_n12039_ | ~new_n9456_;
  assign new_n12075_ = ~new_n9444_ | ~new_n12056_;
  assign new_n12076_ = ~pi0679 | ~new_n12051_;
  assign new_n12077_ = ~new_n12040_ | ~new_n9464_;
  assign new_n12078_ = ~new_n9528_ | ~new_n9455_;
  assign new_n12079_ = ~new_n12039_ | ~new_n9454_;
  assign new_n12080_ = ~new_n9443_ | ~new_n12056_;
  assign new_n12081_ = ~pi0680 | ~new_n12051_;
  assign new_n12082_ = ~new_n12040_ | ~new_n9473_;
  assign new_n12083_ = ~new_n9528_ | ~new_n9453_;
  assign new_n12084_ = ~new_n12039_ | ~new_n9452_;
  assign new_n12085_ = ~new_n9442_ | ~new_n12056_;
  assign new_n12086_ = ~pi0681 | ~new_n12051_;
  assign new_n12087_ = ~new_n12040_ | ~new_n9469_;
  assign new_n12088_ = ~new_n9528_ | ~new_n9451_;
  assign new_n12089_ = ~new_n12039_ | ~new_n9450_;
  assign new_n12090_ = ~new_n9441_ | ~new_n12056_;
  assign new_n12091_ = ~pi0682 | ~new_n12051_;
  assign new_n12092_ = ~new_n12040_ | ~new_n9472_;
  assign new_n12093_ = ~new_n9528_ | ~new_n9449_;
  assign new_n12094_ = ~new_n12039_ | ~new_n9448_;
  assign new_n12095_ = ~new_n9440_ | ~new_n12056_;
  assign new_n12096_ = ~pi0683 | ~new_n12051_;
  assign new_n12097_ = ~new_n10455_;
  assign new_n12098_ = ~new_n10454_;
  assign new_n12099_ = ~new_n10289_;
  assign new_n12100_ = ~new_n10604_;
  assign new_n12101_ = ~new_n10456_;
  assign new_n12102_ = ~new_n11679_ | ~new_n9517_;
  assign new_n12103_ = ~new_n9531_ | ~new_n9403_;
  assign new_n12104_ = ~new_n11486_ | ~new_n12103_;
  assign new_n12105_ = ~new_n12104_ | ~new_n10289_;
  assign new_n12106_ = ~new_n12101_ | ~pi0625;
  assign new_n12107_ = ~pi0624 | ~new_n10454_;
  assign new_n12108_ = ~new_n12105_ | ~new_n10826_;
  assign new_n12109_ = ~new_n9531_ | ~new_n9439_;
  assign new_n12110_ = ~new_n11486_ | ~new_n12109_;
  assign new_n12111_ = ~new_n12110_ | ~new_n12099_;
  assign new_n12112_ = ~pi0625 | ~new_n10456_;
  assign new_n12113_ = ~new_n12112_ | ~new_n12111_;
  assign new_n12114_ = ~new_n12098_ | ~new_n9466_;
  assign new_n12115_ = ~new_n9530_ | ~new_n9463_;
  assign new_n12116_ = ~new_n12097_ | ~new_n9462_;
  assign new_n12117_ = ~new_n9447_ | ~new_n12113_;
  assign new_n12118_ = ~pi0684 | ~new_n12108_;
  assign new_n12119_ = ~new_n12098_ | ~new_n9467_;
  assign new_n12120_ = ~new_n9530_ | ~new_n9461_;
  assign new_n12121_ = ~new_n12097_ | ~new_n9460_;
  assign new_n12122_ = ~new_n9446_ | ~new_n12113_;
  assign new_n12123_ = ~pi0685 | ~new_n12108_;
  assign new_n12124_ = ~new_n12098_ | ~new_n9470_;
  assign new_n12125_ = ~new_n9530_ | ~new_n9459_;
  assign new_n12126_ = ~new_n12097_ | ~new_n9458_;
  assign new_n12127_ = ~new_n9445_ | ~new_n12113_;
  assign new_n12128_ = ~pi0686 | ~new_n12108_;
  assign new_n12129_ = ~new_n12098_ | ~new_n9465_;
  assign new_n12130_ = ~new_n9530_ | ~new_n9457_;
  assign new_n12131_ = ~new_n12097_ | ~new_n9456_;
  assign new_n12132_ = ~new_n9444_ | ~new_n12113_;
  assign new_n12133_ = ~pi0687 | ~new_n12108_;
  assign new_n12134_ = ~new_n12098_ | ~new_n9464_;
  assign new_n12135_ = ~new_n9530_ | ~new_n9455_;
  assign new_n12136_ = ~new_n12097_ | ~new_n9454_;
  assign new_n12137_ = ~new_n9443_ | ~new_n12113_;
  assign new_n12138_ = ~pi0688 | ~new_n12108_;
  assign new_n12139_ = ~new_n12098_ | ~new_n9473_;
  assign new_n12140_ = ~new_n9530_ | ~new_n9453_;
  assign new_n12141_ = ~new_n12097_ | ~new_n9452_;
  assign new_n12142_ = ~new_n9442_ | ~new_n12113_;
  assign new_n12143_ = ~pi0689 | ~new_n12108_;
  assign new_n12144_ = ~new_n12098_ | ~new_n9469_;
  assign new_n12145_ = ~new_n9530_ | ~new_n9451_;
  assign new_n12146_ = ~new_n12097_ | ~new_n9450_;
  assign new_n12147_ = ~new_n9441_ | ~new_n12113_;
  assign new_n12148_ = ~pi0690 | ~new_n12108_;
  assign new_n12149_ = ~new_n12098_ | ~new_n9472_;
  assign new_n12150_ = ~new_n9530_ | ~new_n9449_;
  assign new_n12151_ = ~new_n12097_ | ~new_n9448_;
  assign new_n12152_ = ~new_n9440_ | ~new_n12113_;
  assign new_n12153_ = ~pi0691 | ~new_n12108_;
  assign new_n12154_ = ~new_n10468_;
  assign new_n12155_ = ~new_n9482_ | ~new_n9485_;
  assign new_n12156_ = ~new_n10470_;
  assign new_n12157_ = ~new_n10603_;
  assign new_n12158_ = ~new_n10471_;
  assign new_n12159_ = ~new_n9534_ | ~new_n9403_;
  assign new_n12160_ = ~new_n11486_ | ~new_n12159_;
  assign new_n12161_ = ~new_n12156_ | ~new_n12160_;
  assign new_n12162_ = ~new_n12158_ | ~pi0625;
  assign new_n12163_ = ~pi0624 | ~new_n10465_;
  assign new_n12164_ = ~new_n12161_ | ~new_n10835_;
  assign new_n12165_ = ~new_n9534_ | ~new_n9439_;
  assign new_n12166_ = ~new_n11486_ | ~new_n12165_;
  assign new_n12167_ = ~new_n12166_ | ~new_n10470_;
  assign new_n12168_ = ~pi0625 | ~new_n10471_;
  assign new_n12169_ = ~new_n12168_ | ~new_n12167_;
  assign new_n12170_ = ~new_n11685_ | ~new_n9466_;
  assign new_n12171_ = ~new_n11492_ | ~new_n9463_;
  assign new_n12172_ = ~new_n12154_ | ~new_n9462_;
  assign new_n12173_ = ~new_n9447_ | ~new_n12169_;
  assign new_n12174_ = ~pi0692 | ~new_n12164_;
  assign new_n12175_ = ~new_n11685_ | ~new_n9467_;
  assign new_n12176_ = ~new_n11492_ | ~new_n9461_;
  assign new_n12177_ = ~new_n12154_ | ~new_n9460_;
  assign new_n12178_ = ~new_n9446_ | ~new_n12169_;
  assign new_n12179_ = ~pi0693 | ~new_n12164_;
  assign new_n12180_ = ~new_n11685_ | ~new_n9470_;
  assign new_n12181_ = ~new_n11492_ | ~new_n9459_;
  assign new_n12182_ = ~new_n12154_ | ~new_n9458_;
  assign new_n12183_ = ~new_n9445_ | ~new_n12169_;
  assign new_n12184_ = ~pi0694 | ~new_n12164_;
  assign new_n12185_ = ~new_n11685_ | ~new_n9465_;
  assign new_n12186_ = ~new_n11492_ | ~new_n9457_;
  assign new_n12187_ = ~new_n12154_ | ~new_n9456_;
  assign new_n12188_ = ~new_n9444_ | ~new_n12169_;
  assign new_n12189_ = ~pi0695 | ~new_n12164_;
  assign new_n12190_ = ~new_n11685_ | ~new_n9464_;
  assign new_n12191_ = ~new_n11492_ | ~new_n9455_;
  assign new_n12192_ = ~new_n12154_ | ~new_n9454_;
  assign new_n12193_ = ~new_n9443_ | ~new_n12169_;
  assign new_n12194_ = ~pi0696 | ~new_n12164_;
  assign new_n12195_ = ~new_n11685_ | ~new_n9473_;
  assign new_n12196_ = ~new_n11492_ | ~new_n9453_;
  assign new_n12197_ = ~new_n12154_ | ~new_n9452_;
  assign new_n12198_ = ~new_n9442_ | ~new_n12169_;
  assign new_n12199_ = ~pi0697 | ~new_n12164_;
  assign new_n12200_ = ~new_n11685_ | ~new_n9469_;
  assign new_n12201_ = ~new_n11492_ | ~new_n9451_;
  assign new_n12202_ = ~new_n12154_ | ~new_n9450_;
  assign new_n12203_ = ~new_n9441_ | ~new_n12169_;
  assign new_n12204_ = ~pi0698 | ~new_n12164_;
  assign new_n12205_ = ~new_n11685_ | ~new_n9472_;
  assign new_n12206_ = ~new_n11492_ | ~new_n9449_;
  assign new_n12207_ = ~new_n12154_ | ~new_n9448_;
  assign new_n12208_ = ~new_n9440_ | ~new_n12169_;
  assign new_n12209_ = ~pi0699 | ~new_n12164_;
  assign new_n12210_ = ~new_n10481_;
  assign new_n12211_ = ~new_n10480_;
  assign new_n12212_ = ~new_n10290_;
  assign new_n12213_ = ~new_n10602_;
  assign new_n12214_ = ~new_n10482_;
  assign new_n12215_ = ~new_n11674_ | ~new_n9501_;
  assign new_n12216_ = ~new_n9536_ | ~new_n9403_;
  assign new_n12217_ = ~new_n11486_ | ~new_n12216_;
  assign new_n12218_ = ~new_n12217_ | ~new_n10290_;
  assign new_n12219_ = ~new_n12214_ | ~pi0625;
  assign new_n12220_ = ~pi0624 | ~new_n10480_;
  assign new_n12221_ = ~new_n12218_ | ~new_n10844_;
  assign new_n12222_ = ~new_n9536_ | ~new_n9439_;
  assign new_n12223_ = ~new_n11486_ | ~new_n12222_;
  assign new_n12224_ = ~new_n12223_ | ~new_n12212_;
  assign new_n12225_ = ~pi0625 | ~new_n10482_;
  assign new_n12226_ = ~new_n12225_ | ~new_n12224_;
  assign new_n12227_ = ~new_n12211_ | ~new_n9466_;
  assign new_n12228_ = ~new_n9535_ | ~new_n9463_;
  assign new_n12229_ = ~new_n12210_ | ~new_n9462_;
  assign new_n12230_ = ~new_n9447_ | ~new_n12226_;
  assign new_n12231_ = ~pi0700 | ~new_n12221_;
  assign new_n12232_ = ~new_n12211_ | ~new_n9467_;
  assign new_n12233_ = ~new_n9535_ | ~new_n9461_;
  assign new_n12234_ = ~new_n12210_ | ~new_n9460_;
  assign new_n12235_ = ~new_n9446_ | ~new_n12226_;
  assign new_n12236_ = ~pi0701 | ~new_n12221_;
  assign new_n12237_ = ~new_n12211_ | ~new_n9470_;
  assign new_n12238_ = ~new_n9535_ | ~new_n9459_;
  assign new_n12239_ = ~new_n12210_ | ~new_n9458_;
  assign new_n12240_ = ~new_n9445_ | ~new_n12226_;
  assign new_n12241_ = ~pi0702 | ~new_n12221_;
  assign new_n12242_ = ~new_n12211_ | ~new_n9465_;
  assign new_n12243_ = ~new_n9535_ | ~new_n9457_;
  assign new_n12244_ = ~new_n12210_ | ~new_n9456_;
  assign new_n12245_ = ~new_n9444_ | ~new_n12226_;
  assign new_n12246_ = ~pi0703 | ~new_n12221_;
  assign new_n12247_ = ~new_n12211_ | ~new_n9464_;
  assign new_n12248_ = ~new_n9535_ | ~new_n9455_;
  assign new_n12249_ = ~new_n12210_ | ~new_n9454_;
  assign new_n12250_ = ~new_n9443_ | ~new_n12226_;
  assign new_n12251_ = ~pi0704 | ~new_n12221_;
  assign new_n12252_ = ~new_n12211_ | ~new_n9473_;
  assign new_n12253_ = ~new_n9535_ | ~new_n9453_;
  assign new_n12254_ = ~new_n12210_ | ~new_n9452_;
  assign new_n12255_ = ~new_n9442_ | ~new_n12226_;
  assign new_n12256_ = ~pi0705 | ~new_n12221_;
  assign new_n12257_ = ~new_n12211_ | ~new_n9469_;
  assign new_n12258_ = ~new_n9535_ | ~new_n9451_;
  assign new_n12259_ = ~new_n12210_ | ~new_n9450_;
  assign new_n12260_ = ~new_n9441_ | ~new_n12226_;
  assign new_n12261_ = ~pi0706 | ~new_n12221_;
  assign new_n12262_ = ~new_n12211_ | ~new_n9472_;
  assign new_n12263_ = ~new_n9535_ | ~new_n9449_;
  assign new_n12264_ = ~new_n12210_ | ~new_n9448_;
  assign new_n12265_ = ~new_n9440_ | ~new_n12226_;
  assign new_n12266_ = ~pi0707 | ~new_n12221_;
  assign new_n12267_ = ~new_n10492_;
  assign new_n12268_ = ~new_n10491_;
  assign new_n12269_ = ~new_n9482_ | ~new_n9486_;
  assign new_n12270_ = ~new_n10493_;
  assign new_n12271_ = ~new_n10601_;
  assign new_n12272_ = ~new_n10494_;
  assign new_n12273_ = ~new_n11675_ | ~new_n9501_;
  assign new_n12274_ = ~new_n9538_ | ~new_n9403_;
  assign new_n12275_ = ~new_n11486_ | ~new_n12274_;
  assign new_n12276_ = ~new_n12270_ | ~new_n12275_;
  assign new_n12277_ = ~new_n12272_ | ~pi0625;
  assign new_n12278_ = ~pi0624 | ~new_n10491_;
  assign new_n12279_ = ~new_n12276_ | ~new_n10853_;
  assign new_n12280_ = ~new_n9538_ | ~new_n9439_;
  assign new_n12281_ = ~new_n11486_ | ~new_n12280_;
  assign new_n12282_ = ~new_n12281_ | ~new_n10493_;
  assign new_n12283_ = ~pi0625 | ~new_n10494_;
  assign new_n12284_ = ~new_n12283_ | ~new_n12282_;
  assign new_n12285_ = ~new_n12268_ | ~new_n9466_;
  assign new_n12286_ = ~new_n9537_ | ~new_n9463_;
  assign new_n12287_ = ~new_n12267_ | ~new_n9462_;
  assign new_n12288_ = ~new_n9447_ | ~new_n12284_;
  assign new_n12289_ = ~pi0708 | ~new_n12279_;
  assign new_n12290_ = ~new_n12268_ | ~new_n9467_;
  assign new_n12291_ = ~new_n9537_ | ~new_n9461_;
  assign new_n12292_ = ~new_n12267_ | ~new_n9460_;
  assign new_n12293_ = ~new_n9446_ | ~new_n12284_;
  assign new_n12294_ = ~pi0709 | ~new_n12279_;
  assign new_n12295_ = ~new_n12268_ | ~new_n9470_;
  assign new_n12296_ = ~new_n9537_ | ~new_n9459_;
  assign new_n12297_ = ~new_n12267_ | ~new_n9458_;
  assign new_n12298_ = ~new_n9445_ | ~new_n12284_;
  assign new_n12299_ = ~pi0710 | ~new_n12279_;
  assign new_n12300_ = ~new_n12268_ | ~new_n9465_;
  assign new_n12301_ = ~new_n9537_ | ~new_n9457_;
  assign new_n12302_ = ~new_n12267_ | ~new_n9456_;
  assign new_n12303_ = ~new_n9444_ | ~new_n12284_;
  assign new_n12304_ = ~pi0711 | ~new_n12279_;
  assign new_n12305_ = ~new_n12268_ | ~new_n9464_;
  assign new_n12306_ = ~new_n9537_ | ~new_n9455_;
  assign new_n12307_ = ~new_n12267_ | ~new_n9454_;
  assign new_n12308_ = ~new_n9443_ | ~new_n12284_;
  assign new_n12309_ = ~pi0712 | ~new_n12279_;
  assign new_n12310_ = ~new_n12268_ | ~new_n9473_;
  assign new_n12311_ = ~new_n9537_ | ~new_n9453_;
  assign new_n12312_ = ~new_n12267_ | ~new_n9452_;
  assign new_n12313_ = ~new_n9442_ | ~new_n12284_;
  assign new_n12314_ = ~pi0713 | ~new_n12279_;
  assign new_n12315_ = ~new_n12268_ | ~new_n9469_;
  assign new_n12316_ = ~new_n9537_ | ~new_n9451_;
  assign new_n12317_ = ~new_n12267_ | ~new_n9450_;
  assign new_n12318_ = ~new_n9441_ | ~new_n12284_;
  assign new_n12319_ = ~pi0714 | ~new_n12279_;
  assign new_n12320_ = ~new_n12268_ | ~new_n9472_;
  assign new_n12321_ = ~new_n9537_ | ~new_n9449_;
  assign new_n12322_ = ~new_n12267_ | ~new_n9448_;
  assign new_n12323_ = ~new_n9440_ | ~new_n12284_;
  assign new_n12324_ = ~pi0715 | ~new_n12279_;
  assign new_n12325_ = ~new_n10504_;
  assign new_n12326_ = ~new_n10503_;
  assign new_n12327_ = ~new_n10291_;
  assign new_n12328_ = ~new_n10600_;
  assign new_n12329_ = ~new_n10505_;
  assign new_n12330_ = ~new_n9517_ | ~new_n9501_;
  assign new_n12331_ = ~new_n9540_ | ~new_n9403_;
  assign new_n12332_ = ~new_n11486_ | ~new_n12331_;
  assign new_n12333_ = ~new_n12332_ | ~new_n10291_;
  assign new_n12334_ = ~new_n12329_ | ~pi0625;
  assign new_n12335_ = ~pi0624 | ~new_n10503_;
  assign new_n12336_ = ~new_n12333_ | ~new_n10862_;
  assign new_n12337_ = ~new_n9540_ | ~new_n9439_;
  assign new_n12338_ = ~new_n11486_ | ~new_n12337_;
  assign new_n12339_ = ~new_n12338_ | ~new_n12327_;
  assign new_n12340_ = ~pi0625 | ~new_n10505_;
  assign new_n12341_ = ~new_n12340_ | ~new_n12339_;
  assign new_n12342_ = ~new_n12326_ | ~new_n9466_;
  assign new_n12343_ = ~new_n9539_ | ~new_n9463_;
  assign new_n12344_ = ~new_n12325_ | ~new_n9462_;
  assign new_n12345_ = ~new_n9447_ | ~new_n12341_;
  assign new_n12346_ = ~pi0716 | ~new_n12336_;
  assign new_n12347_ = ~new_n12326_ | ~new_n9467_;
  assign new_n12348_ = ~new_n9539_ | ~new_n9461_;
  assign new_n12349_ = ~new_n12325_ | ~new_n9460_;
  assign new_n12350_ = ~new_n9446_ | ~new_n12341_;
  assign new_n12351_ = ~pi0717 | ~new_n12336_;
  assign new_n12352_ = ~new_n12326_ | ~new_n9470_;
  assign new_n12353_ = ~new_n9539_ | ~new_n9459_;
  assign new_n12354_ = ~new_n12325_ | ~new_n9458_;
  assign new_n12355_ = ~new_n9445_ | ~new_n12341_;
  assign new_n12356_ = ~pi0718 | ~new_n12336_;
  assign new_n12357_ = ~new_n12326_ | ~new_n9465_;
  assign new_n12358_ = ~new_n9539_ | ~new_n9457_;
  assign new_n12359_ = ~new_n12325_ | ~new_n9456_;
  assign new_n12360_ = ~new_n9444_ | ~new_n12341_;
  assign new_n12361_ = ~pi0719 | ~new_n12336_;
  assign new_n12362_ = ~new_n12326_ | ~new_n9464_;
  assign new_n12363_ = ~new_n9539_ | ~new_n9455_;
  assign new_n12364_ = ~new_n12325_ | ~new_n9454_;
  assign new_n12365_ = ~new_n9443_ | ~new_n12341_;
  assign new_n12366_ = ~pi0720 | ~new_n12336_;
  assign new_n12367_ = ~new_n12326_ | ~new_n9473_;
  assign new_n12368_ = ~new_n9539_ | ~new_n9453_;
  assign new_n12369_ = ~new_n12325_ | ~new_n9452_;
  assign new_n12370_ = ~new_n9442_ | ~new_n12341_;
  assign new_n12371_ = ~pi0721 | ~new_n12336_;
  assign new_n12372_ = ~new_n12326_ | ~new_n9469_;
  assign new_n12373_ = ~new_n9539_ | ~new_n9451_;
  assign new_n12374_ = ~new_n12325_ | ~new_n9450_;
  assign new_n12375_ = ~new_n9441_ | ~new_n12341_;
  assign new_n12376_ = ~pi0722 | ~new_n12336_;
  assign new_n12377_ = ~new_n12326_ | ~new_n9472_;
  assign new_n12378_ = ~new_n9539_ | ~new_n9449_;
  assign new_n12379_ = ~new_n12325_ | ~new_n9448_;
  assign new_n12380_ = ~new_n9440_ | ~new_n12341_;
  assign new_n12381_ = ~pi0723 | ~new_n12336_;
  assign new_n12382_ = ~new_n10515_;
  assign new_n12383_ = ~new_n10514_;
  assign new_n12384_ = ~new_n9484_ | ~new_n9485_;
  assign new_n12385_ = ~new_n10516_;
  assign new_n12386_ = ~new_n10599_;
  assign new_n12387_ = ~new_n10517_;
  assign new_n12388_ = ~new_n9542_ | ~new_n11678_;
  assign new_n12389_ = ~new_n9546_ | ~new_n9403_;
  assign new_n12390_ = ~new_n11486_ | ~new_n12389_;
  assign new_n12391_ = ~new_n12385_ | ~new_n12390_;
  assign new_n12392_ = ~new_n12387_ | ~pi0625;
  assign new_n12393_ = ~pi0624 | ~new_n10514_;
  assign new_n12394_ = ~new_n12391_ | ~new_n10871_;
  assign new_n12395_ = ~new_n9546_ | ~new_n9439_;
  assign new_n12396_ = ~new_n11486_ | ~new_n12395_;
  assign new_n12397_ = ~new_n12396_ | ~new_n10516_;
  assign new_n12398_ = ~pi0625 | ~new_n10517_;
  assign new_n12399_ = ~new_n12398_ | ~new_n12397_;
  assign new_n12400_ = ~new_n12383_ | ~new_n9466_;
  assign new_n12401_ = ~new_n9543_ | ~new_n9463_;
  assign new_n12402_ = ~new_n12382_ | ~new_n9462_;
  assign new_n12403_ = ~new_n9447_ | ~new_n12399_;
  assign new_n12404_ = ~pi0724 | ~new_n12394_;
  assign new_n12405_ = ~new_n12383_ | ~new_n9467_;
  assign new_n12406_ = ~new_n9543_ | ~new_n9461_;
  assign new_n12407_ = ~new_n12382_ | ~new_n9460_;
  assign new_n12408_ = ~new_n9446_ | ~new_n12399_;
  assign new_n12409_ = ~pi0725 | ~new_n12394_;
  assign new_n12410_ = ~new_n12383_ | ~new_n9470_;
  assign new_n12411_ = ~new_n9543_ | ~new_n9459_;
  assign new_n12412_ = ~new_n12382_ | ~new_n9458_;
  assign new_n12413_ = ~new_n9445_ | ~new_n12399_;
  assign new_n12414_ = ~pi0726 | ~new_n12394_;
  assign new_n12415_ = ~new_n12383_ | ~new_n9465_;
  assign new_n12416_ = ~new_n9543_ | ~new_n9457_;
  assign new_n12417_ = ~new_n12382_ | ~new_n9456_;
  assign new_n12418_ = ~new_n9444_ | ~new_n12399_;
  assign new_n12419_ = ~pi0727 | ~new_n12394_;
  assign new_n12420_ = ~new_n12383_ | ~new_n9464_;
  assign new_n12421_ = ~new_n9543_ | ~new_n9455_;
  assign new_n12422_ = ~new_n12382_ | ~new_n9454_;
  assign new_n12423_ = ~new_n9443_ | ~new_n12399_;
  assign new_n12424_ = ~pi0728 | ~new_n12394_;
  assign new_n12425_ = ~new_n12383_ | ~new_n9473_;
  assign new_n12426_ = ~new_n9543_ | ~new_n9453_;
  assign new_n12427_ = ~new_n12382_ | ~new_n9452_;
  assign new_n12428_ = ~new_n9442_ | ~new_n12399_;
  assign new_n12429_ = ~pi0729 | ~new_n12394_;
  assign new_n12430_ = ~new_n12383_ | ~new_n9469_;
  assign new_n12431_ = ~new_n9543_ | ~new_n9451_;
  assign new_n12432_ = ~new_n12382_ | ~new_n9450_;
  assign new_n12433_ = ~new_n9441_ | ~new_n12399_;
  assign new_n12434_ = ~pi0730 | ~new_n12394_;
  assign new_n12435_ = ~new_n12383_ | ~new_n9472_;
  assign new_n12436_ = ~new_n9543_ | ~new_n9449_;
  assign new_n12437_ = ~new_n12382_ | ~new_n9448_;
  assign new_n12438_ = ~new_n9440_ | ~new_n12399_;
  assign new_n12439_ = ~pi0731 | ~new_n12394_;
  assign new_n12440_ = ~new_n10527_;
  assign new_n12441_ = ~new_n10526_;
  assign new_n12442_ = ~new_n10292_;
  assign new_n12443_ = ~new_n10598_;
  assign new_n12444_ = ~new_n10528_;
  assign new_n12445_ = ~new_n9542_ | ~new_n11674_;
  assign new_n12446_ = ~new_n9548_ | ~new_n9403_;
  assign new_n12447_ = ~new_n11486_ | ~new_n12446_;
  assign new_n12448_ = ~new_n12447_ | ~new_n10292_;
  assign new_n12449_ = ~new_n12444_ | ~pi0625;
  assign new_n12450_ = ~pi0624 | ~new_n10526_;
  assign new_n12451_ = ~new_n12448_ | ~new_n10880_;
  assign new_n12452_ = ~new_n9548_ | ~new_n9439_;
  assign new_n12453_ = ~new_n11486_ | ~new_n12452_;
  assign new_n12454_ = ~new_n12453_ | ~new_n12442_;
  assign new_n12455_ = ~pi0625 | ~new_n10528_;
  assign new_n12456_ = ~new_n12455_ | ~new_n12454_;
  assign new_n12457_ = ~new_n12441_ | ~new_n9466_;
  assign new_n12458_ = ~new_n9547_ | ~new_n9463_;
  assign new_n12459_ = ~new_n12440_ | ~new_n9462_;
  assign new_n12460_ = ~new_n9447_ | ~new_n12456_;
  assign new_n12461_ = ~pi0732 | ~new_n12451_;
  assign new_n12462_ = ~new_n12441_ | ~new_n9467_;
  assign new_n12463_ = ~new_n9547_ | ~new_n9461_;
  assign new_n12464_ = ~new_n12440_ | ~new_n9460_;
  assign new_n12465_ = ~new_n9446_ | ~new_n12456_;
  assign new_n12466_ = ~pi0733 | ~new_n12451_;
  assign new_n12467_ = ~new_n12441_ | ~new_n9470_;
  assign new_n12468_ = ~new_n9547_ | ~new_n9459_;
  assign new_n12469_ = ~new_n12440_ | ~new_n9458_;
  assign new_n12470_ = ~new_n9445_ | ~new_n12456_;
  assign new_n12471_ = ~pi0734 | ~new_n12451_;
  assign new_n12472_ = ~new_n12441_ | ~new_n9465_;
  assign new_n12473_ = ~new_n9547_ | ~new_n9457_;
  assign new_n12474_ = ~new_n12440_ | ~new_n9456_;
  assign new_n12475_ = ~new_n9444_ | ~new_n12456_;
  assign new_n12476_ = ~pi0735 | ~new_n12451_;
  assign new_n12477_ = ~new_n12441_ | ~new_n9464_;
  assign new_n12478_ = ~new_n9547_ | ~new_n9455_;
  assign new_n12479_ = ~new_n12440_ | ~new_n9454_;
  assign new_n12480_ = ~new_n9443_ | ~new_n12456_;
  assign new_n12481_ = ~pi0736 | ~new_n12451_;
  assign new_n12482_ = ~new_n12441_ | ~new_n9473_;
  assign new_n12483_ = ~new_n9547_ | ~new_n9453_;
  assign new_n12484_ = ~new_n12440_ | ~new_n9452_;
  assign new_n12485_ = ~new_n9442_ | ~new_n12456_;
  assign new_n12486_ = ~pi0737 | ~new_n12451_;
  assign new_n12487_ = ~new_n12441_ | ~new_n9469_;
  assign new_n12488_ = ~new_n9547_ | ~new_n9451_;
  assign new_n12489_ = ~new_n12440_ | ~new_n9450_;
  assign new_n12490_ = ~new_n9441_ | ~new_n12456_;
  assign new_n12491_ = ~pi0738 | ~new_n12451_;
  assign new_n12492_ = ~new_n12441_ | ~new_n9472_;
  assign new_n12493_ = ~new_n9547_ | ~new_n9449_;
  assign new_n12494_ = ~new_n12440_ | ~new_n9448_;
  assign new_n12495_ = ~new_n9440_ | ~new_n12456_;
  assign new_n12496_ = ~pi0739 | ~new_n12451_;
  assign new_n12497_ = ~new_n10538_;
  assign new_n12498_ = ~new_n10537_;
  assign new_n12499_ = ~new_n9484_ | ~new_n9486_;
  assign new_n12500_ = ~new_n10539_;
  assign new_n12501_ = ~new_n10597_;
  assign new_n12502_ = ~new_n10540_;
  assign new_n12503_ = ~new_n9542_ | ~new_n11675_;
  assign new_n12504_ = ~new_n9550_ | ~new_n9403_;
  assign new_n12505_ = ~new_n11486_ | ~new_n12504_;
  assign new_n12506_ = ~new_n12500_ | ~new_n12505_;
  assign new_n12507_ = ~new_n12502_ | ~pi0625;
  assign new_n12508_ = ~pi0624 | ~new_n10537_;
  assign new_n12509_ = ~new_n12506_ | ~new_n10889_;
  assign new_n12510_ = ~new_n9550_ | ~new_n9439_;
  assign new_n12511_ = ~new_n11486_ | ~new_n12510_;
  assign new_n12512_ = ~new_n12511_ | ~new_n10539_;
  assign new_n12513_ = ~pi0625 | ~new_n10540_;
  assign new_n12514_ = ~new_n12513_ | ~new_n12512_;
  assign new_n12515_ = ~new_n12498_ | ~new_n9466_;
  assign new_n12516_ = ~new_n9549_ | ~new_n9463_;
  assign new_n12517_ = ~new_n12497_ | ~new_n9462_;
  assign new_n12518_ = ~new_n9447_ | ~new_n12514_;
  assign new_n12519_ = ~pi0740 | ~new_n12509_;
  assign new_n12520_ = ~new_n12498_ | ~new_n9467_;
  assign new_n12521_ = ~new_n9549_ | ~new_n9461_;
  assign new_n12522_ = ~new_n12497_ | ~new_n9460_;
  assign new_n12523_ = ~new_n9446_ | ~new_n12514_;
  assign new_n12524_ = ~pi0741 | ~new_n12509_;
  assign new_n12525_ = ~new_n12498_ | ~new_n9470_;
  assign new_n12526_ = ~new_n9549_ | ~new_n9459_;
  assign new_n12527_ = ~new_n12497_ | ~new_n9458_;
  assign new_n12528_ = ~new_n9445_ | ~new_n12514_;
  assign new_n12529_ = ~pi0742 | ~new_n12509_;
  assign new_n12530_ = ~new_n12498_ | ~new_n9465_;
  assign new_n12531_ = ~new_n9549_ | ~new_n9457_;
  assign new_n12532_ = ~new_n12497_ | ~new_n9456_;
  assign new_n12533_ = ~new_n9444_ | ~new_n12514_;
  assign new_n12534_ = ~pi0743 | ~new_n12509_;
  assign new_n12535_ = ~new_n12498_ | ~new_n9464_;
  assign new_n12536_ = ~new_n9549_ | ~new_n9455_;
  assign new_n12537_ = ~new_n12497_ | ~new_n9454_;
  assign new_n12538_ = ~new_n9443_ | ~new_n12514_;
  assign new_n12539_ = ~pi0744 | ~new_n12509_;
  assign new_n12540_ = ~new_n12498_ | ~new_n9473_;
  assign new_n12541_ = ~new_n9549_ | ~new_n9453_;
  assign new_n12542_ = ~new_n12497_ | ~new_n9452_;
  assign new_n12543_ = ~new_n9442_ | ~new_n12514_;
  assign new_n12544_ = ~pi0745 | ~new_n12509_;
  assign new_n12545_ = ~new_n12498_ | ~new_n9469_;
  assign new_n12546_ = ~new_n9549_ | ~new_n9451_;
  assign new_n12547_ = ~new_n12497_ | ~new_n9450_;
  assign new_n12548_ = ~new_n9441_ | ~new_n12514_;
  assign new_n12549_ = ~pi0746 | ~new_n12509_;
  assign new_n12550_ = ~new_n12498_ | ~new_n9472_;
  assign new_n12551_ = ~new_n9549_ | ~new_n9449_;
  assign new_n12552_ = ~new_n12497_ | ~new_n9448_;
  assign new_n12553_ = ~new_n9440_ | ~new_n12514_;
  assign new_n12554_ = ~pi0747 | ~new_n12509_;
  assign new_n12555_ = ~new_n10550_;
  assign new_n12556_ = ~new_n10549_;
  assign new_n12557_ = ~new_n10293_;
  assign new_n12558_ = ~new_n10596_;
  assign new_n12559_ = ~new_n10551_;
  assign new_n12560_ = ~new_n9542_ | ~new_n9517_;
  assign new_n12561_ = ~new_n9552_ | ~new_n9403_;
  assign new_n12562_ = ~new_n11486_ | ~new_n12561_;
  assign new_n12563_ = ~new_n12562_ | ~new_n10293_;
  assign new_n12564_ = ~new_n12559_ | ~pi0625;
  assign new_n12565_ = ~pi0624 | ~new_n10549_;
  assign new_n12566_ = ~new_n12563_ | ~new_n10898_;
  assign new_n12567_ = ~new_n9552_ | ~new_n9439_;
  assign new_n12568_ = ~new_n11486_ | ~new_n12567_;
  assign new_n12569_ = ~new_n12568_ | ~new_n12557_;
  assign new_n12570_ = ~pi0625 | ~new_n10551_;
  assign new_n12571_ = ~new_n12570_ | ~new_n12569_;
  assign new_n12572_ = ~new_n12556_ | ~new_n9466_;
  assign new_n12573_ = ~new_n9551_ | ~new_n9463_;
  assign new_n12574_ = ~new_n12555_ | ~new_n9462_;
  assign new_n12575_ = ~new_n9447_ | ~new_n12571_;
  assign new_n12576_ = ~pi0748 | ~new_n12566_;
  assign new_n12577_ = ~new_n12556_ | ~new_n9467_;
  assign new_n12578_ = ~new_n9551_ | ~new_n9461_;
  assign new_n12579_ = ~new_n12555_ | ~new_n9460_;
  assign new_n12580_ = ~new_n9446_ | ~new_n12571_;
  assign new_n12581_ = ~pi0749 | ~new_n12566_;
  assign new_n12582_ = ~new_n12556_ | ~new_n9470_;
  assign new_n12583_ = ~new_n9551_ | ~new_n9459_;
  assign new_n12584_ = ~new_n12555_ | ~new_n9458_;
  assign new_n12585_ = ~new_n9445_ | ~new_n12571_;
  assign new_n12586_ = ~pi0750 | ~new_n12566_;
  assign new_n12587_ = ~new_n12556_ | ~new_n9465_;
  assign new_n12588_ = ~new_n9551_ | ~new_n9457_;
  assign new_n12589_ = ~new_n12555_ | ~new_n9456_;
  assign new_n12590_ = ~new_n9444_ | ~new_n12571_;
  assign new_n12591_ = ~pi0751 | ~new_n12566_;
  assign new_n12592_ = ~new_n12556_ | ~new_n9464_;
  assign new_n12593_ = ~new_n9551_ | ~new_n9455_;
  assign new_n12594_ = ~new_n12555_ | ~new_n9454_;
  assign new_n12595_ = ~new_n9443_ | ~new_n12571_;
  assign new_n12596_ = ~pi0752 | ~new_n12566_;
  assign new_n12597_ = ~new_n12556_ | ~new_n9473_;
  assign new_n12598_ = ~new_n9551_ | ~new_n9453_;
  assign new_n12599_ = ~new_n12555_ | ~new_n9452_;
  assign new_n12600_ = ~new_n9442_ | ~new_n12571_;
  assign new_n12601_ = ~pi0753 | ~new_n12566_;
  assign new_n12602_ = ~new_n12556_ | ~new_n9469_;
  assign new_n12603_ = ~new_n9551_ | ~new_n9451_;
  assign new_n12604_ = ~new_n12555_ | ~new_n9450_;
  assign new_n12605_ = ~new_n9441_ | ~new_n12571_;
  assign new_n12606_ = ~pi0754 | ~new_n12566_;
  assign new_n12607_ = ~new_n12556_ | ~new_n9472_;
  assign new_n12608_ = ~new_n9551_ | ~new_n9449_;
  assign new_n12609_ = ~new_n12555_ | ~new_n9448_;
  assign new_n12610_ = ~new_n9440_ | ~new_n12571_;
  assign new_n12611_ = ~pi0755 | ~new_n12566_;
  assign new_n12612_ = ~new_n10320_ | ~new_n14910_;
  assign new_n12613_ = ~new_n10615_;
  assign new_n12614_ = ~new_n14902_ | ~new_n14904_ | ~new_n9658_;
  assign new_n12615_ = ~new_n10562_ | ~new_n10330_ | ~new_n10296_ | ~new_n14936_;
  assign new_n12616_ = ~new_n9398_ | ~new_n14912_;
  assign new_n12617_ = ~new_n11458_ | ~new_n10615_;
  assign new_n12618_ = ~new_n11469_ | ~new_n11465_;
  assign new_n12619_ = ~new_n10565_ | ~new_n12618_;
  assign new_n12620_ = ~new_n30327_ | ~new_n12619_ | ~new_n10306_;
  assign new_n12621_ = ~new_n11477_ | ~new_n28599_;
  assign new_n12622_ = ~new_n11447_;
  assign new_n12623_ = ~new_n9415_ | ~new_n11447_;
  assign new_n12624_ = ~pi0624 | ~new_n10325_;
  assign new_n12625_ = ~new_n11435_;
  assign new_n12626_ = ~new_n11632_ | ~new_n10317_;
  assign new_n12627_ = ~new_n10919_ | ~new_n9658_ | ~new_n10336_;
  assign new_n12628_ = ~new_n10336_ | ~new_n10296_;
  assign new_n12629_ = ~new_n14906_ | ~new_n10319_;
  assign new_n12630_ = ~new_n10920_ | ~new_n15116_ | ~new_n15115_;
  assign new_n12631_ = ~new_n10566_;
  assign new_n12632_ = ~new_n14779_ | ~new_n10319_;
  assign new_n12633_ = ~new_n12632_ | ~new_n12612_ | ~new_n12614_ | ~new_n10562_;
  assign new_n12634_ = ~new_n11458_ | ~new_n10615_;
  assign new_n12635_ = ~new_n12633_ | ~new_n9657_;
  assign new_n12636_ = ~new_n10918_ | ~new_n12635_;
  assign new_n12637_ = ~new_n10336_ | ~new_n14914_;
  assign new_n12638_ = ~new_n10320_ | ~new_n14912_;
  assign new_n12639_ = ~new_n9658_ | ~new_n10562_;
  assign new_n12640_ = ~new_n11468_ | ~new_n12639_;
  assign new_n12641_ = ~new_n12638_ | ~new_n10321_;
  assign new_n12642_ = ~new_n9477_ | ~new_n14925_;
  assign new_n12643_ = ~new_n10568_ | ~new_n10319_;
  assign new_n12644_ = ~new_n9555_ | ~new_n10329_;
  assign new_n12645_ = ~new_n11511_ | ~new_n15118_ | ~new_n15117_;
  assign new_n12646_ = ~new_n10337_ | ~new_n10563_;
  assign new_n12647_ = ~new_n10619_ | ~new_n11478_;
  assign new_n12648_ = ~new_n11436_ | ~new_n12646_;
  assign new_n12649_ = ~new_n10622_ | ~new_n12647_;
  assign new_n12650_ = ~new_n29006_ | ~new_n12645_;
  assign new_n12651_ = ~new_n27643_ | ~new_n12644_;
  assign new_n12652_ = ~new_n10925_ | ~new_n12651_;
  assign new_n12653_ = ~new_n28369_ | ~new_n11510_;
  assign new_n12654_ = ~new_n11507_ | ~new_n12652_;
  assign new_n12655_ = ~new_n12654_ | ~new_n12653_;
  assign new_n12656_ = ~pi0758 | ~new_n11632_;
  assign new_n12657_ = ~new_n10571_;
  assign new_n12658_ = ~new_n29007_ | ~new_n12645_;
  assign new_n12659_ = ~new_n27644_ | ~new_n12644_;
  assign new_n12660_ = ~new_n10926_ | ~new_n12659_;
  assign new_n12661_ = ~pi0626 | ~new_n10639_ | ~new_n10638_;
  assign new_n12662_ = ~new_n28333_ | ~new_n11510_;
  assign new_n12663_ = ~new_n11507_ | ~new_n12660_;
  assign new_n12664_ = ~new_n12661_ | ~new_n12662_ | ~new_n12663_;
  assign new_n12665_ = ~new_n11470_ | ~new_n9490_ | ~new_n14902_;
  assign new_n12666_ = ~new_n14923_ | ~new_n12665_;
  assign new_n12667_ = ~new_n10928_ | ~new_n15138_;
  assign new_n12668_ = ~new_n29002_ | ~new_n12645_;
  assign new_n12669_ = ~new_n27553_ | ~new_n12644_;
  assign new_n12670_ = ~new_n10929_ | ~new_n12669_;
  assign new_n12671_ = ~new_n10638_ | ~pi0626 | ~new_n15131_;
  assign new_n12672_ = ~new_n28361_ | ~new_n11510_;
  assign new_n12673_ = ~new_n11507_ | ~new_n12670_;
  assign new_n12674_ = ~new_n12671_ | ~new_n12672_ | ~new_n12673_;
  assign new_n12675_ = ~new_n10930_ | ~new_n15138_;
  assign new_n12676_ = ~pi0760 | ~new_n12645_;
  assign new_n12677_ = ~new_n27642_ | ~new_n12644_;
  assign new_n12678_ = ~new_n10931_ | ~new_n12677_;
  assign new_n12679_ = ~new_n28362_ | ~new_n11510_;
  assign new_n12680_ = ~new_n11507_ | ~new_n12678_;
  assign new_n12681_ = ~new_n15128_ | ~pi0626;
  assign new_n12682_ = ~new_n12681_ | ~new_n12680_ | ~new_n12679_;
  assign new_n12683_ = ~new_n29132_ | ~new_n9489_ | ~pi0627;
  assign new_n12684_ = ~new_n10574_;
  assign new_n12685_ = ~new_n11486_ | ~new_n10344_;
  assign new_n12686_ = ~new_n11677_ | ~new_n10620_;
  assign new_n12687_ = ~new_n10467_ | ~new_n12686_;
  assign new_n12688_ = ~new_n10468_ | ~new_n12687_;
  assign new_n12689_ = ~new_n9439_ | ~new_n12688_;
  assign new_n12690_ = ~new_n28369_ | ~new_n12685_;
  assign new_n12691_ = ~new_n29211_ | ~pi0624;
  assign new_n12692_ = ~new_n10932_ | ~new_n12689_;
  assign new_n12693_ = ~new_n9439_ | ~new_n15150_;
  assign new_n12694_ = ~new_n28333_ | ~new_n12685_;
  assign new_n12695_ = ~new_n29213_ | ~pi0624;
  assign new_n12696_ = ~new_n10933_ | ~new_n12693_;
  assign new_n12697_ = ~new_n10379_ | ~new_n10394_;
  assign new_n12698_ = ~new_n9439_ | ~new_n12697_;
  assign new_n12699_ = ~new_n28361_ | ~new_n12685_;
  assign new_n12700_ = ~new_n29187_ | ~pi0624;
  assign new_n12701_ = ~new_n10934_ | ~new_n12698_;
  assign new_n12702_ = ~new_n10354_ | ~new_n10344_;
  assign new_n12703_ = ~new_n28362_ | ~new_n12702_;
  assign new_n12704_ = ~new_n29204_ | ~pi0624;
  assign new_n12705_ = ~new_n11505_ | ~new_n12703_ | ~new_n12704_;
  assign new_n12706_ = ~new_n9657_ | ~new_n10333_;
  assign new_n12707_ = ~new_n29402_ | ~new_n11458_;
  assign new_n12708_ = ~new_n12707_ | ~new_n12706_;
  assign new_n12709_ = ~new_n15162_ | ~new_n30327_ | ~new_n10306_ | ~new_n15163_;
  assign new_n12710_ = ~new_n11461_ | ~new_n12708_;
  assign new_n12711_ = ~new_n10935_ | ~new_n12710_ | ~new_n11438_ | ~new_n9553_;
  assign new_n12712_ = ~new_n9415_ | ~new_n12711_;
  assign new_n12713_ = ~new_n11502_ | ~new_n10325_;
  assign new_n12714_ = ~new_n10576_;
  assign new_n12715_ = ~new_n11468_ | ~new_n11461_;
  assign new_n12716_ = ~new_n10936_ | ~new_n9555_;
  assign new_n12717_ = ~new_n11458_ | ~new_n11465_;
  assign new_n12718_ = ~new_n11511_ | ~new_n10565_ | ~new_n11478_ | ~new_n12717_;
  assign new_n12719_ = ~new_n11469_ | ~new_n11465_;
  assign new_n12720_ = ~new_n10564_ | ~new_n10337_ | ~new_n12719_;
  assign new_n12721_ = ~new_n9431_ | ~new_n29204_;
  assign new_n12722_ = ~new_n9430_ | ~new_n27642_;
  assign new_n12723_ = ~new_n28636_ | ~new_n9429_;
  assign new_n12724_ = ~new_n30329_ | ~new_n9427_;
  assign new_n12725_ = ~new_n29789_ | ~new_n9426_;
  assign new_n12726_ = ~new_n30737_ | ~new_n9425_;
  assign new_n12727_ = ~pi0957 | ~new_n9422_;
  assign new_n12728_ = ~new_n12714_ | ~pi0766;
  assign new_n12729_ = ~new_n9431_ | ~new_n29187_;
  assign new_n12730_ = ~new_n9430_ | ~new_n27553_;
  assign new_n12731_ = ~new_n28716_ | ~new_n9429_;
  assign new_n12732_ = ~new_n30410_ | ~new_n9427_;
  assign new_n12733_ = ~new_n29712_ | ~new_n9426_;
  assign new_n12734_ = ~new_n30694_ | ~new_n9425_;
  assign new_n12735_ = ~new_n9422_ | ~pi0958;
  assign new_n12736_ = ~new_n12714_ | ~pi0767;
  assign new_n12737_ = ~new_n9431_ | ~new_n29213_;
  assign new_n12738_ = ~new_n9430_ | ~new_n27644_;
  assign new_n12739_ = ~new_n28705_ | ~new_n9429_;
  assign new_n12740_ = ~new_n30330_ | ~new_n9427_;
  assign new_n12741_ = ~new_n29798_ | ~new_n9426_;
  assign new_n12742_ = ~new_n30748_ | ~new_n9425_;
  assign new_n12743_ = ~new_n9422_ | ~pi0959;
  assign new_n12744_ = ~pi0768 | ~new_n12714_;
  assign new_n12745_ = ~new_n9431_ | ~new_n29211_;
  assign new_n12746_ = ~new_n9430_ | ~new_n27643_;
  assign new_n12747_ = ~new_n28702_ | ~new_n9429_;
  assign new_n12748_ = ~new_n30420_ | ~new_n9427_;
  assign new_n12749_ = ~new_n29796_ | ~new_n9426_;
  assign new_n12750_ = ~new_n30753_ | ~new_n9425_;
  assign new_n12751_ = ~new_n9422_ | ~pi0960;
  assign new_n12752_ = ~pi0769 | ~new_n12714_;
  assign new_n12753_ = ~new_n29210_ | ~new_n9431_;
  assign new_n12754_ = ~new_n27646_ | ~new_n9430_;
  assign new_n12755_ = ~new_n28701_ | ~new_n9429_;
  assign new_n12756_ = ~new_n30401_ | ~new_n9427_;
  assign new_n12757_ = ~new_n29795_ | ~new_n9426_;
  assign new_n12758_ = ~new_n30749_ | ~new_n9425_;
  assign new_n12759_ = ~new_n9422_ | ~pi0961;
  assign new_n12760_ = ~pi0770 | ~new_n12714_;
  assign new_n12761_ = ~new_n29209_ | ~new_n9431_;
  assign new_n12762_ = ~new_n27619_ | ~new_n9430_;
  assign new_n12763_ = ~new_n28700_ | ~new_n9429_;
  assign new_n12764_ = ~new_n30404_ | ~new_n9427_;
  assign new_n12765_ = ~new_n29794_ | ~new_n9426_;
  assign new_n12766_ = ~new_n30750_ | ~new_n9425_;
  assign new_n12767_ = ~new_n9422_ | ~pi0962;
  assign new_n12768_ = ~pi0771 | ~new_n12714_;
  assign new_n12769_ = ~new_n29208_ | ~new_n9431_;
  assign new_n12770_ = ~new_n27618_ | ~new_n9430_;
  assign new_n12771_ = ~new_n28699_ | ~new_n9429_;
  assign new_n12772_ = ~new_n30388_ | ~new_n9427_;
  assign new_n12773_ = ~new_n29793_ | ~new_n9426_;
  assign new_n12774_ = ~new_n30747_ | ~new_n9425_;
  assign new_n12775_ = ~new_n9422_ | ~pi0963;
  assign new_n12776_ = ~pi0772 | ~new_n12714_;
  assign new_n12777_ = ~new_n29207_ | ~new_n9431_;
  assign new_n12778_ = ~new_n27617_ | ~new_n9430_;
  assign new_n12779_ = ~new_n28698_ | ~new_n9429_;
  assign new_n12780_ = ~new_n30414_ | ~new_n9427_;
  assign new_n12781_ = ~new_n29792_ | ~new_n9426_;
  assign new_n12782_ = ~new_n30754_ | ~new_n9425_;
  assign new_n12783_ = ~new_n9422_ | ~pi0964;
  assign new_n12784_ = ~pi0773 | ~new_n12714_;
  assign new_n12785_ = ~new_n29206_ | ~new_n9431_;
  assign new_n12786_ = ~new_n27616_ | ~new_n9430_;
  assign new_n12787_ = ~new_n28697_ | ~new_n9429_;
  assign new_n12788_ = ~new_n30405_ | ~new_n9427_;
  assign new_n12789_ = ~new_n29791_ | ~new_n9426_;
  assign new_n12790_ = ~new_n30751_ | ~new_n9425_;
  assign new_n12791_ = ~new_n9422_ | ~pi0965;
  assign new_n12792_ = ~pi0774 | ~new_n12714_;
  assign new_n12793_ = ~new_n29205_ | ~new_n9431_;
  assign new_n12794_ = ~new_n27615_ | ~new_n9430_;
  assign new_n12795_ = ~new_n28696_ | ~new_n9429_;
  assign new_n12796_ = ~new_n30395_ | ~new_n9427_;
  assign new_n12797_ = ~new_n29790_ | ~new_n9426_;
  assign new_n12798_ = ~new_n30787_ | ~new_n9425_;
  assign new_n12799_ = ~new_n9422_ | ~pi0966;
  assign new_n12800_ = ~pi0775 | ~new_n12714_;
  assign new_n12801_ = ~new_n29233_ | ~new_n9431_;
  assign new_n12802_ = ~new_n27641_ | ~new_n9430_;
  assign new_n12803_ = ~new_n28726_ | ~new_n9429_;
  assign new_n12804_ = ~new_n30408_ | ~new_n9427_;
  assign new_n12805_ = ~new_n29818_ | ~new_n9426_;
  assign new_n12806_ = ~new_n30682_ | ~new_n9425_;
  assign new_n12807_ = ~new_n9422_ | ~pi0967;
  assign new_n12808_ = ~pi0776 | ~new_n12714_;
  assign new_n12809_ = ~new_n29232_ | ~new_n9431_;
  assign new_n12810_ = ~new_n27640_ | ~new_n9430_;
  assign new_n12811_ = ~new_n28725_ | ~new_n9429_;
  assign new_n12812_ = ~new_n30398_ | ~new_n9427_;
  assign new_n12813_ = ~new_n29817_ | ~new_n9426_;
  assign new_n12814_ = ~new_n30683_ | ~new_n9425_;
  assign new_n12815_ = ~new_n9422_ | ~pi0968;
  assign new_n12816_ = ~pi0777 | ~new_n12714_;
  assign new_n12817_ = ~new_n29231_ | ~new_n9431_;
  assign new_n12818_ = ~new_n27639_ | ~new_n9430_;
  assign new_n12819_ = ~new_n28724_ | ~new_n9429_;
  assign new_n12820_ = ~new_n30413_ | ~new_n9427_;
  assign new_n12821_ = ~new_n29816_ | ~new_n9426_;
  assign new_n12822_ = ~new_n30745_ | ~new_n9425_;
  assign new_n12823_ = ~new_n9422_ | ~pi0969;
  assign new_n12824_ = ~pi0778 | ~new_n12714_;
  assign new_n12825_ = ~new_n29230_ | ~new_n9431_;
  assign new_n12826_ = ~new_n27638_ | ~new_n9430_;
  assign new_n12827_ = ~new_n28723_ | ~new_n9429_;
  assign new_n12828_ = ~new_n30394_ | ~new_n9427_;
  assign new_n12829_ = ~new_n29815_ | ~new_n9426_;
  assign new_n12830_ = ~new_n30684_ | ~new_n9425_;
  assign new_n12831_ = ~new_n9422_ | ~pi0970;
  assign new_n12832_ = ~pi0779 | ~new_n12714_;
  assign new_n12833_ = ~new_n29229_ | ~new_n9431_;
  assign new_n12834_ = ~new_n27637_ | ~new_n9430_;
  assign new_n12835_ = ~new_n28722_ | ~new_n9429_;
  assign new_n12836_ = ~new_n30403_ | ~new_n9427_;
  assign new_n12837_ = ~new_n29814_ | ~new_n9426_;
  assign new_n12838_ = ~new_n30685_ | ~new_n9425_;
  assign new_n12839_ = ~new_n9422_ | ~pi0971;
  assign new_n12840_ = ~pi0780 | ~new_n12714_;
  assign new_n12841_ = ~new_n29228_ | ~new_n9431_;
  assign new_n12842_ = ~new_n27636_ | ~new_n9430_;
  assign new_n12843_ = ~new_n28721_ | ~new_n9429_;
  assign new_n12844_ = ~new_n30400_ | ~new_n9427_;
  assign new_n12845_ = ~new_n29813_ | ~new_n9426_;
  assign new_n12846_ = ~new_n30742_ | ~new_n9425_;
  assign new_n12847_ = ~new_n9422_ | ~pi0972;
  assign new_n12848_ = ~pi0781 | ~new_n12714_;
  assign new_n12849_ = ~new_n29227_ | ~new_n9431_;
  assign new_n12850_ = ~new_n27635_ | ~new_n9430_;
  assign new_n12851_ = ~new_n28720_ | ~new_n9429_;
  assign new_n12852_ = ~new_n30416_ | ~new_n9427_;
  assign new_n12853_ = ~new_n29812_ | ~new_n9426_;
  assign new_n12854_ = ~new_n30686_ | ~new_n9425_;
  assign new_n12855_ = ~new_n9422_ | ~pi0973;
  assign new_n12856_ = ~pi0782 | ~new_n12714_;
  assign new_n12857_ = ~new_n29226_ | ~new_n9431_;
  assign new_n12858_ = ~new_n27634_ | ~new_n9430_;
  assign new_n12859_ = ~new_n28719_ | ~new_n9429_;
  assign new_n12860_ = ~new_n30392_ | ~new_n9427_;
  assign new_n12861_ = ~new_n29811_ | ~new_n9426_;
  assign new_n12862_ = ~new_n30740_ | ~new_n9425_;
  assign new_n12863_ = ~new_n9422_ | ~pi0974;
  assign new_n12864_ = ~pi0783 | ~new_n12714_;
  assign new_n12865_ = ~new_n29225_ | ~new_n9431_;
  assign new_n12866_ = ~new_n27633_ | ~new_n9430_;
  assign new_n12867_ = ~new_n28718_ | ~new_n9429_;
  assign new_n12868_ = ~new_n30397_ | ~new_n9427_;
  assign new_n12869_ = ~new_n29810_ | ~new_n9426_;
  assign new_n12870_ = ~new_n30741_ | ~new_n9425_;
  assign new_n12871_ = ~new_n9422_ | ~pi0975;
  assign new_n12872_ = ~pi0784 | ~new_n12714_;
  assign new_n12873_ = ~new_n29224_ | ~new_n9431_;
  assign new_n12874_ = ~new_n27632_ | ~new_n9430_;
  assign new_n12875_ = ~new_n28717_ | ~new_n9429_;
  assign new_n12876_ = ~new_n30407_ | ~new_n9427_;
  assign new_n12877_ = ~new_n29809_ | ~new_n9426_;
  assign new_n12878_ = ~new_n30687_ | ~new_n9425_;
  assign new_n12879_ = ~new_n9422_ | ~pi0976;
  assign new_n12880_ = ~pi0785 | ~new_n12714_;
  assign new_n12881_ = ~new_n29223_ | ~new_n9431_;
  assign new_n12882_ = ~new_n27631_ | ~new_n9430_;
  assign new_n12883_ = ~new_n28715_ | ~new_n9429_;
  assign new_n12884_ = ~new_n30393_ | ~new_n9427_;
  assign new_n12885_ = ~new_n29808_ | ~new_n9426_;
  assign new_n12886_ = ~new_n30688_ | ~new_n9425_;
  assign new_n12887_ = ~new_n9422_ | ~pi0977;
  assign new_n12888_ = ~pi0786 | ~new_n12714_;
  assign new_n12889_ = ~new_n29222_ | ~new_n9431_;
  assign new_n12890_ = ~new_n27630_ | ~new_n9430_;
  assign new_n12891_ = ~new_n28714_ | ~new_n9429_;
  assign new_n12892_ = ~new_n30412_ | ~new_n9427_;
  assign new_n12893_ = ~new_n29807_ | ~new_n9426_;
  assign new_n12894_ = ~new_n30744_ | ~new_n9425_;
  assign new_n12895_ = ~new_n9422_ | ~pi0978;
  assign new_n12896_ = ~pi0787 | ~new_n12714_;
  assign new_n12897_ = ~new_n29221_ | ~new_n9431_;
  assign new_n12898_ = ~new_n27629_ | ~new_n9430_;
  assign new_n12899_ = ~new_n28713_ | ~new_n9429_;
  assign new_n12900_ = ~new_n30396_ | ~new_n9427_;
  assign new_n12901_ = ~new_n29806_ | ~new_n9426_;
  assign new_n12902_ = ~new_n30689_ | ~new_n9425_;
  assign new_n12903_ = ~new_n9422_ | ~pi0979;
  assign new_n12904_ = ~pi0788 | ~new_n12714_;
  assign new_n12905_ = ~new_n29220_ | ~new_n9431_;
  assign new_n12906_ = ~new_n27628_ | ~new_n9430_;
  assign new_n12907_ = ~new_n28712_ | ~new_n9429_;
  assign new_n12908_ = ~new_n30406_ | ~new_n9427_;
  assign new_n12909_ = ~new_n29805_ | ~new_n9426_;
  assign new_n12910_ = ~new_n30690_ | ~new_n9425_;
  assign new_n12911_ = ~new_n9422_ | ~pi0980;
  assign new_n12912_ = ~pi0789 | ~new_n12714_;
  assign new_n12913_ = ~new_n29219_ | ~new_n9431_;
  assign new_n12914_ = ~new_n27627_ | ~new_n9430_;
  assign new_n12915_ = ~new_n28711_ | ~new_n9429_;
  assign new_n12916_ = ~new_n30391_ | ~new_n9427_;
  assign new_n12917_ = ~new_n29804_ | ~new_n9426_;
  assign new_n12918_ = ~new_n30739_ | ~new_n9425_;
  assign new_n12919_ = ~new_n9422_ | ~pi0981;
  assign new_n12920_ = ~pi0790 | ~new_n12714_;
  assign new_n12921_ = ~new_n29218_ | ~new_n9431_;
  assign new_n12922_ = ~new_n27626_ | ~new_n9430_;
  assign new_n12923_ = ~new_n28710_ | ~new_n9429_;
  assign new_n12924_ = ~new_n30415_ | ~new_n9427_;
  assign new_n12925_ = ~new_n29803_ | ~new_n9426_;
  assign new_n12926_ = ~new_n30746_ | ~new_n9425_;
  assign new_n12927_ = ~new_n9422_ | ~pi0982;
  assign new_n12928_ = ~pi0791 | ~new_n12714_;
  assign new_n12929_ = ~new_n29217_ | ~new_n9431_;
  assign new_n12930_ = ~new_n27625_ | ~new_n9430_;
  assign new_n12931_ = ~new_n28709_ | ~new_n9429_;
  assign new_n12932_ = ~new_n30399_ | ~new_n9427_;
  assign new_n12933_ = ~new_n29802_ | ~new_n9426_;
  assign new_n12934_ = ~new_n30691_ | ~new_n9425_;
  assign new_n12935_ = ~new_n9422_ | ~pi0983;
  assign new_n12936_ = ~pi0792 | ~new_n12714_;
  assign new_n12937_ = ~new_n29216_ | ~new_n9431_;
  assign new_n12938_ = ~new_n27624_ | ~new_n9430_;
  assign new_n12939_ = ~new_n28708_ | ~new_n9429_;
  assign new_n12940_ = ~new_n30402_ | ~new_n9427_;
  assign new_n12941_ = ~new_n29801_ | ~new_n9426_;
  assign new_n12942_ = ~new_n30743_ | ~new_n9425_;
  assign new_n12943_ = ~new_n9422_ | ~pi0984;
  assign new_n12944_ = ~pi0793 | ~new_n12714_;
  assign new_n12945_ = ~new_n29215_ | ~new_n9431_;
  assign new_n12946_ = ~new_n27623_ | ~new_n9430_;
  assign new_n12947_ = ~new_n28707_ | ~new_n9429_;
  assign new_n12948_ = ~new_n30411_ | ~new_n9427_;
  assign new_n12949_ = ~new_n29800_ | ~new_n9426_;
  assign new_n12950_ = ~new_n30692_ | ~new_n9425_;
  assign new_n12951_ = ~new_n9422_ | ~pi0985;
  assign new_n12952_ = ~pi0794 | ~new_n12714_;
  assign new_n12953_ = ~new_n29214_ | ~new_n9431_;
  assign new_n12954_ = ~new_n27622_ | ~new_n9430_;
  assign new_n12955_ = ~new_n28706_ | ~new_n9429_;
  assign new_n12956_ = ~new_n30390_ | ~new_n9427_;
  assign new_n12957_ = ~new_n29799_ | ~new_n9426_;
  assign new_n12958_ = ~new_n30693_ | ~new_n9425_;
  assign new_n12959_ = ~new_n9422_ | ~pi0986;
  assign new_n12960_ = ~pi0795 | ~new_n12714_;
  assign new_n12961_ = ~new_n29212_ | ~new_n9431_;
  assign new_n12962_ = ~new_n27621_ | ~new_n9430_;
  assign new_n12963_ = ~new_n28704_ | ~new_n9429_;
  assign new_n12964_ = ~new_n30389_ | ~new_n9427_;
  assign new_n12965_ = ~new_n29797_ | ~new_n9426_;
  assign new_n12966_ = ~new_n30738_ | ~new_n9425_;
  assign new_n12967_ = ~new_n9422_ | ~pi0987;
  assign new_n12968_ = ~pi0796 | ~new_n12714_;
  assign new_n12969_ = ~new_n29186_ | ~new_n9431_;
  assign new_n12970_ = ~new_n27620_ | ~new_n9430_;
  assign new_n12971_ = ~new_n28703_ | ~new_n9429_;
  assign new_n12972_ = ~new_n30409_ | ~new_n9427_;
  assign new_n12973_ = ~new_n29711_ | ~new_n9426_;
  assign new_n12974_ = ~new_n30752_ | ~new_n9425_;
  assign new_n12975_ = ~new_n9422_ | ~pi0988;
  assign new_n12976_ = ~pi0797 | ~new_n12714_;
  assign new_n12977_ = ~new_n11654_ | ~new_n11461_ | ~new_n9415_;
  assign new_n12978_ = ~new_n12702_ | ~new_n10325_;
  assign new_n12979_ = ~new_n10578_;
  assign new_n12980_ = ~pi0626 | ~new_n10343_;
  assign new_n12981_ = ~new_n10581_ | ~new_n12980_;
  assign new_n12982_ = ~pi0798 | ~new_n9428_;
  assign new_n12983_ = ~new_n9414_ | ~new_n30737_;
  assign new_n12984_ = ~new_n9413_ | ~new_n27642_;
  assign new_n12985_ = ~new_n9412_ | ~pi0957;
  assign new_n12986_ = ~new_n9411_ | ~new_n29789_;
  assign new_n12987_ = ~pi0798 | ~new_n12979_;
  assign new_n12988_ = ~new_n28823_ | ~new_n9428_;
  assign new_n12989_ = ~new_n9414_ | ~new_n30694_;
  assign new_n12990_ = ~new_n9413_ | ~new_n27553_;
  assign new_n12991_ = ~new_n9412_ | ~pi0958;
  assign new_n12992_ = ~new_n9411_ | ~new_n29712_;
  assign new_n12993_ = ~pi0799 | ~new_n12979_;
  assign new_n12994_ = ~new_n28889_ | ~new_n9428_;
  assign new_n12995_ = ~new_n9414_ | ~new_n30748_;
  assign new_n12996_ = ~new_n9413_ | ~new_n27644_;
  assign new_n12997_ = ~new_n9412_ | ~pi0959;
  assign new_n12998_ = ~new_n9411_ | ~new_n29798_;
  assign new_n12999_ = ~pi0800 | ~new_n12979_;
  assign new_n13000_ = ~new_n28886_ | ~new_n9428_;
  assign new_n13001_ = ~new_n9414_ | ~new_n30753_;
  assign new_n13002_ = ~new_n9413_ | ~new_n27643_;
  assign new_n13003_ = ~new_n9412_ | ~pi0960;
  assign new_n13004_ = ~new_n9411_ | ~new_n29796_;
  assign new_n13005_ = ~pi0801 | ~new_n12979_;
  assign new_n13006_ = ~new_n28885_ | ~new_n9428_;
  assign new_n13007_ = ~new_n9414_ | ~new_n30749_;
  assign new_n13008_ = ~new_n9413_ | ~new_n27646_;
  assign new_n13009_ = ~new_n9412_ | ~pi0961;
  assign new_n13010_ = ~new_n9411_ | ~new_n29795_;
  assign new_n13011_ = ~pi0802 | ~new_n12979_;
  assign new_n13012_ = ~new_n28884_ | ~new_n9428_;
  assign new_n13013_ = ~new_n9414_ | ~new_n30750_;
  assign new_n13014_ = ~new_n9413_ | ~new_n27619_;
  assign new_n13015_ = ~new_n9412_ | ~pi0962;
  assign new_n13016_ = ~new_n9411_ | ~new_n29794_;
  assign new_n13017_ = ~pi0803 | ~new_n12979_;
  assign new_n13018_ = ~new_n28883_ | ~new_n9428_;
  assign new_n13019_ = ~new_n9414_ | ~new_n30747_;
  assign new_n13020_ = ~new_n9413_ | ~new_n27618_;
  assign new_n13021_ = ~new_n9412_ | ~pi0963;
  assign new_n13022_ = ~new_n9411_ | ~new_n29793_;
  assign new_n13023_ = ~pi0804 | ~new_n12979_;
  assign new_n13024_ = ~new_n28882_ | ~new_n9428_;
  assign new_n13025_ = ~new_n9414_ | ~new_n30754_;
  assign new_n13026_ = ~new_n9413_ | ~new_n27617_;
  assign new_n13027_ = ~new_n9412_ | ~pi0964;
  assign new_n13028_ = ~new_n9411_ | ~new_n29792_;
  assign new_n13029_ = ~pi0805 | ~new_n12979_;
  assign new_n13030_ = ~new_n28881_ | ~new_n9428_;
  assign new_n13031_ = ~new_n9414_ | ~new_n30751_;
  assign new_n13032_ = ~new_n9413_ | ~new_n27616_;
  assign new_n13033_ = ~new_n9412_ | ~pi0965;
  assign new_n13034_ = ~new_n9411_ | ~new_n29791_;
  assign new_n13035_ = ~pi0806 | ~new_n12979_;
  assign new_n13036_ = ~new_n28880_ | ~new_n9428_;
  assign new_n13037_ = ~new_n9414_ | ~new_n30787_;
  assign new_n13038_ = ~new_n9413_ | ~new_n27615_;
  assign new_n13039_ = ~new_n9412_ | ~pi0966;
  assign new_n13040_ = ~new_n9411_ | ~new_n29790_;
  assign new_n13041_ = ~pi0807 | ~new_n12979_;
  assign new_n13042_ = ~new_n28909_ | ~new_n9428_;
  assign new_n13043_ = ~new_n9414_ | ~new_n30682_;
  assign new_n13044_ = ~new_n9413_ | ~new_n27641_;
  assign new_n13045_ = ~new_n9412_ | ~pi0967;
  assign new_n13046_ = ~new_n9411_ | ~new_n29818_;
  assign new_n13047_ = ~pi0808 | ~new_n12979_;
  assign new_n13048_ = ~new_n28908_ | ~new_n9428_;
  assign new_n13049_ = ~new_n9414_ | ~new_n30683_;
  assign new_n13050_ = ~new_n9413_ | ~new_n27640_;
  assign new_n13051_ = ~new_n9412_ | ~pi0968;
  assign new_n13052_ = ~new_n9411_ | ~new_n29817_;
  assign new_n13053_ = ~pi0809 | ~new_n12979_;
  assign new_n13054_ = ~new_n28907_ | ~new_n9428_;
  assign new_n13055_ = ~new_n9414_ | ~new_n30745_;
  assign new_n13056_ = ~new_n9413_ | ~new_n27639_;
  assign new_n13057_ = ~new_n9412_ | ~pi0969;
  assign new_n13058_ = ~new_n9411_ | ~new_n29816_;
  assign new_n13059_ = ~pi0810 | ~new_n12979_;
  assign new_n13060_ = ~new_n28906_ | ~new_n9428_;
  assign new_n13061_ = ~new_n9414_ | ~new_n30684_;
  assign new_n13062_ = ~new_n9413_ | ~new_n27638_;
  assign new_n13063_ = ~new_n9412_ | ~pi0970;
  assign new_n13064_ = ~new_n9411_ | ~new_n29815_;
  assign new_n13065_ = ~pi0811 | ~new_n12979_;
  assign new_n13066_ = ~new_n28905_ | ~new_n9428_;
  assign new_n13067_ = ~new_n9414_ | ~new_n30685_;
  assign new_n13068_ = ~new_n9413_ | ~new_n27637_;
  assign new_n13069_ = ~new_n9412_ | ~pi0971;
  assign new_n13070_ = ~new_n9411_ | ~new_n29814_;
  assign new_n13071_ = ~pi0812 | ~new_n12979_;
  assign new_n13072_ = ~new_n28904_ | ~new_n9428_;
  assign new_n13073_ = ~new_n9414_ | ~new_n30742_;
  assign new_n13074_ = ~new_n9413_ | ~new_n27636_;
  assign new_n13075_ = ~new_n9412_ | ~pi0972;
  assign new_n13076_ = ~new_n9411_ | ~new_n29813_;
  assign new_n13077_ = ~pi0813 | ~new_n12979_;
  assign new_n13078_ = ~new_n28903_ | ~new_n9428_;
  assign new_n13079_ = ~new_n9414_ | ~new_n30686_;
  assign new_n13080_ = ~new_n9413_ | ~new_n27635_;
  assign new_n13081_ = ~new_n9412_ | ~pi0973;
  assign new_n13082_ = ~new_n9411_ | ~new_n29812_;
  assign new_n13083_ = ~pi0814 | ~new_n12979_;
  assign new_n13084_ = ~new_n28902_ | ~new_n9428_;
  assign new_n13085_ = ~new_n9414_ | ~new_n30740_;
  assign new_n13086_ = ~new_n9413_ | ~new_n27634_;
  assign new_n13087_ = ~new_n9412_ | ~pi0974;
  assign new_n13088_ = ~new_n9411_ | ~new_n29811_;
  assign new_n13089_ = ~pi0815 | ~new_n12979_;
  assign new_n13090_ = ~new_n28901_ | ~new_n9428_;
  assign new_n13091_ = ~new_n9414_ | ~new_n30741_;
  assign new_n13092_ = ~new_n9413_ | ~new_n27633_;
  assign new_n13093_ = ~new_n9412_ | ~pi0975;
  assign new_n13094_ = ~new_n9411_ | ~new_n29810_;
  assign new_n13095_ = ~pi0816 | ~new_n12979_;
  assign new_n13096_ = ~new_n28900_ | ~new_n9428_;
  assign new_n13097_ = ~new_n9414_ | ~new_n30687_;
  assign new_n13098_ = ~new_n9413_ | ~new_n27632_;
  assign new_n13099_ = ~new_n9412_ | ~pi0976;
  assign new_n13100_ = ~new_n9411_ | ~new_n29809_;
  assign new_n13101_ = ~pi0817 | ~new_n12979_;
  assign new_n13102_ = ~new_n28899_ | ~new_n9428_;
  assign new_n13103_ = ~new_n9414_ | ~new_n30688_;
  assign new_n13104_ = ~new_n9413_ | ~new_n27631_;
  assign new_n13105_ = ~new_n9412_ | ~pi0977;
  assign new_n13106_ = ~new_n9411_ | ~new_n29808_;
  assign new_n13107_ = ~pi0818 | ~new_n12979_;
  assign new_n13108_ = ~new_n28898_ | ~new_n9428_;
  assign new_n13109_ = ~new_n9414_ | ~new_n30744_;
  assign new_n13110_ = ~new_n9413_ | ~new_n27630_;
  assign new_n13111_ = ~new_n9412_ | ~pi0978;
  assign new_n13112_ = ~new_n9411_ | ~new_n29807_;
  assign new_n13113_ = ~pi0819 | ~new_n12979_;
  assign new_n13114_ = ~new_n28897_ | ~new_n9428_;
  assign new_n13115_ = ~new_n9414_ | ~new_n30689_;
  assign new_n13116_ = ~new_n9413_ | ~new_n27629_;
  assign new_n13117_ = ~new_n9412_ | ~pi0979;
  assign new_n13118_ = ~new_n9411_ | ~new_n29806_;
  assign new_n13119_ = ~pi0820 | ~new_n12979_;
  assign new_n13120_ = ~new_n28896_ | ~new_n9428_;
  assign new_n13121_ = ~new_n9414_ | ~new_n30690_;
  assign new_n13122_ = ~new_n9413_ | ~new_n27628_;
  assign new_n13123_ = ~new_n9412_ | ~pi0980;
  assign new_n13124_ = ~new_n9411_ | ~new_n29805_;
  assign new_n13125_ = ~pi0821 | ~new_n12979_;
  assign new_n13126_ = ~new_n28895_ | ~new_n9428_;
  assign new_n13127_ = ~new_n9414_ | ~new_n30739_;
  assign new_n13128_ = ~new_n9413_ | ~new_n27627_;
  assign new_n13129_ = ~new_n9412_ | ~pi0981;
  assign new_n13130_ = ~new_n9411_ | ~new_n29804_;
  assign new_n13131_ = ~pi0822 | ~new_n12979_;
  assign new_n13132_ = ~new_n28894_ | ~new_n9428_;
  assign new_n13133_ = ~new_n9414_ | ~new_n30746_;
  assign new_n13134_ = ~new_n9413_ | ~new_n27626_;
  assign new_n13135_ = ~new_n9412_ | ~pi0982;
  assign new_n13136_ = ~new_n9411_ | ~new_n29803_;
  assign new_n13137_ = ~pi0823 | ~new_n12979_;
  assign new_n13138_ = ~new_n28893_ | ~new_n9428_;
  assign new_n13139_ = ~new_n9414_ | ~new_n30691_;
  assign new_n13140_ = ~new_n9413_ | ~new_n27625_;
  assign new_n13141_ = ~new_n9412_ | ~pi0983;
  assign new_n13142_ = ~new_n9411_ | ~new_n29802_;
  assign new_n13143_ = ~pi0824 | ~new_n12979_;
  assign new_n13144_ = ~new_n28892_ | ~new_n9428_;
  assign new_n13145_ = ~new_n9414_ | ~new_n30743_;
  assign new_n13146_ = ~new_n9413_ | ~new_n27624_;
  assign new_n13147_ = ~new_n9412_ | ~pi0984;
  assign new_n13148_ = ~new_n9411_ | ~new_n29801_;
  assign new_n13149_ = ~pi0825 | ~new_n12979_;
  assign new_n13150_ = ~new_n28891_ | ~new_n9428_;
  assign new_n13151_ = ~new_n9414_ | ~new_n30692_;
  assign new_n13152_ = ~new_n9413_ | ~new_n27623_;
  assign new_n13153_ = ~new_n9412_ | ~pi0985;
  assign new_n13154_ = ~new_n9411_ | ~new_n29800_;
  assign new_n13155_ = ~pi0826 | ~new_n12979_;
  assign new_n13156_ = ~new_n28890_ | ~new_n9428_;
  assign new_n13157_ = ~new_n9414_ | ~new_n30693_;
  assign new_n13158_ = ~new_n9413_ | ~new_n27622_;
  assign new_n13159_ = ~new_n9412_ | ~pi0986;
  assign new_n13160_ = ~new_n9411_ | ~new_n29799_;
  assign new_n13161_ = ~pi0827 | ~new_n12979_;
  assign new_n13162_ = ~new_n28888_ | ~new_n9428_;
  assign new_n13163_ = ~new_n9414_ | ~new_n30738_;
  assign new_n13164_ = ~new_n9413_ | ~new_n27621_;
  assign new_n13165_ = ~new_n9412_ | ~pi0987;
  assign new_n13166_ = ~new_n9411_ | ~new_n29797_;
  assign new_n13167_ = ~pi0828 | ~new_n12979_;
  assign new_n13168_ = ~new_n28887_ | ~new_n9428_;
  assign new_n13169_ = ~new_n9414_ | ~new_n30752_;
  assign new_n13170_ = ~new_n9413_ | ~new_n27620_;
  assign new_n13171_ = ~new_n9412_ | ~pi0988;
  assign new_n13172_ = ~new_n9411_ | ~new_n29711_;
  assign new_n13173_ = ~pi0829 | ~new_n12979_;
  assign new_n13174_ = ~new_n2973_ | ~new_n9657_;
  assign new_n13175_ = ~pi0908 | ~new_n9436_;
  assign new_n13176_ = ~new_n3070_ | ~new_n9435_;
  assign new_n13177_ = ~pi0830 | ~new_n10579_;
  assign new_n13178_ = ~pi0907 | ~new_n9436_;
  assign new_n13179_ = ~new_n3071_ | ~new_n9435_;
  assign new_n13180_ = ~pi0831 | ~new_n10579_;
  assign new_n13181_ = ~pi0906 | ~new_n9436_;
  assign new_n13182_ = ~new_n3072_ | ~new_n9435_;
  assign new_n13183_ = ~pi0832 | ~new_n10579_;
  assign new_n13184_ = ~pi0905 | ~new_n9436_;
  assign new_n13185_ = ~new_n3073_ | ~new_n9435_;
  assign new_n13186_ = ~pi0833 | ~new_n10579_;
  assign new_n13187_ = ~pi0904 | ~new_n9436_;
  assign new_n13188_ = ~new_n3074_ | ~new_n9435_;
  assign new_n13189_ = ~pi0834 | ~new_n10579_;
  assign new_n13190_ = ~pi0903 | ~new_n9436_;
  assign new_n13191_ = ~new_n3075_ | ~new_n9435_;
  assign new_n13192_ = ~pi0835 | ~new_n10579_;
  assign new_n13193_ = ~pi0902 | ~new_n9436_;
  assign new_n13194_ = ~new_n3045_ | ~new_n9435_;
  assign new_n13195_ = ~pi0836 | ~new_n10579_;
  assign new_n13196_ = ~pi0901 | ~new_n9436_;
  assign new_n13197_ = ~new_n3046_ | ~new_n9435_;
  assign new_n13198_ = ~pi0837 | ~new_n10579_;
  assign new_n13199_ = ~pi0900 | ~new_n9436_;
  assign new_n13200_ = ~new_n9435_ | ~new_n3047_;
  assign new_n13201_ = ~pi0838 | ~new_n10579_;
  assign new_n13202_ = ~pi0899 | ~new_n9436_;
  assign new_n13203_ = ~new_n9435_ | ~new_n3048_;
  assign new_n13204_ = ~pi0839 | ~new_n10579_;
  assign new_n13205_ = ~pi0898 | ~new_n9436_;
  assign new_n13206_ = ~new_n9435_ | ~new_n3049_;
  assign new_n13207_ = ~pi0840 | ~new_n10579_;
  assign new_n13208_ = ~pi0897 | ~new_n9436_;
  assign new_n13209_ = ~new_n9435_ | ~new_n3050_;
  assign new_n13210_ = ~pi0841 | ~new_n10579_;
  assign new_n13211_ = ~pi0896 | ~new_n9436_;
  assign new_n13212_ = ~new_n9435_ | ~new_n3051_;
  assign new_n13213_ = ~pi0842 | ~new_n10579_;
  assign new_n13214_ = ~pi0895 | ~new_n9436_;
  assign new_n13215_ = ~new_n9435_ | ~new_n3054_;
  assign new_n13216_ = ~pi0843 | ~new_n10579_;
  assign new_n13217_ = ~pi0894 | ~new_n9436_;
  assign new_n13218_ = ~new_n9435_ | ~new_n3065_;
  assign new_n13219_ = ~pi0844 | ~new_n10579_;
  assign new_n13220_ = ~pi0893 | ~new_n9436_;
  assign new_n13221_ = ~new_n9435_ | ~new_n3076_;
  assign new_n13222_ = ~pi0845 | ~new_n10579_;
  assign new_n13223_ = ~pi0923 | ~new_n9436_;
  assign new_n13224_ = ~new_n3071_ | ~new_n9435_;
  assign new_n13225_ = ~pi0846 | ~new_n10579_;
  assign new_n13226_ = ~pi0922 | ~new_n9436_;
  assign new_n13227_ = ~new_n3072_ | ~new_n9435_;
  assign new_n13228_ = ~pi0847 | ~new_n10579_;
  assign new_n13229_ = ~pi0921 | ~new_n9436_;
  assign new_n13230_ = ~new_n3073_ | ~new_n9435_;
  assign new_n13231_ = ~pi0848 | ~new_n10579_;
  assign new_n13232_ = ~pi0920 | ~new_n9436_;
  assign new_n13233_ = ~new_n3074_ | ~new_n9435_;
  assign new_n13234_ = ~pi0849 | ~new_n10579_;
  assign new_n13235_ = ~pi0919 | ~new_n9436_;
  assign new_n13236_ = ~new_n3075_ | ~new_n9435_;
  assign new_n13237_ = ~pi0850 | ~new_n10579_;
  assign new_n13238_ = ~pi0918 | ~new_n9436_;
  assign new_n13239_ = ~new_n3045_ | ~new_n9435_;
  assign new_n13240_ = ~pi0851 | ~new_n10579_;
  assign new_n13241_ = ~pi0917 | ~new_n9436_;
  assign new_n13242_ = ~new_n3046_ | ~new_n9435_;
  assign new_n13243_ = ~pi0852 | ~new_n10579_;
  assign new_n13244_ = ~pi0916 | ~new_n9436_;
  assign new_n13245_ = ~new_n9435_ | ~new_n3047_;
  assign new_n13246_ = ~pi0853 | ~new_n10579_;
  assign new_n13247_ = ~pi0915 | ~new_n9436_;
  assign new_n13248_ = ~new_n9435_ | ~new_n3048_;
  assign new_n13249_ = ~pi0854 | ~new_n10579_;
  assign new_n13250_ = ~pi0914 | ~new_n9436_;
  assign new_n13251_ = ~new_n9435_ | ~new_n3049_;
  assign new_n13252_ = ~pi0855 | ~new_n10579_;
  assign new_n13253_ = ~pi0913 | ~new_n9436_;
  assign new_n13254_ = ~new_n9435_ | ~new_n3050_;
  assign new_n13255_ = ~pi0856 | ~new_n10579_;
  assign new_n13256_ = ~pi0912 | ~new_n9436_;
  assign new_n13257_ = ~new_n9435_ | ~new_n3051_;
  assign new_n13258_ = ~pi0857 | ~new_n10579_;
  assign new_n13259_ = ~pi0911 | ~new_n9436_;
  assign new_n13260_ = ~new_n9435_ | ~new_n3054_;
  assign new_n13261_ = ~pi0858 | ~new_n10579_;
  assign new_n13262_ = ~pi0910 | ~new_n9436_;
  assign new_n13263_ = ~new_n9435_ | ~new_n3065_;
  assign new_n13264_ = ~pi0859 | ~new_n10579_;
  assign new_n13265_ = ~pi0909 | ~new_n9436_;
  assign new_n13266_ = ~new_n9435_ | ~new_n3076_;
  assign new_n13267_ = ~pi0860 | ~new_n10579_;
  assign new_n13268_ = ~new_n28599_ | ~new_n11098_ | ~new_n11462_;
  assign new_n13269_ = ~new_n11099_ | ~new_n9487_;
  assign new_n13270_ = ~new_n13269_ | ~new_n13268_;
  assign new_n13271_ = ~new_n11452_ | ~new_n13270_;
  assign new_n13272_ = ~new_n11508_ | ~pi0626;
  assign new_n13273_ = ~new_n10582_;
  assign new_n13274_ = ~new_n9471_ | ~pi0893;
  assign new_n13275_ = ~new_n9437_ | ~pi0845;
  assign new_n13276_ = ~pi0861 | ~new_n13273_;
  assign new_n13277_ = ~new_n9471_ | ~pi0894;
  assign new_n13278_ = ~new_n9437_ | ~pi0844;
  assign new_n13279_ = ~pi0862 | ~new_n13273_;
  assign new_n13280_ = ~new_n9471_ | ~pi0895;
  assign new_n13281_ = ~new_n9437_ | ~pi0843;
  assign new_n13282_ = ~pi0863 | ~new_n13273_;
  assign new_n13283_ = ~new_n9471_ | ~pi0896;
  assign new_n13284_ = ~new_n9437_ | ~pi0842;
  assign new_n13285_ = ~pi0864 | ~new_n13273_;
  assign new_n13286_ = ~new_n9471_ | ~pi0897;
  assign new_n13287_ = ~new_n9437_ | ~pi0841;
  assign new_n13288_ = ~pi0865 | ~new_n13273_;
  assign new_n13289_ = ~new_n9471_ | ~pi0898;
  assign new_n13290_ = ~new_n9437_ | ~pi0840;
  assign new_n13291_ = ~pi0866 | ~new_n13273_;
  assign new_n13292_ = ~new_n9471_ | ~pi0899;
  assign new_n13293_ = ~new_n9437_ | ~pi0839;
  assign new_n13294_ = ~pi0867 | ~new_n13273_;
  assign new_n13295_ = ~new_n9471_ | ~pi0900;
  assign new_n13296_ = ~new_n9437_ | ~pi0838;
  assign new_n13297_ = ~pi0868 | ~new_n13273_;
  assign new_n13298_ = ~new_n9471_ | ~pi0901;
  assign new_n13299_ = ~new_n9437_ | ~pi0837;
  assign new_n13300_ = ~pi0869 | ~new_n13273_;
  assign new_n13301_ = ~new_n9471_ | ~pi0902;
  assign new_n13302_ = ~new_n9437_ | ~pi0836;
  assign new_n13303_ = ~pi0870 | ~new_n13273_;
  assign new_n13304_ = ~new_n9471_ | ~pi0903;
  assign new_n13305_ = ~new_n9437_ | ~pi0835;
  assign new_n13306_ = ~pi0871 | ~new_n13273_;
  assign new_n13307_ = ~new_n9471_ | ~pi0904;
  assign new_n13308_ = ~new_n9437_ | ~pi0834;
  assign new_n13309_ = ~pi0872 | ~new_n13273_;
  assign new_n13310_ = ~new_n9471_ | ~pi0905;
  assign new_n13311_ = ~new_n9437_ | ~pi0833;
  assign new_n13312_ = ~pi0873 | ~new_n13273_;
  assign new_n13313_ = ~new_n9471_ | ~pi0906;
  assign new_n13314_ = ~new_n9437_ | ~pi0832;
  assign new_n13315_ = ~pi0874 | ~new_n13273_;
  assign new_n13316_ = ~new_n9471_ | ~pi0907;
  assign new_n13317_ = ~new_n9437_ | ~pi0831;
  assign new_n13318_ = ~pi0875 | ~new_n13273_;
  assign new_n13319_ = ~new_n9471_ | ~pi0908;
  assign new_n13320_ = ~new_n9437_ | ~pi0830;
  assign new_n13321_ = ~pi0876 | ~new_n13273_;
  assign new_n13322_ = ~new_n9476_ | ~pi0909;
  assign new_n13323_ = ~new_n9437_ | ~pi0860;
  assign new_n13324_ = ~pi0877 | ~new_n13273_;
  assign new_n13325_ = ~new_n9476_ | ~pi0910;
  assign new_n13326_ = ~new_n9437_ | ~pi0859;
  assign new_n13327_ = ~pi0878 | ~new_n13273_;
  assign new_n13328_ = ~new_n9476_ | ~pi0911;
  assign new_n13329_ = ~new_n9437_ | ~pi0858;
  assign new_n13330_ = ~pi0879 | ~new_n13273_;
  assign new_n13331_ = ~new_n9476_ | ~pi0912;
  assign new_n13332_ = ~new_n9437_ | ~pi0857;
  assign new_n13333_ = ~pi0880 | ~new_n13273_;
  assign new_n13334_ = ~new_n9476_ | ~pi0913;
  assign new_n13335_ = ~new_n9437_ | ~pi0856;
  assign new_n13336_ = ~pi0881 | ~new_n13273_;
  assign new_n13337_ = ~new_n9476_ | ~pi0914;
  assign new_n13338_ = ~new_n9437_ | ~pi0855;
  assign new_n13339_ = ~pi0882 | ~new_n13273_;
  assign new_n13340_ = ~new_n9476_ | ~pi0915;
  assign new_n13341_ = ~new_n9437_ | ~pi0854;
  assign new_n13342_ = ~pi0883 | ~new_n13273_;
  assign new_n13343_ = ~new_n9476_ | ~pi0916;
  assign new_n13344_ = ~new_n9437_ | ~pi0853;
  assign new_n13345_ = ~pi0884 | ~new_n13273_;
  assign new_n13346_ = ~new_n9476_ | ~pi0917;
  assign new_n13347_ = ~new_n9437_ | ~pi0852;
  assign new_n13348_ = ~pi0885 | ~new_n13273_;
  assign new_n13349_ = ~new_n9476_ | ~pi0918;
  assign new_n13350_ = ~new_n9437_ | ~pi0851;
  assign new_n13351_ = ~pi0886 | ~new_n13273_;
  assign new_n13352_ = ~new_n9476_ | ~pi0919;
  assign new_n13353_ = ~new_n9437_ | ~pi0850;
  assign new_n13354_ = ~pi0887 | ~new_n13273_;
  assign new_n13355_ = ~new_n9476_ | ~pi0920;
  assign new_n13356_ = ~new_n9437_ | ~pi0849;
  assign new_n13357_ = ~pi0888 | ~new_n13273_;
  assign new_n13358_ = ~new_n9476_ | ~pi0921;
  assign new_n13359_ = ~new_n9437_ | ~pi0848;
  assign new_n13360_ = ~pi0889 | ~new_n13273_;
  assign new_n13361_ = ~new_n9476_ | ~pi0922;
  assign new_n13362_ = ~new_n9437_ | ~pi0847;
  assign new_n13363_ = ~pi0890 | ~new_n13273_;
  assign new_n13364_ = ~new_n9476_ | ~pi0923;
  assign new_n13365_ = ~new_n9437_ | ~pi0846;
  assign new_n13366_ = ~pi0891 | ~new_n13273_;
  assign new_n13367_ = ~new_n9554_ | ~new_n10295_;
  assign new_n13368_ = ~new_n9474_ | ~new_n3076_;
  assign new_n13369_ = ~new_n27856_ | ~new_n9438_;
  assign new_n13370_ = ~new_n9421_ | ~new_n29204_;
  assign new_n13371_ = ~pi0893 | ~new_n10583_;
  assign new_n13372_ = ~new_n9474_ | ~new_n3065_;
  assign new_n13373_ = ~new_n27781_ | ~new_n9438_;
  assign new_n13374_ = ~new_n9421_ | ~new_n29187_;
  assign new_n13375_ = ~pi0894 | ~new_n10583_;
  assign new_n13376_ = ~new_n9474_ | ~new_n3054_;
  assign new_n13377_ = ~new_n27861_ | ~new_n9438_;
  assign new_n13378_ = ~new_n9421_ | ~new_n29213_;
  assign new_n13379_ = ~pi0895 | ~new_n10583_;
  assign new_n13380_ = ~new_n9474_ | ~new_n3051_;
  assign new_n13381_ = ~new_n27860_ | ~new_n9438_;
  assign new_n13382_ = ~new_n9421_ | ~new_n29211_;
  assign new_n13383_ = ~pi0896 | ~new_n10583_;
  assign new_n13384_ = ~new_n9474_ | ~new_n3050_;
  assign new_n13385_ = ~new_n27859_ | ~new_n9438_;
  assign new_n13386_ = ~new_n9421_ | ~new_n29210_;
  assign new_n13387_ = ~pi0897 | ~new_n10583_;
  assign new_n13388_ = ~new_n9474_ | ~new_n3049_;
  assign new_n13389_ = ~new_n27778_ | ~new_n9438_;
  assign new_n13390_ = ~new_n9421_ | ~new_n29209_;
  assign new_n13391_ = ~pi0898 | ~new_n10583_;
  assign new_n13392_ = ~new_n9474_ | ~new_n3048_;
  assign new_n13393_ = ~new_n27858_ | ~new_n9438_;
  assign new_n13394_ = ~new_n9421_ | ~new_n29208_;
  assign new_n13395_ = ~pi0899 | ~new_n10583_;
  assign new_n13396_ = ~new_n9474_ | ~new_n3047_;
  assign new_n13397_ = ~new_n27779_ | ~new_n9438_;
  assign new_n13398_ = ~new_n9421_ | ~new_n29207_;
  assign new_n13399_ = ~pi0900 | ~new_n10583_;
  assign new_n13400_ = ~new_n9474_ | ~new_n3046_;
  assign new_n13401_ = ~new_n27857_ | ~new_n9438_;
  assign new_n13402_ = ~new_n9421_ | ~new_n29206_;
  assign new_n13403_ = ~pi0901 | ~new_n10583_;
  assign new_n13404_ = ~new_n9474_ | ~new_n3045_;
  assign new_n13405_ = ~new_n27780_ | ~new_n9438_;
  assign new_n13406_ = ~new_n9421_ | ~new_n29205_;
  assign new_n13407_ = ~pi0902 | ~new_n10583_;
  assign new_n13408_ = ~new_n9474_ | ~new_n3075_;
  assign new_n13409_ = ~new_n27878_ | ~new_n9438_;
  assign new_n13410_ = ~new_n9421_ | ~new_n29233_;
  assign new_n13411_ = ~pi0903 | ~new_n10583_;
  assign new_n13412_ = ~new_n9474_ | ~new_n3074_;
  assign new_n13413_ = ~new_n27774_ | ~new_n9438_;
  assign new_n13414_ = ~new_n9421_ | ~new_n29232_;
  assign new_n13415_ = ~pi0904 | ~new_n10583_;
  assign new_n13416_ = ~new_n9474_ | ~new_n3073_;
  assign new_n13417_ = ~new_n27877_ | ~new_n9438_;
  assign new_n13418_ = ~new_n9421_ | ~new_n29231_;
  assign new_n13419_ = ~pi0905 | ~new_n10583_;
  assign new_n13420_ = ~new_n9474_ | ~new_n3072_;
  assign new_n13421_ = ~new_n27775_ | ~new_n9438_;
  assign new_n13422_ = ~new_n9421_ | ~new_n29230_;
  assign new_n13423_ = ~pi0906 | ~new_n10583_;
  assign new_n13424_ = ~new_n9474_ | ~new_n3071_;
  assign new_n13425_ = ~new_n27876_ | ~new_n9438_;
  assign new_n13426_ = ~new_n9421_ | ~new_n29229_;
  assign new_n13427_ = ~pi0907 | ~new_n10583_;
  assign new_n13428_ = ~new_n9474_ | ~new_n3070_;
  assign new_n13429_ = ~new_n27776_ | ~new_n9438_;
  assign new_n13430_ = ~new_n9421_ | ~new_n29228_;
  assign new_n13431_ = ~pi0908 | ~new_n10583_;
  assign new_n13432_ = ~new_n9475_ | ~new_n3076_;
  assign new_n13433_ = ~new_n9468_ | ~new_n3069_;
  assign new_n13434_ = ~new_n27875_ | ~new_n9438_;
  assign new_n13435_ = ~new_n9421_ | ~new_n29227_;
  assign new_n13436_ = ~pi0909 | ~new_n10583_;
  assign new_n13437_ = ~new_n9475_ | ~new_n3065_;
  assign new_n13438_ = ~new_n9468_ | ~new_n3068_;
  assign new_n13439_ = ~new_n27874_ | ~new_n9438_;
  assign new_n13440_ = ~new_n9421_ | ~new_n29226_;
  assign new_n13441_ = ~pi0910 | ~new_n10583_;
  assign new_n13442_ = ~new_n9475_ | ~new_n3054_;
  assign new_n13443_ = ~new_n9468_ | ~new_n3067_;
  assign new_n13444_ = ~new_n27873_ | ~new_n9438_;
  assign new_n13445_ = ~new_n9421_ | ~new_n29225_;
  assign new_n13446_ = ~pi0911 | ~new_n10583_;
  assign new_n13447_ = ~new_n9475_ | ~new_n3051_;
  assign new_n13448_ = ~new_n9468_ | ~new_n3066_;
  assign new_n13449_ = ~new_n27872_ | ~new_n9438_;
  assign new_n13450_ = ~new_n9421_ | ~new_n29224_;
  assign new_n13451_ = ~pi0912 | ~new_n10583_;
  assign new_n13452_ = ~new_n9475_ | ~new_n3050_;
  assign new_n13453_ = ~new_n9468_ | ~new_n3064_;
  assign new_n13454_ = ~new_n27871_ | ~new_n9438_;
  assign new_n13455_ = ~new_n9421_ | ~new_n29223_;
  assign new_n13456_ = ~pi0913 | ~new_n10583_;
  assign new_n13457_ = ~new_n9475_ | ~new_n3049_;
  assign new_n13458_ = ~new_n9468_ | ~new_n3063_;
  assign new_n13459_ = ~new_n27870_ | ~new_n9438_;
  assign new_n13460_ = ~new_n9421_ | ~new_n29222_;
  assign new_n13461_ = ~pi0914 | ~new_n10583_;
  assign new_n13462_ = ~new_n9475_ | ~new_n3048_;
  assign new_n13463_ = ~new_n9468_ | ~new_n3062_;
  assign new_n13464_ = ~new_n27869_ | ~new_n9438_;
  assign new_n13465_ = ~new_n9421_ | ~new_n29221_;
  assign new_n13466_ = ~pi0915 | ~new_n10583_;
  assign new_n13467_ = ~new_n9475_ | ~new_n3047_;
  assign new_n13468_ = ~new_n9468_ | ~new_n3061_;
  assign new_n13469_ = ~new_n27868_ | ~new_n9438_;
  assign new_n13470_ = ~new_n9421_ | ~new_n29220_;
  assign new_n13471_ = ~pi0916 | ~new_n10583_;
  assign new_n13472_ = ~new_n9475_ | ~new_n3046_;
  assign new_n13473_ = ~new_n9468_ | ~new_n3060_;
  assign new_n13474_ = ~new_n27867_ | ~new_n9438_;
  assign new_n13475_ = ~new_n9421_ | ~new_n29219_;
  assign new_n13476_ = ~pi0917 | ~new_n10583_;
  assign new_n13477_ = ~new_n9475_ | ~new_n3045_;
  assign new_n13478_ = ~new_n9468_ | ~new_n3059_;
  assign new_n13479_ = ~new_n27866_ | ~new_n9438_;
  assign new_n13480_ = ~new_n9421_ | ~new_n29218_;
  assign new_n13481_ = ~pi0918 | ~new_n10583_;
  assign new_n13482_ = ~new_n9475_ | ~new_n3075_;
  assign new_n13483_ = ~new_n9468_ | ~new_n3058_;
  assign new_n13484_ = ~new_n27865_ | ~new_n9438_;
  assign new_n13485_ = ~new_n9421_ | ~new_n29217_;
  assign new_n13486_ = ~pi0919 | ~new_n10583_;
  assign new_n13487_ = ~new_n9475_ | ~new_n3074_;
  assign new_n13488_ = ~new_n9468_ | ~new_n3057_;
  assign new_n13489_ = ~new_n27864_ | ~new_n9438_;
  assign new_n13490_ = ~new_n9421_ | ~new_n29216_;
  assign new_n13491_ = ~pi0920 | ~new_n10583_;
  assign new_n13492_ = ~new_n9475_ | ~new_n3073_;
  assign new_n13493_ = ~new_n9468_ | ~new_n3056_;
  assign new_n13494_ = ~new_n27863_ | ~new_n9438_;
  assign new_n13495_ = ~new_n9421_ | ~new_n29215_;
  assign new_n13496_ = ~pi0921 | ~new_n10583_;
  assign new_n13497_ = ~new_n9475_ | ~new_n3072_;
  assign new_n13498_ = ~new_n9468_ | ~new_n3055_;
  assign new_n13499_ = ~new_n27862_ | ~new_n9438_;
  assign new_n13500_ = ~new_n9421_ | ~new_n29214_;
  assign new_n13501_ = ~pi0922 | ~new_n10583_;
  assign new_n13502_ = ~new_n9475_ | ~new_n3071_;
  assign new_n13503_ = ~new_n9468_ | ~new_n3053_;
  assign new_n13504_ = ~new_n27777_ | ~new_n9438_;
  assign new_n13505_ = ~new_n9421_ | ~new_n29212_;
  assign new_n13506_ = ~pi0923 | ~new_n10583_;
  assign new_n13507_ = ~new_n9468_ | ~new_n3052_;
  assign new_n13508_ = ~new_n9421_ | ~new_n29186_;
  assign new_n13509_ = ~pi0924 | ~new_n10583_;
  assign new_n13510_ = ~new_n11476_ | ~new_n10338_;
  assign new_n13511_ = ~new_n10619_ | ~new_n13510_;
  assign new_n13512_ = ~new_n9434_ | ~new_n28362_;
  assign new_n13513_ = ~new_n9420_ | ~new_n27642_;
  assign new_n13514_ = ~pi0925 | ~new_n10584_;
  assign new_n13515_ = ~new_n9434_ | ~new_n28361_;
  assign new_n13516_ = ~new_n9420_ | ~new_n27553_;
  assign new_n13517_ = ~pi0926 | ~new_n10584_;
  assign new_n13518_ = ~new_n9434_ | ~new_n28333_;
  assign new_n13519_ = ~new_n9420_ | ~new_n27644_;
  assign new_n13520_ = ~pi0927 | ~new_n10584_;
  assign new_n13521_ = ~new_n9434_ | ~new_n28369_;
  assign new_n13522_ = ~new_n9420_ | ~new_n27643_;
  assign new_n13523_ = ~pi0928 | ~new_n10584_;
  assign new_n13524_ = ~new_n28368_ | ~new_n9434_;
  assign new_n13525_ = ~new_n9420_ | ~new_n27646_;
  assign new_n13526_ = ~pi0929 | ~new_n10584_;
  assign new_n13527_ = ~new_n28367_ | ~new_n9434_;
  assign new_n13528_ = ~new_n9420_ | ~new_n27619_;
  assign new_n13529_ = ~pi0930 | ~new_n10584_;
  assign new_n13530_ = ~new_n28366_ | ~new_n9434_;
  assign new_n13531_ = ~new_n9420_ | ~new_n27618_;
  assign new_n13532_ = ~pi0931 | ~new_n10584_;
  assign new_n13533_ = ~new_n28365_ | ~new_n9434_;
  assign new_n13534_ = ~new_n9420_ | ~new_n27617_;
  assign new_n13535_ = ~pi0932 | ~new_n10584_;
  assign new_n13536_ = ~new_n28364_ | ~new_n9434_;
  assign new_n13537_ = ~new_n9420_ | ~new_n27616_;
  assign new_n13538_ = ~pi0933 | ~new_n10584_;
  assign new_n13539_ = ~new_n28363_ | ~new_n9434_;
  assign new_n13540_ = ~new_n9420_ | ~new_n27615_;
  assign new_n13541_ = ~pi0934 | ~new_n10584_;
  assign new_n13542_ = ~new_n28389_ | ~new_n9434_;
  assign new_n13543_ = ~new_n9420_ | ~new_n27641_;
  assign new_n13544_ = ~pi0935 | ~new_n10584_;
  assign new_n13545_ = ~new_n28388_ | ~new_n9434_;
  assign new_n13546_ = ~new_n9420_ | ~new_n27640_;
  assign new_n13547_ = ~pi0936 | ~new_n10584_;
  assign new_n13548_ = ~new_n28387_ | ~new_n9434_;
  assign new_n13549_ = ~new_n9420_ | ~new_n27639_;
  assign new_n13550_ = ~pi0937 | ~new_n10584_;
  assign new_n13551_ = ~new_n28386_ | ~new_n9434_;
  assign new_n13552_ = ~new_n9420_ | ~new_n27638_;
  assign new_n13553_ = ~pi0938 | ~new_n10584_;
  assign new_n13554_ = ~new_n28385_ | ~new_n9434_;
  assign new_n13555_ = ~new_n9420_ | ~new_n27637_;
  assign new_n13556_ = ~pi0939 | ~new_n10584_;
  assign new_n13557_ = ~new_n28384_ | ~new_n9434_;
  assign new_n13558_ = ~new_n9420_ | ~new_n27636_;
  assign new_n13559_ = ~pi0940 | ~new_n10584_;
  assign new_n13560_ = ~new_n28383_ | ~new_n9434_;
  assign new_n13561_ = ~new_n9420_ | ~new_n27635_;
  assign new_n13562_ = ~pi0941 | ~new_n10584_;
  assign new_n13563_ = ~new_n28382_ | ~new_n9434_;
  assign new_n13564_ = ~new_n9420_ | ~new_n27634_;
  assign new_n13565_ = ~pi0942 | ~new_n10584_;
  assign new_n13566_ = ~new_n28381_ | ~new_n9434_;
  assign new_n13567_ = ~new_n9420_ | ~new_n27633_;
  assign new_n13568_ = ~pi0943 | ~new_n10584_;
  assign new_n13569_ = ~new_n28380_ | ~new_n9434_;
  assign new_n13570_ = ~new_n9420_ | ~new_n27632_;
  assign new_n13571_ = ~pi0944 | ~new_n10584_;
  assign new_n13572_ = ~new_n28379_ | ~new_n9434_;
  assign new_n13573_ = ~new_n9420_ | ~new_n27631_;
  assign new_n13574_ = ~pi0945 | ~new_n10584_;
  assign new_n13575_ = ~new_n28378_ | ~new_n9434_;
  assign new_n13576_ = ~new_n9420_ | ~new_n27630_;
  assign new_n13577_ = ~pi0946 | ~new_n10584_;
  assign new_n13578_ = ~new_n28377_ | ~new_n9434_;
  assign new_n13579_ = ~new_n9420_ | ~new_n27629_;
  assign new_n13580_ = ~pi0947 | ~new_n10584_;
  assign new_n13581_ = ~new_n28376_ | ~new_n9434_;
  assign new_n13582_ = ~new_n9420_ | ~new_n27628_;
  assign new_n13583_ = ~pi0948 | ~new_n10584_;
  assign new_n13584_ = ~new_n28375_ | ~new_n9434_;
  assign new_n13585_ = ~new_n9420_ | ~new_n27627_;
  assign new_n13586_ = ~pi0949 | ~new_n10584_;
  assign new_n13587_ = ~new_n28374_ | ~new_n9434_;
  assign new_n13588_ = ~new_n9420_ | ~new_n27626_;
  assign new_n13589_ = ~pi0950 | ~new_n10584_;
  assign new_n13590_ = ~new_n28373_ | ~new_n9434_;
  assign new_n13591_ = ~new_n9420_ | ~new_n27625_;
  assign new_n13592_ = ~pi0951 | ~new_n10584_;
  assign new_n13593_ = ~new_n28372_ | ~new_n9434_;
  assign new_n13594_ = ~new_n9420_ | ~new_n27624_;
  assign new_n13595_ = ~pi0952 | ~new_n10584_;
  assign new_n13596_ = ~new_n28371_ | ~new_n9434_;
  assign new_n13597_ = ~new_n9420_ | ~new_n27623_;
  assign new_n13598_ = ~pi0953 | ~new_n10584_;
  assign new_n13599_ = ~new_n28370_ | ~new_n9434_;
  assign new_n13600_ = ~new_n9420_ | ~new_n27622_;
  assign new_n13601_ = ~pi0954 | ~new_n10584_;
  assign new_n13602_ = ~new_n28334_ | ~new_n9434_;
  assign new_n13603_ = ~new_n9420_ | ~new_n27621_;
  assign new_n13604_ = ~pi0955 | ~new_n10584_;
  assign new_n13605_ = ~new_n9420_ | ~new_n27620_;
  assign new_n13606_ = ~pi0956 | ~new_n10584_;
  assign new_n13607_ = ~new_n30327_ | ~new_n11644_;
  assign new_n13608_ = ~new_n11474_ | ~new_n28599_;
  assign new_n13609_ = ~new_n13608_ | ~new_n13607_;
  assign new_n13610_ = ~new_n11502_ | ~new_n10325_;
  assign new_n13611_ = ~new_n10587_;
  assign new_n13612_ = ~new_n10586_;
  assign new_n13613_ = pi0996 | new_n2973_;
  assign new_n13614_ = ~new_n30527_ | ~new_n9628_;
  assign new_n13615_ = ~new_n9629_ | ~new_n29204_;
  assign new_n13616_ = ~pi0925 | ~new_n14784_;
  assign new_n13617_ = ~new_n9478_ | ~new_n28362_;
  assign new_n13618_ = ~new_n9433_ | ~new_n27642_;
  assign new_n13619_ = ~new_n9424_ | ~pi0798;
  assign new_n13620_ = ~new_n9423_ | ~new_n10724_;
  assign new_n13621_ = ~new_n9419_ | ~pi0798;
  assign new_n13622_ = ~new_n13611_ | ~pi0957;
  assign new_n13623_ = ~new_n30549_ | ~new_n9628_;
  assign new_n13624_ = ~new_n9629_ | ~new_n29187_;
  assign new_n13625_ = ~pi0926 | ~new_n14784_;
  assign new_n13626_ = ~new_n9478_ | ~new_n28361_;
  assign new_n13627_ = ~new_n9433_ | ~new_n27553_;
  assign new_n13628_ = ~new_n9424_ | ~new_n28823_;
  assign new_n13629_ = ~new_n9423_ | ~new_n29599_;
  assign new_n13630_ = ~new_n9419_ | ~pi0799;
  assign new_n13631_ = ~new_n13611_ | ~pi0958;
  assign new_n13632_ = ~new_n30571_ | ~new_n9628_;
  assign new_n13633_ = ~new_n9629_ | ~new_n29213_;
  assign new_n13634_ = ~pi0927 | ~new_n14784_;
  assign new_n13635_ = ~new_n9478_ | ~new_n28333_;
  assign new_n13636_ = ~new_n9433_ | ~new_n27644_;
  assign new_n13637_ = ~new_n9424_ | ~new_n28889_;
  assign new_n13638_ = ~new_n29567_ | ~new_n9423_;
  assign new_n13639_ = ~new_n9419_ | ~pi0800;
  assign new_n13640_ = ~new_n13611_ | ~pi0959;
  assign new_n13641_ = ~new_n30523_ | ~new_n9628_;
  assign new_n13642_ = ~new_n9629_ | ~new_n29211_;
  assign new_n13643_ = ~pi0928 | ~new_n14784_;
  assign new_n13644_ = ~new_n9478_ | ~new_n28369_;
  assign new_n13645_ = ~new_n9433_ | ~new_n27643_;
  assign new_n13646_ = ~new_n9424_ | ~new_n28886_;
  assign new_n13647_ = ~new_n29609_ | ~new_n9423_;
  assign new_n13648_ = ~new_n9419_ | ~pi0801;
  assign new_n13649_ = ~new_n13611_ | ~pi0960;
  assign new_n13650_ = ~new_n30566_ | ~new_n9628_;
  assign new_n13651_ = ~new_n9629_ | ~new_n29210_;
  assign new_n13652_ = ~pi0929 | ~new_n14784_;
  assign new_n13653_ = ~new_n9478_ | ~new_n28368_;
  assign new_n13654_ = ~new_n9433_ | ~new_n27646_;
  assign new_n13655_ = ~new_n9424_ | ~new_n28885_;
  assign new_n13656_ = ~new_n29568_ | ~new_n9423_;
  assign new_n13657_ = ~new_n9419_ | ~pi0802;
  assign new_n13658_ = ~new_n13611_ | ~pi0961;
  assign new_n13659_ = ~new_n30524_ | ~new_n9628_;
  assign new_n13660_ = ~new_n9629_ | ~new_n29209_;
  assign new_n13661_ = ~pi0930 | ~new_n14784_;
  assign new_n13662_ = ~new_n9478_ | ~new_n28367_;
  assign new_n13663_ = ~new_n9433_ | ~new_n27619_;
  assign new_n13664_ = ~new_n9424_ | ~new_n28884_;
  assign new_n13665_ = ~new_n29607_ | ~new_n9423_;
  assign new_n13666_ = ~new_n9419_ | ~pi0803;
  assign new_n13667_ = ~new_n13611_ | ~pi0962;
  assign new_n13668_ = ~new_n30564_ | ~new_n9628_;
  assign new_n13669_ = ~new_n9629_ | ~new_n29208_;
  assign new_n13670_ = ~pi0931 | ~new_n14784_;
  assign new_n13671_ = ~new_n9433_ | ~new_n27618_;
  assign new_n13672_ = ~new_n9424_ | ~new_n28883_;
  assign new_n13673_ = ~new_n29569_ | ~new_n9423_;
  assign new_n13674_ = ~new_n9419_ | ~pi0804;
  assign new_n13675_ = ~new_n13611_ | ~pi0963;
  assign new_n13676_ = ~new_n30525_ | ~new_n9628_;
  assign new_n13677_ = ~new_n9629_ | ~new_n29207_;
  assign new_n13678_ = ~pi0932 | ~new_n14784_;
  assign new_n13679_ = ~new_n9433_ | ~new_n27617_;
  assign new_n13680_ = ~new_n9424_ | ~new_n28882_;
  assign new_n13681_ = ~new_n29605_ | ~new_n9423_;
  assign new_n13682_ = ~new_n9419_ | ~pi0805;
  assign new_n13683_ = ~new_n13611_ | ~pi0964;
  assign new_n13684_ = ~new_n30562_ | ~new_n9628_;
  assign new_n13685_ = ~new_n9629_ | ~new_n29206_;
  assign new_n13686_ = ~pi0933 | ~new_n14784_;
  assign new_n13687_ = ~new_n9433_ | ~new_n27616_;
  assign new_n13688_ = ~new_n9424_ | ~new_n28881_;
  assign new_n13689_ = ~new_n29570_ | ~new_n9423_;
  assign new_n13690_ = ~new_n9419_ | ~pi0806;
  assign new_n13691_ = ~new_n13611_ | ~pi0965;
  assign new_n13692_ = ~new_n30526_ | ~new_n9628_;
  assign new_n13693_ = ~new_n9629_ | ~new_n29205_;
  assign new_n13694_ = ~pi0934 | ~new_n14784_;
  assign new_n13695_ = ~new_n9433_ | ~new_n27615_;
  assign new_n13696_ = ~new_n9424_ | ~new_n28880_;
  assign new_n13697_ = ~new_n29603_ | ~new_n9423_;
  assign new_n13698_ = ~new_n9419_ | ~pi0807;
  assign new_n13699_ = ~new_n13611_ | ~pi0966;
  assign new_n13700_ = ~new_n30593_ | ~new_n9628_;
  assign new_n13701_ = ~new_n9629_ | ~new_n29233_;
  assign new_n13702_ = ~pi0935 | ~new_n14784_;
  assign new_n13703_ = ~new_n9433_ | ~new_n27641_;
  assign new_n13704_ = ~new_n9424_ | ~new_n28909_;
  assign new_n13705_ = ~new_n29556_ | ~new_n9423_;
  assign new_n13706_ = ~new_n9419_ | ~pi0808;
  assign new_n13707_ = ~new_n13611_ | ~pi0967;
  assign new_n13708_ = ~new_n30512_ | ~new_n9628_;
  assign new_n13709_ = ~new_n9629_ | ~new_n29232_;
  assign new_n13710_ = ~pi0936 | ~new_n14784_;
  assign new_n13711_ = ~new_n9433_ | ~new_n27640_;
  assign new_n13712_ = ~new_n9424_ | ~new_n28908_;
  assign new_n13713_ = ~new_n29632_ | ~new_n9423_;
  assign new_n13714_ = ~new_n9419_ | ~pi0809;
  assign new_n13715_ = ~new_n13611_ | ~pi0968;
  assign new_n13716_ = ~new_n30591_ | ~new_n9628_;
  assign new_n13717_ = ~new_n9629_ | ~new_n29231_;
  assign new_n13718_ = ~pi0937 | ~new_n14784_;
  assign new_n13719_ = ~new_n9433_ | ~new_n27639_;
  assign new_n13720_ = ~new_n9424_ | ~new_n28907_;
  assign new_n13721_ = ~new_n29557_ | ~new_n9423_;
  assign new_n13722_ = ~new_n9419_ | ~pi0810;
  assign new_n13723_ = ~new_n13611_ | ~pi0969;
  assign new_n13724_ = ~new_n30513_ | ~new_n9628_;
  assign new_n13725_ = ~new_n9629_ | ~new_n29230_;
  assign new_n13726_ = ~pi0938 | ~new_n14784_;
  assign new_n13727_ = ~new_n9433_ | ~new_n27638_;
  assign new_n13728_ = ~new_n9424_ | ~new_n28906_;
  assign new_n13729_ = ~new_n29630_ | ~new_n9423_;
  assign new_n13730_ = ~new_n9419_ | ~pi0811;
  assign new_n13731_ = ~new_n13611_ | ~pi0970;
  assign new_n13732_ = ~new_n30589_ | ~new_n9628_;
  assign new_n13733_ = ~new_n9629_ | ~new_n29229_;
  assign new_n13734_ = ~pi0939 | ~new_n14784_;
  assign new_n13735_ = ~new_n9433_ | ~new_n27637_;
  assign new_n13736_ = ~new_n9424_ | ~new_n28905_;
  assign new_n13737_ = ~new_n29558_ | ~new_n9423_;
  assign new_n13738_ = ~new_n9419_ | ~pi0812;
  assign new_n13739_ = ~new_n13611_ | ~pi0971;
  assign new_n13740_ = ~new_n30514_ | ~new_n9628_;
  assign new_n13741_ = ~new_n9629_ | ~new_n29228_;
  assign new_n13742_ = ~pi0940 | ~new_n14784_;
  assign new_n13743_ = ~new_n9433_ | ~new_n27636_;
  assign new_n13744_ = ~new_n9424_ | ~new_n28904_;
  assign new_n13745_ = ~new_n29628_ | ~new_n9423_;
  assign new_n13746_ = ~new_n9419_ | ~pi0813;
  assign new_n13747_ = ~new_n13611_ | ~pi0972;
  assign new_n13748_ = ~new_n30587_ | ~new_n9628_;
  assign new_n13749_ = ~new_n9629_ | ~new_n29227_;
  assign new_n13750_ = ~pi0941 | ~new_n14784_;
  assign new_n13751_ = ~new_n9433_ | ~new_n27635_;
  assign new_n13752_ = ~new_n9424_ | ~new_n28903_;
  assign new_n13753_ = ~new_n29559_ | ~new_n9423_;
  assign new_n13754_ = ~new_n9419_ | ~pi0814;
  assign new_n13755_ = ~new_n13611_ | ~pi0973;
  assign new_n13756_ = ~new_n30515_ | ~new_n9628_;
  assign new_n13757_ = ~new_n9629_ | ~new_n29226_;
  assign new_n13758_ = ~pi0942 | ~new_n14784_;
  assign new_n13759_ = ~new_n9433_ | ~new_n27634_;
  assign new_n13760_ = ~new_n9424_ | ~new_n28902_;
  assign new_n13761_ = ~new_n29626_ | ~new_n9423_;
  assign new_n13762_ = ~new_n9419_ | ~pi0815;
  assign new_n13763_ = ~new_n13611_ | ~pi0974;
  assign new_n13764_ = ~new_n30585_ | ~new_n9628_;
  assign new_n13765_ = ~new_n9629_ | ~new_n29225_;
  assign new_n13766_ = ~pi0943 | ~new_n14784_;
  assign new_n13767_ = ~new_n9433_ | ~new_n27633_;
  assign new_n13768_ = ~new_n9424_ | ~new_n28901_;
  assign new_n13769_ = ~new_n29560_ | ~new_n9423_;
  assign new_n13770_ = ~new_n9419_ | ~pi0816;
  assign new_n13771_ = ~new_n13611_ | ~pi0975;
  assign new_n13772_ = ~new_n30516_ | ~new_n9628_;
  assign new_n13773_ = ~new_n9629_ | ~new_n29224_;
  assign new_n13774_ = ~pi0944 | ~new_n14784_;
  assign new_n13775_ = ~new_n9433_ | ~new_n27632_;
  assign new_n13776_ = ~new_n9424_ | ~new_n28900_;
  assign new_n13777_ = ~new_n29624_ | ~new_n9423_;
  assign new_n13778_ = ~new_n9419_ | ~pi0817;
  assign new_n13779_ = ~new_n13611_ | ~pi0976;
  assign new_n13780_ = ~new_n30581_ | ~new_n9628_;
  assign new_n13781_ = ~new_n9629_ | ~new_n29223_;
  assign new_n13782_ = ~pi0945 | ~new_n14784_;
  assign new_n13783_ = ~new_n9433_ | ~new_n27631_;
  assign new_n13784_ = ~new_n9424_ | ~new_n28899_;
  assign new_n13785_ = ~new_n29561_ | ~new_n9423_;
  assign new_n13786_ = ~new_n9419_ | ~pi0818;
  assign new_n13787_ = ~new_n13611_ | ~pi0977;
  assign new_n13788_ = ~new_n30517_ | ~new_n9628_;
  assign new_n13789_ = ~new_n9629_ | ~new_n29222_;
  assign new_n13790_ = ~pi0946 | ~new_n14784_;
  assign new_n13791_ = ~new_n9433_ | ~new_n27630_;
  assign new_n13792_ = ~new_n9424_ | ~new_n28898_;
  assign new_n13793_ = ~new_n29620_ | ~new_n9423_;
  assign new_n13794_ = ~new_n9419_ | ~pi0819;
  assign new_n13795_ = ~new_n13611_ | ~pi0978;
  assign new_n13796_ = ~new_n30579_ | ~new_n9628_;
  assign new_n13797_ = ~new_n9629_ | ~new_n29221_;
  assign new_n13798_ = ~pi0947 | ~new_n14784_;
  assign new_n13799_ = ~new_n9433_ | ~new_n27629_;
  assign new_n13800_ = ~new_n9424_ | ~new_n28897_;
  assign new_n13801_ = ~new_n29562_ | ~new_n9423_;
  assign new_n13802_ = ~new_n9419_ | ~pi0820;
  assign new_n13803_ = ~new_n13611_ | ~pi0979;
  assign new_n13804_ = ~new_n30518_ | ~new_n9628_;
  assign new_n13805_ = ~new_n9629_ | ~new_n29220_;
  assign new_n13806_ = ~pi0948 | ~new_n14784_;
  assign new_n13807_ = ~new_n9433_ | ~new_n27628_;
  assign new_n13808_ = ~new_n9424_ | ~new_n28896_;
  assign new_n13809_ = ~new_n29618_ | ~new_n9423_;
  assign new_n13810_ = ~new_n9419_ | ~pi0821;
  assign new_n13811_ = ~new_n13611_ | ~pi0980;
  assign new_n13812_ = ~new_n30577_ | ~new_n9628_;
  assign new_n13813_ = ~new_n9629_ | ~new_n29219_;
  assign new_n13814_ = ~pi0949 | ~new_n14784_;
  assign new_n13815_ = ~new_n9433_ | ~new_n27627_;
  assign new_n13816_ = ~new_n9424_ | ~new_n28895_;
  assign new_n13817_ = ~new_n29563_ | ~new_n9423_;
  assign new_n13818_ = ~new_n9419_ | ~pi0822;
  assign new_n13819_ = ~new_n13611_ | ~pi0981;
  assign new_n13820_ = ~new_n30519_ | ~new_n9628_;
  assign new_n13821_ = ~new_n9629_ | ~new_n29218_;
  assign new_n13822_ = ~pi0950 | ~new_n14784_;
  assign new_n13823_ = ~new_n9433_ | ~new_n27626_;
  assign new_n13824_ = ~new_n9424_ | ~new_n28894_;
  assign new_n13825_ = ~new_n29616_ | ~new_n9423_;
  assign new_n13826_ = ~new_n9419_ | ~pi0823;
  assign new_n13827_ = ~new_n13611_ | ~pi0982;
  assign new_n13828_ = ~new_n30575_ | ~new_n9628_;
  assign new_n13829_ = ~new_n9629_ | ~new_n29217_;
  assign new_n13830_ = ~pi0951 | ~new_n14784_;
  assign new_n13831_ = ~new_n9433_ | ~new_n27625_;
  assign new_n13832_ = ~new_n9424_ | ~new_n28893_;
  assign new_n13833_ = ~new_n29564_ | ~new_n9423_;
  assign new_n13834_ = ~new_n9419_ | ~pi0824;
  assign new_n13835_ = ~new_n13611_ | ~pi0983;
  assign new_n13836_ = ~new_n30520_ | ~new_n9628_;
  assign new_n13837_ = ~new_n9629_ | ~new_n29216_;
  assign new_n13838_ = ~pi0952 | ~new_n14784_;
  assign new_n13839_ = ~new_n9433_ | ~new_n27624_;
  assign new_n13840_ = ~new_n9424_ | ~new_n28892_;
  assign new_n13841_ = ~new_n29614_ | ~new_n9423_;
  assign new_n13842_ = ~new_n9419_ | ~pi0825;
  assign new_n13843_ = ~new_n13611_ | ~pi0984;
  assign new_n13844_ = ~new_n30573_ | ~new_n9628_;
  assign new_n13845_ = ~new_n9629_ | ~new_n29215_;
  assign new_n13846_ = ~pi0953 | ~new_n14784_;
  assign new_n13847_ = ~new_n9433_ | ~new_n27623_;
  assign new_n13848_ = ~new_n9424_ | ~new_n28891_;
  assign new_n13849_ = ~new_n29565_ | ~new_n9423_;
  assign new_n13850_ = ~new_n9419_ | ~pi0826;
  assign new_n13851_ = ~new_n13611_ | ~pi0985;
  assign new_n13852_ = ~new_n30521_ | ~new_n9628_;
  assign new_n13853_ = ~new_n9629_ | ~new_n29214_;
  assign new_n13854_ = ~pi0954 | ~new_n14784_;
  assign new_n13855_ = ~new_n9433_ | ~new_n27622_;
  assign new_n13856_ = ~new_n9424_ | ~new_n28890_;
  assign new_n13857_ = ~new_n29566_ | ~new_n9423_;
  assign new_n13858_ = ~new_n9419_ | ~pi0827;
  assign new_n13859_ = ~new_n13611_ | ~pi0986;
  assign new_n13860_ = ~new_n30522_ | ~new_n9628_;
  assign new_n13861_ = ~new_n9629_ | ~new_n29212_;
  assign new_n13862_ = ~pi0955 | ~new_n14784_;
  assign new_n13863_ = ~new_n9433_ | ~new_n27621_;
  assign new_n13864_ = ~new_n9424_ | ~new_n28888_;
  assign new_n13865_ = ~new_n29612_ | ~new_n9423_;
  assign new_n13866_ = ~new_n9419_ | ~pi0828;
  assign new_n13867_ = ~new_n13611_ | ~pi0987;
  assign new_n13868_ = ~new_n30569_ | ~new_n9628_;
  assign new_n13869_ = ~new_n9629_ | ~new_n29186_;
  assign new_n13870_ = ~pi0956 | ~new_n14784_;
  assign new_n13871_ = ~new_n9433_ | ~new_n27620_;
  assign new_n13872_ = ~new_n9424_ | ~new_n28887_;
  assign new_n13873_ = ~new_n29600_ | ~new_n9423_;
  assign new_n13874_ = ~new_n9419_ | ~pi0829;
  assign new_n13875_ = ~new_n13611_ | ~pi0988;
  assign new_n13876_ = ~pi0593 | ~pi0592;
  assign new_n13877_ = ~new_n11518_ | ~pi0957;
  assign new_n13878_ = ~pi0991 | ~new_n10588_;
  assign new_n13879_ = ~new_n11441_;
  assign new_n13880_ = ~new_n11440_ | ~new_n11467_ | ~new_n11509_;
  assign new_n13881_ = ~pi0994 | ~new_n11441_;
  assign new_n13882_ = ~new_n11228_ | ~new_n11508_;
  assign new_n13883_ = ~new_n11507_ | ~new_n10325_;
  assign new_n13884_ = ~new_n11443_;
  assign new_n13885_ = ~new_n11452_ | ~pi0996;
  assign new_n13886_ = ~new_n9756_;
  assign new_n13887_ = ~new_n9756_ | ~new_n10577_;
  assign new_n13888_ = ~new_n11452_ | ~new_n10306_;
  assign new_n13889_ = ~new_n11225_ | ~new_n9397_;
  assign new_n13890_ = ~new_n11459_ | ~new_n13888_;
  assign new_n13891_ = ~new_n2973_ | ~new_n13887_;
  assign new_n13892_ = pi0625 | pi0626;
  assign new_n13893_ = ~new_n11227_ | ~new_n13892_ | ~new_n13891_;
  assign new_n13894_ = ~new_n9415_ | ~new_n9500_;
  assign new_n13895_ = ~pi1000 | ~new_n13894_;
  assign new_n13896_ = ~new_n11502_ | ~pi0627;
  assign new_n13897_ = ~pi1001 | ~pi0591;
  assign new_n13898_ = ~new_n11444_;
  assign new_n13899_ = ~new_n10335_ | ~pi0625 | ~new_n10327_;
  assign new_n13900_ = ~new_n11445_ | ~new_n11462_ | ~new_n11509_;
  assign new_n13901_ = ~new_n11230_ | ~new_n9487_;
  assign new_n13902_ = ~pi1003 | ~new_n13900_;
  assign new_n13903_ = ~new_n9579_ | ~pi0684;
  assign new_n13904_ = ~new_n9578_ | ~pi0676;
  assign new_n13905_ = ~new_n9577_ | ~pi0668;
  assign new_n13906_ = ~new_n9576_ | ~pi0660;
  assign new_n13907_ = ~new_n9575_ | ~pi0652;
  assign new_n13908_ = ~new_n9574_ | ~pi0644;
  assign new_n13909_ = ~new_n9572_ | ~pi0636;
  assign new_n13910_ = ~new_n9571_ | ~pi0628;
  assign new_n13911_ = ~new_n9569_ | ~pi0692;
  assign new_n13912_ = ~new_n9568_ | ~pi0700;
  assign new_n13913_ = ~new_n9567_ | ~pi0708;
  assign new_n13914_ = ~new_n9565_ | ~pi0716;
  assign new_n13915_ = ~new_n9563_ | ~pi0724;
  assign new_n13916_ = ~new_n9562_ | ~pi0732;
  assign new_n13917_ = ~new_n9560_ | ~pi0740;
  assign new_n13918_ = ~new_n9558_ | ~pi0748;
  assign new_n13919_ = ~new_n9603_ | ~pi0628;
  assign new_n13920_ = ~new_n9602_ | ~pi0636;
  assign new_n13921_ = ~new_n9601_ | ~pi0644;
  assign new_n13922_ = ~new_n9600_ | ~pi0652;
  assign new_n13923_ = ~new_n9599_ | ~pi0660;
  assign new_n13924_ = ~new_n9598_ | ~pi0668;
  assign new_n13925_ = ~new_n9596_ | ~pi0676;
  assign new_n13926_ = ~new_n9595_ | ~pi0684;
  assign new_n13927_ = ~new_n9593_ | ~pi0692;
  assign new_n13928_ = ~new_n9592_ | ~pi0700;
  assign new_n13929_ = ~new_n9591_ | ~pi0708;
  assign new_n13930_ = ~new_n9589_ | ~pi0716;
  assign new_n13931_ = ~new_n9587_ | ~pi0724;
  assign new_n13932_ = ~new_n9586_ | ~pi0732;
  assign new_n13933_ = ~new_n9584_ | ~pi0740;
  assign new_n13934_ = ~new_n9582_ | ~pi0748;
  assign new_n13935_ = ~new_n9603_ | ~pi0629;
  assign new_n13936_ = ~new_n9602_ | ~pi0637;
  assign new_n13937_ = ~new_n9601_ | ~pi0645;
  assign new_n13938_ = ~new_n9600_ | ~pi0653;
  assign new_n13939_ = ~new_n9599_ | ~pi0661;
  assign new_n13940_ = ~new_n9598_ | ~pi0669;
  assign new_n13941_ = ~new_n9596_ | ~pi0677;
  assign new_n13942_ = ~new_n9595_ | ~pi0685;
  assign new_n13943_ = ~new_n9593_ | ~pi0693;
  assign new_n13944_ = ~new_n9592_ | ~pi0701;
  assign new_n13945_ = ~new_n9591_ | ~pi0709;
  assign new_n13946_ = ~new_n9589_ | ~pi0717;
  assign new_n13947_ = ~new_n9587_ | ~pi0725;
  assign new_n13948_ = ~new_n9586_ | ~pi0733;
  assign new_n13949_ = ~new_n9584_ | ~pi0741;
  assign new_n13950_ = ~new_n9582_ | ~pi0749;
  assign new_n13951_ = ~new_n9603_ | ~pi0630;
  assign new_n13952_ = ~new_n9602_ | ~pi0638;
  assign new_n13953_ = ~new_n9601_ | ~pi0646;
  assign new_n13954_ = ~new_n9600_ | ~pi0654;
  assign new_n13955_ = ~new_n9599_ | ~pi0662;
  assign new_n13956_ = ~new_n9598_ | ~pi0670;
  assign new_n13957_ = ~new_n9596_ | ~pi0678;
  assign new_n13958_ = ~new_n9595_ | ~pi0686;
  assign new_n13959_ = ~new_n9593_ | ~pi0694;
  assign new_n13960_ = ~new_n9592_ | ~pi0702;
  assign new_n13961_ = ~new_n9591_ | ~pi0710;
  assign new_n13962_ = ~new_n9589_ | ~pi0718;
  assign new_n13963_ = ~new_n9587_ | ~pi0726;
  assign new_n13964_ = ~new_n9586_ | ~pi0734;
  assign new_n13965_ = ~new_n9584_ | ~pi0742;
  assign new_n13966_ = ~new_n9582_ | ~pi0750;
  assign new_n13967_ = ~new_n9603_ | ~pi0631;
  assign new_n13968_ = ~new_n9602_ | ~pi0639;
  assign new_n13969_ = ~new_n9601_ | ~pi0647;
  assign new_n13970_ = ~new_n9600_ | ~pi0655;
  assign new_n13971_ = ~new_n9599_ | ~pi0663;
  assign new_n13972_ = ~new_n9598_ | ~pi0671;
  assign new_n13973_ = ~new_n9596_ | ~pi0679;
  assign new_n13974_ = ~new_n9595_ | ~pi0687;
  assign new_n13975_ = ~new_n9593_ | ~pi0695;
  assign new_n13976_ = ~new_n9592_ | ~pi0703;
  assign new_n13977_ = ~new_n9591_ | ~pi0711;
  assign new_n13978_ = ~new_n9589_ | ~pi0719;
  assign new_n13979_ = ~new_n9587_ | ~pi0727;
  assign new_n13980_ = ~new_n9586_ | ~pi0735;
  assign new_n13981_ = ~new_n9584_ | ~pi0743;
  assign new_n13982_ = ~new_n9582_ | ~pi0751;
  assign new_n13983_ = ~new_n9603_ | ~pi0632;
  assign new_n13984_ = ~new_n9602_ | ~pi0640;
  assign new_n13985_ = ~new_n9601_ | ~pi0648;
  assign new_n13986_ = ~new_n9600_ | ~pi0656;
  assign new_n13987_ = ~new_n9599_ | ~pi0664;
  assign new_n13988_ = ~new_n9598_ | ~pi0672;
  assign new_n13989_ = ~new_n9596_ | ~pi0680;
  assign new_n13990_ = ~new_n9595_ | ~pi0688;
  assign new_n13991_ = ~new_n9593_ | ~pi0696;
  assign new_n13992_ = ~new_n9592_ | ~pi0704;
  assign new_n13993_ = ~new_n9591_ | ~pi0712;
  assign new_n13994_ = ~new_n9589_ | ~pi0720;
  assign new_n13995_ = ~new_n9587_ | ~pi0728;
  assign new_n13996_ = ~new_n9586_ | ~pi0736;
  assign new_n13997_ = ~new_n9584_ | ~pi0744;
  assign new_n13998_ = ~new_n9582_ | ~pi0752;
  assign new_n13999_ = ~new_n9603_ | ~pi0633;
  assign new_n14000_ = ~new_n9602_ | ~pi0641;
  assign new_n14001_ = ~new_n9601_ | ~pi0649;
  assign new_n14002_ = ~new_n9600_ | ~pi0657;
  assign new_n14003_ = ~new_n9599_ | ~pi0665;
  assign new_n14004_ = ~new_n9598_ | ~pi0673;
  assign new_n14005_ = ~new_n9596_ | ~pi0681;
  assign new_n14006_ = ~new_n9595_ | ~pi0689;
  assign new_n14007_ = ~new_n9593_ | ~pi0697;
  assign new_n14008_ = ~new_n9592_ | ~pi0705;
  assign new_n14009_ = ~new_n9591_ | ~pi0713;
  assign new_n14010_ = ~new_n9589_ | ~pi0721;
  assign new_n14011_ = ~new_n9587_ | ~pi0729;
  assign new_n14012_ = ~new_n9586_ | ~pi0737;
  assign new_n14013_ = ~new_n9584_ | ~pi0745;
  assign new_n14014_ = ~new_n9582_ | ~pi0753;
  assign new_n14015_ = ~new_n9603_ | ~pi0634;
  assign new_n14016_ = ~new_n9602_ | ~pi0642;
  assign new_n14017_ = ~new_n9601_ | ~pi0650;
  assign new_n14018_ = ~new_n9600_ | ~pi0658;
  assign new_n14019_ = ~new_n9599_ | ~pi0666;
  assign new_n14020_ = ~new_n9598_ | ~pi0674;
  assign new_n14021_ = ~new_n9596_ | ~pi0682;
  assign new_n14022_ = ~new_n9595_ | ~pi0690;
  assign new_n14023_ = ~new_n9593_ | ~pi0698;
  assign new_n14024_ = ~new_n9592_ | ~pi0706;
  assign new_n14025_ = ~new_n9591_ | ~pi0714;
  assign new_n14026_ = ~new_n9589_ | ~pi0722;
  assign new_n14027_ = ~new_n9587_ | ~pi0730;
  assign new_n14028_ = ~new_n9586_ | ~pi0738;
  assign new_n14029_ = ~new_n9584_ | ~pi0746;
  assign new_n14030_ = ~new_n9582_ | ~pi0754;
  assign new_n14031_ = ~new_n9603_ | ~pi0635;
  assign new_n14032_ = ~new_n9602_ | ~pi0643;
  assign new_n14033_ = ~new_n9601_ | ~pi0651;
  assign new_n14034_ = ~new_n9600_ | ~pi0659;
  assign new_n14035_ = ~new_n9599_ | ~pi0667;
  assign new_n14036_ = ~new_n9598_ | ~pi0675;
  assign new_n14037_ = ~new_n9596_ | ~pi0683;
  assign new_n14038_ = ~new_n9595_ | ~pi0691;
  assign new_n14039_ = ~new_n9593_ | ~pi0699;
  assign new_n14040_ = ~new_n9592_ | ~pi0707;
  assign new_n14041_ = ~new_n9591_ | ~pi0715;
  assign new_n14042_ = ~new_n9589_ | ~pi0723;
  assign new_n14043_ = ~new_n9587_ | ~pi0731;
  assign new_n14044_ = ~new_n9586_ | ~pi0739;
  assign new_n14045_ = ~new_n9584_ | ~pi0747;
  assign new_n14046_ = ~new_n9582_ | ~pi0755;
  assign new_n14047_ = pi0760 | pi0759;
  assign new_n14048_ = ~new_n11446_;
  assign new_n14049_ = ~new_n9627_ | ~pi0748;
  assign new_n14050_ = ~new_n9626_ | ~pi0740;
  assign new_n14051_ = ~new_n9625_ | ~pi0732;
  assign new_n14052_ = ~new_n9624_ | ~pi0724;
  assign new_n14053_ = ~new_n9622_ | ~pi0716;
  assign new_n14054_ = ~new_n9621_ | ~pi0708;
  assign new_n14055_ = ~new_n9620_ | ~pi0700;
  assign new_n14056_ = ~new_n9619_ | ~pi0692;
  assign new_n14057_ = ~new_n9617_ | ~pi0684;
  assign new_n14058_ = ~new_n9616_ | ~pi0676;
  assign new_n14059_ = ~new_n9615_ | ~pi0668;
  assign new_n14060_ = ~new_n9614_ | ~pi0660;
  assign new_n14061_ = ~new_n9612_ | ~pi0652;
  assign new_n14062_ = ~new_n9610_ | ~pi0644;
  assign new_n14063_ = ~new_n9608_ | ~pi0636;
  assign new_n14064_ = ~new_n9606_ | ~pi0628;
  assign new_n14065_ = ~new_n9627_ | ~pi0749;
  assign new_n14066_ = ~new_n9626_ | ~pi0741;
  assign new_n14067_ = ~new_n9625_ | ~pi0733;
  assign new_n14068_ = ~new_n9624_ | ~pi0725;
  assign new_n14069_ = ~new_n9622_ | ~pi0717;
  assign new_n14070_ = ~new_n9621_ | ~pi0709;
  assign new_n14071_ = ~new_n9620_ | ~pi0701;
  assign new_n14072_ = ~new_n9619_ | ~pi0693;
  assign new_n14073_ = ~new_n9617_ | ~pi0685;
  assign new_n14074_ = ~new_n9616_ | ~pi0677;
  assign new_n14075_ = ~new_n9615_ | ~pi0669;
  assign new_n14076_ = ~new_n9614_ | ~pi0661;
  assign new_n14077_ = ~new_n9612_ | ~pi0653;
  assign new_n14078_ = ~new_n9610_ | ~pi0645;
  assign new_n14079_ = ~new_n9608_ | ~pi0637;
  assign new_n14080_ = ~new_n9606_ | ~pi0629;
  assign new_n14081_ = ~new_n9627_ | ~pi0750;
  assign new_n14082_ = ~new_n9626_ | ~pi0742;
  assign new_n14083_ = ~new_n9625_ | ~pi0734;
  assign new_n14084_ = ~new_n9624_ | ~pi0726;
  assign new_n14085_ = ~new_n9622_ | ~pi0718;
  assign new_n14086_ = ~new_n9621_ | ~pi0710;
  assign new_n14087_ = ~new_n9620_ | ~pi0702;
  assign new_n14088_ = ~new_n9619_ | ~pi0694;
  assign new_n14089_ = ~new_n9617_ | ~pi0686;
  assign new_n14090_ = ~new_n9616_ | ~pi0678;
  assign new_n14091_ = ~new_n9615_ | ~pi0670;
  assign new_n14092_ = ~new_n9614_ | ~pi0662;
  assign new_n14093_ = ~new_n9612_ | ~pi0654;
  assign new_n14094_ = ~new_n9610_ | ~pi0646;
  assign new_n14095_ = ~new_n9608_ | ~pi0638;
  assign new_n14096_ = ~new_n9606_ | ~pi0630;
  assign new_n14097_ = ~new_n9627_ | ~pi0751;
  assign new_n14098_ = ~new_n9626_ | ~pi0743;
  assign new_n14099_ = ~new_n9625_ | ~pi0735;
  assign new_n14100_ = ~new_n9624_ | ~pi0727;
  assign new_n14101_ = ~new_n9622_ | ~pi0719;
  assign new_n14102_ = ~new_n9621_ | ~pi0711;
  assign new_n14103_ = ~new_n9620_ | ~pi0703;
  assign new_n14104_ = ~new_n9619_ | ~pi0695;
  assign new_n14105_ = ~new_n9617_ | ~pi0687;
  assign new_n14106_ = ~new_n9616_ | ~pi0679;
  assign new_n14107_ = ~new_n9615_ | ~pi0671;
  assign new_n14108_ = ~new_n9614_ | ~pi0663;
  assign new_n14109_ = ~new_n9612_ | ~pi0655;
  assign new_n14110_ = ~new_n9610_ | ~pi0647;
  assign new_n14111_ = ~new_n9608_ | ~pi0639;
  assign new_n14112_ = ~new_n9606_ | ~pi0631;
  assign new_n14113_ = ~new_n9627_ | ~pi0752;
  assign new_n14114_ = ~new_n9626_ | ~pi0744;
  assign new_n14115_ = ~new_n9625_ | ~pi0736;
  assign new_n14116_ = ~new_n9624_ | ~pi0728;
  assign new_n14117_ = ~new_n9622_ | ~pi0720;
  assign new_n14118_ = ~new_n9621_ | ~pi0712;
  assign new_n14119_ = ~new_n9620_ | ~pi0704;
  assign new_n14120_ = ~new_n9619_ | ~pi0696;
  assign new_n14121_ = ~new_n9617_ | ~pi0688;
  assign new_n14122_ = ~new_n9616_ | ~pi0680;
  assign new_n14123_ = ~new_n9615_ | ~pi0672;
  assign new_n14124_ = ~new_n9614_ | ~pi0664;
  assign new_n14125_ = ~new_n9612_ | ~pi0656;
  assign new_n14126_ = ~new_n9610_ | ~pi0648;
  assign new_n14127_ = ~new_n9608_ | ~pi0640;
  assign new_n14128_ = ~new_n9606_ | ~pi0632;
  assign new_n14129_ = ~new_n9627_ | ~pi0753;
  assign new_n14130_ = ~new_n9626_ | ~pi0745;
  assign new_n14131_ = ~new_n9625_ | ~pi0737;
  assign new_n14132_ = ~new_n9624_ | ~pi0729;
  assign new_n14133_ = ~new_n9622_ | ~pi0721;
  assign new_n14134_ = ~new_n9621_ | ~pi0713;
  assign new_n14135_ = ~new_n9620_ | ~pi0705;
  assign new_n14136_ = ~new_n9619_ | ~pi0697;
  assign new_n14137_ = ~new_n9617_ | ~pi0689;
  assign new_n14138_ = ~new_n9616_ | ~pi0681;
  assign new_n14139_ = ~new_n9615_ | ~pi0673;
  assign new_n14140_ = ~new_n9614_ | ~pi0665;
  assign new_n14141_ = ~new_n9612_ | ~pi0657;
  assign new_n14142_ = ~new_n9610_ | ~pi0649;
  assign new_n14143_ = ~new_n9608_ | ~pi0641;
  assign new_n14144_ = ~new_n9606_ | ~pi0633;
  assign new_n14145_ = ~new_n9627_ | ~pi0754;
  assign new_n14146_ = ~new_n9626_ | ~pi0746;
  assign new_n14147_ = ~new_n9625_ | ~pi0738;
  assign new_n14148_ = ~new_n9624_ | ~pi0730;
  assign new_n14149_ = ~new_n9622_ | ~pi0722;
  assign new_n14150_ = ~new_n9621_ | ~pi0714;
  assign new_n14151_ = ~new_n9620_ | ~pi0706;
  assign new_n14152_ = ~new_n9619_ | ~pi0698;
  assign new_n14153_ = ~new_n9617_ | ~pi0690;
  assign new_n14154_ = ~new_n9616_ | ~pi0682;
  assign new_n14155_ = ~new_n9615_ | ~pi0674;
  assign new_n14156_ = ~new_n9614_ | ~pi0666;
  assign new_n14157_ = ~new_n9612_ | ~pi0658;
  assign new_n14158_ = ~new_n9610_ | ~pi0650;
  assign new_n14159_ = ~new_n9608_ | ~pi0642;
  assign new_n14160_ = ~new_n9606_ | ~pi0634;
  assign new_n14161_ = ~new_n9627_ | ~pi0755;
  assign new_n14162_ = ~new_n9626_ | ~pi0747;
  assign new_n14163_ = ~new_n9625_ | ~pi0739;
  assign new_n14164_ = ~new_n9624_ | ~pi0731;
  assign new_n14165_ = ~new_n9622_ | ~pi0723;
  assign new_n14166_ = ~new_n9621_ | ~pi0715;
  assign new_n14167_ = ~new_n9620_ | ~pi0707;
  assign new_n14168_ = ~new_n9619_ | ~pi0699;
  assign new_n14169_ = ~new_n9617_ | ~pi0691;
  assign new_n14170_ = ~new_n9616_ | ~pi0683;
  assign new_n14171_ = ~new_n9615_ | ~pi0675;
  assign new_n14172_ = ~new_n9614_ | ~pi0667;
  assign new_n14173_ = ~new_n9612_ | ~pi0659;
  assign new_n14174_ = ~new_n9610_ | ~pi0651;
  assign new_n14175_ = ~new_n9608_ | ~pi0643;
  assign new_n14176_ = ~new_n9606_ | ~pi0635;
  assign new_n14177_ = ~new_n10595_;
  assign new_n14178_ = ~new_n14177_ | ~new_n10341_;
  assign new_n14179_ = ~new_n11508_ | ~new_n27643_;
  assign new_n14180_ = ~pi0757 | ~new_n14178_;
  assign new_n14181_ = ~new_n11471_ | ~new_n10469_;
  assign new_n14182_ = ~new_n28267_ | ~new_n9396_;
  assign new_n14183_ = ~new_n9395_ | ~new_n9647_;
  assign new_n14184_ = ~new_n9646_ | ~new_n9396_;
  assign new_n14185_ = ~new_n9395_ | ~new_n9646_;
  assign new_n14186_ = ~new_n9645_ | ~new_n9396_;
  assign new_n14187_ = ~new_n9395_ | ~new_n9645_;
  assign new_n14188_ = ~new_n9644_ | ~new_n9396_;
  assign new_n14189_ = ~new_n9395_ | ~new_n9644_;
  assign new_n14190_ = ~new_n11508_ | ~new_n27644_;
  assign new_n14191_ = ~pi0758 | ~new_n14178_;
  assign new_n14192_ = ~new_n11471_ | ~new_n10621_;
  assign new_n14193_ = ~new_n9643_ | ~new_n9396_;
  assign new_n14194_ = ~new_n9395_ | ~new_n9643_;
  assign new_n14195_ = ~new_n9642_ | ~new_n9396_;
  assign new_n14196_ = ~new_n9395_ | ~new_n9642_;
  assign new_n14197_ = ~new_n9641_ | ~new_n9396_;
  assign new_n14198_ = ~new_n9395_ | ~new_n9641_;
  assign new_n14199_ = ~new_n9640_ | ~new_n9396_;
  assign new_n14200_ = ~new_n9395_ | ~new_n9640_;
  assign new_n14201_ = ~new_n11508_ | ~new_n27553_;
  assign new_n14202_ = ~pi0759 | ~new_n14178_;
  assign new_n14203_ = ~new_n11471_ | ~new_n10284_;
  assign new_n14204_ = ~new_n11508_ | ~new_n27642_;
  assign new_n14205_ = ~pi0760 | ~new_n14178_;
  assign new_n14206_ = ~new_n11471_ | ~new_n10348_;
  assign new_n14207_ = ~pi0755 | ~new_n9396_;
  assign new_n14208_ = ~new_n12558_ | ~pi0748;
  assign new_n14209_ = ~new_n12501_ | ~pi0740;
  assign new_n14210_ = ~new_n12443_ | ~pi0732;
  assign new_n14211_ = ~new_n12386_ | ~pi0724;
  assign new_n14212_ = ~new_n12328_ | ~pi0716;
  assign new_n14213_ = ~new_n12271_ | ~pi0708;
  assign new_n14214_ = ~new_n12213_ | ~pi0700;
  assign new_n14215_ = ~new_n12157_ | ~pi0692;
  assign new_n14216_ = ~new_n12100_ | ~pi0684;
  assign new_n14217_ = ~new_n12043_ | ~pi0676;
  assign new_n14218_ = ~new_n11985_ | ~pi0668;
  assign new_n14219_ = ~new_n11928_ | ~pi0660;
  assign new_n14220_ = ~new_n11870_ | ~pi0652;
  assign new_n14221_ = ~new_n11813_ | ~pi0644;
  assign new_n14222_ = ~new_n11754_ | ~pi0636;
  assign new_n14223_ = ~new_n11694_ | ~pi0628;
  assign new_n14224_ = ~new_n11320_ | ~new_n11318_ | ~new_n11319_ | ~new_n11321_;
  assign new_n14225_ = ~new_n12558_ | ~pi0749;
  assign new_n14226_ = ~new_n12501_ | ~pi0741;
  assign new_n14227_ = ~new_n12443_ | ~pi0733;
  assign new_n14228_ = ~new_n12386_ | ~pi0725;
  assign new_n14229_ = ~new_n12328_ | ~pi0717;
  assign new_n14230_ = ~new_n12271_ | ~pi0709;
  assign new_n14231_ = ~new_n12213_ | ~pi0701;
  assign new_n14232_ = ~new_n12157_ | ~pi0693;
  assign new_n14233_ = ~new_n12100_ | ~pi0685;
  assign new_n14234_ = ~new_n12043_ | ~pi0677;
  assign new_n14235_ = ~new_n11985_ | ~pi0669;
  assign new_n14236_ = ~new_n11928_ | ~pi0661;
  assign new_n14237_ = ~new_n11870_ | ~pi0653;
  assign new_n14238_ = ~new_n11813_ | ~pi0645;
  assign new_n14239_ = ~new_n11754_ | ~pi0637;
  assign new_n14240_ = ~new_n11694_ | ~pi0629;
  assign new_n14241_ = ~new_n11324_ | ~new_n11322_ | ~new_n11323_ | ~new_n11325_;
  assign new_n14242_ = ~new_n9579_ | ~pi0685;
  assign new_n14243_ = ~new_n9578_ | ~pi0677;
  assign new_n14244_ = ~new_n9577_ | ~pi0669;
  assign new_n14245_ = ~new_n9576_ | ~pi0661;
  assign new_n14246_ = ~new_n9575_ | ~pi0653;
  assign new_n14247_ = ~new_n9574_ | ~pi0645;
  assign new_n14248_ = ~new_n9572_ | ~pi0637;
  assign new_n14249_ = ~new_n9571_ | ~pi0629;
  assign new_n14250_ = ~new_n9569_ | ~pi0693;
  assign new_n14251_ = ~new_n9568_ | ~pi0701;
  assign new_n14252_ = ~new_n9567_ | ~pi0709;
  assign new_n14253_ = ~new_n9565_ | ~pi0717;
  assign new_n14254_ = ~new_n9563_ | ~pi0725;
  assign new_n14255_ = ~new_n9562_ | ~pi0733;
  assign new_n14256_ = ~new_n9560_ | ~pi0741;
  assign new_n14257_ = ~new_n9558_ | ~pi0749;
  assign new_n14258_ = ~new_n11328_ | ~new_n11326_ | ~new_n11327_ | ~new_n11329_;
  assign new_n14259_ = ~new_n12558_ | ~pi0750;
  assign new_n14260_ = ~new_n12501_ | ~pi0742;
  assign new_n14261_ = ~new_n12443_ | ~pi0734;
  assign new_n14262_ = ~new_n12386_ | ~pi0726;
  assign new_n14263_ = ~new_n12328_ | ~pi0718;
  assign new_n14264_ = ~new_n12271_ | ~pi0710;
  assign new_n14265_ = ~new_n12213_ | ~pi0702;
  assign new_n14266_ = ~new_n12157_ | ~pi0694;
  assign new_n14267_ = ~new_n12100_ | ~pi0686;
  assign new_n14268_ = ~new_n12043_ | ~pi0678;
  assign new_n14269_ = ~new_n11985_ | ~pi0670;
  assign new_n14270_ = ~new_n11928_ | ~pi0662;
  assign new_n14271_ = ~new_n11870_ | ~pi0654;
  assign new_n14272_ = ~new_n11813_ | ~pi0646;
  assign new_n14273_ = ~new_n11754_ | ~pi0638;
  assign new_n14274_ = ~new_n11694_ | ~pi0630;
  assign new_n14275_ = ~new_n11332_ | ~new_n11330_ | ~new_n11331_ | ~new_n11333_;
  assign new_n14276_ = ~new_n9579_ | ~pi0686;
  assign new_n14277_ = ~new_n9578_ | ~pi0678;
  assign new_n14278_ = ~new_n9577_ | ~pi0670;
  assign new_n14279_ = ~new_n9576_ | ~pi0662;
  assign new_n14280_ = ~new_n9575_ | ~pi0654;
  assign new_n14281_ = ~new_n9574_ | ~pi0646;
  assign new_n14282_ = ~new_n9572_ | ~pi0638;
  assign new_n14283_ = ~new_n9571_ | ~pi0630;
  assign new_n14284_ = ~new_n9569_ | ~pi0694;
  assign new_n14285_ = ~new_n9568_ | ~pi0702;
  assign new_n14286_ = ~new_n9567_ | ~pi0710;
  assign new_n14287_ = ~new_n9565_ | ~pi0718;
  assign new_n14288_ = ~new_n9563_ | ~pi0726;
  assign new_n14289_ = ~new_n9562_ | ~pi0734;
  assign new_n14290_ = ~new_n9560_ | ~pi0742;
  assign new_n14291_ = ~new_n9558_ | ~pi0750;
  assign new_n14292_ = ~new_n11336_ | ~new_n11334_ | ~new_n11335_ | ~new_n11337_;
  assign new_n14293_ = ~new_n12558_ | ~pi0751;
  assign new_n14294_ = ~new_n12501_ | ~pi0743;
  assign new_n14295_ = ~new_n12443_ | ~pi0735;
  assign new_n14296_ = ~new_n12386_ | ~pi0727;
  assign new_n14297_ = ~new_n12328_ | ~pi0719;
  assign new_n14298_ = ~new_n12271_ | ~pi0711;
  assign new_n14299_ = ~new_n12213_ | ~pi0703;
  assign new_n14300_ = ~new_n12157_ | ~pi0695;
  assign new_n14301_ = ~new_n12100_ | ~pi0687;
  assign new_n14302_ = ~new_n12043_ | ~pi0679;
  assign new_n14303_ = ~new_n11985_ | ~pi0671;
  assign new_n14304_ = ~new_n11928_ | ~pi0663;
  assign new_n14305_ = ~new_n11870_ | ~pi0655;
  assign new_n14306_ = ~new_n11813_ | ~pi0647;
  assign new_n14307_ = ~new_n11754_ | ~pi0639;
  assign new_n14308_ = ~new_n11694_ | ~pi0631;
  assign new_n14309_ = ~new_n11340_ | ~new_n11338_ | ~new_n11339_ | ~new_n11341_;
  assign new_n14310_ = ~new_n9579_ | ~pi0687;
  assign new_n14311_ = ~new_n9578_ | ~pi0679;
  assign new_n14312_ = ~new_n9577_ | ~pi0671;
  assign new_n14313_ = ~new_n9576_ | ~pi0663;
  assign new_n14314_ = ~new_n9575_ | ~pi0655;
  assign new_n14315_ = ~new_n9574_ | ~pi0647;
  assign new_n14316_ = ~new_n9572_ | ~pi0639;
  assign new_n14317_ = ~new_n9571_ | ~pi0631;
  assign new_n14318_ = ~new_n9569_ | ~pi0695;
  assign new_n14319_ = ~new_n9568_ | ~pi0703;
  assign new_n14320_ = ~new_n9567_ | ~pi0711;
  assign new_n14321_ = ~new_n9565_ | ~pi0719;
  assign new_n14322_ = ~new_n9563_ | ~pi0727;
  assign new_n14323_ = ~new_n9562_ | ~pi0735;
  assign new_n14324_ = ~new_n9560_ | ~pi0743;
  assign new_n14325_ = ~new_n9558_ | ~pi0751;
  assign new_n14326_ = ~new_n11344_ | ~new_n11342_ | ~new_n11343_ | ~new_n11345_;
  assign new_n14327_ = ~new_n12558_ | ~pi0752;
  assign new_n14328_ = ~new_n12501_ | ~pi0744;
  assign new_n14329_ = ~new_n12443_ | ~pi0736;
  assign new_n14330_ = ~new_n12386_ | ~pi0728;
  assign new_n14331_ = ~new_n12328_ | ~pi0720;
  assign new_n14332_ = ~new_n12271_ | ~pi0712;
  assign new_n14333_ = ~new_n12213_ | ~pi0704;
  assign new_n14334_ = ~new_n12157_ | ~pi0696;
  assign new_n14335_ = ~new_n12100_ | ~pi0688;
  assign new_n14336_ = ~new_n12043_ | ~pi0680;
  assign new_n14337_ = ~new_n11985_ | ~pi0672;
  assign new_n14338_ = ~new_n11928_ | ~pi0664;
  assign new_n14339_ = ~new_n11870_ | ~pi0656;
  assign new_n14340_ = ~new_n11813_ | ~pi0648;
  assign new_n14341_ = ~new_n11754_ | ~pi0640;
  assign new_n14342_ = ~new_n11694_ | ~pi0632;
  assign new_n14343_ = ~new_n11348_ | ~new_n11346_ | ~new_n11347_ | ~new_n11349_;
  assign new_n14344_ = ~new_n9579_ | ~pi0688;
  assign new_n14345_ = ~new_n9578_ | ~pi0680;
  assign new_n14346_ = ~new_n9577_ | ~pi0672;
  assign new_n14347_ = ~new_n9576_ | ~pi0664;
  assign new_n14348_ = ~new_n9575_ | ~pi0656;
  assign new_n14349_ = ~new_n9574_ | ~pi0648;
  assign new_n14350_ = ~new_n9572_ | ~pi0640;
  assign new_n14351_ = ~new_n9571_ | ~pi0632;
  assign new_n14352_ = ~new_n9569_ | ~pi0696;
  assign new_n14353_ = ~new_n9568_ | ~pi0704;
  assign new_n14354_ = ~new_n9567_ | ~pi0712;
  assign new_n14355_ = ~new_n9565_ | ~pi0720;
  assign new_n14356_ = ~new_n9563_ | ~pi0728;
  assign new_n14357_ = ~new_n9562_ | ~pi0736;
  assign new_n14358_ = ~new_n9560_ | ~pi0744;
  assign new_n14359_ = ~new_n9558_ | ~pi0752;
  assign new_n14360_ = ~new_n11352_ | ~new_n11350_ | ~new_n11351_ | ~new_n11353_;
  assign new_n14361_ = ~new_n12558_ | ~pi0753;
  assign new_n14362_ = ~new_n12501_ | ~pi0745;
  assign new_n14363_ = ~new_n12443_ | ~pi0737;
  assign new_n14364_ = ~new_n12386_ | ~pi0729;
  assign new_n14365_ = ~new_n12328_ | ~pi0721;
  assign new_n14366_ = ~new_n12271_ | ~pi0713;
  assign new_n14367_ = ~new_n12213_ | ~pi0705;
  assign new_n14368_ = ~new_n12157_ | ~pi0697;
  assign new_n14369_ = ~new_n12100_ | ~pi0689;
  assign new_n14370_ = ~new_n12043_ | ~pi0681;
  assign new_n14371_ = ~new_n11985_ | ~pi0673;
  assign new_n14372_ = ~new_n11928_ | ~pi0665;
  assign new_n14373_ = ~new_n11870_ | ~pi0657;
  assign new_n14374_ = ~new_n11813_ | ~pi0649;
  assign new_n14375_ = ~new_n11754_ | ~pi0641;
  assign new_n14376_ = ~new_n11694_ | ~pi0633;
  assign new_n14377_ = ~new_n11356_ | ~new_n11354_ | ~new_n11355_ | ~new_n11357_;
  assign new_n14378_ = ~new_n9579_ | ~pi0689;
  assign new_n14379_ = ~new_n9578_ | ~pi0681;
  assign new_n14380_ = ~new_n9577_ | ~pi0673;
  assign new_n14381_ = ~new_n9576_ | ~pi0665;
  assign new_n14382_ = ~new_n9575_ | ~pi0657;
  assign new_n14383_ = ~new_n9574_ | ~pi0649;
  assign new_n14384_ = ~new_n9572_ | ~pi0641;
  assign new_n14385_ = ~new_n9571_ | ~pi0633;
  assign new_n14386_ = ~new_n9569_ | ~pi0697;
  assign new_n14387_ = ~new_n9568_ | ~pi0705;
  assign new_n14388_ = ~new_n9567_ | ~pi0713;
  assign new_n14389_ = ~new_n9565_ | ~pi0721;
  assign new_n14390_ = ~new_n9563_ | ~pi0729;
  assign new_n14391_ = ~new_n9562_ | ~pi0737;
  assign new_n14392_ = ~new_n9560_ | ~pi0745;
  assign new_n14393_ = ~new_n9558_ | ~pi0753;
  assign new_n14394_ = ~new_n11360_ | ~new_n11358_ | ~new_n11359_ | ~new_n11361_;
  assign new_n14395_ = ~new_n12558_ | ~pi0754;
  assign new_n14396_ = ~new_n12501_ | ~pi0746;
  assign new_n14397_ = ~new_n12443_ | ~pi0738;
  assign new_n14398_ = ~new_n12386_ | ~pi0730;
  assign new_n14399_ = ~new_n12328_ | ~pi0722;
  assign new_n14400_ = ~new_n12271_ | ~pi0714;
  assign new_n14401_ = ~new_n12213_ | ~pi0706;
  assign new_n14402_ = ~new_n12157_ | ~pi0698;
  assign new_n14403_ = ~new_n12100_ | ~pi0690;
  assign new_n14404_ = ~new_n12043_ | ~pi0682;
  assign new_n14405_ = ~new_n11985_ | ~pi0674;
  assign new_n14406_ = ~new_n11928_ | ~pi0666;
  assign new_n14407_ = ~new_n11870_ | ~pi0658;
  assign new_n14408_ = ~new_n11813_ | ~pi0650;
  assign new_n14409_ = ~new_n11754_ | ~pi0642;
  assign new_n14410_ = ~new_n11694_ | ~pi0634;
  assign new_n14411_ = ~new_n11364_ | ~new_n11362_ | ~new_n11363_ | ~new_n11365_;
  assign new_n14412_ = ~new_n9579_ | ~pi0690;
  assign new_n14413_ = ~new_n9578_ | ~pi0682;
  assign new_n14414_ = ~new_n9577_ | ~pi0674;
  assign new_n14415_ = ~new_n9576_ | ~pi0666;
  assign new_n14416_ = ~new_n9575_ | ~pi0658;
  assign new_n14417_ = ~new_n9574_ | ~pi0650;
  assign new_n14418_ = ~new_n9572_ | ~pi0642;
  assign new_n14419_ = ~new_n9571_ | ~pi0634;
  assign new_n14420_ = ~new_n9569_ | ~pi0698;
  assign new_n14421_ = ~new_n9568_ | ~pi0706;
  assign new_n14422_ = ~new_n9567_ | ~pi0714;
  assign new_n14423_ = ~new_n9565_ | ~pi0722;
  assign new_n14424_ = ~new_n9563_ | ~pi0730;
  assign new_n14425_ = ~new_n9562_ | ~pi0738;
  assign new_n14426_ = ~new_n9560_ | ~pi0746;
  assign new_n14427_ = ~new_n9558_ | ~pi0754;
  assign new_n14428_ = ~new_n11368_ | ~new_n11366_ | ~new_n11367_ | ~new_n11369_;
  assign new_n14429_ = ~new_n12558_ | ~pi0755;
  assign new_n14430_ = ~new_n12501_ | ~pi0747;
  assign new_n14431_ = ~new_n12443_ | ~pi0739;
  assign new_n14432_ = ~new_n12386_ | ~pi0731;
  assign new_n14433_ = ~new_n12328_ | ~pi0723;
  assign new_n14434_ = ~new_n12271_ | ~pi0715;
  assign new_n14435_ = ~new_n12213_ | ~pi0707;
  assign new_n14436_ = ~new_n12157_ | ~pi0699;
  assign new_n14437_ = ~new_n12100_ | ~pi0691;
  assign new_n14438_ = ~new_n12043_ | ~pi0683;
  assign new_n14439_ = ~new_n11985_ | ~pi0675;
  assign new_n14440_ = ~new_n11928_ | ~pi0667;
  assign new_n14441_ = ~new_n11870_ | ~pi0659;
  assign new_n14442_ = ~new_n11813_ | ~pi0651;
  assign new_n14443_ = ~new_n11754_ | ~pi0643;
  assign new_n14444_ = ~new_n11694_ | ~pi0635;
  assign new_n14445_ = ~new_n11372_ | ~new_n11370_ | ~new_n11371_ | ~new_n11373_;
  assign new_n14446_ = ~new_n9579_ | ~pi0691;
  assign new_n14447_ = ~new_n9578_ | ~pi0683;
  assign new_n14448_ = ~new_n9577_ | ~pi0675;
  assign new_n14449_ = ~new_n9576_ | ~pi0667;
  assign new_n14450_ = ~new_n9575_ | ~pi0659;
  assign new_n14451_ = ~new_n9574_ | ~pi0651;
  assign new_n14452_ = ~new_n9572_ | ~pi0643;
  assign new_n14453_ = ~new_n9571_ | ~pi0635;
  assign new_n14454_ = ~new_n9569_ | ~pi0699;
  assign new_n14455_ = ~new_n9568_ | ~pi0707;
  assign new_n14456_ = ~new_n9567_ | ~pi0715;
  assign new_n14457_ = ~new_n9565_ | ~pi0723;
  assign new_n14458_ = ~new_n9563_ | ~pi0731;
  assign new_n14459_ = ~new_n9562_ | ~pi0739;
  assign new_n14460_ = ~new_n9560_ | ~pi0747;
  assign new_n14461_ = ~new_n9558_ | ~pi0755;
  assign new_n14462_ = ~new_n11376_ | ~new_n11374_ | ~new_n11375_ | ~new_n11377_;
  assign new_n14463_ = ~new_n9393_ | ~new_n14360_;
  assign new_n14464_ = ~pi0762 | ~pi0624;
  assign new_n14465_ = ~new_n9393_ | ~new_n14394_;
  assign new_n14466_ = ~pi0763 | ~pi0624;
  assign new_n14467_ = ~new_n9480_ | ~new_n10336_;
  assign new_n14468_ = ~new_n9393_ | ~new_n14428_;
  assign new_n14469_ = ~pi0764 | ~pi0624;
  assign new_n14470_ = ~new_n9393_ | ~new_n14462_;
  assign new_n14471_ = ~pi0765 | ~pi0624;
  assign new_n14472_ = ~new_n9480_ | ~new_n10320_;
  assign new_n14473_ = ~new_n11454_ | ~new_n11455_ | ~new_n14472_;
  assign new_n14474_ = ~pi0775 | ~new_n14473_;
  assign new_n14475_ = ~new_n9394_ | ~pi0966;
  assign new_n14476_ = ~new_n11453_ | ~pi0902;
  assign new_n14477_ = ~new_n9393_ | ~new_n9649_;
  assign new_n14478_ = ~pi0774 | ~new_n14473_;
  assign new_n14479_ = ~new_n9394_ | ~pi0965;
  assign new_n14480_ = ~new_n11453_ | ~pi0901;
  assign new_n14481_ = ~new_n9393_ | ~new_n9648_;
  assign new_n14482_ = ~pi0773 | ~new_n14473_;
  assign new_n14483_ = ~new_n9394_ | ~pi0964;
  assign new_n14484_ = ~new_n11453_ | ~pi0900;
  assign new_n14485_ = ~pi0772 | ~new_n14473_;
  assign new_n14486_ = ~new_n9394_ | ~pi0963;
  assign new_n14487_ = ~new_n11453_ | ~pi0899;
  assign new_n14488_ = ~pi0771 | ~new_n14473_;
  assign new_n14489_ = ~new_n9394_ | ~pi0962;
  assign new_n14490_ = ~new_n11453_ | ~pi0898;
  assign new_n14491_ = ~pi0770 | ~new_n14473_;
  assign new_n14492_ = ~new_n9394_ | ~pi0961;
  assign new_n14493_ = ~new_n11453_ | ~pi0897;
  assign new_n14494_ = ~pi0797 | ~new_n14473_;
  assign new_n14495_ = ~new_n9394_ | ~pi0988;
  assign new_n14496_ = ~new_n11453_ | ~pi0924;
  assign new_n14497_ = ~pi0796 | ~new_n14473_;
  assign new_n14498_ = ~new_n9394_ | ~pi0987;
  assign new_n14499_ = ~new_n11453_ | ~pi0923;
  assign new_n14500_ = ~pi0769 | ~new_n14473_;
  assign new_n14501_ = ~new_n9394_ | ~pi0960;
  assign new_n14502_ = ~new_n11453_ | ~pi0896;
  assign new_n14503_ = ~pi0795 | ~new_n14473_;
  assign new_n14504_ = ~new_n9394_ | ~pi0986;
  assign new_n14505_ = ~new_n11453_ | ~pi0922;
  assign new_n14506_ = ~pi0794 | ~new_n14473_;
  assign new_n14507_ = ~new_n9394_ | ~pi0985;
  assign new_n14508_ = ~new_n11453_ | ~pi0921;
  assign new_n14509_ = ~pi0793 | ~new_n14473_;
  assign new_n14510_ = ~new_n9394_ | ~pi0984;
  assign new_n14511_ = ~new_n11453_ | ~pi0920;
  assign new_n14512_ = ~pi0792 | ~new_n14473_;
  assign new_n14513_ = ~new_n9394_ | ~pi0983;
  assign new_n14514_ = ~new_n11453_ | ~pi0919;
  assign new_n14515_ = ~pi0791 | ~new_n14473_;
  assign new_n14516_ = ~new_n9394_ | ~pi0982;
  assign new_n14517_ = ~new_n11453_ | ~pi0918;
  assign new_n14518_ = ~pi0790 | ~new_n14473_;
  assign new_n14519_ = ~new_n9394_ | ~pi0981;
  assign new_n14520_ = ~new_n11453_ | ~pi0917;
  assign new_n14521_ = ~pi0789 | ~new_n14473_;
  assign new_n14522_ = ~new_n9394_ | ~pi0980;
  assign new_n14523_ = ~new_n11453_ | ~pi0916;
  assign new_n14524_ = ~pi0788 | ~new_n14473_;
  assign new_n14525_ = ~new_n9394_ | ~pi0979;
  assign new_n14526_ = ~new_n11453_ | ~pi0915;
  assign new_n14527_ = ~pi0787 | ~new_n14473_;
  assign new_n14528_ = ~new_n9394_ | ~pi0978;
  assign new_n14529_ = ~new_n11453_ | ~pi0914;
  assign new_n14530_ = ~pi0786 | ~new_n14473_;
  assign new_n14531_ = ~new_n9394_ | ~pi0977;
  assign new_n14532_ = ~new_n11453_ | ~pi0913;
  assign new_n14533_ = ~pi0768 | ~new_n14473_;
  assign new_n14534_ = ~new_n9394_ | ~pi0959;
  assign new_n14535_ = ~new_n11453_ | ~pi0895;
  assign new_n14536_ = ~pi0785 | ~new_n14473_;
  assign new_n14537_ = ~new_n9394_ | ~pi0976;
  assign new_n14538_ = ~new_n11453_ | ~pi0912;
  assign new_n14539_ = ~pi0784 | ~new_n14473_;
  assign new_n14540_ = ~new_n9394_ | ~pi0975;
  assign new_n14541_ = ~new_n11453_ | ~pi0911;
  assign new_n14542_ = ~pi0783 | ~new_n14473_;
  assign new_n14543_ = ~new_n9394_ | ~pi0974;
  assign new_n14544_ = ~new_n11453_ | ~pi0910;
  assign new_n14545_ = ~pi0782 | ~new_n14473_;
  assign new_n14546_ = ~new_n9394_ | ~pi0973;
  assign new_n14547_ = ~new_n11453_ | ~pi0909;
  assign new_n14548_ = ~pi0781 | ~new_n14473_;
  assign new_n14549_ = ~new_n9394_ | ~pi0972;
  assign new_n14550_ = ~new_n11453_ | ~pi0908;
  assign new_n14551_ = ~new_n9393_ | ~new_n9655_;
  assign new_n14552_ = ~pi0780 | ~new_n14473_;
  assign new_n14553_ = ~new_n9394_ | ~pi0971;
  assign new_n14554_ = ~new_n11453_ | ~pi0907;
  assign new_n14555_ = ~new_n9393_ | ~new_n9654_;
  assign new_n14556_ = ~pi0779 | ~new_n14473_;
  assign new_n14557_ = ~new_n9394_ | ~pi0970;
  assign new_n14558_ = ~new_n11453_ | ~pi0906;
  assign new_n14559_ = ~new_n9393_ | ~new_n9653_;
  assign new_n14560_ = ~pi0778 | ~new_n14473_;
  assign new_n14561_ = ~new_n9394_ | ~pi0969;
  assign new_n14562_ = ~new_n11453_ | ~pi0905;
  assign new_n14563_ = ~new_n9393_ | ~new_n9652_;
  assign new_n14564_ = ~pi0777 | ~new_n14473_;
  assign new_n14565_ = ~new_n9394_ | ~pi0968;
  assign new_n14566_ = ~new_n11453_ | ~pi0904;
  assign new_n14567_ = ~new_n9393_ | ~new_n9651_;
  assign new_n14568_ = ~pi0776 | ~new_n14473_;
  assign new_n14569_ = ~new_n9394_ | ~pi0967;
  assign new_n14570_ = ~new_n11453_ | ~pi0903;
  assign new_n14571_ = ~new_n9393_ | ~new_n9650_;
  assign new_n14572_ = ~pi0767 | ~new_n14473_;
  assign new_n14573_ = ~new_n9394_ | ~pi0958;
  assign new_n14574_ = ~new_n11453_ | ~pi0894;
  assign new_n14575_ = ~pi0766 | ~new_n14473_;
  assign new_n14576_ = ~new_n9394_ | ~pi0957;
  assign new_n14577_ = ~new_n11453_ | ~pi0893;
  assign new_n14578_ = ~pi0934 | ~new_n14910_;
  assign new_n14579_ = ~pi0933 | ~new_n14910_;
  assign new_n14580_ = ~pi0956 | ~new_n14910_;
  assign new_n14581_ = ~pi0955 | ~new_n14910_;
  assign new_n14582_ = ~pi0954 | ~new_n14910_;
  assign new_n14583_ = ~pi0953 | ~new_n14910_;
  assign new_n14584_ = ~pi0952 | ~new_n14910_;
  assign new_n14585_ = ~pi0951 | ~new_n14910_;
  assign new_n14586_ = ~pi0950 | ~new_n14910_;
  assign new_n14587_ = ~pi0949 | ~new_n14910_;
  assign new_n14588_ = ~pi0948 | ~new_n14910_;
  assign new_n14589_ = ~pi0947 | ~new_n14910_;
  assign new_n14590_ = ~pi0946 | ~new_n14910_;
  assign new_n14591_ = ~pi0945 | ~new_n14910_;
  assign new_n14592_ = ~pi0944 | ~new_n14910_;
  assign new_n14593_ = ~pi0943 | ~new_n14910_;
  assign new_n14594_ = ~pi0942 | ~new_n14910_;
  assign new_n14595_ = ~pi0941 | ~new_n14910_;
  assign new_n14596_ = ~pi0940 | ~new_n14910_;
  assign new_n14597_ = ~pi0939 | ~new_n14910_;
  assign new_n14598_ = ~pi0938 | ~new_n14910_;
  assign new_n14599_ = ~pi0937 | ~new_n14910_;
  assign new_n14600_ = ~pi0936 | ~new_n14910_;
  assign new_n14601_ = ~pi0935 | ~new_n14910_;
  assign new_n14602_ = ~new_n11637_ | ~new_n10335_;
  assign new_n14603_ = ~new_n11469_ | ~new_n14326_;
  assign new_n14604_ = ~pi0756 | ~new_n14602_;
  assign new_n14605_ = ~new_n11469_ | ~new_n14360_;
  assign new_n14606_ = ~pi0757 | ~new_n14602_;
  assign new_n14607_ = ~new_n11469_ | ~new_n14394_;
  assign new_n14608_ = ~pi0758 | ~new_n14602_;
  assign new_n14609_ = ~new_n11469_ | ~new_n14428_;
  assign new_n14610_ = ~pi0759 | ~new_n14602_;
  assign new_n14611_ = ~new_n11469_ | ~new_n14462_;
  assign new_n14612_ = ~pi0760 | ~new_n14602_;
  assign new_n14613_ = ~pi0761 | ~new_n14602_;
  assign new_n14614_ = ~pi0762 | ~new_n14602_;
  assign new_n14615_ = ~pi0763 | ~new_n14602_;
  assign new_n14616_ = ~pi0764 | ~new_n14602_;
  assign new_n14617_ = ~pi0765 | ~new_n14602_;
  assign new_n14618_ = ~new_n11418_ | ~new_n12613_;
  assign new_n14619_ = ~pi0627 | ~new_n11473_;
  assign new_n14620_ = ~new_n9658_ | ~new_n9491_;
  assign new_n14621_ = ~new_n11417_ | ~new_n12633_;
  assign new_n14622_ = ~new_n14908_ | ~new_n10566_ | ~new_n13886_;
  assign new_n14623_ = ~new_n11512_ | ~pi0762;
  assign new_n14624_ = ~pi0757 | ~new_n14931_;
  assign new_n14625_ = ~pi0758 | ~new_n14931_;
  assign new_n14626_ = ~pi0763 | ~new_n10325_;
  assign new_n14627_ = ~new_n11422_ | ~new_n11465_;
  assign new_n14628_ = ~new_n11512_ | ~pi0764;
  assign new_n14629_ = ~pi0759 | ~new_n14931_;
  assign new_n14630_ = ~new_n9631_ | ~new_n13886_;
  assign new_n14631_ = ~new_n11512_ | ~pi0765;
  assign new_n14632_ = ~new_n11457_ | ~new_n9417_ | ~new_n14912_;
  assign new_n14633_ = ~new_n10326_ | ~new_n10580_ | ~new_n11463_ | ~new_n14632_;
  assign new_n14634_ = ~pi0775 | ~new_n14633_;
  assign new_n14635_ = ~pi0807 | ~pi0626;
  assign new_n14636_ = ~new_n11464_ | ~pi0966;
  assign new_n14637_ = ~new_n9399_ | ~pi0934;
  assign new_n14638_ = ~pi0774 | ~new_n14633_;
  assign new_n14639_ = ~pi0806 | ~pi0626;
  assign new_n14640_ = ~new_n11464_ | ~pi0965;
  assign new_n14641_ = ~new_n9399_ | ~pi0933;
  assign new_n14642_ = ~pi0773 | ~new_n14633_;
  assign new_n14643_ = ~pi0805 | ~pi0626;
  assign new_n14644_ = ~new_n11464_ | ~pi0964;
  assign new_n14645_ = ~new_n9399_ | ~pi0932;
  assign new_n14646_ = ~pi0772 | ~new_n14633_;
  assign new_n14647_ = ~pi0804 | ~pi0626;
  assign new_n14648_ = ~new_n11464_ | ~pi0963;
  assign new_n14649_ = ~new_n9399_ | ~pi0931;
  assign new_n14650_ = ~pi0771 | ~new_n14633_;
  assign new_n14651_ = ~pi0803 | ~pi0626;
  assign new_n14652_ = ~new_n11464_ | ~pi0962;
  assign new_n14653_ = ~new_n9399_ | ~pi0930;
  assign new_n14654_ = ~pi0770 | ~new_n14633_;
  assign new_n14655_ = ~pi0802 | ~pi0626;
  assign new_n14656_ = ~new_n11464_ | ~pi0961;
  assign new_n14657_ = ~new_n9399_ | ~pi0929;
  assign new_n14658_ = ~pi0797 | ~new_n14633_;
  assign new_n14659_ = ~pi0829 | ~pi0626;
  assign new_n14660_ = ~new_n11464_ | ~pi0988;
  assign new_n14661_ = ~new_n9399_ | ~pi0956;
  assign new_n14662_ = ~pi0796 | ~new_n14633_;
  assign new_n14663_ = ~pi0828 | ~pi0626;
  assign new_n14664_ = ~new_n11464_ | ~pi0987;
  assign new_n14665_ = ~new_n9399_ | ~pi0955;
  assign new_n14666_ = ~pi0769 | ~new_n14633_;
  assign new_n14667_ = ~pi0801 | ~pi0626;
  assign new_n14668_ = ~new_n11464_ | ~pi0960;
  assign new_n14669_ = ~new_n9399_ | ~pi0928;
  assign new_n14670_ = ~pi0795 | ~new_n14633_;
  assign new_n14671_ = ~pi0827 | ~pi0626;
  assign new_n14672_ = ~new_n11464_ | ~pi0986;
  assign new_n14673_ = ~new_n9399_ | ~pi0954;
  assign new_n14674_ = ~pi0794 | ~new_n14633_;
  assign new_n14675_ = ~pi0826 | ~pi0626;
  assign new_n14676_ = ~new_n11464_ | ~pi0985;
  assign new_n14677_ = ~new_n9399_ | ~pi0953;
  assign new_n14678_ = ~pi0793 | ~new_n14633_;
  assign new_n14679_ = ~pi0825 | ~pi0626;
  assign new_n14680_ = ~new_n11464_ | ~pi0984;
  assign new_n14681_ = ~new_n9399_ | ~pi0952;
  assign new_n14682_ = ~pi0792 | ~new_n14633_;
  assign new_n14683_ = ~pi0824 | ~pi0626;
  assign new_n14684_ = ~new_n11464_ | ~pi0983;
  assign new_n14685_ = ~new_n9399_ | ~pi0951;
  assign new_n14686_ = ~pi0791 | ~new_n14633_;
  assign new_n14687_ = ~pi0823 | ~pi0626;
  assign new_n14688_ = ~new_n11464_ | ~pi0982;
  assign new_n14689_ = ~new_n9399_ | ~pi0950;
  assign new_n14690_ = ~pi0790 | ~new_n14633_;
  assign new_n14691_ = ~pi0822 | ~pi0626;
  assign new_n14692_ = ~new_n11464_ | ~pi0981;
  assign new_n14693_ = ~new_n9399_ | ~pi0949;
  assign new_n14694_ = ~pi0789 | ~new_n14633_;
  assign new_n14695_ = ~pi0821 | ~pi0626;
  assign new_n14696_ = ~new_n11464_ | ~pi0980;
  assign new_n14697_ = ~new_n9399_ | ~pi0948;
  assign new_n14698_ = ~pi0788 | ~new_n14633_;
  assign new_n14699_ = ~pi0820 | ~pi0626;
  assign new_n14700_ = ~new_n11464_ | ~pi0979;
  assign new_n14701_ = ~new_n9399_ | ~pi0947;
  assign new_n14702_ = ~pi0787 | ~new_n14633_;
  assign new_n14703_ = ~pi0819 | ~pi0626;
  assign new_n14704_ = ~new_n11464_ | ~pi0978;
  assign new_n14705_ = ~new_n9399_ | ~pi0946;
  assign new_n14706_ = ~pi0786 | ~new_n14633_;
  assign new_n14707_ = ~pi0818 | ~pi0626;
  assign new_n14708_ = ~new_n11464_ | ~pi0977;
  assign new_n14709_ = ~new_n9399_ | ~pi0945;
  assign new_n14710_ = ~pi0768 | ~new_n14633_;
  assign new_n14711_ = ~pi0800 | ~pi0626;
  assign new_n14712_ = ~new_n11464_ | ~pi0959;
  assign new_n14713_ = ~new_n9399_ | ~pi0927;
  assign new_n14714_ = ~pi0785 | ~new_n14633_;
  assign new_n14715_ = ~pi0817 | ~pi0626;
  assign new_n14716_ = ~new_n11464_ | ~pi0976;
  assign new_n14717_ = ~new_n9399_ | ~pi0944;
  assign new_n14718_ = ~pi0784 | ~new_n14633_;
  assign new_n14719_ = ~pi0816 | ~pi0626;
  assign new_n14720_ = ~new_n11464_ | ~pi0975;
  assign new_n14721_ = ~new_n9399_ | ~pi0943;
  assign new_n14722_ = ~pi0783 | ~new_n14633_;
  assign new_n14723_ = ~pi0815 | ~pi0626;
  assign new_n14724_ = ~new_n11464_ | ~pi0974;
  assign new_n14725_ = ~new_n9399_ | ~pi0942;
  assign new_n14726_ = ~pi0782 | ~new_n14633_;
  assign new_n14727_ = ~pi0814 | ~pi0626;
  assign new_n14728_ = ~new_n11464_ | ~pi0973;
  assign new_n14729_ = ~new_n9399_ | ~pi0941;
  assign new_n14730_ = ~pi0781 | ~new_n14633_;
  assign new_n14731_ = ~pi0813 | ~pi0626;
  assign new_n14732_ = ~new_n11464_ | ~pi0972;
  assign new_n14733_ = ~new_n9399_ | ~pi0940;
  assign new_n14734_ = ~pi0780 | ~new_n14633_;
  assign new_n14735_ = ~pi0812 | ~pi0626;
  assign new_n14736_ = ~new_n11464_ | ~pi0971;
  assign new_n14737_ = ~new_n9399_ | ~pi0939;
  assign new_n14738_ = ~pi0779 | ~new_n14633_;
  assign new_n14739_ = ~pi0811 | ~pi0626;
  assign new_n14740_ = ~new_n11464_ | ~pi0970;
  assign new_n14741_ = ~new_n9399_ | ~pi0938;
  assign new_n14742_ = ~pi0778 | ~new_n14633_;
  assign new_n14743_ = ~pi0810 | ~pi0626;
  assign new_n14744_ = ~new_n11464_ | ~pi0969;
  assign new_n14745_ = ~new_n9399_ | ~pi0937;
  assign new_n14746_ = ~pi0777 | ~new_n14633_;
  assign new_n14747_ = ~pi0809 | ~pi0626;
  assign new_n14748_ = ~new_n11464_ | ~pi0968;
  assign new_n14749_ = ~new_n9399_ | ~pi0936;
  assign new_n14750_ = ~pi0776 | ~new_n14633_;
  assign new_n14751_ = ~pi0808 | ~pi0626;
  assign new_n14752_ = ~new_n11464_ | ~pi0967;
  assign new_n14753_ = ~new_n9399_ | ~pi0935;
  assign new_n14754_ = ~pi0767 | ~new_n14633_;
  assign new_n14755_ = ~pi0799 | ~pi0626;
  assign new_n14756_ = ~new_n11464_ | ~pi0958;
  assign new_n14757_ = ~new_n9399_ | ~pi0926;
  assign new_n14758_ = ~new_n11428_ | ~new_n14926_;
  assign new_n14759_ = ~pi0766 | ~new_n14780_;
  assign new_n14760_ = ~pi0798 | ~pi0626;
  assign new_n14761_ = ~new_n11464_ | ~pi0957;
  assign new_n14762_ = ~new_n9399_ | ~pi0925;
  assign new_n14763_ = ~new_n14761_ | ~new_n10616_;
  assign new_n14764_ = ~new_n10591_ | ~new_n10577_;
  assign new_n14765_ = ~new_n29041_ | ~new_n14764_;
  assign new_n14766_ = ~new_n29043_ | ~new_n14764_;
  assign new_n14767_ = ~new_n29508_ | ~new_n9397_;
  assign new_n14768_ = ~pi0756 | ~new_n10325_;
  assign new_n14769_ = ~new_n29509_ | ~new_n9397_;
  assign new_n14770_ = ~pi0757 | ~new_n10325_;
  assign new_n14771_ = ~new_n29510_ | ~new_n9397_;
  assign new_n14772_ = ~pi0758 | ~new_n10325_;
  assign new_n14773_ = ~new_n29511_ | ~new_n9397_;
  assign new_n14774_ = ~pi0759 | ~new_n10325_;
  assign new_n14775_ = ~new_n29496_ | ~new_n9397_;
  assign new_n14776_ = ~pi0760 | ~new_n10325_;
  assign new_n14777_ = ~new_n10566_ | ~new_n10336_ | ~new_n14914_;
  assign new_n14778_ = ~new_n14630_ | ~new_n10313_ | ~new_n11463_ | ~new_n14631_;
  assign new_n14779_ = ~new_n14902_ | ~new_n9658_;
  assign new_n14780_ = ~new_n10326_ | ~new_n10580_ | ~new_n11463_ | ~new_n14632_;
  assign new_n14781_ = ~new_n14785_ | ~new_n12612_ | ~new_n12614_ | ~new_n10562_;
  assign new_n14782_ = ~new_n9432_ | ~new_n10585_;
  assign new_n14783_ = ~new_n9418_ | ~new_n13613_;
  assign new_n14784_ = ~new_n14783_ | ~new_n14782_ | ~new_n11489_;
  assign new_n14785_ = ~new_n14786_ | ~new_n10319_;
  assign new_n14786_ = ~new_n14902_ | ~new_n9658_;
  assign new_n14787_ = ~new_n11633_ | ~new_n15044_ | ~new_n15043_;
  assign new_n14788_ = ~new_n11633_ | ~new_n15012_ | ~new_n15011_;
  assign new_n14789_ = ~new_n11633_ | ~new_n14996_ | ~new_n14995_;
  assign new_n14790_ = ~new_n11633_ | ~new_n15076_ | ~new_n15075_;
  assign new_n14791_ = ~new_n11633_ | ~new_n15060_ | ~new_n15059_;
  assign new_n14792_ = ~new_n11633_ | ~new_n15028_ | ~new_n15027_;
  assign new_n14793_ = ~new_n11633_ | ~new_n14980_ | ~new_n14979_;
  assign new_n14794_ = ~new_n11633_ | ~new_n14964_ | ~new_n14963_;
  assign new_n14795_ = ~new_n11633_ | ~new_n15195_ | ~new_n15194_;
  assign new_n14796_ = ~new_n11633_ | ~new_n15211_ | ~new_n15210_;
  assign new_n14797_ = ~new_n11633_ | ~new_n15227_ | ~new_n15226_;
  assign new_n14798_ = ~new_n11633_ | ~new_n15243_ | ~new_n15242_;
  assign new_n14799_ = ~new_n11633_ | ~new_n15259_ | ~new_n15258_;
  assign new_n14800_ = ~new_n11633_ | ~new_n15275_ | ~new_n15274_;
  assign new_n14801_ = ~new_n11633_ | ~new_n15291_ | ~new_n15290_;
  assign new_n14802_ = ~new_n11633_ | ~new_n15307_ | ~new_n15306_;
  assign new_n14803_ = ~new_n11634_ | ~new_n15046_ | ~new_n15045_;
  assign new_n14804_ = ~new_n11634_ | ~new_n15014_ | ~new_n15013_;
  assign new_n14805_ = ~new_n11634_ | ~new_n14998_ | ~new_n14997_;
  assign new_n14806_ = ~new_n11634_ | ~new_n15078_ | ~new_n15077_;
  assign new_n14807_ = ~new_n11634_ | ~new_n15062_ | ~new_n15061_;
  assign new_n14808_ = ~new_n11634_ | ~new_n15030_ | ~new_n15029_;
  assign new_n14809_ = ~new_n11634_ | ~new_n14982_ | ~new_n14981_;
  assign new_n14810_ = ~new_n11634_ | ~new_n14966_ | ~new_n14965_;
  assign new_n14811_ = ~new_n11634_ | ~new_n15197_ | ~new_n15196_;
  assign new_n14812_ = ~new_n11634_ | ~new_n15213_ | ~new_n15212_;
  assign new_n14813_ = ~new_n11634_ | ~new_n15229_ | ~new_n15228_;
  assign new_n14814_ = ~new_n11634_ | ~new_n15245_ | ~new_n15244_;
  assign new_n14815_ = ~new_n11634_ | ~new_n15261_ | ~new_n15260_;
  assign new_n14816_ = ~new_n11634_ | ~new_n15277_ | ~new_n15276_;
  assign new_n14817_ = ~new_n11634_ | ~new_n15293_ | ~new_n15292_;
  assign new_n14818_ = ~new_n11634_ | ~new_n15309_ | ~new_n15308_;
  assign new_n14819_ = ~new_n9497_ | ~new_n15048_ | ~new_n15047_;
  assign new_n14820_ = ~new_n9497_ | ~new_n15016_ | ~new_n15015_;
  assign new_n14821_ = ~new_n9497_ | ~new_n15000_ | ~new_n14999_;
  assign new_n14822_ = ~new_n9497_ | ~new_n15080_ | ~new_n15079_;
  assign new_n14823_ = ~new_n9497_ | ~new_n15064_ | ~new_n15063_;
  assign new_n14824_ = ~new_n9497_ | ~new_n15032_ | ~new_n15031_;
  assign new_n14825_ = ~new_n9497_ | ~new_n14984_ | ~new_n14983_;
  assign new_n14826_ = ~new_n9497_ | ~new_n14968_ | ~new_n14967_;
  assign new_n14827_ = ~new_n9497_ | ~new_n15199_ | ~new_n15198_;
  assign new_n14828_ = ~new_n9497_ | ~new_n15215_ | ~new_n15214_;
  assign new_n14829_ = ~new_n9497_ | ~new_n15231_ | ~new_n15230_;
  assign new_n14830_ = ~new_n9497_ | ~new_n15247_ | ~new_n15246_;
  assign new_n14831_ = ~new_n9497_ | ~new_n15263_ | ~new_n15262_;
  assign new_n14832_ = ~new_n9497_ | ~new_n15279_ | ~new_n15278_;
  assign new_n14833_ = ~new_n9497_ | ~new_n15295_ | ~new_n15294_;
  assign new_n14834_ = ~new_n9497_ | ~new_n15311_ | ~new_n15310_;
  assign new_n14835_ = ~new_n9495_ | ~new_n15050_ | ~new_n15049_;
  assign new_n14836_ = ~new_n9495_ | ~new_n15018_ | ~new_n15017_;
  assign new_n14837_ = ~new_n9495_ | ~new_n15002_ | ~new_n15001_;
  assign new_n14838_ = ~new_n9495_ | ~new_n15082_ | ~new_n15081_;
  assign new_n14839_ = ~new_n9495_ | ~new_n15066_ | ~new_n15065_;
  assign new_n14840_ = ~new_n9495_ | ~new_n15034_ | ~new_n15033_;
  assign new_n14841_ = ~new_n9495_ | ~new_n14986_ | ~new_n14985_;
  assign new_n14842_ = ~new_n9495_ | ~new_n14970_ | ~new_n14969_;
  assign new_n14843_ = ~new_n9495_ | ~new_n15201_ | ~new_n15200_;
  assign new_n14844_ = ~new_n9495_ | ~new_n15217_ | ~new_n15216_;
  assign new_n14845_ = ~new_n9495_ | ~new_n15233_ | ~new_n15232_;
  assign new_n14846_ = ~new_n9495_ | ~new_n15249_ | ~new_n15248_;
  assign new_n14847_ = ~new_n9495_ | ~new_n15265_ | ~new_n15264_;
  assign new_n14848_ = ~new_n9495_ | ~new_n15281_ | ~new_n15280_;
  assign new_n14849_ = ~new_n9495_ | ~new_n15297_ | ~new_n15296_;
  assign new_n14850_ = ~new_n9495_ | ~new_n15313_ | ~new_n15312_;
  assign new_n14851_ = ~new_n11631_ | ~new_n15052_ | ~new_n15051_;
  assign new_n14852_ = ~new_n11631_ | ~new_n15020_ | ~new_n15019_;
  assign new_n14853_ = ~new_n11631_ | ~new_n15004_ | ~new_n15003_;
  assign new_n14854_ = ~new_n11631_ | ~new_n15084_ | ~new_n15083_;
  assign new_n14855_ = ~new_n11631_ | ~new_n15068_ | ~new_n15067_;
  assign new_n14856_ = ~new_n11631_ | ~new_n15036_ | ~new_n15035_;
  assign new_n14857_ = ~new_n11631_ | ~new_n14988_ | ~new_n14987_;
  assign new_n14858_ = ~new_n11631_ | ~new_n14972_ | ~new_n14971_;
  assign new_n14859_ = ~new_n11631_ | ~new_n15203_ | ~new_n15202_;
  assign new_n14860_ = ~new_n11631_ | ~new_n15219_ | ~new_n15218_;
  assign new_n14861_ = ~new_n11631_ | ~new_n15235_ | ~new_n15234_;
  assign new_n14862_ = ~new_n11631_ | ~new_n15251_ | ~new_n15250_;
  assign new_n14863_ = ~new_n11631_ | ~new_n15267_ | ~new_n15266_;
  assign new_n14864_ = ~new_n11631_ | ~new_n15283_ | ~new_n15282_;
  assign new_n14865_ = ~new_n11631_ | ~new_n15299_ | ~new_n15298_;
  assign new_n14866_ = ~new_n11631_ | ~new_n15315_ | ~new_n15314_;
  assign new_n14867_ = ~new_n9494_ | ~new_n15054_ | ~new_n15053_;
  assign new_n14868_ = ~new_n9494_ | ~new_n15022_ | ~new_n15021_;
  assign new_n14869_ = ~new_n9494_ | ~new_n15006_ | ~new_n15005_;
  assign new_n14870_ = ~new_n9494_ | ~new_n15086_ | ~new_n15085_;
  assign new_n14871_ = ~new_n9494_ | ~new_n15070_ | ~new_n15069_;
  assign new_n14872_ = ~new_n9494_ | ~new_n15038_ | ~new_n15037_;
  assign new_n14873_ = ~new_n9494_ | ~new_n14990_ | ~new_n14989_;
  assign new_n14874_ = ~new_n9494_ | ~new_n14974_ | ~new_n14973_;
  assign new_n14875_ = ~new_n9494_ | ~new_n15205_ | ~new_n15204_;
  assign new_n14876_ = ~new_n9494_ | ~new_n15221_ | ~new_n15220_;
  assign new_n14877_ = ~new_n9494_ | ~new_n15237_ | ~new_n15236_;
  assign new_n14878_ = ~new_n9494_ | ~new_n15253_ | ~new_n15252_;
  assign new_n14879_ = ~new_n9494_ | ~new_n15269_ | ~new_n15268_;
  assign new_n14880_ = ~new_n9494_ | ~new_n15285_ | ~new_n15284_;
  assign new_n14881_ = ~new_n9494_ | ~new_n15301_ | ~new_n15300_;
  assign new_n14882_ = ~new_n9494_ | ~new_n15317_ | ~new_n15316_;
  assign new_n14883_ = ~new_n9493_ | ~new_n15056_ | ~new_n15055_;
  assign new_n14884_ = ~new_n9493_ | ~new_n15024_ | ~new_n15023_;
  assign new_n14885_ = ~new_n9493_ | ~new_n15008_ | ~new_n15007_;
  assign new_n14886_ = ~new_n9493_ | ~new_n15088_ | ~new_n15087_;
  assign new_n14887_ = ~new_n9493_ | ~new_n15072_ | ~new_n15071_;
  assign new_n14888_ = ~new_n9493_ | ~new_n15040_ | ~new_n15039_;
  assign new_n14889_ = ~new_n9493_ | ~new_n14992_ | ~new_n14991_;
  assign new_n14890_ = ~new_n9493_ | ~new_n14976_ | ~new_n14975_;
  assign new_n14891_ = ~new_n9493_ | ~new_n15207_ | ~new_n15206_;
  assign new_n14892_ = ~new_n9493_ | ~new_n15223_ | ~new_n15222_;
  assign new_n14893_ = ~new_n9493_ | ~new_n15239_ | ~new_n15238_;
  assign new_n14894_ = ~new_n9493_ | ~new_n15255_ | ~new_n15254_;
  assign new_n14895_ = ~new_n9493_ | ~new_n15271_ | ~new_n15270_;
  assign new_n14896_ = ~new_n9493_ | ~new_n15287_ | ~new_n15286_;
  assign new_n14897_ = ~new_n9493_ | ~new_n15303_ | ~new_n15302_;
  assign new_n14898_ = ~new_n9493_ | ~new_n15319_ | ~new_n15318_;
  assign new_n14899_ = ~new_n9496_ | ~new_n15058_ | ~new_n15057_;
  assign new_n14900_ = ~new_n10321_;
  assign new_n14901_ = ~new_n9496_ | ~new_n15026_ | ~new_n15025_;
  assign new_n14902_ = ~new_n10320_;
  assign new_n14903_ = ~new_n9496_ | ~new_n15010_ | ~new_n15009_;
  assign new_n14904_ = ~new_n10319_;
  assign new_n14905_ = ~new_n9496_ | ~new_n15090_ | ~new_n15089_;
  assign new_n14906_ = ~new_n10562_;
  assign new_n14907_ = ~new_n9496_ | ~new_n15074_ | ~new_n15073_;
  assign new_n14908_ = ~new_n10296_;
  assign new_n14909_ = ~new_n9496_ | ~new_n15042_ | ~new_n15041_;
  assign new_n14910_ = ~new_n9658_;
  assign new_n14911_ = ~new_n9496_ | ~new_n14994_ | ~new_n14993_;
  assign new_n14912_ = ~new_n10294_;
  assign new_n14913_ = ~new_n9496_ | ~new_n14978_ | ~new_n14977_;
  assign new_n14914_ = ~new_n9657_;
  assign new_n14915_ = ~new_n9496_ | ~new_n15209_ | ~new_n15208_;
  assign new_n14916_ = ~new_n9496_ | ~new_n15225_ | ~new_n15224_;
  assign new_n14917_ = ~new_n9496_ | ~new_n15241_ | ~new_n15240_;
  assign new_n14918_ = ~new_n9496_ | ~new_n15257_ | ~new_n15256_;
  assign new_n14919_ = ~new_n9496_ | ~new_n15273_ | ~new_n15272_;
  assign new_n14920_ = ~new_n9496_ | ~new_n15289_ | ~new_n15288_;
  assign new_n14921_ = ~new_n9496_ | ~new_n15305_ | ~new_n15304_;
  assign new_n14922_ = ~new_n9496_ | ~new_n15321_ | ~new_n15320_;
  assign new_n14923_ = ~new_n12631_ | ~new_n11469_;
  assign new_n14924_ = ~new_n12637_ | ~new_n10566_;
  assign new_n14925_ = ~new_n11637_ | ~new_n14924_;
  assign new_n14926_ = ~new_n10294_ | ~new_n15389_ | ~new_n15388_;
  assign new_n14927_ = ~new_n14763_ | ~new_n12630_;
  assign new_n14928_ = ~new_n11500_ | ~new_n12630_;
  assign new_n14929_ = ~new_n11427_ | ~new_n11425_ | ~new_n11426_ | ~new_n9630_ | ~new_n14928_;
  assign new_n14930_ = ~new_n11500_ | ~new_n12630_;
  assign new_n14931_ = ~new_n11499_ | ~new_n11420_ | ~new_n9630_ | ~new_n14930_;
  assign new_n14932_ = ~new_n11610_ | ~new_n11613_ | ~pi0590;
  assign new_n14933_ = ~pi0591 | ~pi0997 | ~new_n10285_;
  assign new_n14934_ = ~pi0590 | ~new_n11610_;
  assign new_n14935_ = ~new_n11641_ | ~new_n11656_;
  assign new_n14936_ = ~new_n14904_ | ~new_n14912_;
  assign new_n14937_ = ~new_n10296_ | ~new_n12636_;
  assign new_n14938_ = ~new_n11470_ | ~new_n12630_;
  assign new_n14939_ = ~pi0957 | ~pi0592;
  assign new_n14940_ = ~pi0555 | ~new_n10300_;
  assign new_n14941_ = ~pi0989 | ~new_n11480_;
  assign new_n14942_ = ~pi0556 | ~new_n10300_;
  assign new_n14943_ = ~pi0990 | ~new_n11480_;
  assign new_n14944_ = ~pi0557 | ~new_n10300_;
  assign new_n14945_ = ~pi0991 | ~new_n11480_;
  assign new_n14946_ = ~pi0558 | ~new_n10300_;
  assign new_n14947_ = ~pi0992 | ~new_n11480_;
  assign new_n14948_ = ~pi0591 | ~new_n10309_ | ~new_n10308_;
  assign new_n14949_ = pi0034 | pi0591;
  assign new_n14950_ = ~pi0589 | ~new_n10307_;
  assign new_n14951_ = ~new_n11609_ | ~pi0591;
  assign new_n14952_ = ~pi0590 | ~new_n11622_ | ~new_n11613_;
  assign new_n14953_ = ~new_n11623_ | ~new_n10299_;
  assign new_n14954_ = ~pi0589 | ~pi0591 | ~new_n10308_;
  assign new_n14955_ = ~new_n11625_ | ~new_n10285_;
  assign new_n14956_ = pi0591 | pi0590;
  assign new_n14957_ = ~pi0591 | ~new_n11514_;
  assign new_n14958_ = ~new_n10630_;
  assign new_n14959_ = ~new_n14958_ | ~pi0592;
  assign new_n14960_ = ~new_n10631_ | ~new_n10630_;
  assign new_n14961_ = ~new_n10630_ | ~new_n11630_;
  assign new_n14962_ = ~new_n14958_ | ~pi0593;
  assign new_n14963_ = ~pi0757 | ~new_n10429_;
  assign new_n14964_ = pi0757 | pi0730;
  assign new_n14965_ = pi0757 | pi0754;
  assign new_n14966_ = ~pi0757 | ~new_n10463_;
  assign new_n14967_ = pi0757 | pi0746;
  assign new_n14968_ = ~pi0757 | ~new_n10452_;
  assign new_n14969_ = ~pi0757 | ~new_n10415_;
  assign new_n14970_ = pi0757 | pi0722;
  assign new_n14971_ = ~pi0757 | ~new_n10374_;
  assign new_n14972_ = pi0757 | pi0698;
  assign new_n14973_ = ~pi0757 | ~new_n10404_;
  assign new_n14974_ = pi0757 | pi0714;
  assign new_n14975_ = ~pi0757 | ~new_n10388_;
  assign new_n14976_ = pi0757 | pi0706;
  assign new_n14977_ = ~pi0757 | ~new_n10440_;
  assign new_n14978_ = pi0757 | pi0738;
  assign new_n14979_ = ~pi0757 | ~new_n10430_;
  assign new_n14980_ = pi0757 | pi0731;
  assign new_n14981_ = pi0757 | pi0755;
  assign new_n14982_ = ~pi0757 | ~new_n10464_;
  assign new_n14983_ = pi0757 | pi0747;
  assign new_n14984_ = ~pi0757 | ~new_n10453_;
  assign new_n14985_ = ~pi0757 | ~new_n10416_;
  assign new_n14986_ = pi0757 | pi0723;
  assign new_n14987_ = ~pi0757 | ~new_n10375_;
  assign new_n14988_ = pi0757 | pi0699;
  assign new_n14989_ = ~pi0757 | ~new_n10405_;
  assign new_n14990_ = pi0757 | pi0715;
  assign new_n14991_ = ~pi0757 | ~new_n10389_;
  assign new_n14992_ = pi0757 | pi0707;
  assign new_n14993_ = ~pi0757 | ~new_n10441_;
  assign new_n14994_ = pi0757 | pi0739;
  assign new_n14995_ = ~pi0757 | ~new_n10426_;
  assign new_n14996_ = pi0757 | pi0727;
  assign new_n14997_ = pi0757 | pi0751;
  assign new_n14998_ = ~pi0757 | ~new_n10460_;
  assign new_n14999_ = pi0757 | pi0743;
  assign new_n15000_ = ~pi0757 | ~new_n10449_;
  assign new_n15001_ = ~pi0757 | ~new_n10412_;
  assign new_n15002_ = pi0757 | pi0719;
  assign new_n15003_ = ~pi0757 | ~new_n10371_;
  assign new_n15004_ = pi0757 | pi0695;
  assign new_n15005_ = ~pi0757 | ~new_n10401_;
  assign new_n15006_ = pi0757 | pi0711;
  assign new_n15007_ = ~pi0757 | ~new_n10385_;
  assign new_n15008_ = pi0757 | pi0703;
  assign new_n15009_ = ~pi0757 | ~new_n10437_;
  assign new_n15010_ = pi0757 | pi0735;
  assign new_n15011_ = ~pi0757 | ~new_n10424_;
  assign new_n15012_ = pi0757 | pi0725;
  assign new_n15013_ = pi0757 | pi0749;
  assign new_n15014_ = ~pi0757 | ~new_n10458_;
  assign new_n15015_ = pi0757 | pi0741;
  assign new_n15016_ = ~pi0757 | ~new_n10447_;
  assign new_n15017_ = ~pi0757 | ~new_n10410_;
  assign new_n15018_ = pi0757 | pi0717;
  assign new_n15019_ = ~pi0757 | ~new_n10369_;
  assign new_n15020_ = pi0757 | pi0693;
  assign new_n15021_ = ~pi0757 | ~new_n10399_;
  assign new_n15022_ = pi0757 | pi0709;
  assign new_n15023_ = ~pi0757 | ~new_n10383_;
  assign new_n15024_ = pi0757 | pi0701;
  assign new_n15025_ = ~pi0757 | ~new_n10435_;
  assign new_n15026_ = pi0757 | pi0733;
  assign new_n15027_ = ~pi0757 | ~new_n10425_;
  assign new_n15028_ = pi0757 | pi0726;
  assign new_n15029_ = pi0757 | pi0750;
  assign new_n15030_ = ~pi0757 | ~new_n10459_;
  assign new_n15031_ = pi0757 | pi0742;
  assign new_n15032_ = ~pi0757 | ~new_n10448_;
  assign new_n15033_ = ~pi0757 | ~new_n10411_;
  assign new_n15034_ = pi0757 | pi0718;
  assign new_n15035_ = ~pi0757 | ~new_n10370_;
  assign new_n15036_ = pi0757 | pi0694;
  assign new_n15037_ = ~pi0757 | ~new_n10400_;
  assign new_n15038_ = pi0757 | pi0710;
  assign new_n15039_ = ~pi0757 | ~new_n10384_;
  assign new_n15040_ = pi0757 | pi0702;
  assign new_n15041_ = ~pi0757 | ~new_n10436_;
  assign new_n15042_ = pi0757 | pi0734;
  assign new_n15043_ = ~pi0757 | ~new_n10428_;
  assign new_n15044_ = pi0757 | pi0729;
  assign new_n15045_ = pi0757 | pi0753;
  assign new_n15046_ = ~pi0757 | ~new_n10462_;
  assign new_n15047_ = pi0757 | pi0745;
  assign new_n15048_ = ~pi0757 | ~new_n10451_;
  assign new_n15049_ = ~pi0757 | ~new_n10414_;
  assign new_n15050_ = pi0757 | pi0721;
  assign new_n15051_ = ~pi0757 | ~new_n10373_;
  assign new_n15052_ = pi0757 | pi0697;
  assign new_n15053_ = ~pi0757 | ~new_n10403_;
  assign new_n15054_ = pi0757 | pi0713;
  assign new_n15055_ = ~pi0757 | ~new_n10387_;
  assign new_n15056_ = pi0757 | pi0705;
  assign new_n15057_ = ~pi0757 | ~new_n10439_;
  assign new_n15058_ = pi0757 | pi0737;
  assign new_n15059_ = ~pi0757 | ~new_n10427_;
  assign new_n15060_ = pi0757 | pi0728;
  assign new_n15061_ = pi0757 | pi0752;
  assign new_n15062_ = ~pi0757 | ~new_n10461_;
  assign new_n15063_ = pi0757 | pi0744;
  assign new_n15064_ = ~pi0757 | ~new_n10450_;
  assign new_n15065_ = ~pi0757 | ~new_n10413_;
  assign new_n15066_ = pi0757 | pi0720;
  assign new_n15067_ = ~pi0757 | ~new_n10372_;
  assign new_n15068_ = pi0757 | pi0696;
  assign new_n15069_ = ~pi0757 | ~new_n10402_;
  assign new_n15070_ = pi0757 | pi0712;
  assign new_n15071_ = ~pi0757 | ~new_n10386_;
  assign new_n15072_ = pi0757 | pi0704;
  assign new_n15073_ = ~pi0757 | ~new_n10438_;
  assign new_n15074_ = pi0757 | pi0736;
  assign new_n15075_ = ~pi0757 | ~new_n10423_;
  assign new_n15076_ = pi0757 | pi0724;
  assign new_n15077_ = pi0757 | pi0748;
  assign new_n15078_ = ~pi0757 | ~new_n10457_;
  assign new_n15079_ = pi0757 | pi0740;
  assign new_n15080_ = ~pi0757 | ~new_n10446_;
  assign new_n15081_ = ~pi0757 | ~new_n10409_;
  assign new_n15082_ = pi0757 | pi0716;
  assign new_n15083_ = ~pi0757 | ~new_n10368_;
  assign new_n15084_ = pi0757 | pi0692;
  assign new_n15085_ = ~pi0757 | ~new_n10398_;
  assign new_n15086_ = pi0757 | pi0708;
  assign new_n15087_ = ~pi0757 | ~new_n10382_;
  assign new_n15088_ = pi0757 | pi0700;
  assign new_n15089_ = ~pi0757 | ~new_n10434_;
  assign new_n15090_ = pi0757 | pi0732;
  assign new_n15091_ = ~new_n28599_ | ~new_n11476_;
  assign new_n15092_ = ~new_n11645_ | ~new_n10338_;
  assign new_n15093_ = ~new_n14912_ | ~new_n10334_;
  assign new_n15094_ = ~new_n10294_ | ~new_n10323_;
  assign new_n15095_ = ~new_n11468_ | ~new_n10338_;
  assign new_n15096_ = ~new_n10330_ | ~new_n10561_;
  assign new_n15097_ = new_n2973_ | pi0627;
  assign new_n15098_ = ~pi0627 | ~new_n11658_;
  assign new_n15099_ = ~pi0624 | ~new_n10340_;
  assign new_n15100_ = ~new_n9489_ | ~new_n11661_;
  assign new_n15101_ = ~pi0627 | ~new_n11672_;
  assign new_n15102_ = ~new_n10325_ | ~new_n11671_ | ~new_n11660_;
  assign new_n15103_ = ~new_n28333_ | ~new_n10359_;
  assign new_n15104_ = ~new_n11678_ | ~new_n10357_;
  assign new_n15105_ = ~new_n10620_;
  assign new_n15106_ = ~pi0763 | ~new_n10352_;
  assign new_n15107_ = ~new_n11683_ | ~new_n10351_;
  assign new_n15108_ = ~new_n10621_;
  assign new_n15109_ = ~new_n14900_ | ~new_n12615_;
  assign new_n15110_ = ~new_n10321_ | ~new_n12616_;
  assign new_n15111_ = ~new_n11476_ | ~new_n10338_;
  assign new_n15112_ = ~new_n28599_ | ~new_n11474_ | ~new_n9400_;
  assign new_n15113_ = ~new_n10635_ | ~new_n11435_;
  assign new_n15114_ = ~new_n12625_ | ~pi0756;
  assign new_n15115_ = ~new_n10321_ | ~new_n12627_;
  assign new_n15116_ = ~new_n14900_ | ~new_n9658_ | ~new_n10320_;
  assign new_n15117_ = ~new_n11465_ | ~new_n10294_;
  assign new_n15118_ = ~new_n11516_ | ~new_n14912_;
  assign new_n15119_ = ~pi0757 | ~new_n12626_;
  assign new_n15120_ = ~new_n10314_ | ~new_n11632_ | ~new_n10317_;
  assign new_n15121_ = ~pi0757 | ~new_n10318_;
  assign new_n15122_ = ~new_n11631_ | ~new_n10314_;
  assign new_n15123_ = ~new_n10622_;
  assign new_n15124_ = ~new_n12625_ | ~pi0757;
  assign new_n15125_ = ~new_n12655_ | ~new_n11435_;
  assign new_n15126_ = ~pi0766 | ~new_n10569_;
  assign new_n15127_ = ~new_n10688_ | ~new_n10724_;
  assign new_n15128_ = ~new_n10638_;
  assign new_n15129_ = ~pi0767 | ~new_n10569_;
  assign new_n15130_ = ~new_n29599_ | ~new_n10688_;
  assign new_n15131_ = ~new_n10639_;
  assign new_n15132_ = ~new_n12657_ | ~new_n12646_;
  assign new_n15133_ = ~new_n10571_ | ~new_n12647_;
  assign new_n15134_ = ~new_n12625_ | ~pi0758;
  assign new_n15135_ = ~new_n12664_ | ~new_n11435_;
  assign new_n15136_ = ~new_n10296_ | ~new_n10927_ | ~new_n11638_;
  assign new_n15137_ = ~new_n14908_ | ~new_n14910_ | ~new_n12666_;
  assign new_n15138_ = ~new_n15137_ | ~new_n15136_;
  assign new_n15139_ = ~pi0760 | ~new_n10312_;
  assign new_n15140_ = ~pi0759 | ~new_n10313_;
  assign new_n15141_ = ~new_n10623_;
  assign new_n15142_ = ~new_n12625_ | ~pi0759;
  assign new_n15143_ = ~new_n12674_ | ~new_n11435_;
  assign new_n15144_ = ~new_n12625_ | ~pi0760;
  assign new_n15145_ = ~new_n12682_ | ~new_n11435_;
  assign new_n15146_ = ~new_n12684_ | ~pi0762;
  assign new_n15147_ = ~new_n12692_ | ~new_n10574_;
  assign new_n15148_ = ~new_n15105_ | ~new_n11677_;
  assign new_n15149_ = ~new_n10620_ | ~new_n10360_;
  assign new_n15150_ = ~new_n15149_ | ~new_n15148_;
  assign new_n15151_ = ~new_n12684_ | ~pi0763;
  assign new_n15152_ = ~new_n12696_ | ~new_n10574_;
  assign new_n15153_ = ~new_n12684_ | ~pi0764;
  assign new_n15154_ = ~new_n12701_ | ~new_n10574_;
  assign new_n15155_ = ~new_n12684_ | ~pi0765;
  assign new_n15156_ = ~new_n12705_ | ~new_n10574_;
  assign new_n15157_ = ~new_n9657_ | ~new_n9400_ | ~new_n10321_;
  assign new_n15158_ = ~new_n9479_ | ~new_n14914_;
  assign new_n15159_ = ~new_n15158_ | ~new_n15157_;
  assign new_n15160_ = ~new_n10338_ | ~new_n10294_ | ~new_n10319_;
  assign new_n15161_ = ~new_n15159_ | ~new_n28599_;
  assign new_n15162_ = ~new_n14900_ | ~new_n14914_;
  assign new_n15163_ = ~new_n9657_ | ~new_n10323_;
  assign new_n15164_ = ~pi0989 | ~new_n10588_;
  assign new_n15165_ = ~new_n10647_ | ~new_n11479_;
  assign new_n15166_ = ~pi0990 | ~new_n10588_;
  assign new_n15167_ = ~new_n10648_ | ~new_n11479_;
  assign new_n15168_ = ~pi0992 | ~new_n10588_;
  assign new_n15169_ = ~new_n11479_ | ~pi0957;
  assign new_n15170_ = ~new_n11480_ | ~new_n10593_;
  assign new_n15171_ = ~pi0993 | ~new_n10300_;
  assign new_n15172_ = ~new_n10328_ | ~new_n14914_;
  assign new_n15173_ = ~new_n29132_ | ~new_n9657_;
  assign new_n15174_ = ~new_n13879_ | ~new_n10298_;
  assign new_n15175_ = ~pi0995 | ~new_n11441_;
  assign new_n15176_ = ~new_n14958_ | ~pi0996;
  assign new_n15177_ = ~pi0035 | ~new_n10630_;
  assign new_n15178_ = ~new_n13884_ | ~pi0997;
  assign new_n15179_ = ~new_n13893_ | ~new_n11443_;
  assign new_n15180_ = ~new_n11480_ | ~new_n10592_;
  assign new_n15181_ = ~pi0998 | ~new_n10300_;
  assign new_n15182_ = ~pi0999 | ~new_n10300_;
  assign new_n15183_ = ~pi1003 | ~new_n11480_;
  assign new_n15184_ = ~new_n13898_ | ~pi1002;
  assign new_n15185_ = ~new_n13899_ | ~new_n11444_;
  assign new_n15186_ = ~new_n14914_ | ~new_n10561_;
  assign new_n15187_ = ~new_n9657_ | ~new_n10338_;
  assign new_n15188_ = ~pi0757 | ~new_n11446_;
  assign new_n15189_ = ~new_n14048_ | ~new_n10314_;
  assign new_n15190_ = ~new_n10624_;
  assign new_n15191_ = ~pi0758 | ~new_n10314_;
  assign new_n15192_ = ~pi0757 | ~new_n10317_;
  assign new_n15193_ = ~new_n10625_;
  assign new_n15194_ = ~new_n10625_ | ~new_n10368_;
  assign new_n15195_ = ~new_n15193_ | ~new_n10472_;
  assign new_n15196_ = ~new_n10625_ | ~new_n10409_;
  assign new_n15197_ = ~new_n15193_ | ~new_n10506_;
  assign new_n15198_ = ~new_n10625_ | ~new_n10398_;
  assign new_n15199_ = ~new_n15193_ | ~new_n10495_;
  assign new_n15200_ = ~new_n10625_ | ~new_n10457_;
  assign new_n15201_ = ~new_n15193_ | ~new_n10552_;
  assign new_n15202_ = ~new_n10625_ | ~new_n10423_;
  assign new_n15203_ = ~new_n15193_ | ~new_n10518_;
  assign new_n15204_ = ~new_n10625_ | ~new_n10446_;
  assign new_n15205_ = ~new_n15193_ | ~new_n10541_;
  assign new_n15206_ = ~new_n10625_ | ~new_n10434_;
  assign new_n15207_ = ~new_n15193_ | ~new_n10529_;
  assign new_n15208_ = ~new_n10625_ | ~new_n10382_;
  assign new_n15209_ = ~new_n15193_ | ~new_n10483_;
  assign new_n15210_ = ~new_n10625_ | ~new_n10369_;
  assign new_n15211_ = ~new_n15193_ | ~new_n10473_;
  assign new_n15212_ = ~new_n10625_ | ~new_n10410_;
  assign new_n15213_ = ~new_n15193_ | ~new_n10507_;
  assign new_n15214_ = ~new_n10625_ | ~new_n10399_;
  assign new_n15215_ = ~new_n15193_ | ~new_n10496_;
  assign new_n15216_ = ~new_n10625_ | ~new_n10458_;
  assign new_n15217_ = ~new_n15193_ | ~new_n10553_;
  assign new_n15218_ = ~new_n10625_ | ~new_n10424_;
  assign new_n15219_ = ~new_n15193_ | ~new_n10519_;
  assign new_n15220_ = ~new_n10625_ | ~new_n10447_;
  assign new_n15221_ = ~new_n15193_ | ~new_n10542_;
  assign new_n15222_ = ~new_n10625_ | ~new_n10435_;
  assign new_n15223_ = ~new_n15193_ | ~new_n10530_;
  assign new_n15224_ = ~new_n10625_ | ~new_n10383_;
  assign new_n15225_ = ~new_n15193_ | ~new_n10484_;
  assign new_n15226_ = ~new_n10625_ | ~new_n10370_;
  assign new_n15227_ = ~new_n15193_ | ~new_n10474_;
  assign new_n15228_ = ~new_n10625_ | ~new_n10411_;
  assign new_n15229_ = ~new_n15193_ | ~new_n10508_;
  assign new_n15230_ = ~new_n10625_ | ~new_n10400_;
  assign new_n15231_ = ~new_n15193_ | ~new_n10497_;
  assign new_n15232_ = ~new_n10625_ | ~new_n10459_;
  assign new_n15233_ = ~new_n15193_ | ~new_n10554_;
  assign new_n15234_ = ~new_n10625_ | ~new_n10425_;
  assign new_n15235_ = ~new_n15193_ | ~new_n10520_;
  assign new_n15236_ = ~new_n10625_ | ~new_n10448_;
  assign new_n15237_ = ~new_n15193_ | ~new_n10543_;
  assign new_n15238_ = ~new_n10625_ | ~new_n10436_;
  assign new_n15239_ = ~new_n15193_ | ~new_n10531_;
  assign new_n15240_ = ~new_n10625_ | ~new_n10384_;
  assign new_n15241_ = ~new_n15193_ | ~new_n10485_;
  assign new_n15242_ = ~new_n10625_ | ~new_n10371_;
  assign new_n15243_ = ~new_n15193_ | ~new_n10475_;
  assign new_n15244_ = ~new_n10625_ | ~new_n10412_;
  assign new_n15245_ = ~new_n15193_ | ~new_n10509_;
  assign new_n15246_ = ~new_n10625_ | ~new_n10401_;
  assign new_n15247_ = ~new_n15193_ | ~new_n10498_;
  assign new_n15248_ = ~new_n10625_ | ~new_n10460_;
  assign new_n15249_ = ~new_n15193_ | ~new_n10555_;
  assign new_n15250_ = ~new_n10625_ | ~new_n10426_;
  assign new_n15251_ = ~new_n15193_ | ~new_n10521_;
  assign new_n15252_ = ~new_n10625_ | ~new_n10449_;
  assign new_n15253_ = ~new_n15193_ | ~new_n10544_;
  assign new_n15254_ = ~new_n10625_ | ~new_n10437_;
  assign new_n15255_ = ~new_n15193_ | ~new_n10532_;
  assign new_n15256_ = ~new_n10625_ | ~new_n10385_;
  assign new_n15257_ = ~new_n15193_ | ~new_n10486_;
  assign new_n15258_ = ~new_n10625_ | ~new_n10372_;
  assign new_n15259_ = ~new_n15193_ | ~new_n10476_;
  assign new_n15260_ = ~new_n10625_ | ~new_n10413_;
  assign new_n15261_ = ~new_n15193_ | ~new_n10510_;
  assign new_n15262_ = ~new_n10625_ | ~new_n10402_;
  assign new_n15263_ = ~new_n15193_ | ~new_n10499_;
  assign new_n15264_ = ~new_n10625_ | ~new_n10461_;
  assign new_n15265_ = ~new_n15193_ | ~new_n10556_;
  assign new_n15266_ = ~new_n10625_ | ~new_n10427_;
  assign new_n15267_ = ~new_n15193_ | ~new_n10522_;
  assign new_n15268_ = ~new_n10625_ | ~new_n10450_;
  assign new_n15269_ = ~new_n15193_ | ~new_n10545_;
  assign new_n15270_ = ~new_n10625_ | ~new_n10438_;
  assign new_n15271_ = ~new_n15193_ | ~new_n10533_;
  assign new_n15272_ = ~new_n10625_ | ~new_n10386_;
  assign new_n15273_ = ~new_n15193_ | ~new_n10487_;
  assign new_n15274_ = ~new_n10625_ | ~new_n10373_;
  assign new_n15275_ = ~new_n15193_ | ~new_n10477_;
  assign new_n15276_ = ~new_n10625_ | ~new_n10414_;
  assign new_n15277_ = ~new_n15193_ | ~new_n10511_;
  assign new_n15278_ = ~new_n10625_ | ~new_n10403_;
  assign new_n15279_ = ~new_n15193_ | ~new_n10500_;
  assign new_n15280_ = ~new_n10625_ | ~new_n10462_;
  assign new_n15281_ = ~new_n15193_ | ~new_n10557_;
  assign new_n15282_ = ~new_n10625_ | ~new_n10428_;
  assign new_n15283_ = ~new_n15193_ | ~new_n10523_;
  assign new_n15284_ = ~new_n10625_ | ~new_n10451_;
  assign new_n15285_ = ~new_n15193_ | ~new_n10546_;
  assign new_n15286_ = ~new_n10625_ | ~new_n10439_;
  assign new_n15287_ = ~new_n15193_ | ~new_n10534_;
  assign new_n15288_ = ~new_n10625_ | ~new_n10387_;
  assign new_n15289_ = ~new_n15193_ | ~new_n10488_;
  assign new_n15290_ = ~new_n10625_ | ~new_n10374_;
  assign new_n15291_ = ~new_n15193_ | ~new_n10478_;
  assign new_n15292_ = ~new_n10625_ | ~new_n10415_;
  assign new_n15293_ = ~new_n15193_ | ~new_n10512_;
  assign new_n15294_ = ~new_n10625_ | ~new_n10404_;
  assign new_n15295_ = ~new_n15193_ | ~new_n10501_;
  assign new_n15296_ = ~new_n10625_ | ~new_n10463_;
  assign new_n15297_ = ~new_n15193_ | ~new_n10558_;
  assign new_n15298_ = ~new_n10625_ | ~new_n10429_;
  assign new_n15299_ = ~new_n15193_ | ~new_n10524_;
  assign new_n15300_ = ~new_n10625_ | ~new_n10452_;
  assign new_n15301_ = ~new_n15193_ | ~new_n10547_;
  assign new_n15302_ = ~new_n10625_ | ~new_n10440_;
  assign new_n15303_ = ~new_n15193_ | ~new_n10535_;
  assign new_n15304_ = ~new_n10625_ | ~new_n10388_;
  assign new_n15305_ = ~new_n15193_ | ~new_n10489_;
  assign new_n15306_ = ~new_n10625_ | ~new_n10375_;
  assign new_n15307_ = ~new_n15193_ | ~new_n10479_;
  assign new_n15308_ = ~new_n10625_ | ~new_n10416_;
  assign new_n15309_ = ~new_n15193_ | ~new_n10513_;
  assign new_n15310_ = ~new_n10625_ | ~new_n10405_;
  assign new_n15311_ = ~new_n15193_ | ~new_n10502_;
  assign new_n15312_ = ~new_n10625_ | ~new_n10464_;
  assign new_n15313_ = ~new_n15193_ | ~new_n10559_;
  assign new_n15314_ = ~new_n10625_ | ~new_n10430_;
  assign new_n15315_ = ~new_n15193_ | ~new_n10525_;
  assign new_n15316_ = ~new_n10625_ | ~new_n10453_;
  assign new_n15317_ = ~new_n15193_ | ~new_n10548_;
  assign new_n15318_ = ~new_n10625_ | ~new_n10441_;
  assign new_n15319_ = ~new_n15193_ | ~new_n10536_;
  assign new_n15320_ = ~new_n10625_ | ~new_n10389_;
  assign new_n15321_ = ~new_n15193_ | ~new_n10490_;
  assign new_n15322_ = ~pi0758 | ~new_n10560_;
  assign new_n15323_ = ~pi0994 | ~new_n10639_ | ~new_n10638_;
  assign new_n15324_ = ~pi0759 | ~new_n10560_;
  assign new_n15325_ = ~pi0994 | ~new_n10638_ | ~new_n15131_;
  assign new_n15326_ = ~pi0760 | ~new_n10560_;
  assign new_n15327_ = ~new_n15128_ | ~pi0994;
  assign new_n15328_ = ~new_n10657_ | ~new_n11447_;
  assign new_n15329_ = ~new_n12622_ | ~pi0756;
  assign new_n15330_ = ~new_n12622_ | ~pi0757;
  assign new_n15331_ = ~new_n12652_ | ~new_n11447_;
  assign new_n15332_ = ~new_n12622_ | ~pi0758;
  assign new_n15333_ = ~new_n12660_ | ~new_n11447_;
  assign new_n15334_ = ~new_n12622_ | ~pi0759;
  assign new_n15335_ = ~new_n12670_ | ~new_n11447_;
  assign new_n15336_ = ~new_n12622_ | ~pi0760;
  assign new_n15337_ = ~new_n12678_ | ~new_n11447_;
  assign new_n15338_ = ~new_n10283_ | ~new_n14914_;
  assign new_n15339_ = ~new_n9657_ | ~new_n14224_;
  assign new_n15340_ = ~new_n14258_ | ~new_n14914_;
  assign new_n15341_ = ~new_n9657_ | ~new_n14241_;
  assign new_n15342_ = ~new_n14292_ | ~new_n14914_;
  assign new_n15343_ = ~new_n9657_ | ~new_n14275_;
  assign new_n15344_ = ~new_n14326_ | ~new_n14914_;
  assign new_n15345_ = ~new_n9657_ | ~new_n14309_;
  assign new_n15346_ = ~new_n14360_ | ~new_n14914_;
  assign new_n15347_ = ~new_n9657_ | ~new_n14343_;
  assign new_n15348_ = ~new_n14394_ | ~new_n14914_;
  assign new_n15349_ = ~new_n9657_ | ~new_n14377_;
  assign new_n15350_ = ~new_n14428_ | ~new_n14914_;
  assign new_n15351_ = ~new_n9657_ | ~new_n14411_;
  assign new_n15352_ = ~new_n14462_ | ~new_n14914_;
  assign new_n15353_ = ~new_n9657_ | ~new_n14445_;
  assign new_n15354_ = ~new_n29429_ | ~new_n10613_;
  assign new_n15355_ = ~new_n10283_ | ~new_n30562_;
  assign new_n15356_ = ~new_n29441_ | ~new_n10613_;
  assign new_n15357_ = ~new_n10283_ | ~new_n30525_;
  assign new_n15358_ = ~new_n29442_ | ~new_n10613_;
  assign new_n15359_ = ~new_n10283_ | ~new_n30564_;
  assign new_n15360_ = ~new_n29443_ | ~new_n10613_;
  assign new_n15361_ = ~new_n10283_ | ~new_n30524_;
  assign new_n15362_ = ~new_n29444_ | ~new_n10613_;
  assign new_n15363_ = ~new_n10283_ | ~new_n30566_;
  assign new_n15364_ = ~new_n29450_ | ~new_n10613_;
  assign new_n15365_ = ~new_n10283_ | ~new_n30523_;
  assign new_n15366_ = ~new_n29446_ | ~new_n10613_;
  assign new_n15367_ = ~new_n10283_ | ~new_n30571_;
  assign new_n15368_ = ~new_n29428_ | ~new_n10613_;
  assign new_n15369_ = ~new_n10283_ | ~new_n30549_;
  assign new_n15370_ = ~new_n29445_ | ~new_n10613_;
  assign new_n15371_ = ~new_n10283_ | ~new_n30527_;
  assign new_n15372_ = ~new_n29037_ | ~new_n9658_;
  assign new_n15373_ = ~pi0932 | ~new_n14910_;
  assign new_n15374_ = ~new_n29038_ | ~new_n9658_;
  assign new_n15375_ = ~pi0931 | ~new_n14910_;
  assign new_n15376_ = ~new_n29039_ | ~new_n9658_;
  assign new_n15377_ = ~pi0930 | ~new_n14910_;
  assign new_n15378_ = ~new_n29040_ | ~new_n9658_;
  assign new_n15379_ = ~pi0929 | ~new_n14910_;
  assign new_n15380_ = ~new_n29041_ | ~new_n9658_;
  assign new_n15381_ = ~pi0928 | ~new_n14910_;
  assign new_n15382_ = ~new_n29042_ | ~new_n9658_;
  assign new_n15383_ = ~pi0927 | ~new_n14910_;
  assign new_n15384_ = ~new_n29043_ | ~new_n9658_;
  assign new_n15385_ = ~pi0926 | ~new_n14910_;
  assign new_n15386_ = ~new_n29021_ | ~new_n9658_;
  assign new_n15387_ = ~pi0925 | ~new_n14910_;
  assign new_n15388_ = ~new_n10296_ | ~new_n14781_;
  assign new_n15389_ = ~new_n14908_ | ~new_n10566_;
  assign new_n15390_ = ~new_n28887_ | ~new_n10325_;
  assign new_n15391_ = ~pi0797 | ~pi0627;
  assign new_n15392_ = ~new_n29495_ | ~new_n10324_;
  assign new_n15393_ = ~new_n30269_ | ~new_n11458_;
  assign new_n15394_ = ~new_n29508_ | ~new_n10324_;
  assign new_n15395_ = ~new_n30280_ | ~new_n11458_;
  assign new_n15396_ = ~new_n29509_ | ~new_n10324_;
  assign new_n15397_ = ~new_n30281_ | ~new_n11458_;
  assign new_n15398_ = ~new_n29510_ | ~new_n10324_;
  assign new_n15399_ = ~new_n30282_ | ~new_n11458_;
  assign new_n15400_ = ~new_n29511_ | ~new_n10324_;
  assign new_n15401_ = ~new_n30283_ | ~new_n11458_;
  assign new_n15402_ = ~new_n28880_ | ~new_n10325_;
  assign new_n15403_ = ~pi0775 | ~pi0627;
  assign new_n15404_ = ~new_n28881_ | ~new_n10325_;
  assign new_n15405_ = ~pi0774 | ~pi0627;
  assign new_n15406_ = ~new_n28882_ | ~new_n10325_;
  assign new_n15407_ = ~pi0773 | ~pi0627;
  assign new_n15408_ = ~new_n28883_ | ~new_n10325_;
  assign new_n15409_ = ~pi0772 | ~pi0627;
  assign new_n15410_ = ~new_n28884_ | ~new_n10325_;
  assign new_n15411_ = ~pi0771 | ~pi0627;
  assign new_n15412_ = ~new_n28885_ | ~new_n10325_;
  assign new_n15413_ = ~pi0770 | ~pi0627;
  assign new_n15414_ = ~new_n28888_ | ~new_n10325_;
  assign new_n15415_ = ~pi0796 | ~pi0627;
  assign new_n15416_ = ~new_n28886_ | ~new_n10325_;
  assign new_n15417_ = ~pi0769 | ~pi0627;
  assign new_n15418_ = ~new_n28890_ | ~new_n10325_;
  assign new_n15419_ = ~pi0795 | ~pi0627;
  assign new_n15420_ = ~new_n28891_ | ~new_n10325_;
  assign new_n15421_ = ~pi0794 | ~pi0627;
  assign new_n15422_ = ~new_n28892_ | ~new_n10325_;
  assign new_n15423_ = ~pi0793 | ~pi0627;
  assign new_n15424_ = ~new_n28893_ | ~new_n10325_;
  assign new_n15425_ = ~pi0792 | ~pi0627;
  assign new_n15426_ = ~new_n28894_ | ~new_n10325_;
  assign new_n15427_ = ~pi0791 | ~pi0627;
  assign new_n15428_ = ~new_n28895_ | ~new_n10325_;
  assign new_n15429_ = ~pi0790 | ~pi0627;
  assign new_n15430_ = ~new_n28896_ | ~new_n10325_;
  assign new_n15431_ = ~pi0789 | ~pi0627;
  assign new_n15432_ = ~new_n28897_ | ~new_n10325_;
  assign new_n15433_ = ~pi0788 | ~pi0627;
  assign new_n15434_ = ~new_n28898_ | ~new_n10325_;
  assign new_n15435_ = ~pi0787 | ~pi0627;
  assign new_n15436_ = ~new_n28899_ | ~new_n10325_;
  assign new_n15437_ = ~pi0786 | ~pi0627;
  assign new_n15438_ = ~new_n28889_ | ~new_n10325_;
  assign new_n15439_ = ~pi0768 | ~pi0627;
  assign new_n15440_ = ~new_n28900_ | ~new_n10325_;
  assign new_n15441_ = ~pi0785 | ~pi0627;
  assign new_n15442_ = ~new_n28901_ | ~new_n10325_;
  assign new_n15443_ = ~pi0784 | ~pi0627;
  assign new_n15444_ = ~new_n28902_ | ~new_n10325_;
  assign new_n15445_ = ~pi0783 | ~pi0627;
  assign new_n15446_ = ~new_n28903_ | ~new_n10325_;
  assign new_n15447_ = ~pi0782 | ~pi0627;
  assign new_n15448_ = ~new_n28904_ | ~new_n10325_;
  assign new_n15449_ = ~pi0781 | ~pi0627;
  assign new_n15450_ = ~new_n28905_ | ~new_n10325_;
  assign new_n15451_ = ~pi0780 | ~pi0627;
  assign new_n15452_ = ~new_n28906_ | ~new_n10325_;
  assign new_n15453_ = ~pi0779 | ~pi0627;
  assign new_n15454_ = ~new_n28907_ | ~new_n10325_;
  assign new_n15455_ = ~pi0778 | ~pi0627;
  assign new_n15456_ = ~new_n28908_ | ~new_n10325_;
  assign new_n15457_ = ~pi0777 | ~pi0627;
  assign new_n15458_ = ~new_n28909_ | ~new_n10325_;
  assign new_n15459_ = ~pi0776 | ~pi0627;
  assign new_n15460_ = ~new_n28823_ | ~new_n10325_;
  assign new_n15461_ = ~pi0767 | ~pi0627;
  assign new_n15462_ = ~pi0798 | ~new_n10325_;
  assign new_n15463_ = ~pi0766 | ~pi0627;
  assign new_n15464_ = ~new_n29495_ | ~new_n10310_;
  assign new_n15465_ = ~new_n9656_ | ~pi0626;
  assign new_n15466_ = ~new_n29508_ | ~new_n10310_;
  assign new_n15467_ = ~new_n9656_ | ~pi0626;
  assign new_n15468_ = ~new_n29509_ | ~new_n10310_;
  assign new_n15469_ = ~new_n29138_ | ~pi0626;
  assign new_n15470_ = ~new_n29510_ | ~new_n10310_;
  assign new_n15471_ = ~new_n29139_ | ~pi0626;
  assign new_n15472_ = ~new_n29511_ | ~new_n10310_;
  assign new_n15473_ = ~new_n29136_ | ~pi0626;
  assign new_n15474_ = ~new_n29496_ | ~new_n10310_;
  assign new_n15475_ = ~new_n29137_ | ~pi0626;
  assign new_n15476_ = ~pi1218 | ~new_n20995_;
  assign new_n15477_ = ~new_n15521_ | ~new_n20997_;
  assign new_n15478_ = ~pi1246 | ~new_n20996_;
  assign new_n15479_ = ~new_n20985_ | ~new_n33677_;
  assign new_n15480_ = ~pi1225 | ~new_n33676_;
  assign new_n15481_ = ~new_n20976_ | ~new_n33695_;
  assign new_n15482_ = ~pi1234 | ~new_n33694_;
  assign new_n15483_ = ~new_n15530_ | ~new_n33703_;
  assign new_n15484_ = ~pi1238 | ~new_n33702_;
  assign new_n15485_ = ~new_n20987_ | ~new_n33673_;
  assign new_n15486_ = ~pi1223 | ~new_n33672_;
  assign new_n15487_ = ~new_n20990_ | ~new_n33667_;
  assign new_n15488_ = ~pi1220 | ~new_n33666_;
  assign new_n15489_ = ~new_n20981_ | ~new_n33685_;
  assign new_n15490_ = ~pi1229 | ~new_n33684_;
  assign new_n15491_ = ~new_n15526_ | ~new_n33711_;
  assign new_n15492_ = ~pi1242 | ~new_n33710_;
  assign new_n15493_ = ~new_n20991_ | ~new_n33665_;
  assign new_n15494_ = ~pi1219 | ~new_n33664_;
  assign new_n15495_ = ~new_n20980_ | ~new_n33687_;
  assign new_n15496_ = ~pi1230 | ~new_n33686_;
  assign new_n15497_ = ~new_n15527_ | ~new_n33709_;
  assign new_n15498_ = ~pi1241 | ~new_n33708_;
  assign new_n15499_ = ~new_n20984_ | ~new_n33679_;
  assign new_n15500_ = ~pi1226 | ~new_n33678_;
  assign new_n15501_ = ~new_n20977_ | ~new_n33693_;
  assign new_n15502_ = ~pi1233 | ~new_n33692_;
  assign new_n15503_ = ~new_n15531_ | ~new_n33701_;
  assign new_n15504_ = ~pi1237 | ~new_n33700_;
  assign new_n15505_ = ~new_n20986_ | ~new_n33675_;
  assign new_n15506_ = ~pi1224 | ~new_n33674_;
  assign new_n15507_ = ~new_n20982_ | ~new_n33683_;
  assign new_n15508_ = ~pi1228 | ~new_n33682_;
  assign new_n15509_ = ~new_n15800_ | ~new_n33697_;
  assign new_n15510_ = ~pi1235 | ~new_n33696_;
  assign new_n15511_ = ~new_n20978_ | ~new_n33691_;
  assign new_n15512_ = ~pi1232 | ~new_n33690_;
  assign new_n15513_ = ~new_n15529_ | ~new_n33705_;
  assign new_n15514_ = ~pi1239 | ~new_n33704_;
  assign new_n15515_ = ~new_n15524_ | ~new_n33715_;
  assign new_n15516_ = ~pi1244 | ~new_n33714_;
  assign new_n15517_ = ~new_n15523_ | ~new_n33716_;
  assign new_n15518_ = ~pi1245 | ~new_n33717_;
  assign new_n15519_ = ~new_n20989_ | ~new_n33668_;
  assign new_n15520_ = ~pi1221 | ~new_n33669_;
  assign new_n15521_ = ~new_n20996_;
  assign new_n15522_ = ~pi1217 | ~pi1216 | ~pi1215;
  assign new_n15523_ = ~new_n33717_;
  assign new_n15524_ = ~new_n33714_;
  assign new_n15525_ = ~new_n33712_;
  assign new_n15526_ = ~new_n33710_;
  assign new_n15527_ = ~new_n33708_;
  assign new_n15528_ = ~new_n33706_;
  assign new_n15529_ = ~new_n33704_;
  assign new_n15530_ = ~new_n33702_;
  assign new_n15531_ = ~new_n33700_;
  assign new_n15532_ = ~new_n33698_;
  assign new_n15533_ = ~pi1445 & ~pi1074;
  assign new_n15534_ = new_n17412_ & pi1074;
  assign new_n15535_ = new_n17446_ & new_n17658_;
  assign new_n15536_ = new_n16415_ & new_n15631_;
  assign new_n15537_ = new_n33497_ & new_n17373_;
  assign new_n15538_ = new_n33065_ & new_n19140_ & new_n17046_;
  assign new_n15539_ = new_n15569_ & new_n17405_;
  assign new_n15540_ = pi1074 & new_n16612_;
  assign new_n15541_ = pi1074 & new_n16595_;
  assign new_n15542_ = new_n17405_ & pi1073;
  assign new_n15543_ = new_n15540_ & new_n17389_;
  assign new_n15544_ = new_n15540_ & new_n17391_;
  assign new_n15545_ = new_n17045_ & new_n16597_;
  assign new_n15546_ = new_n17442_ & new_n16597_;
  assign new_n15547_ = new_n16611_ & new_n16612_ & pi1075;
  assign new_n15548_ = new_n33164_ & pi1075 & new_n16612_;
  assign new_n15549_ = new_n17416_ & pi1076;
  assign new_n15550_ = new_n15543_ & new_n17678_;
  assign new_n15551_ = new_n16595_ & new_n16444_;
  assign new_n15552_ = new_n17403_ & new_n17630_;
  assign new_n15553_ = pi1076 & new_n16597_;
  assign new_n15554_ = pi1073 & new_n16612_;
  assign new_n15555_ = new_n15541_ & new_n17395_;
  assign new_n15556_ = new_n15541_ & new_n17397_;
  assign new_n15557_ = new_n18979_ & new_n16597_;
  assign new_n15558_ = new_n16943_ & new_n16595_;
  assign new_n15559_ = new_n15541_ & new_n18750_;
  assign new_n15560_ = new_n15544_ & new_n16461_;
  assign new_n15561_ = new_n15541_ & new_n20789_;
  assign new_n15562_ = new_n15538_ & new_n16452_;
  assign new_n15563_ = new_n15538_ & new_n17658_;
  assign new_n15564_ = new_n17403_ & new_n16572_;
  assign new_n15565_ = pi1076 & new_n16598_;
  assign new_n15566_ = new_n16598_ & new_n16475_;
  assign new_n15567_ = new_n17404_ & new_n16604_;
  assign new_n15568_ = new_n17065_ & new_n17404_;
  assign new_n15569_ = pi1445 & new_n17390_;
  assign new_n15570_ = new_n15633_ & new_n20675_;
  assign new_n15571_ = new_n3108_ & new_n17405_;
  assign new_n15572_ = new_n3097_ & new_n17405_;
  assign new_n15573_ = new_n3086_ & new_n17405_;
  assign new_n15574_ = new_n3083_ & new_n17405_;
  assign new_n15575_ = new_n3082_ & new_n17405_;
  assign new_n15576_ = new_n3081_ & new_n17405_;
  assign new_n15577_ = new_n3080_ & new_n17405_;
  assign new_n15578_ = new_n3079_ & new_n17405_;
  assign new_n15579_ = new_n3092_ & new_n15539_;
  assign new_n15580_ = new_n3101_ & new_n15539_;
  assign new_n15581_ = new_n3091_ & new_n15539_;
  assign new_n15582_ = new_n3100_ & new_n15539_;
  assign new_n15583_ = new_n3090_ & new_n15539_;
  assign new_n15584_ = new_n3099_ & new_n15539_;
  assign new_n15585_ = new_n3089_ & new_n15539_;
  assign new_n15586_ = new_n3098_ & new_n15539_;
  assign new_n15587_ = new_n3088_ & new_n15539_;
  assign new_n15588_ = new_n3096_ & new_n15539_;
  assign new_n15589_ = new_n3087_ & new_n15539_;
  assign new_n15590_ = new_n3095_ & new_n15539_;
  assign new_n15591_ = new_n3085_ & new_n15539_;
  assign new_n15592_ = new_n3094_ & new_n15539_;
  assign new_n15593_ = new_n3084_ & new_n15539_;
  assign new_n15594_ = new_n3093_ & new_n15539_;
  assign new_n15595_ = new_n15542_ & new_n16452_;
  assign new_n15596_ = new_n15542_ & new_n16572_;
  assign new_n15597_ = new_n15542_ & new_n16458_;
  assign new_n15598_ = new_n15542_ & new_n16465_;
  assign new_n15599_ = new_n15542_ & new_n16464_;
  assign new_n15600_ = new_n15542_ & new_n16459_;
  assign new_n15601_ = new_n15542_ & new_n17354_;
  assign new_n15602_ = new_n15542_ & new_n17352_;
  assign new_n15603_ = new_n17404_ & new_n18642_;
  assign new_n15604_ = new_n17404_ & new_n17412_;
  assign new_n15605_ = new_n15565_ & new_n16465_;
  assign new_n15606_ = new_n15549_ & new_n15629_;
  assign new_n15607_ = new_n17070_ & new_n16612_;
  assign new_n15608_ = ~pi1075 & ~pi1073;
  assign new_n15609_ = pi1074 & pi1075;
  assign new_n15610_ = new_n19547_ & new_n16612_;
  assign new_n15611_ = pi1075 & new_n16568_;
  assign new_n15612_ = new_n17380_ & new_n20675_;
  assign new_n15613_ = new_n16636_ & new_n16541_;
  assign new_n15614_ = new_n17721_ & new_n16636_;
  assign new_n15615_ = new_n20877_ & new_n16541_;
  assign new_n15616_ = new_n17721_ & new_n20877_;
  assign new_n15617_ = new_n16416_ & new_n16482_;
  assign new_n15618_ = new_n17724_ & new_n16482_;
  assign new_n15619_ = new_n31187_ & new_n31170_;
  assign new_n15620_ = new_n31187_ & new_n16497_;
  assign new_n15621_ = new_n31170_ & new_n16498_;
  assign new_n15622_ = ~new_n31187_ & ~new_n31170_;
  assign new_n15623_ = new_n31178_ & new_n31179_;
  assign new_n15624_ = new_n31178_ & new_n16499_;
  assign new_n15625_ = new_n31179_ & new_n16500_;
  assign new_n15626_ = ~new_n31178_ & ~new_n31179_;
  assign new_n15627_ = pi1075 & new_n16652_;
  assign new_n15628_ = new_n16758_ & new_n15633_;
  assign new_n15629_ = new_n33065_ & new_n16465_;
  assign new_n15630_ = new_n17675_ & new_n16452_;
  assign new_n15631_ = pi1076 & new_n17581_;
  assign new_n15632_ = new_n17432_ & pi1076;
  assign new_n15633_ = new_n16458_ & new_n17354_ & new_n16572_ & new_n17581_;
  assign new_n15634_ = pi1209 & pi1207 & pi1208 & pi1206;
  assign new_n15635_ = pi1208 & new_n16447_;
  assign new_n15636_ = pi1208 & new_n16447_ & pi1207 & pi1206;
  assign new_n15637_ = pi1209 & new_n16446_;
  assign new_n15638_ = pi1209 & new_n16446_ & pi1207 & pi1206;
  assign new_n15639_ = new_n16688_ & new_n17559_;
  assign new_n15640_ = pi1209 & new_n16445_ & pi1208 & pi1206;
  assign new_n15641_ = pi1208 & new_n16445_ & new_n16447_;
  assign new_n15642_ = new_n16687_ & new_n16686_;
  assign new_n15643_ = pi1209 & new_n16445_ & new_n16446_;
  assign new_n15644_ = new_n16685_ & new_n16684_;
  assign new_n15645_ = pi1206 & new_n17561_;
  assign new_n15646_ = new_n16683_ & new_n16682_;
  assign new_n15647_ = new_n16681_ & new_n16680_;
  assign new_n15648_ = new_n17559_ & pi1207 & new_n16451_;
  assign new_n15649_ = new_n16679_ & new_n16678_;
  assign new_n15650_ = ~pi1206 & ~pi1207;
  assign new_n15651_ = new_n15650_ & pi1208 & new_n16447_;
  assign new_n15652_ = new_n15650_ & pi1209 & new_n16446_;
  assign new_n15653_ = new_n17561_ & new_n16451_;
  assign new_n15654_ = new_n16587_ & new_n20861_ & new_n20860_;
  assign new_n15655_ = new_n31276_ & new_n16493_;
  assign new_n15656_ = new_n16635_ & new_n16539_;
  assign new_n15657_ = new_n31235_ & new_n31276_;
  assign new_n15658_ = new_n17709_ & new_n15657_;
  assign new_n15659_ = pi1212 & pi1211;
  assign new_n15660_ = pi1212 & new_n16484_;
  assign new_n15661_ = new_n16496_ & new_n17729_;
  assign new_n15662_ = new_n17705_ & new_n15657_;
  assign new_n15663_ = new_n16508_ & new_n17787_;
  assign new_n15664_ = new_n17706_ & new_n15657_;
  assign new_n15665_ = new_n16515_ & new_n17846_;
  assign new_n15666_ = new_n17707_ & new_n31270_;
  assign new_n15667_ = ~new_n31270_ & ~new_n31277_;
  assign new_n15668_ = new_n15667_ & new_n15657_;
  assign new_n15669_ = ~pi1214 & ~pi1213;
  assign new_n15670_ = new_n16519_ & new_n17903_;
  assign new_n15671_ = new_n20874_ & new_n16539_;
  assign new_n15672_ = new_n17710_ & new_n17709_;
  assign new_n15673_ = new_n16524_ & new_n17961_;
  assign new_n15674_ = new_n17710_ & new_n17705_;
  assign new_n15675_ = new_n16528_ & new_n18018_;
  assign new_n15676_ = new_n17710_ & new_n17706_;
  assign new_n15677_ = new_n16531_ & new_n18076_;
  assign new_n15678_ = new_n17710_ & new_n15667_;
  assign new_n15679_ = new_n16535_ & new_n18133_;
  assign new_n15680_ = new_n17712_ & new_n16635_;
  assign new_n15681_ = new_n16540_ & new_n16538_;
  assign new_n15682_ = new_n17705_ & new_n15655_;
  assign new_n15683_ = new_n16545_ & new_n18246_;
  assign new_n15684_ = new_n17706_ & new_n15655_;
  assign new_n15685_ = new_n16548_ & new_n18304_;
  assign new_n15686_ = new_n15667_ & new_n15655_;
  assign new_n15687_ = new_n16552_ & new_n18361_;
  assign new_n15688_ = new_n17712_ & new_n20874_;
  assign new_n15689_ = ~new_n31276_ & ~new_n31235_;
  assign new_n15690_ = new_n15689_ & new_n17709_;
  assign new_n15691_ = ~pi1211 & ~pi1212;
  assign new_n15692_ = new_n16555_ & new_n18419_;
  assign new_n15693_ = new_n15689_ & new_n17705_;
  assign new_n15694_ = new_n16559_ & new_n18476_;
  assign new_n15695_ = new_n15689_ & new_n17706_;
  assign new_n15696_ = new_n16562_ & new_n18534_;
  assign new_n15697_ = new_n15689_ & new_n15667_;
  assign new_n15698_ = new_n16566_ & new_n18591_;
  assign new_n15699_ = new_n18649_ & new_n20881_ & new_n20880_;
  assign new_n15700_ = new_n16925_ & new_n18680_;
  assign new_n15701_ = new_n17400_ & new_n16627_;
  assign new_n15702_ = pi1209 & new_n16583_;
  assign new_n15703_ = new_n18664_ & new_n18692_;
  assign new_n15704_ = new_n15703_ & new_n15702_;
  assign new_n15705_ = new_n16447_ & new_n16583_;
  assign new_n15706_ = new_n15703_ & new_n15705_;
  assign new_n15707_ = new_n18700_ & pi1209;
  assign new_n15708_ = new_n15703_ & new_n15707_;
  assign new_n15709_ = new_n18700_ & new_n16447_;
  assign new_n15710_ = new_n15703_ & new_n15709_;
  assign new_n15711_ = new_n18664_ & new_n16582_;
  assign new_n15712_ = new_n15711_ & new_n15702_;
  assign new_n15713_ = new_n15711_ & new_n15705_;
  assign new_n15714_ = new_n15711_ & new_n15707_;
  assign new_n15715_ = new_n15711_ & new_n15709_;
  assign new_n15716_ = new_n18692_ & new_n16619_;
  assign new_n15717_ = new_n15716_ & new_n15702_;
  assign new_n15718_ = new_n15716_ & new_n15705_;
  assign new_n15719_ = new_n15716_ & new_n15707_;
  assign new_n15720_ = new_n15716_ & new_n15709_;
  assign new_n15721_ = new_n16619_ & new_n16582_;
  assign new_n15722_ = new_n15702_ & new_n15721_;
  assign new_n15723_ = new_n15705_ & new_n15721_;
  assign new_n15724_ = new_n15707_ & new_n15721_;
  assign new_n15725_ = new_n15709_ & new_n15721_;
  assign new_n15726_ = new_n18661_ & new_n20901_;
  assign new_n15727_ = new_n15726_ & new_n15635_;
  assign new_n15728_ = new_n15726_ & new_n16679_;
  assign new_n15729_ = new_n15726_ & new_n17559_;
  assign new_n15730_ = new_n15726_ & new_n15637_;
  assign new_n15731_ = new_n18661_ & new_n16637_;
  assign new_n15732_ = new_n15731_ & new_n15635_;
  assign new_n15733_ = new_n15731_ & new_n16679_;
  assign new_n15734_ = new_n15731_ & new_n17559_;
  assign new_n15735_ = new_n15731_ & new_n15637_;
  assign new_n15736_ = new_n20901_ & new_n16623_;
  assign new_n15737_ = new_n15736_ & new_n15635_;
  assign new_n15738_ = new_n15736_ & new_n16679_;
  assign new_n15739_ = new_n15736_ & new_n17559_;
  assign new_n15740_ = new_n15736_ & new_n15637_;
  assign new_n15741_ = new_n16637_ & new_n16623_;
  assign new_n15742_ = new_n15741_ & new_n15635_;
  assign new_n15743_ = new_n15741_ & new_n16679_;
  assign new_n15744_ = new_n15741_ & new_n17559_;
  assign new_n15745_ = new_n15741_ & new_n15637_;
  assign new_n15746_ = new_n20246_ & new_n17560_;
  assign new_n15747_ = new_n20246_ & new_n15641_;
  assign new_n15748_ = new_n20246_ & new_n15643_;
  assign new_n15749_ = new_n20246_ & new_n17561_;
  assign new_n15750_ = new_n20246_ & pi1207;
  assign new_n15751_ = new_n15750_ & new_n16679_;
  assign new_n15752_ = new_n15750_ & new_n15635_;
  assign new_n15753_ = new_n15750_ & new_n15637_;
  assign new_n15754_ = new_n15750_ & new_n17559_;
  assign new_n15755_ = new_n17560_ & new_n16626_;
  assign new_n15756_ = new_n15641_ & new_n16626_;
  assign new_n15757_ = new_n15643_ & new_n16626_;
  assign new_n15758_ = new_n17561_ & new_n16626_;
  assign new_n15759_ = pi1207 & new_n16626_;
  assign new_n15760_ = new_n15759_ & new_n16679_;
  assign new_n15761_ = new_n15759_ & new_n15635_;
  assign new_n15762_ = new_n15759_ & new_n15637_;
  assign new_n15763_ = new_n15759_ & new_n17559_;
  assign new_n15764_ = new_n20971_ & new_n17365_;
  assign new_n15765_ = new_n15764_ & new_n15705_;
  assign new_n15766_ = new_n15764_ & new_n15702_;
  assign new_n15767_ = new_n15764_ & new_n15709_;
  assign new_n15768_ = new_n15764_ & new_n15707_;
  assign new_n15769_ = new_n20971_ & new_n16633_;
  assign new_n15770_ = new_n15769_ & new_n15705_;
  assign new_n15771_ = new_n15769_ & new_n15702_;
  assign new_n15772_ = new_n15769_ & new_n15709_;
  assign new_n15773_ = new_n15769_ & new_n15707_;
  assign new_n15774_ = new_n17365_ & new_n16638_;
  assign new_n15775_ = new_n15774_ & new_n15705_;
  assign new_n15776_ = new_n15774_ & new_n15702_;
  assign new_n15777_ = new_n15774_ & new_n15709_;
  assign new_n15778_ = new_n15774_ & new_n15707_;
  assign new_n15779_ = new_n16638_ & new_n16633_;
  assign new_n15780_ = new_n15779_ & new_n15705_;
  assign new_n15781_ = new_n15779_ & new_n15702_;
  assign new_n15782_ = new_n15779_ & new_n15709_;
  assign new_n15783_ = new_n15779_ & new_n15707_;
  assign new_n15784_ = pi1076 & new_n16570_;
  assign new_n15785_ = pi1405 & new_n15560_;
  assign new_n15786_ = new_n16714_ & new_n16711_ & new_n16712_ & new_n16713_ & new_n15788_;
  assign new_n15787_ = new_n20685_ & new_n16608_;
  assign new_n15788_ = new_n20853_ & new_n20852_;
  assign new_n15789_ = new_n20968_ & new_n20967_;
  assign new_n15790_ = ~new_n20036_ | ~new_n20034_ | ~new_n20035_;
  assign new_n15791_ = ~new_n20037_ | ~new_n17207_;
  assign new_n15792_ = ~new_n20024_ | ~new_n20022_ | ~new_n20023_;
  assign new_n15793_ = ~new_n20027_ | ~new_n20025_ | ~new_n20026_;
  assign new_n15794_ = ~new_n20030_ | ~new_n20028_ | ~new_n20029_;
  assign new_n15795_ = ~new_n19937_ | ~new_n17186_;
  assign new_n15796_ = ~new_n19934_ | ~new_n17185_;
  assign new_n15797_ = ~new_n20033_ | ~new_n20031_ | ~new_n20032_;
  assign new_n15798_ = ~new_n19931_ | ~new_n17184_;
  assign new_n15799_ = ~new_n19928_ | ~new_n17183_;
  assign new_n15800_ = ~new_n33696_;
  assign new_n15801_ = new_n31372_ & new_n19927_;
  assign new_n15802_ = new_n31372_ & new_n19927_;
  assign new_n15803_ = new_n31372_ & new_n19927_;
  assign new_n15804_ = new_n31372_ & new_n19927_;
  assign new_n15805_ = new_n31372_ & new_n19927_;
  assign new_n15806_ = new_n31372_ & new_n19927_;
  assign new_n15807_ = new_n31372_ & new_n19927_;
  assign new_n15808_ = new_n31372_ & new_n19927_;
  assign new_n15809_ = new_n31372_ & new_n19927_;
  assign new_n15810_ = new_n31372_ & new_n19927_;
  assign new_n15811_ = new_n31372_ & new_n19927_;
  assign new_n15812_ = new_n31372_ & new_n19927_;
  assign new_n15813_ = new_n31372_ & new_n19927_;
  assign new_n15814_ = new_n31372_ & new_n19927_;
  assign new_n15815_ = new_n31238_ & new_n19927_;
  assign new_n15816_ = new_n31264_ & new_n19927_;
  assign new_n15817_ = new_n31265_ & new_n19927_;
  assign new_n15818_ = new_n31266_ & new_n19927_;
  assign new_n15819_ = new_n31267_ & new_n19927_;
  assign new_n15820_ = new_n31268_ & new_n19927_;
  assign new_n15821_ = new_n31269_ & new_n19927_;
  assign new_n15822_ = new_n31257_ & new_n19927_;
  assign new_n15823_ = new_n31307_ & new_n19927_;
  assign new_n15824_ = new_n31237_ & new_n19927_;
  assign new_n15825_ = new_n31236_ & new_n19927_;
  assign new_n15826_ = new_n31272_ & new_n19927_;
  assign new_n15827_ = new_n31274_ & new_n19927_;
  assign new_n15828_ = new_n31235_ & new_n19927_;
  assign new_n15829_ = ~new_n16621_ | ~new_n20050_;
  assign new_n15830_ = new_n31277_ & new_n19927_;
  assign new_n15831_ = pi1074 & new_n20051_;
  assign new_n15832_ = ~new_n19951_ | ~new_n19950_ | ~new_n19949_;
  assign new_n15833_ = ~new_n19952_ | ~new_n17190_;
  assign new_n15834_ = ~new_n19961_ | ~new_n17192_;
  assign new_n15835_ = ~new_n19965_ | ~new_n17193_;
  assign new_n15836_ = ~new_n19969_ | ~new_n17194_;
  assign new_n15837_ = ~new_n19973_ | ~new_n17195_;
  assign new_n15838_ = ~new_n19977_ | ~new_n17196_;
  assign new_n15839_ = ~new_n19981_ | ~new_n17197_;
  assign new_n15840_ = ~new_n19985_ | ~new_n17198_;
  assign new_n15841_ = ~new_n19989_ | ~new_n17199_;
  assign new_n15842_ = ~new_n19993_ | ~new_n17200_;
  assign new_n15843_ = ~new_n19997_ | ~new_n17201_;
  assign new_n15844_ = ~new_n20006_ | ~new_n17203_;
  assign new_n15845_ = ~new_n20010_ | ~new_n17204_;
  assign new_n15846_ = ~new_n20014_ | ~new_n17205_;
  assign new_n15847_ = ~new_n20018_ | ~new_n17206_;
  assign new_n15848_ = ~new_n19940_ | ~new_n17187_;
  assign new_n15849_ = ~new_n19947_ | ~new_n19944_ | ~new_n17189_ | ~new_n19948_;
  assign new_n15850_ = ~new_n19959_ | ~new_n19956_ | ~new_n17191_ | ~new_n19960_;
  assign new_n15851_ = ~new_n20004_ | ~new_n20001_ | ~new_n17202_ | ~new_n20005_;
  assign new_n15852_ = ~new_n20043_ | ~new_n20040_ | ~new_n17208_ | ~new_n20044_;
  assign new_n15853_ = ~new_n20047_ | ~new_n20048_ | ~new_n20049_ | ~new_n20046_ | ~new_n20045_;
  assign new_n15854_ = ~new_n20639_ | ~new_n20638_;
  assign new_n15855_ = ~new_n20641_ | ~new_n20640_;
  assign new_n15856_ = ~new_n17349_ | ~new_n20644_;
  assign new_n15857_ = ~new_n17350_ | ~new_n20647_;
  assign new_n15858_ = ~new_n20648_ | ~new_n20975_ | ~new_n20974_;
  assign new_n15859_ = ~new_n20637_ | ~new_n16465_;
  assign new_n15860_ = ~new_n20586_ | ~new_n20585_;
  assign new_n15861_ = ~new_n20588_ | ~new_n20587_;
  assign new_n15862_ = ~new_n20592_ | ~new_n20591_;
  assign new_n15863_ = ~new_n20594_ | ~new_n20593_;
  assign new_n15864_ = ~new_n20596_ | ~new_n20595_;
  assign new_n15865_ = ~new_n20598_ | ~new_n20597_;
  assign new_n15866_ = ~new_n20600_ | ~new_n20599_;
  assign new_n15867_ = ~new_n20602_ | ~new_n20601_;
  assign new_n15868_ = ~new_n20604_ | ~new_n20603_;
  assign new_n15869_ = ~new_n20606_ | ~new_n20605_;
  assign new_n15870_ = ~new_n20608_ | ~new_n20607_;
  assign new_n15871_ = ~new_n20610_ | ~new_n20609_;
  assign new_n15872_ = ~new_n20614_ | ~new_n20613_;
  assign new_n15873_ = ~new_n20616_ | ~new_n20615_;
  assign new_n15874_ = ~new_n20618_ | ~new_n20617_;
  assign new_n15875_ = ~new_n20620_ | ~new_n20619_;
  assign new_n15876_ = ~new_n20622_ | ~new_n20621_;
  assign new_n15877_ = ~new_n20624_ | ~new_n20623_;
  assign new_n15878_ = ~new_n20626_ | ~new_n20625_;
  assign new_n15879_ = ~new_n20628_ | ~new_n20627_;
  assign new_n15880_ = ~new_n20630_ | ~new_n20629_;
  assign new_n15881_ = ~new_n20632_ | ~new_n20631_;
  assign new_n15882_ = ~new_n20574_ | ~new_n20573_;
  assign new_n15883_ = ~new_n20576_ | ~new_n20575_;
  assign new_n15884_ = ~new_n20578_ | ~new_n20577_;
  assign new_n15885_ = ~new_n20580_ | ~new_n20579_;
  assign new_n15886_ = ~new_n20582_ | ~new_n20581_;
  assign new_n15887_ = ~new_n20584_ | ~new_n20583_;
  assign new_n15888_ = ~new_n20590_ | ~new_n20589_;
  assign new_n15889_ = ~new_n20612_ | ~new_n20611_;
  assign new_n15890_ = ~new_n20634_ | ~new_n20633_;
  assign new_n15891_ = ~new_n20636_ | ~new_n20635_;
  assign new_n15892_ = ~new_n20558_ | ~new_n20557_;
  assign new_n15893_ = ~new_n20560_ | ~new_n20559_;
  assign new_n15894_ = ~new_n17346_ | ~new_n17420_;
  assign new_n15895_ = ~new_n20566_ | ~new_n16615_ | ~new_n17347_ | ~new_n20567_;
  assign new_n15896_ = ~new_n17420_ | ~new_n17348_;
  assign new_n15897_ = ~new_n20546_ | ~new_n20545_;
  assign new_n15898_ = ~new_n20548_ | ~new_n20547_;
  assign new_n15899_ = ~new_n17342_ | ~new_n20549_;
  assign new_n15900_ = ~new_n17343_ | ~new_n20551_;
  assign new_n15901_ = ~new_n17344_ | ~new_n20553_;
  assign new_n15902_ = ~new_n17345_ | ~new_n20555_;
  assign new_n15903_ = ~new_n17340_ | ~new_n17373_;
  assign new_n15904_ = new_n20417_ & new_n20264_;
  assign new_n15905_ = new_n20434_ & new_n20264_;
  assign new_n15906_ = new_n20451_ & new_n20264_;
  assign new_n15907_ = new_n20801_ & new_n20264_;
  assign new_n15908_ = new_n20483_ & new_n20264_;
  assign new_n15909_ = new_n20500_ & new_n20264_;
  assign new_n15910_ = new_n20517_ & new_n20264_;
  assign new_n15911_ = new_n20534_ & new_n20264_;
  assign new_n15912_ = ~new_n15787_ | ~new_n20535_;
  assign new_n15913_ = new_n20264_ & new_n20263_;
  assign new_n15914_ = new_n20295_ & new_n20264_;
  assign new_n15915_ = new_n20312_ & new_n20264_;
  assign new_n15916_ = new_n20799_ & new_n20264_;
  assign new_n15917_ = new_n20344_ & new_n20264_;
  assign new_n15918_ = new_n20361_ & new_n20264_;
  assign new_n15919_ = new_n20378_ & new_n20264_;
  assign new_n15920_ = new_n20395_ & new_n20264_;
  assign new_n15921_ = pi1205 & new_n20244_;
  assign new_n15922_ = ~new_n17259_ | ~new_n20277_;
  assign new_n15923_ = new_n20673_ & new_n20672_;
  assign new_n15924_ = new_n20687_ & new_n20651_;
  assign new_n15925_ = new_n20660_ & new_n20659_;
  assign new_n15926_ = ~new_n20229_ | ~new_n20228_;
  assign new_n15927_ = ~new_n20231_ | ~new_n20230_;
  assign new_n15928_ = ~new_n20233_ | ~new_n20232_;
  assign new_n15929_ = ~new_n20797_ | ~new_n20234_;
  assign new_n15930_ = ~new_n20236_ | ~new_n20235_;
  assign new_n15931_ = ~new_n20238_ | ~new_n20237_;
  assign new_n15932_ = ~new_n17242_ | ~new_n20239_;
  assign new_n15933_ = ~new_n20242_ | ~new_n17243_ | ~new_n20241_;
  assign new_n15934_ = new_n20138_ & new_n20090_;
  assign new_n15935_ = new_n20155_ & new_n20090_;
  assign new_n15936_ = new_n20172_ & new_n20090_;
  assign new_n15937_ = new_n20796_ & new_n20090_;
  assign new_n15938_ = new_n20204_ & new_n20090_;
  assign new_n15939_ = new_n20221_ & new_n20090_;
  assign new_n15940_ = new_n20090_ & new_n20089_;
  assign new_n15941_ = new_n20107_ & new_n20090_;
  assign new_n15942_ = ~new_n20109_ | ~new_n20108_;
  assign new_n15943_ = ~new_n20111_ | ~new_n20110_;
  assign new_n15944_ = ~new_n20113_ | ~new_n20112_;
  assign new_n15945_ = ~new_n20115_ | ~new_n20114_;
  assign new_n15946_ = ~new_n20118_ | ~new_n20117_ | ~new_n20116_;
  assign new_n15947_ = ~new_n20121_ | ~new_n20120_ | ~new_n20119_;
  assign new_n15948_ = ~new_n20223_ | ~new_n20224_ | ~new_n20222_;
  assign new_n15949_ = ~new_n20226_ | ~new_n20227_ | ~new_n20225_;
  assign new_n15950_ = new_n31372_ & new_n17340_;
  assign new_n15951_ = new_n17340_ & new_n31372_;
  assign new_n15952_ = new_n17340_ & new_n31372_;
  assign new_n15953_ = new_n17340_ & new_n31372_;
  assign new_n15954_ = new_n17340_ & new_n31372_;
  assign new_n15955_ = new_n17340_ & new_n31372_;
  assign new_n15956_ = new_n17340_ & new_n31372_;
  assign new_n15957_ = new_n17340_ & new_n31372_;
  assign new_n15958_ = new_n17340_ & new_n31372_;
  assign new_n15959_ = new_n17340_ & new_n31372_;
  assign new_n15960_ = new_n17340_ & new_n31372_;
  assign new_n15961_ = new_n17340_ & new_n31372_;
  assign new_n15962_ = new_n17340_ & new_n31372_;
  assign new_n15963_ = new_n17340_ & new_n31372_;
  assign new_n15964_ = new_n17340_ & new_n31372_;
  assign new_n15965_ = new_n17340_ & new_n31238_;
  assign new_n15966_ = new_n17340_ & new_n31264_;
  assign new_n15967_ = new_n17340_ & new_n31265_;
  assign new_n15968_ = new_n17340_ & new_n31266_;
  assign new_n15969_ = new_n17340_ & new_n31267_;
  assign new_n15970_ = new_n17340_ & new_n31268_;
  assign new_n15971_ = new_n17340_ & new_n31269_;
  assign new_n15972_ = new_n17340_ & new_n31257_;
  assign new_n15973_ = ~new_n20053_ | ~new_n20052_;
  assign new_n15974_ = ~new_n20055_ | ~new_n20054_;
  assign new_n15975_ = ~new_n20057_ | ~new_n20056_;
  assign new_n15976_ = ~new_n20059_ | ~new_n20058_;
  assign new_n15977_ = ~new_n20061_ | ~new_n20060_;
  assign new_n15978_ = ~new_n20063_ | ~new_n20062_;
  assign new_n15979_ = ~new_n20064_ | ~new_n20065_ | ~new_n20066_;
  assign new_n15980_ = ~new_n20067_ | ~new_n17209_ | ~new_n20068_;
  assign new_n15981_ = ~new_n20070_ | ~new_n20071_ | ~new_n20072_;
  assign po1511 = ~new_n20679_ | ~new_n19798_ | ~new_n16613_;
  assign po1509 = ~new_n20831_ | ~new_n19794_;
  assign po1508 = ~new_n19793_ | ~new_n19792_;
  assign po1506 = ~new_n17424_ | ~new_n20950_ | ~new_n20949_;
  assign po1504 = ~new_n17424_ | ~new_n20946_ | ~new_n20945_;
  assign po1502 = ~new_n19782_ | ~new_n17429_;
  assign po1499 = ~new_n17421_ | ~new_n20938_ | ~new_n20937_;
  assign po1497 = ~new_n17421_ | ~new_n20928_ | ~new_n20927_;
  assign po1496 = ~new_n19774_ | ~new_n19776_ | ~new_n19772_ | ~new_n17130_ | ~new_n17129_;
  assign po1495 = ~new_n19767_ | ~new_n19769_ | ~new_n19765_ | ~new_n17128_ | ~new_n17127_;
  assign po1494 = ~new_n19760_ | ~new_n19762_ | ~new_n19758_ | ~new_n17126_ | ~new_n17125_;
  assign po1493 = ~new_n19753_ | ~new_n19755_ | ~new_n19751_ | ~new_n17124_ | ~new_n17123_;
  assign po1492 = ~new_n19746_ | ~new_n19748_ | ~new_n19744_ | ~new_n17122_ | ~new_n17121_;
  assign po1491 = ~new_n19739_ | ~new_n19741_ | ~new_n19737_ | ~new_n17120_ | ~new_n17119_;
  assign po1490 = ~new_n19732_ | ~new_n19734_ | ~new_n19730_ | ~new_n17118_ | ~new_n17117_;
  assign po1489 = ~new_n19725_ | ~new_n19727_ | ~new_n19723_ | ~new_n17116_ | ~new_n17115_;
  assign po1488 = ~new_n19718_ | ~new_n19720_ | ~new_n19716_ | ~new_n17114_ | ~new_n17113_;
  assign po1487 = ~new_n19711_ | ~new_n19713_ | ~new_n19709_ | ~new_n17112_ | ~new_n17111_;
  assign po1486 = ~new_n19704_ | ~new_n19706_ | ~new_n19702_ | ~new_n17110_ | ~new_n17109_;
  assign po1485 = ~new_n19697_ | ~new_n19699_ | ~new_n19695_ | ~new_n17108_ | ~new_n17107_;
  assign po1484 = ~new_n17105_ | ~new_n19692_ | ~new_n19688_ | ~new_n17106_ | ~new_n19690_;
  assign po1483 = ~new_n17103_ | ~new_n19685_ | ~new_n19681_ | ~new_n17104_ | ~new_n19683_;
  assign po1482 = ~new_n17101_ | ~new_n19678_ | ~new_n19674_ | ~new_n17102_ | ~new_n19676_;
  assign po1481 = ~new_n19669_ | ~new_n19671_ | ~new_n17099_ | ~new_n17100_ | ~new_n19668_;
  assign po1480 = ~new_n19662_ | ~new_n19664_ | ~new_n17097_ | ~new_n17098_ | ~new_n19661_;
  assign po1479 = ~new_n17096_ | ~new_n19657_ | ~new_n19654_ | ~new_n17095_ | ~new_n19655_;
  assign po1478 = ~new_n17094_ | ~new_n19650_ | ~new_n19647_ | ~new_n17093_ | ~new_n19648_;
  assign po1477 = ~new_n17092_ | ~new_n19643_ | ~new_n19640_ | ~new_n17091_ | ~new_n19641_;
  assign po1476 = ~new_n17090_ | ~new_n19636_ | ~new_n19633_ | ~new_n17089_ | ~new_n19634_;
  assign po1475 = ~new_n17088_ | ~new_n19629_ | ~new_n19626_ | ~new_n17087_ | ~new_n19627_;
  assign po1474 = ~new_n17086_ | ~new_n19622_ | ~new_n19619_ | ~new_n17085_ | ~new_n19620_;
  assign po1473 = ~new_n17084_ | ~new_n19615_ | ~new_n19612_ | ~new_n17083_ | ~new_n19613_;
  assign po1472 = ~new_n17082_ | ~new_n19608_ | ~new_n19605_ | ~new_n17081_ | ~new_n19606_;
  assign po1471 = ~new_n17080_ | ~new_n19601_ | ~new_n19598_ | ~new_n17079_ | ~new_n19599_;
  assign po1470 = ~new_n19590_ | ~new_n17078_ | ~new_n19591_ | ~new_n17077_;
  assign po1469 = ~new_n17075_ | ~new_n19583_ | ~new_n19584_ | ~new_n17076_ | ~new_n19582_;
  assign po1468 = ~new_n19573_ | ~new_n17074_ | ~new_n19575_ | ~new_n19574_;
  assign po1467 = ~new_n19565_ | ~new_n17073_ | ~new_n19567_ | ~new_n19566_;
  assign po1466 = ~new_n19557_ | ~new_n17072_ | ~new_n19559_ | ~new_n19558_;
  assign po1465 = ~new_n19549_ | ~new_n17071_ | ~new_n19551_ | ~new_n19550_;
  assign po1464 = ~new_n19540_ | ~new_n19539_;
  assign po1463 = ~new_n19536_ | ~new_n19537_ | ~new_n19538_;
  assign po1462 = ~new_n19533_ | ~new_n19534_ | ~new_n19535_;
  assign po1461 = ~new_n19530_ | ~new_n19531_ | ~new_n19532_;
  assign po1460 = ~new_n19527_ | ~new_n19528_ | ~new_n19529_;
  assign po1459 = ~new_n19524_ | ~new_n19525_ | ~new_n19526_;
  assign po1458 = ~new_n19521_ | ~new_n19522_ | ~new_n19523_;
  assign po1457 = ~new_n19518_ | ~new_n19519_ | ~new_n19520_;
  assign po1456 = ~new_n19515_ | ~new_n19516_ | ~new_n19517_;
  assign po1455 = ~new_n19512_ | ~new_n19513_ | ~new_n19514_;
  assign po1454 = ~new_n19509_ | ~new_n19510_ | ~new_n19511_;
  assign po1453 = ~new_n19506_ | ~new_n19507_ | ~new_n19508_;
  assign po1452 = ~new_n19503_ | ~new_n19504_ | ~new_n19505_;
  assign po1451 = ~new_n19500_ | ~new_n19501_ | ~new_n19502_;
  assign po1450 = ~new_n19497_ | ~new_n19498_ | ~new_n19499_;
  assign po1449 = ~new_n19494_ | ~new_n19495_ | ~new_n19496_;
  assign po1448 = ~new_n19491_ | ~new_n19492_ | ~new_n19493_;
  assign po1447 = ~new_n19488_ | ~new_n19489_ | ~new_n19490_;
  assign po1446 = ~new_n19485_ | ~new_n19486_ | ~new_n19487_;
  assign po1445 = ~new_n19482_ | ~new_n19483_ | ~new_n19484_;
  assign po1444 = ~new_n19479_ | ~new_n19480_ | ~new_n19481_;
  assign po1443 = ~new_n19476_ | ~new_n19477_ | ~new_n19478_;
  assign po1442 = ~new_n19473_ | ~new_n19474_ | ~new_n19475_;
  assign po1441 = ~new_n19470_ | ~new_n19471_ | ~new_n19472_;
  assign po1440 = ~new_n19467_ | ~new_n19468_ | ~new_n19469_;
  assign po1439 = ~new_n19464_ | ~new_n19465_ | ~new_n19466_;
  assign po1438 = ~new_n19461_ | ~new_n19462_ | ~new_n19463_;
  assign po1437 = ~new_n19458_ | ~new_n19459_ | ~new_n19460_;
  assign po1436 = ~new_n19455_ | ~new_n19456_ | ~new_n19457_;
  assign po1435 = ~new_n19452_ | ~new_n19453_ | ~new_n19454_;
  assign po1434 = ~new_n19449_ | ~new_n19450_ | ~new_n19451_;
  assign po1433 = ~new_n19448_ | ~new_n19447_ | ~new_n19446_;
  assign po1432 = ~new_n17357_ | ~new_n19443_;
  assign po1431 = ~new_n19439_ | ~new_n19441_ | ~new_n19442_ | ~new_n19440_;
  assign po1430 = ~new_n19435_ | ~new_n19437_ | ~new_n19438_ | ~new_n19436_;
  assign po1429 = ~new_n19431_ | ~new_n19433_ | ~new_n19434_ | ~new_n19432_;
  assign po1428 = ~new_n19427_ | ~new_n19429_ | ~new_n19430_ | ~new_n19428_;
  assign po1427 = ~new_n19423_ | ~new_n19425_ | ~new_n19426_ | ~new_n19424_;
  assign po1426 = ~new_n19419_ | ~new_n19421_ | ~new_n19422_ | ~new_n19420_;
  assign po1425 = ~new_n19415_ | ~new_n19417_ | ~new_n19418_ | ~new_n19416_;
  assign po1424 = ~new_n19411_ | ~new_n19413_ | ~new_n19414_ | ~new_n19412_;
  assign po1423 = ~new_n19407_ | ~new_n19409_ | ~new_n19410_ | ~new_n19408_;
  assign po1422 = ~new_n19403_ | ~new_n19405_ | ~new_n19406_ | ~new_n19404_;
  assign po1421 = ~new_n19399_ | ~new_n19401_ | ~new_n19402_ | ~new_n19400_;
  assign po1420 = ~new_n19395_ | ~new_n19397_ | ~new_n19398_ | ~new_n19396_;
  assign po1419 = ~new_n19391_ | ~new_n19393_ | ~new_n19394_ | ~new_n19392_;
  assign po1418 = ~new_n19387_ | ~new_n19389_ | ~new_n19390_ | ~new_n19388_;
  assign po1417 = ~new_n19383_ | ~new_n19385_ | ~new_n19386_ | ~new_n19384_;
  assign po1416 = ~new_n19381_ | ~new_n19382_ | ~new_n19380_;
  assign po1415 = ~new_n19378_ | ~new_n19379_ | ~new_n19377_;
  assign po1414 = ~new_n19375_ | ~new_n19376_ | ~new_n19374_;
  assign po1413 = ~new_n19372_ | ~new_n19373_ | ~new_n19371_;
  assign po1412 = ~new_n19369_ | ~new_n19370_ | ~new_n19368_;
  assign po1411 = ~new_n19366_ | ~new_n19367_ | ~new_n19365_;
  assign po1410 = ~new_n19363_ | ~new_n19364_ | ~new_n19362_;
  assign po1409 = ~new_n19360_ | ~new_n19361_ | ~new_n19359_;
  assign po1408 = ~new_n19357_ | ~new_n19358_ | ~new_n19356_;
  assign po1407 = ~new_n19354_ | ~new_n19355_ | ~new_n19353_;
  assign po1406 = ~new_n19351_ | ~new_n19352_ | ~new_n19350_;
  assign po1405 = ~new_n19348_ | ~new_n19349_ | ~new_n19347_;
  assign po1404 = ~new_n19345_ | ~new_n19346_ | ~new_n19344_;
  assign po1403 = ~new_n19342_ | ~new_n19343_ | ~new_n19341_;
  assign po1402 = ~new_n19340_ | ~new_n19339_ | ~new_n19338_;
  assign po1401 = ~new_n19337_ | ~new_n19336_ | ~new_n19335_;
  assign po1400 = pi1341 & new_n19236_;
  assign po1399 = ~new_n17063_ | ~new_n19327_;
  assign po1398 = ~new_n17062_ | ~new_n19324_;
  assign po1397 = ~new_n17061_ | ~new_n19321_;
  assign po1396 = ~new_n17060_ | ~new_n19318_;
  assign po1395 = ~new_n17059_ | ~new_n19315_;
  assign po1394 = ~new_n17058_ | ~new_n19312_;
  assign po1393 = ~new_n17057_ | ~new_n19309_;
  assign po1392 = ~new_n17056_ | ~new_n19306_;
  assign po1391 = ~new_n17055_ | ~new_n19303_;
  assign po1390 = ~new_n17054_ | ~new_n19300_;
  assign po1389 = ~new_n17053_ | ~new_n19297_;
  assign po1388 = ~new_n17052_ | ~new_n19294_;
  assign po1387 = ~new_n17051_ | ~new_n19291_;
  assign po1386 = ~new_n17050_ | ~new_n19288_;
  assign po1385 = ~new_n17049_ | ~new_n19285_;
  assign po1384 = ~new_n19284_ | ~new_n19283_ | ~new_n19282_;
  assign po1383 = ~new_n19281_ | ~new_n19280_ | ~new_n19279_;
  assign po1382 = ~new_n19278_ | ~new_n19277_ | ~new_n19276_;
  assign po1381 = ~new_n19275_ | ~new_n19274_ | ~new_n19273_;
  assign po1380 = ~new_n19272_ | ~new_n19271_ | ~new_n19270_;
  assign po1379 = ~new_n19269_ | ~new_n19268_ | ~new_n19267_;
  assign po1378 = ~new_n19266_ | ~new_n19265_ | ~new_n19264_;
  assign po1377 = ~new_n19263_ | ~new_n19262_ | ~new_n19261_;
  assign po1376 = ~new_n19260_ | ~new_n19259_ | ~new_n19258_;
  assign po1375 = ~new_n19257_ | ~new_n19256_ | ~new_n19255_;
  assign po1374 = ~new_n19254_ | ~new_n19253_ | ~new_n19252_;
  assign po1373 = ~new_n19251_ | ~new_n19250_ | ~new_n19249_;
  assign po1372 = ~new_n19248_ | ~new_n19247_ | ~new_n19246_;
  assign po1371 = ~new_n19245_ | ~new_n19244_ | ~new_n19243_;
  assign po1370 = ~new_n19242_ | ~new_n19241_ | ~new_n19240_;
  assign po1369 = ~new_n19239_ | ~new_n19238_ | ~new_n19237_;
  assign po1368 = ~new_n20721_ | ~new_n20723_;
  assign po1367 = ~new_n20720_ | ~new_n20725_;
  assign po1366 = ~new_n20719_ | ~new_n20727_;
  assign po1365 = ~new_n20718_ | ~new_n20729_;
  assign po1364 = ~new_n20717_ | ~new_n20731_;
  assign po1363 = ~new_n20716_ | ~new_n20733_;
  assign po1362 = ~new_n20715_ | ~new_n20735_;
  assign po1361 = ~new_n20714_ | ~new_n20737_;
  assign po1360 = ~new_n20713_ | ~new_n20739_;
  assign po1359 = ~new_n20712_ | ~new_n20741_;
  assign po1358 = ~new_n20711_ | ~new_n20743_;
  assign po1357 = ~new_n20710_ | ~new_n20745_;
  assign po1356 = ~new_n20709_ | ~new_n20747_;
  assign po1355 = ~new_n20708_ | ~new_n20749_;
  assign po1354 = ~new_n20707_ | ~new_n20751_;
  assign po1353 = ~new_n20706_ | ~new_n20753_;
  assign po1352 = ~new_n20705_ | ~new_n20755_;
  assign po1351 = ~new_n20704_ | ~new_n20757_;
  assign po1350 = ~new_n20703_ | ~new_n20759_;
  assign po1349 = ~new_n20702_ | ~new_n20761_;
  assign po1348 = ~new_n20701_ | ~new_n20763_;
  assign po1347 = ~new_n20700_ | ~new_n20765_;
  assign po1346 = ~new_n20699_ | ~new_n20767_;
  assign po1345 = ~new_n20698_ | ~new_n20769_;
  assign po1344 = ~new_n20697_ | ~new_n20771_;
  assign po1343 = ~new_n20696_ | ~new_n20773_;
  assign po1342 = ~new_n20695_ | ~new_n20775_;
  assign po1341 = ~new_n20694_ | ~new_n20777_;
  assign po1340 = ~new_n20693_ | ~new_n20779_;
  assign po1339 = ~new_n20692_ | ~new_n20781_;
  assign po1338 = ~new_n20691_ | ~new_n20783_;
  assign po1337 = ~new_n19137_ | ~new_n19138_ | ~new_n19136_ | ~new_n19139_ | ~new_n19135_;
  assign po1336 = ~new_n19132_ | ~new_n19133_ | ~new_n19131_ | ~new_n19134_ | ~new_n19130_;
  assign po1335 = ~new_n19127_ | ~new_n19128_ | ~new_n19126_ | ~new_n19129_ | ~new_n19125_;
  assign po1334 = ~new_n19122_ | ~new_n19123_ | ~new_n19121_ | ~new_n19124_ | ~new_n19120_;
  assign po1333 = ~new_n19117_ | ~new_n19118_ | ~new_n19116_ | ~new_n19119_ | ~new_n19115_;
  assign po1332 = ~new_n19112_ | ~new_n19113_ | ~new_n19111_ | ~new_n19114_ | ~new_n19110_;
  assign po1331 = ~new_n19107_ | ~new_n19108_ | ~new_n19106_ | ~new_n19109_ | ~new_n19105_;
  assign po1330 = ~new_n19102_ | ~new_n19103_ | ~new_n19101_ | ~new_n19104_ | ~new_n19100_;
  assign po1329 = ~new_n19097_ | ~new_n19098_ | ~new_n19096_ | ~new_n19099_ | ~new_n19095_;
  assign po1328 = ~new_n19092_ | ~new_n19093_ | ~new_n19091_ | ~new_n19094_ | ~new_n19090_;
  assign po1327 = ~new_n19087_ | ~new_n19088_ | ~new_n19086_ | ~new_n19089_ | ~new_n19085_;
  assign po1326 = ~new_n19082_ | ~new_n19083_ | ~new_n19081_ | ~new_n19084_ | ~new_n19080_;
  assign po1325 = ~new_n19077_ | ~new_n19078_ | ~new_n19076_ | ~new_n19079_ | ~new_n19075_;
  assign po1324 = ~new_n19072_ | ~new_n19073_ | ~new_n19071_ | ~new_n19074_ | ~new_n19070_;
  assign po1323 = ~new_n19067_ | ~new_n19068_ | ~new_n19066_ | ~new_n19069_ | ~new_n19065_;
  assign po1322 = ~new_n19062_ | ~new_n19063_ | ~new_n19061_ | ~new_n19064_ | ~new_n19060_;
  assign po1321 = ~new_n19057_ | ~new_n19058_ | ~new_n19056_ | ~new_n19059_ | ~new_n19055_;
  assign po1320 = ~new_n19052_ | ~new_n19053_ | ~new_n19051_ | ~new_n19054_ | ~new_n19050_;
  assign po1319 = ~new_n19047_ | ~new_n19048_ | ~new_n19046_ | ~new_n19049_ | ~new_n19045_;
  assign po1318 = ~new_n19042_ | ~new_n19043_ | ~new_n19041_ | ~new_n19044_ | ~new_n19040_;
  assign po1317 = ~new_n19037_ | ~new_n19038_ | ~new_n19036_ | ~new_n19039_ | ~new_n19035_;
  assign po1316 = ~new_n19032_ | ~new_n19033_ | ~new_n19031_ | ~new_n19034_ | ~new_n19030_;
  assign po1315 = ~new_n19027_ | ~new_n19028_ | ~new_n19026_ | ~new_n19029_ | ~new_n19025_;
  assign po1314 = ~new_n19022_ | ~new_n19023_ | ~new_n19021_ | ~new_n19024_ | ~new_n19020_;
  assign po1313 = ~new_n19017_ | ~new_n19018_ | ~new_n19019_ | ~new_n19016_ | ~new_n19015_;
  assign po1312 = ~new_n19012_ | ~new_n19013_ | ~new_n19014_ | ~new_n19011_ | ~new_n19010_;
  assign po1311 = ~new_n19007_ | ~new_n19008_ | ~new_n19009_ | ~new_n19006_ | ~new_n19005_;
  assign po1310 = ~new_n19002_ | ~new_n19003_ | ~new_n19004_ | ~new_n19001_ | ~new_n19000_;
  assign po1309 = ~new_n18997_ | ~new_n18998_ | ~new_n18999_ | ~new_n18996_ | ~new_n18995_;
  assign po1308 = ~new_n18992_ | ~new_n18993_ | ~new_n18994_ | ~new_n18991_ | ~new_n18990_;
  assign po1307 = ~new_n18986_ | ~new_n18988_ | ~new_n18989_ | ~new_n18987_ | ~new_n18985_;
  assign po1306 = ~new_n18981_ | ~new_n18983_ | ~new_n18984_ | ~new_n18982_ | ~new_n18980_;
  assign po1305 = ~new_n17040_ | ~new_n18970_ | ~new_n18968_ | ~new_n17042_;
  assign po1304 = ~new_n17037_ | ~new_n18963_ | ~new_n18961_ | ~new_n17039_;
  assign po1303 = ~new_n17034_ | ~new_n18956_ | ~new_n18954_ | ~new_n17036_;
  assign po1302 = ~new_n17031_ | ~new_n18949_ | ~new_n18947_ | ~new_n17033_;
  assign po1301 = ~new_n17028_ | ~new_n18942_ | ~new_n18940_ | ~new_n17030_;
  assign po1300 = ~new_n17025_ | ~new_n18935_ | ~new_n18933_ | ~new_n17027_;
  assign po1299 = ~new_n17022_ | ~new_n18928_ | ~new_n18926_ | ~new_n17024_;
  assign po1298 = ~new_n17019_ | ~new_n18921_ | ~new_n18919_ | ~new_n17021_;
  assign po1297 = ~new_n17016_ | ~new_n18914_ | ~new_n18912_ | ~new_n17018_;
  assign po1296 = ~new_n17013_ | ~new_n18907_ | ~new_n18905_ | ~new_n17015_;
  assign po1295 = ~new_n17010_ | ~new_n18900_ | ~new_n18898_ | ~new_n17012_;
  assign po1294 = ~new_n17007_ | ~new_n18893_ | ~new_n18891_ | ~new_n17009_;
  assign po1293 = ~new_n17004_ | ~new_n18886_ | ~new_n18884_ | ~new_n17006_;
  assign po1292 = ~new_n17001_ | ~new_n18879_ | ~new_n18877_ | ~new_n17003_;
  assign po1291 = ~new_n16998_ | ~new_n18872_ | ~new_n18870_ | ~new_n17000_;
  assign po1290 = ~new_n16995_ | ~new_n18865_ | ~new_n18863_ | ~new_n16997_;
  assign po1289 = ~new_n16992_ | ~new_n18858_ | ~new_n18856_ | ~new_n16994_;
  assign po1288 = ~new_n16989_ | ~new_n18851_ | ~new_n18849_ | ~new_n16991_;
  assign po1287 = ~new_n16986_ | ~new_n18844_ | ~new_n18842_ | ~new_n16988_;
  assign po1286 = ~new_n18837_ | ~new_n16983_ | ~new_n16985_;
  assign po1285 = ~new_n18830_ | ~new_n16980_ | ~new_n16982_;
  assign po1284 = ~new_n18823_ | ~new_n16977_ | ~new_n16979_;
  assign po1283 = ~new_n18816_ | ~new_n16974_ | ~new_n16976_;
  assign po1282 = ~new_n18809_ | ~new_n16971_ | ~new_n16973_;
  assign po1281 = ~new_n18802_ | ~new_n16968_ | ~new_n16970_;
  assign po1280 = ~new_n18795_ | ~new_n16965_ | ~new_n16967_;
  assign po1279 = ~new_n18788_ | ~new_n16962_ | ~new_n16964_;
  assign po1278 = ~new_n18781_ | ~new_n16959_ | ~new_n16961_;
  assign po1277 = ~new_n16956_ | ~new_n16957_;
  assign po1276 = ~new_n16955_ | ~new_n16953_ | ~new_n16952_;
  assign po1275 = ~new_n16951_ | ~new_n16949_ | ~new_n16948_;
  assign po1274 = ~new_n16947_ | ~new_n16945_ | ~new_n16944_;
  assign po1269 = pi1210 & new_n18718_;
  assign po1263 = ~new_n16911_ | ~new_n18641_ | ~new_n18640_;
  assign po1262 = ~new_n16910_ | ~new_n18636_ | ~new_n18635_;
  assign po1261 = ~new_n16909_ | ~new_n18631_ | ~new_n18630_;
  assign po1260 = ~new_n16908_ | ~new_n18626_ | ~new_n18625_;
  assign po1259 = ~new_n16907_ | ~new_n20793_ | ~new_n18621_;
  assign po1258 = ~new_n16906_ | ~new_n18617_ | ~new_n18616_;
  assign po1257 = ~new_n16905_ | ~new_n18612_ | ~new_n18611_;
  assign po1256 = ~new_n16904_ | ~new_n18607_ | ~new_n18606_;
  assign po1255 = ~new_n16902_ | ~new_n18585_ | ~new_n18584_;
  assign po1254 = ~new_n16901_ | ~new_n18580_ | ~new_n18579_;
  assign po1253 = ~new_n16900_ | ~new_n18575_ | ~new_n18574_;
  assign po1252 = ~new_n16899_ | ~new_n18570_ | ~new_n18569_;
  assign po1251 = ~new_n16898_ | ~new_n18565_ | ~new_n18564_;
  assign po1250 = ~new_n16897_ | ~new_n18560_ | ~new_n18559_;
  assign po1249 = ~new_n16896_ | ~new_n18555_ | ~new_n18554_;
  assign po1248 = ~new_n16895_ | ~new_n18550_ | ~new_n18549_;
  assign po1247 = ~new_n16893_ | ~new_n18527_ | ~new_n18526_;
  assign po1246 = ~new_n16892_ | ~new_n18522_ | ~new_n18521_;
  assign po1245 = ~new_n16891_ | ~new_n18517_ | ~new_n18516_;
  assign po1244 = ~new_n16890_ | ~new_n18512_ | ~new_n18511_;
  assign po1243 = ~new_n16889_ | ~new_n18507_ | ~new_n18506_;
  assign po1242 = ~new_n16888_ | ~new_n18502_ | ~new_n18501_;
  assign po1241 = ~new_n16887_ | ~new_n18497_ | ~new_n18496_;
  assign po1240 = ~new_n16886_ | ~new_n18492_ | ~new_n18491_;
  assign po1239 = ~new_n16884_ | ~new_n18470_ | ~new_n18469_;
  assign po1238 = ~new_n16883_ | ~new_n18465_ | ~new_n18464_;
  assign po1237 = ~new_n16882_ | ~new_n18460_ | ~new_n18459_;
  assign po1236 = ~new_n16881_ | ~new_n18455_ | ~new_n18454_;
  assign po1235 = ~new_n16880_ | ~new_n18450_ | ~new_n18449_;
  assign po1234 = ~new_n16879_ | ~new_n18445_ | ~new_n18444_;
  assign po1233 = ~new_n16878_ | ~new_n18440_ | ~new_n18439_;
  assign po1232 = ~new_n16877_ | ~new_n18435_ | ~new_n18434_;
  assign po1231 = ~new_n16875_ | ~new_n18412_ | ~new_n18411_;
  assign po1230 = ~new_n16874_ | ~new_n18407_ | ~new_n18406_;
  assign po1229 = ~new_n16873_ | ~new_n18402_ | ~new_n18401_;
  assign po1228 = ~new_n16872_ | ~new_n18397_ | ~new_n18396_;
  assign po1227 = ~new_n16871_ | ~new_n18392_ | ~new_n18391_;
  assign po1226 = ~new_n16870_ | ~new_n18387_ | ~new_n18386_;
  assign po1225 = ~new_n16869_ | ~new_n18382_ | ~new_n18381_;
  assign po1224 = ~new_n16868_ | ~new_n18377_ | ~new_n18376_;
  assign po1223 = ~new_n16866_ | ~new_n18355_ | ~new_n18354_;
  assign po1222 = ~new_n16865_ | ~new_n18350_ | ~new_n18349_;
  assign po1221 = ~new_n16864_ | ~new_n18345_ | ~new_n18344_;
  assign po1220 = ~new_n16863_ | ~new_n18340_ | ~new_n18339_;
  assign po1219 = ~new_n16862_ | ~new_n18335_ | ~new_n18334_;
  assign po1218 = ~new_n16861_ | ~new_n18330_ | ~new_n18329_;
  assign po1217 = ~new_n16860_ | ~new_n18325_ | ~new_n18324_;
  assign po1216 = ~new_n16859_ | ~new_n18320_ | ~new_n18319_;
  assign po1215 = ~new_n16857_ | ~new_n18297_ | ~new_n18296_;
  assign po1214 = ~new_n16856_ | ~new_n18292_ | ~new_n18291_;
  assign po1213 = ~new_n16855_ | ~new_n18287_ | ~new_n18286_;
  assign po1212 = ~new_n16854_ | ~new_n18282_ | ~new_n18281_;
  assign po1211 = ~new_n16853_ | ~new_n18277_ | ~new_n18276_;
  assign po1210 = ~new_n16852_ | ~new_n18272_ | ~new_n18271_;
  assign po1209 = ~new_n16851_ | ~new_n18267_ | ~new_n18266_;
  assign po1208 = ~new_n16850_ | ~new_n18262_ | ~new_n18261_;
  assign po1207 = ~new_n16848_ | ~new_n18240_ | ~new_n18239_;
  assign po1206 = ~new_n16847_ | ~new_n18235_ | ~new_n18234_;
  assign po1205 = ~new_n16846_ | ~new_n18230_ | ~new_n18229_;
  assign po1204 = ~new_n16845_ | ~new_n18225_ | ~new_n18224_;
  assign po1203 = ~new_n16844_ | ~new_n18220_ | ~new_n18219_;
  assign po1202 = ~new_n16843_ | ~new_n18215_ | ~new_n18214_;
  assign po1201 = ~new_n16842_ | ~new_n18210_ | ~new_n18209_;
  assign po1200 = ~new_n16841_ | ~new_n18205_ | ~new_n18204_;
  assign po1199 = ~new_n16839_ | ~new_n18184_ | ~new_n18183_;
  assign po1198 = ~new_n16838_ | ~new_n18179_ | ~new_n18178_;
  assign po1197 = ~new_n16837_ | ~new_n18174_ | ~new_n18173_;
  assign po1196 = ~new_n16836_ | ~new_n18169_ | ~new_n18168_;
  assign po1195 = ~new_n16835_ | ~new_n18164_ | ~new_n18163_;
  assign po1194 = ~new_n16834_ | ~new_n18159_ | ~new_n18158_;
  assign po1193 = ~new_n16833_ | ~new_n18154_ | ~new_n18153_;
  assign po1192 = ~new_n16832_ | ~new_n18149_ | ~new_n18148_;
  assign po1191 = ~new_n16830_ | ~new_n18127_ | ~new_n18126_;
  assign po1190 = ~new_n16829_ | ~new_n18122_ | ~new_n18121_;
  assign po1189 = ~new_n16828_ | ~new_n18117_ | ~new_n18116_;
  assign po1188 = ~new_n16827_ | ~new_n18112_ | ~new_n18111_;
  assign po1187 = ~new_n16826_ | ~new_n18107_ | ~new_n18106_;
  assign po1186 = ~new_n16825_ | ~new_n18102_ | ~new_n18101_;
  assign po1185 = ~new_n16824_ | ~new_n18097_ | ~new_n18096_;
  assign po1184 = ~new_n16823_ | ~new_n18092_ | ~new_n18091_;
  assign po1183 = ~new_n16821_ | ~new_n18069_ | ~new_n18068_;
  assign po1182 = ~new_n16820_ | ~new_n18064_ | ~new_n18063_;
  assign po1181 = ~new_n16819_ | ~new_n18059_ | ~new_n18058_;
  assign po1180 = ~new_n16818_ | ~new_n18054_ | ~new_n18053_;
  assign po1179 = ~new_n16817_ | ~new_n18049_ | ~new_n18048_;
  assign po1178 = ~new_n16816_ | ~new_n18044_ | ~new_n18043_;
  assign po1177 = ~new_n16815_ | ~new_n18039_ | ~new_n18038_;
  assign po1176 = ~new_n16814_ | ~new_n18034_ | ~new_n18033_;
  assign po1175 = ~new_n16812_ | ~new_n18012_ | ~new_n18011_;
  assign po1174 = ~new_n16811_ | ~new_n18007_ | ~new_n18006_;
  assign po1173 = ~new_n16810_ | ~new_n18002_ | ~new_n18001_;
  assign po1172 = ~new_n16809_ | ~new_n17997_ | ~new_n17996_;
  assign po1171 = ~new_n16808_ | ~new_n17992_ | ~new_n17991_;
  assign po1170 = ~new_n16807_ | ~new_n17987_ | ~new_n17986_;
  assign po1169 = ~new_n16806_ | ~new_n17982_ | ~new_n17981_;
  assign po1168 = ~new_n16805_ | ~new_n17977_ | ~new_n17976_;
  assign po1167 = ~new_n16803_ | ~new_n17954_ | ~new_n17953_;
  assign po1166 = ~new_n16802_ | ~new_n17949_ | ~new_n17948_;
  assign po1165 = ~new_n16801_ | ~new_n17944_ | ~new_n17943_;
  assign po1164 = ~new_n16800_ | ~new_n17939_ | ~new_n17938_;
  assign po1163 = ~new_n16799_ | ~new_n17934_ | ~new_n17933_;
  assign po1162 = ~new_n16798_ | ~new_n17929_ | ~new_n17928_;
  assign po1161 = ~new_n16797_ | ~new_n17924_ | ~new_n17923_;
  assign po1160 = ~new_n16796_ | ~new_n17919_ | ~new_n17918_;
  assign po1159 = ~new_n16794_ | ~new_n17897_ | ~new_n17896_;
  assign po1158 = ~new_n16793_ | ~new_n17892_ | ~new_n17891_;
  assign po1157 = ~new_n16792_ | ~new_n17887_ | ~new_n17886_;
  assign po1156 = ~new_n16791_ | ~new_n17882_ | ~new_n17881_;
  assign po1155 = ~new_n16790_ | ~new_n17877_ | ~new_n17876_;
  assign po1154 = ~new_n16789_ | ~new_n17872_ | ~new_n17871_;
  assign po1153 = ~new_n16788_ | ~new_n17867_ | ~new_n17866_;
  assign po1152 = ~new_n16787_ | ~new_n17862_ | ~new_n17861_;
  assign po1151 = ~new_n16785_ | ~new_n17838_ | ~new_n17837_;
  assign po1150 = ~new_n16784_ | ~new_n17833_ | ~new_n17832_;
  assign po1149 = ~new_n16783_ | ~new_n17828_ | ~new_n17827_;
  assign po1148 = ~new_n16782_ | ~new_n17823_ | ~new_n17822_;
  assign po1147 = ~new_n16781_ | ~new_n17818_ | ~new_n17817_;
  assign po1146 = ~new_n16780_ | ~new_n17813_ | ~new_n17812_;
  assign po1145 = ~new_n16779_ | ~new_n17808_ | ~new_n17807_;
  assign po1144 = ~new_n16778_ | ~new_n17803_ | ~new_n17802_;
  assign po1143 = ~new_n16776_ | ~new_n17780_ | ~new_n17779_;
  assign po1142 = ~new_n16775_ | ~new_n17775_ | ~new_n17774_;
  assign po1141 = ~new_n16774_ | ~new_n17770_ | ~new_n17769_;
  assign po1140 = ~new_n16773_ | ~new_n17765_ | ~new_n17764_;
  assign po1139 = ~new_n16772_ | ~new_n17760_ | ~new_n17759_;
  assign po1138 = ~new_n16771_ | ~new_n17755_ | ~new_n17754_;
  assign po1137 = ~new_n16770_ | ~new_n17750_ | ~new_n17749_;
  assign po1136 = ~new_n16769_ | ~new_n17745_ | ~new_n17744_;
  assign po1135 = ~new_n16767_ | ~new_n20871_ | ~new_n20870_;
  assign po1134 = ~new_n17700_ | ~new_n17425_ | ~new_n17699_ | ~new_n17701_;
  assign po1133 = ~new_n16763_ | ~new_n17697_;
  assign po1131 = pi1072 & new_n20831_;
  assign po1130 = pi1071 & new_n20831_;
  assign po1129 = pi1070 & new_n20831_;
  assign po1128 = pi1069 & new_n20831_;
  assign po1127 = pi1068 & new_n20831_;
  assign po1126 = pi1067 & new_n20831_;
  assign po1125 = pi1066 & new_n20831_;
  assign po1124 = pi1065 & new_n20831_;
  assign po1123 = pi1064 & new_n20831_;
  assign po1122 = pi1063 & new_n20831_;
  assign po1121 = pi1062 & new_n20831_;
  assign po1120 = pi1061 & new_n20831_;
  assign po1119 = pi1060 & new_n20831_;
  assign po1118 = pi1059 & new_n20831_;
  assign po1117 = pi1058 & new_n20831_;
  assign po1116 = pi1057 & new_n20831_;
  assign po1115 = pi1056 & new_n20831_;
  assign po1114 = pi1055 & new_n20831_;
  assign po1113 = pi1054 & new_n20831_;
  assign po1112 = pi1053 & new_n20831_;
  assign po1111 = pi1052 & new_n20831_;
  assign po1110 = pi1051 & new_n20831_;
  assign po1109 = pi1050 & new_n20831_;
  assign po1108 = pi1049 & new_n20831_;
  assign po1107 = pi1048 & new_n20831_;
  assign po1106 = pi1047 & new_n20831_;
  assign po1105 = pi1046 & new_n20831_;
  assign po1104 = pi1045 & new_n20831_;
  assign po1103 = pi1044 & new_n20831_;
  assign po1102 = pi1043 & new_n20831_;
  assign po1099 = ~new_n17556_ | ~new_n20828_ | ~new_n20827_;
  assign po1098 = ~new_n16676_ | ~new_n20826_ | ~new_n20825_;
  assign po1097 = ~new_n16675_ | ~new_n17550_;
  assign po1096 = ~new_n17537_ | ~new_n17536_ | ~new_n17535_;
  assign po1095 = ~new_n17534_ | ~new_n17533_ | ~new_n17532_;
  assign po1094 = ~new_n17531_ | ~new_n17530_ | ~new_n17529_;
  assign po1093 = ~new_n17528_ | ~new_n17527_ | ~new_n17526_;
  assign po1092 = ~new_n17525_ | ~new_n17524_ | ~new_n17523_;
  assign po1091 = ~new_n17522_ | ~new_n17521_ | ~new_n17520_;
  assign po1090 = ~new_n17519_ | ~new_n17518_ | ~new_n17517_;
  assign po1089 = ~new_n17516_ | ~new_n17515_ | ~new_n17514_;
  assign po1088 = ~new_n17513_ | ~new_n17512_ | ~new_n17511_;
  assign po1087 = ~new_n17510_ | ~new_n17509_ | ~new_n17508_;
  assign po1086 = ~new_n17507_ | ~new_n17506_ | ~new_n17505_;
  assign po1085 = ~new_n17504_ | ~new_n17503_ | ~new_n17502_;
  assign po1084 = ~new_n17501_ | ~new_n17500_ | ~new_n17499_;
  assign po1083 = ~new_n17498_ | ~new_n17497_ | ~new_n17496_;
  assign po1082 = ~new_n17495_ | ~new_n17494_ | ~new_n17493_;
  assign po1081 = ~new_n17492_ | ~new_n17491_ | ~new_n17490_;
  assign po1080 = ~new_n17489_ | ~new_n17488_ | ~new_n17487_;
  assign po1079 = ~new_n17486_ | ~new_n17485_ | ~new_n17484_;
  assign po1078 = ~new_n17483_ | ~new_n17482_ | ~new_n17481_;
  assign po1077 = ~new_n17480_ | ~new_n17479_ | ~new_n17478_;
  assign po1076 = ~new_n17477_ | ~new_n17476_ | ~new_n17475_;
  assign po1075 = ~new_n17474_ | ~new_n17473_ | ~new_n17472_;
  assign po1074 = ~new_n17471_ | ~new_n17470_ | ~new_n17469_;
  assign po1073 = ~new_n17468_ | ~new_n17467_ | ~new_n17466_;
  assign po1072 = ~new_n17465_ | ~new_n17464_ | ~new_n17463_;
  assign po1071 = ~new_n17462_ | ~new_n17461_ | ~new_n17460_;
  assign po1070 = ~new_n17459_ | ~new_n17458_ | ~new_n17457_;
  assign po1069 = ~new_n17456_ | ~new_n17455_ | ~new_n17454_;
  assign po1068 = ~new_n17453_ | ~new_n17452_ | ~new_n17451_;
  assign po1067 = ~new_n17450_ | ~new_n17449_ | ~new_n17448_;
  assign new_n16408_ = ~new_n17181_ | ~new_n17179_ | ~new_n17180_ | ~new_n17182_;
  assign new_n16409_ = ~new_n17177_ | ~new_n17175_ | ~new_n17176_ | ~new_n17178_;
  assign new_n16410_ = ~new_n17173_ | ~new_n17171_ | ~new_n17172_ | ~new_n17174_;
  assign new_n16411_ = ~new_n17169_ | ~new_n17167_ | ~new_n17168_ | ~new_n17170_;
  assign new_n16412_ = ~new_n17165_ | ~new_n17163_ | ~new_n17164_ | ~new_n17166_;
  assign new_n16413_ = ~new_n17161_ | ~new_n17159_ | ~new_n17160_ | ~new_n17162_;
  assign new_n16414_ = ~new_n17157_ | ~new_n17155_ | ~new_n17156_ | ~new_n17158_;
  assign new_n16415_ = ~new_n17153_ | ~new_n17151_ | ~new_n17152_ | ~new_n17154_;
  assign new_n16416_ = ~new_n16510_ | ~new_n16504_;
  assign new_n16417_ = ~new_n15613_ | ~new_n16416_;
  assign new_n16418_ = ~new_n15613_ | ~new_n17724_;
  assign new_n16419_ = ~new_n15615_ | ~new_n16416_;
  assign new_n16420_ = ~new_n15615_ | ~new_n17724_;
  assign new_n16421_ = ~new_n15614_ | ~new_n16416_;
  assign new_n16422_ = ~new_n15614_ | ~new_n17724_;
  assign new_n16423_ = ~new_n15616_ | ~new_n16416_;
  assign new_n16424_ = ~new_n15616_ | ~new_n17724_;
  assign new_n16425_ = ~new_n18644_ | ~new_n16572_ | ~new_n16575_;
  assign new_n16426_ = ~new_n20267_ | ~new_n18645_;
  assign new_n16427_ = ~new_n20972_ | ~new_n17337_ | ~new_n17339_ | ~new_n20973_;
  assign new_n16428_ = ~pi1446;
  assign new_n16429_ = ~pi1039;
  assign new_n16430_ = ~pi1039 | ~new_n16439_;
  assign new_n16431_ = ~new_n17402_ | ~new_n16432_;
  assign new_n16432_ = ~pi1038;
  assign new_n16433_ = ~pi1038 | ~new_n17402_;
  assign new_n16434_ = ~pi1407;
  assign new_n16435_ = ~pi1039 | ~new_n16432_;
  assign new_n16436_ = pi1039 | pi1038;
  assign new_n16437_ = ~pi0033;
  assign new_n16438_ = ~new_n2972_;
  assign new_n16439_ = ~pi1040;
  assign new_n16440_ = ~pi1040 | ~new_n16441_;
  assign new_n16441_ = ~pi1446 | ~new_n16437_;
  assign new_n16442_ = pi0033 | pi1446;
  assign new_n16443_ = ~pi1075;
  assign new_n16444_ = ~pi1074;
  assign new_n16445_ = ~pi1207;
  assign new_n16446_ = ~pi1208;
  assign new_n16447_ = ~pi1209;
  assign new_n16448_ = ~pi1208 | ~new_n16451_ | ~pi1207 | ~pi1209;
  assign new_n16449_ = pi1208 | pi1207 | pi1209;
  assign new_n16450_ = pi1208 | pi1209;
  assign new_n16451_ = ~pi1206;
  assign new_n16452_ = ~new_n16747_ | ~new_n16745_ | ~new_n16746_ | ~new_n16748_;
  assign new_n16453_ = ~new_n17677_ | ~new_n16439_;
  assign new_n16454_ = ~new_n33065_;
  assign new_n16455_ = ~pi1207 | ~new_n16451_;
  assign new_n16456_ = ~pi1209 | ~pi1208;
  assign new_n16457_ = ~new_n16699_ | ~new_n16697_ | ~new_n16698_ | ~new_n16700_;
  assign new_n16458_ = ~new_n16720_ | ~new_n16717_ | ~new_n16718_ | ~new_n16719_ | ~new_n17351_;
  assign new_n16459_ = ~new_n16737_ | ~new_n16735_ | ~new_n16736_ | ~new_n16738_;
  assign new_n16460_ = ~new_n16740_ | ~new_n16739_;
  assign new_n16461_ = pi1445 | new_n2972_;
  assign new_n16462_ = ~new_n33065_ | ~new_n17678_;
  assign new_n16463_ = ~new_n17658_ | ~new_n16465_;
  assign new_n16464_ = ~new_n16691_ | ~new_n16689_ | ~new_n16690_ | ~new_n16692_;
  assign new_n16465_ = ~new_n16743_ | ~new_n16741_ | ~new_n16742_ | ~new_n16744_;
  assign new_n16466_ = ~new_n15654_ | ~new_n17682_;
  assign new_n16467_ = ~new_n15570_ | ~new_n16464_;
  assign new_n16468_ = ~new_n17675_ | ~new_n17658_;
  assign new_n16469_ = ~new_n17430_ | ~new_n15628_;
  assign new_n16470_ = ~new_n16572_ | ~new_n16459_ | ~new_n17354_ | ~new_n17641_;
  assign new_n16471_ = ~new_n16452_ | ~new_n16464_;
  assign new_n16472_ = ~new_n17371_ | ~new_n16465_;
  assign new_n16473_ = ~new_n17437_ | ~new_n15612_;
  assign new_n16474_ = ~new_n17359_ | ~new_n33474_ | ~new_n17406_ | ~new_n20807_ | ~new_n17690_;
  assign new_n16475_ = ~pi1076;
  assign new_n16476_ = ~pi1076 | ~new_n20785_;
  assign new_n16477_ = ~pi1073;
  assign new_n16478_ = ~pi1074 | ~new_n16443_;
  assign new_n16479_ = pi1074 | pi1075;
  assign new_n16480_ = ~pi1073 | ~new_n33065_;
  assign new_n16481_ = ~new_n17728_ | ~new_n16475_;
  assign new_n16482_ = ~pi1214;
  assign new_n16483_ = ~pi1213;
  assign new_n16484_ = ~pi1211;
  assign new_n16485_ = ~pi1212;
  assign new_n16486_ = ~pi1213 | ~pi1214;
  assign new_n16487_ = ~new_n17714_ | ~new_n15659_;
  assign new_n16488_ = pi1074 | pi1073;
  assign new_n16489_ = ~pi1445;
  assign new_n16490_ = ~new_n31270_;
  assign new_n16491_ = ~new_n31277_;
  assign new_n16492_ = ~new_n31276_;
  assign new_n16493_ = ~new_n31235_;
  assign new_n16494_ = ~new_n31277_ | ~new_n31270_;
  assign new_n16495_ = ~new_n16513_ | ~new_n16490_;
  assign new_n16496_ = ~new_n17708_ | ~new_n15656_;
  assign new_n16497_ = ~new_n31170_;
  assign new_n16498_ = ~new_n31187_;
  assign new_n16499_ = ~new_n31179_;
  assign new_n16500_ = ~new_n31178_;
  assign new_n16501_ = ~new_n17390_ | ~new_n16489_;
  assign new_n16502_ = ~new_n16487_ | ~new_n17716_;
  assign new_n16503_ = ~new_n16487_ | ~new_n17725_;
  assign new_n16504_ = ~pi1213 | ~new_n16482_;
  assign new_n16505_ = ~new_n17723_ | ~new_n15659_;
  assign new_n16506_ = ~new_n31277_ | ~new_n16490_;
  assign new_n16507_ = ~new_n31270_ | ~new_n16513_;
  assign new_n16508_ = ~new_n17781_ | ~new_n15656_;
  assign new_n16509_ = ~new_n16505_ | ~new_n17784_;
  assign new_n16510_ = ~pi1214 | ~new_n16483_;
  assign new_n16511_ = ~new_n17722_ | ~new_n15659_;
  assign new_n16512_ = ~new_n31270_ | ~new_n16491_;
  assign new_n16513_ = ~new_n16506_ | ~new_n16512_;
  assign new_n16514_ = ~new_n17707_ | ~new_n16490_;
  assign new_n16515_ = ~new_n17839_ | ~new_n15656_;
  assign new_n16516_ = ~new_n16511_ | ~new_n17842_;
  assign new_n16517_ = ~new_n16511_ | ~new_n17844_;
  assign new_n16518_ = ~new_n15669_ | ~new_n15659_;
  assign new_n16519_ = ~new_n15666_ | ~new_n15656_;
  assign new_n16520_ = ~new_n16518_ | ~new_n17900_;
  assign new_n16521_ = ~pi1211 | ~new_n16485_;
  assign new_n16522_ = ~new_n17719_ | ~new_n17714_;
  assign new_n16523_ = ~new_n31235_ | ~new_n16492_;
  assign new_n16524_ = ~new_n15671_ | ~new_n17708_;
  assign new_n16525_ = ~new_n16522_ | ~new_n17957_;
  assign new_n16526_ = ~new_n16522_ | ~new_n17959_;
  assign new_n16527_ = ~new_n17719_ | ~new_n17723_;
  assign new_n16528_ = ~new_n15671_ | ~new_n17781_;
  assign new_n16529_ = ~new_n16527_ | ~new_n18015_;
  assign new_n16530_ = ~new_n17719_ | ~new_n17722_;
  assign new_n16531_ = ~new_n15671_ | ~new_n17839_;
  assign new_n16532_ = ~new_n16530_ | ~new_n18072_;
  assign new_n16533_ = ~new_n16530_ | ~new_n18074_;
  assign new_n16534_ = ~new_n17719_ | ~new_n15669_;
  assign new_n16535_ = ~new_n15671_ | ~new_n15666_;
  assign new_n16536_ = ~new_n16534_ | ~new_n18130_;
  assign new_n16537_ = ~new_n15660_ | ~new_n17714_;
  assign new_n16538_ = ~new_n15655_ | ~new_n17709_;
  assign new_n16539_ = ~new_n16538_ | ~new_n16523_ | ~new_n17711_;
  assign new_n16540_ = ~new_n15680_ | ~new_n17708_;
  assign new_n16541_ = ~new_n16537_ | ~new_n16521_ | ~new_n17720_;
  assign new_n16542_ = ~new_n16537_ | ~new_n18186_;
  assign new_n16543_ = ~new_n16537_ | ~new_n18188_;
  assign new_n16544_ = ~new_n17723_ | ~new_n15660_;
  assign new_n16545_ = ~new_n15680_ | ~new_n17781_;
  assign new_n16546_ = ~new_n16544_ | ~new_n18243_;
  assign new_n16547_ = ~new_n17722_ | ~new_n15660_;
  assign new_n16548_ = ~new_n15680_ | ~new_n17839_;
  assign new_n16549_ = ~new_n16547_ | ~new_n18300_;
  assign new_n16550_ = ~new_n16547_ | ~new_n18302_;
  assign new_n16551_ = ~new_n15669_ | ~new_n15660_;
  assign new_n16552_ = ~new_n15680_ | ~new_n15666_;
  assign new_n16553_ = ~new_n16551_ | ~new_n18358_;
  assign new_n16554_ = ~new_n15691_ | ~new_n17714_;
  assign new_n16555_ = ~new_n15688_ | ~new_n17708_;
  assign new_n16556_ = ~new_n16554_ | ~new_n18415_;
  assign new_n16557_ = ~new_n16554_ | ~new_n18417_;
  assign new_n16558_ = ~new_n15691_ | ~new_n17723_;
  assign new_n16559_ = ~new_n15688_ | ~new_n17781_;
  assign new_n16560_ = ~new_n16558_ | ~new_n18473_;
  assign new_n16561_ = ~new_n15691_ | ~new_n17722_;
  assign new_n16562_ = ~new_n15688_ | ~new_n17839_;
  assign new_n16563_ = ~new_n16561_ | ~new_n18530_;
  assign new_n16564_ = ~new_n16561_ | ~new_n18532_;
  assign new_n16565_ = ~new_n15691_ | ~new_n15669_;
  assign new_n16566_ = ~new_n15688_ | ~new_n15666_;
  assign new_n16567_ = ~new_n16565_ | ~new_n18588_;
  assign new_n16568_ = ~pi1443;
  assign new_n16569_ = ~new_n9378_;
  assign new_n16570_ = ~new_n16465_ | ~new_n16459_;
  assign new_n16571_ = ~new_n16465_ | ~new_n16452_;
  assign new_n16572_ = ~new_n16695_ | ~new_n16693_ | ~new_n16694_ | ~new_n16696_;
  assign new_n16573_ = ~new_n20809_ | ~new_n18671_ | ~new_n18670_;
  assign new_n16574_ = ~new_n17580_ | ~new_n16465_;
  assign new_n16575_ = ~new_n15786_ | ~new_n16458_;
  assign new_n16576_ = ~new_n17675_ | ~new_n17580_ | ~new_n20675_;
  assign new_n16577_ = ~new_n16922_ | ~new_n17428_;
  assign new_n16578_ = ~new_n20675_ | ~new_n17580_ | ~new_n17675_ | ~new_n15786_ | ~new_n17658_;
  assign new_n16579_ = ~new_n15786_ | ~new_n17581_ | ~new_n17630_ | ~new_n17352_ | ~new_n17641_;
  assign new_n16580_ = ~new_n17415_ | ~new_n17380_ | ~new_n17658_;
  assign new_n16581_ = ~new_n15630_ | ~new_n15628_;
  assign new_n16582_ = ~new_n16625_ | ~new_n18691_;
  assign new_n16583_ = ~new_n16450_ | ~new_n16456_;
  assign new_n16584_ = ~new_n32701_;
  assign new_n16585_ = ~new_n18717_ | ~new_n17423_ | ~new_n16481_;
  assign new_n16586_ = ~new_n16465_ | ~pi1076 | ~new_n16459_;
  assign new_n16587_ = ~new_n16452_ | ~new_n16454_;
  assign new_n16588_ = ~new_n16458_ | ~new_n16572_;
  assign new_n16589_ = ~new_n15608_ | ~new_n16475_;
  assign new_n16590_ = ~new_n17641_ | ~new_n16572_;
  assign new_n16591_ = ~new_n17434_ | ~new_n16459_;
  assign new_n16592_ = ~new_n17371_ | ~new_n15633_;
  assign new_n16593_ = ~pi1074 | ~new_n16452_;
  assign new_n16594_ = ~pi1406;
  assign new_n16595_ = ~new_n16937_ | ~new_n18743_;
  assign new_n16596_ = ~new_n17581_ | ~new_n17354_;
  assign new_n16597_ = ~new_n17044_ | ~new_n17429_;
  assign new_n16598_ = ~new_n19235_ | ~new_n19234_;
  assign new_n16599_ = ~pi1076 | ~new_n17675_;
  assign new_n16600_ = ~new_n17580_ | ~new_n20675_;
  assign new_n16601_ = ~new_n17387_ | ~new_n17658_;
  assign new_n16602_ = ~new_n17375_ | ~new_n15612_;
  assign new_n16603_ = ~new_n17391_ | ~pi1076;
  assign new_n16604_ = ~new_n17684_ | ~new_n16572_;
  assign new_n16605_ = ~new_n17416_ | ~new_n19334_;
  assign new_n16606_ = ~pi1076 | ~new_n17397_;
  assign new_n16607_ = ~new_n17416_ | ~new_n19445_;
  assign new_n16608_ = ~new_n17430_ | ~new_n15633_ | ~new_n17067_ | ~pi1076;
  assign new_n16609_ = ~new_n17047_ | ~new_n15628_;
  assign new_n16610_ = ~pi1405;
  assign new_n16611_ = ~new_n33164_;
  assign new_n16612_ = ~new_n17409_ | ~new_n17068_;
  assign new_n16613_ = ~new_n17390_ | ~new_n16443_;
  assign new_n16614_ = ~new_n17139_ | ~new_n17133_ | ~new_n17136_ | ~new_n17143_;
  assign new_n16615_ = ~new_n17387_ | ~new_n16452_;
  assign new_n16616_ = ~pi1449;
  assign new_n16617_ = ~pi1451;
  assign new_n16618_ = ~new_n15628_ | ~new_n17679_;
  assign new_n16619_ = ~new_n16448_ | ~new_n18663_;
  assign new_n16620_ = ~new_n17630_ | ~pi1074;
  assign new_n16621_ = ~pi1445 | ~new_n16444_;
  assign new_n16622_ = ~new_n16415_;
  assign new_n16623_ = ~new_n18660_ | ~new_n18659_;
  assign new_n16624_ = ~new_n15631_ | ~new_n16622_;
  assign new_n16625_ = ~pi1209 | ~pi1208 | ~new_n16445_;
  assign new_n16626_ = ~new_n16455_ | ~new_n20245_;
  assign new_n16627_ = ~new_n17378_ | ~new_n17415_;
  assign new_n16628_ = ~new_n17431_ | ~new_n17412_ | ~new_n17581_;
  assign new_n16629_ = ~new_n17431_ | ~new_n17412_ | ~new_n16459_;
  assign new_n16630_ = ~new_n17658_ | ~new_n17677_;
  assign new_n16631_ = ~new_n20274_ | ~new_n17258_ | ~new_n17256_ | ~new_n17255_;
  assign new_n16632_ = ~new_n17435_ | ~new_n17447_;
  assign new_n16633_ = ~new_n17364_ | ~new_n16449_;
  assign new_n16634_ = ~pi1076 | ~new_n15786_;
  assign new_n16635_ = ~new_n20873_ | ~new_n20872_;
  assign new_n16636_ = ~new_n20876_ | ~new_n20875_;
  assign new_n16637_ = ~new_n20900_ | ~new_n20899_;
  assign new_n16638_ = ~new_n20970_ | ~new_n20969_;
  assign po1063 = ~new_n20815_ | ~new_n20814_;
  assign po1064 = ~new_n20817_ | ~new_n20816_;
  assign po1065 = ~new_n20819_ | ~new_n20818_;
  assign po1066 = ~new_n20821_ | ~new_n20820_;
  assign new_n16643_ = ~new_n20830_ | ~new_n20829_;
  assign new_n16644_ = new_n16436_ & new_n17360_;
  assign po1100 = ~new_n20833_ | ~new_n20832_;
  assign po1101 = ~new_n20835_ | ~new_n20834_;
  assign po1132 = ~new_n20867_ | ~new_n20866_;
  assign new_n16648_ = new_n31169_ & new_n15608_ & new_n17396_;
  assign po1264 = ~new_n20883_ | ~new_n20882_;
  assign po1265 = ~new_n20890_ | ~new_n20889_;
  assign new_n16651_ = ~new_n20892_ | ~new_n20891_;
  assign new_n16652_ = ~new_n20895_ | ~new_n20894_;
  assign po1266 = ~new_n20903_ | ~new_n20902_;
  assign po1267 = ~new_n20905_ | ~new_n20904_;
  assign po1268 = ~new_n20909_ | ~new_n20908_;
  assign po1270 = ~new_n20911_ | ~new_n20910_;
  assign po1271 = ~new_n20916_ | ~new_n20915_;
  assign po1272 = ~new_n20918_ | ~new_n20917_;
  assign po1273 = ~new_n20920_ | ~new_n20919_;
  assign new_n16660_ = new_n32111_ & new_n17630_;
  assign new_n16661_ = ~pi1042 & ~pi1407;
  assign po1498 = ~new_n20936_ | ~new_n20935_;
  assign po1500 = ~new_n20940_ | ~new_n20939_;
  assign po1501 = ~new_n20942_ | ~new_n20941_;
  assign po1503 = ~new_n20944_ | ~new_n20943_;
  assign po1505 = ~new_n20948_ | ~new_n20947_;
  assign po1507 = ~new_n20952_ | ~new_n20951_;
  assign po1510 = ~new_n20954_ | ~new_n20953_;
  assign new_n16669_ = new_n31169_ & new_n17396_;
  assign new_n16670_ = ~new_n20956_ | ~new_n20955_;
  assign new_n16671_ = ~new_n20958_ | ~new_n20957_;
  assign new_n16672_ = ~new_n20960_ | ~new_n20959_;
  assign new_n16673_ = ~new_n20962_ | ~new_n20961_;
  assign new_n16674_ = ~new_n20964_ | ~new_n20963_;
  assign new_n16675_ = new_n17549_ & new_n16433_;
  assign new_n16676_ = new_n17551_ & new_n16431_;
  assign new_n16677_ = pi1446 & pi1040;
  assign new_n16678_ = ~pi1207 & ~pi1206;
  assign new_n16679_ = pi1209 & pi1208;
  assign new_n16680_ = ~pi1208 & ~pi1206;
  assign new_n16681_ = pi1209 & pi1207;
  assign new_n16682_ = ~pi1209 & ~pi1206;
  assign new_n16683_ = pi1208 & pi1207;
  assign new_n16684_ = ~pi1208 & ~pi1207;
  assign new_n16685_ = pi1206 & pi1209;
  assign new_n16686_ = ~pi1209 & ~pi1207;
  assign new_n16687_ = pi1206 & pi1208;
  assign new_n16688_ = pi1206 & pi1207;
  assign new_n16689_ = new_n17566_ & new_n17564_ & new_n17565_ & new_n17567_;
  assign new_n16690_ = new_n17570_ & new_n17568_ & new_n17569_ & new_n17571_;
  assign new_n16691_ = new_n17574_ & new_n17572_ & new_n17573_ & new_n17575_;
  assign new_n16692_ = new_n17578_ & new_n17576_ & new_n17577_ & new_n17579_;
  assign new_n16693_ = new_n17616_ & new_n17614_ & new_n17615_ & new_n17617_;
  assign new_n16694_ = new_n17620_ & new_n17618_ & new_n17619_ & new_n17621_;
  assign new_n16695_ = new_n17624_ & new_n17622_ & new_n17623_ & new_n17625_;
  assign new_n16696_ = new_n17628_ & new_n17626_ & new_n17627_ & new_n17629_;
  assign new_n16697_ = new_n17599_ & new_n17597_ & new_n17598_ & new_n17600_;
  assign new_n16698_ = new_n17603_ & new_n17601_ & new_n17602_ & new_n17604_;
  assign new_n16699_ = new_n17607_ & new_n17605_ & new_n17606_ & new_n17608_;
  assign new_n16700_ = new_n17611_ & new_n17609_ & new_n17610_ & new_n17612_;
  assign new_n16701_ = ~pi1208 & ~pi1206;
  assign new_n16702_ = pi1159 & pi1209;
  assign new_n16703_ = ~pi1209 & ~pi1206;
  assign new_n16704_ = pi1151 & pi1208;
  assign new_n16705_ = pi1206 & pi1135;
  assign new_n16706_ = ~pi1209 & ~pi1207;
  assign new_n16707_ = pi1119 & pi1206;
  assign new_n16708_ = pi1103 & pi1206;
  assign new_n16709_ = ~pi1208 & ~pi1207;
  assign new_n16710_ = pi1127 & pi1209;
  assign new_n16711_ = new_n17584_ & new_n17582_ & new_n17583_ & new_n17585_;
  assign new_n16712_ = new_n17588_ & new_n17586_ & new_n17587_ & new_n17589_;
  assign new_n16713_ = new_n17592_ & new_n17590_ & new_n17591_ & new_n17593_;
  assign new_n16714_ = new_n17595_ & new_n17594_;
  assign new_n16715_ = ~pi1207 & ~pi1206;
  assign new_n16716_ = pi1174 & pi1209;
  assign new_n16717_ = new_n17633_ & new_n17631_ & new_n17632_ & new_n17634_;
  assign new_n16718_ = new_n17637_ & new_n17636_ & new_n17635_;
  assign new_n16719_ = new_n17640_ & new_n17639_ & new_n17638_;
  assign new_n16720_ = new_n20858_ & new_n20856_ & new_n20857_ & new_n20859_;
  assign new_n16721_ = ~pi1207 & ~pi1206;
  assign new_n16722_ = pi1192 & pi1209;
  assign new_n16723_ = ~pi1209 & ~pi1208;
  assign new_n16724_ = pi1168 & pi1207;
  assign new_n16725_ = ~pi1209 & ~pi1208;
  assign new_n16726_ = pi1104 & pi1207;
  assign new_n16727_ = pi1209 & pi1207;
  assign new_n16728_ = pi1096 & pi1206;
  assign new_n16729_ = ~pi1209 & ~pi1206;
  assign new_n16730_ = pi1152 & pi1207;
  assign new_n16731_ = pi1208 & pi1207;
  assign new_n16732_ = pi1088 & pi1206;
  assign new_n16733_ = ~pi1208 & ~pi1207;
  assign new_n16734_ = pi1128 & pi1206;
  assign new_n16735_ = new_n20838_ & new_n20836_ & new_n20837_ & new_n20839_;
  assign new_n16736_ = new_n20842_ & new_n20840_ & new_n20841_ & new_n20843_;
  assign new_n16737_ = new_n20846_ & new_n20844_ & new_n20845_ & new_n20847_;
  assign new_n16738_ = new_n20850_ & new_n20848_ & new_n20849_ & new_n20851_;
  assign new_n16739_ = new_n20675_ & new_n16572_ & new_n16464_;
  assign new_n16740_ = new_n17581_ & new_n17641_ & new_n15786_;
  assign new_n16741_ = new_n17661_ & new_n17659_ & new_n17660_ & new_n17662_;
  assign new_n16742_ = new_n17665_ & new_n17663_ & new_n17664_ & new_n17666_;
  assign new_n16743_ = new_n17669_ & new_n17667_ & new_n17668_ & new_n17670_;
  assign new_n16744_ = new_n17673_ & new_n17671_ & new_n17672_ & new_n17674_;
  assign new_n16745_ = new_n17644_ & new_n17642_ & new_n17643_ & new_n17645_;
  assign new_n16746_ = new_n17648_ & new_n17646_ & new_n17647_ & new_n17649_;
  assign new_n16747_ = new_n17652_ & new_n17650_ & new_n17651_ & new_n17653_;
  assign new_n16748_ = new_n17656_ & new_n17654_ & new_n17655_ & new_n17657_;
  assign new_n16749_ = new_n17558_ & new_n17389_;
  assign new_n16750_ = new_n17599_ & new_n17597_ & new_n17598_ & new_n17600_;
  assign new_n16751_ = new_n17603_ & new_n17601_ & new_n17602_ & new_n17604_;
  assign new_n16752_ = new_n17607_ & new_n17605_ & new_n17606_ & new_n17608_;
  assign new_n16753_ = new_n17611_ & new_n17609_ & new_n17610_ & new_n17612_;
  assign new_n16754_ = new_n17584_ & new_n17582_ & new_n17583_ & new_n17585_;
  assign new_n16755_ = new_n17588_ & new_n17586_ & new_n17587_ & new_n17589_;
  assign new_n16756_ = new_n17592_ & new_n17590_ & new_n17591_ & new_n17593_;
  assign new_n16757_ = new_n17595_ & new_n17594_;
  assign new_n16758_ = new_n17580_ & new_n17352_;
  assign new_n16759_ = new_n17430_ & new_n16464_;
  assign new_n16760_ = new_n16464_ & new_n20675_ & new_n17581_ & new_n16465_;
  assign new_n16761_ = new_n17398_ & new_n16581_;
  assign new_n16762_ = pi1074 & new_n20784_;
  assign new_n16763_ = new_n17696_ & new_n16478_;
  assign new_n16764_ = new_n15608_ & new_n16438_;
  assign new_n16765_ = pi1073 & pi1076;
  assign new_n16766_ = new_n17427_ & new_n17422_;
  assign new_n16767_ = new_n16766_ & new_n17704_;
  assign new_n16768_ = new_n17405_ & new_n17733_ & new_n17734_;
  assign new_n16769_ = new_n17743_ & new_n17742_ & new_n17741_;
  assign new_n16770_ = new_n17748_ & new_n17747_ & new_n17746_;
  assign new_n16771_ = new_n17753_ & new_n17752_ & new_n17751_;
  assign new_n16772_ = new_n17758_ & new_n17757_ & new_n17756_;
  assign new_n16773_ = new_n17763_ & new_n17762_ & new_n17761_;
  assign new_n16774_ = new_n17768_ & new_n17767_ & new_n17766_;
  assign new_n16775_ = new_n17773_ & new_n17772_ & new_n17771_;
  assign new_n16776_ = new_n17778_ & new_n17777_ & new_n17776_;
  assign new_n16777_ = new_n17405_ & new_n17791_ & new_n17792_;
  assign new_n16778_ = new_n17801_ & new_n17800_ & new_n17799_;
  assign new_n16779_ = new_n17806_ & new_n17805_ & new_n17804_;
  assign new_n16780_ = new_n17811_ & new_n17810_ & new_n17809_;
  assign new_n16781_ = new_n17816_ & new_n17815_ & new_n17814_;
  assign new_n16782_ = new_n17821_ & new_n17820_ & new_n17819_;
  assign new_n16783_ = new_n17826_ & new_n17825_ & new_n17824_;
  assign new_n16784_ = new_n17831_ & new_n17830_ & new_n17829_;
  assign new_n16785_ = new_n17836_ & new_n17835_ & new_n17834_;
  assign new_n16786_ = new_n17405_ & new_n17850_ & new_n17851_;
  assign new_n16787_ = new_n17860_ & new_n17859_ & new_n17858_;
  assign new_n16788_ = new_n17865_ & new_n17864_ & new_n17863_;
  assign new_n16789_ = new_n17870_ & new_n17869_ & new_n17868_;
  assign new_n16790_ = new_n17875_ & new_n17874_ & new_n17873_;
  assign new_n16791_ = new_n17880_ & new_n17879_ & new_n17878_;
  assign new_n16792_ = new_n17885_ & new_n17884_ & new_n17883_;
  assign new_n16793_ = new_n17890_ & new_n17889_ & new_n17888_;
  assign new_n16794_ = new_n17895_ & new_n17894_ & new_n17893_;
  assign new_n16795_ = new_n17405_ & new_n17907_ & new_n17908_;
  assign new_n16796_ = new_n17917_ & new_n17916_ & new_n17915_;
  assign new_n16797_ = new_n17922_ & new_n17921_ & new_n17920_;
  assign new_n16798_ = new_n17927_ & new_n17926_ & new_n17925_;
  assign new_n16799_ = new_n17932_ & new_n17931_ & new_n17930_;
  assign new_n16800_ = new_n17937_ & new_n17936_ & new_n17935_;
  assign new_n16801_ = new_n17942_ & new_n17941_ & new_n17940_;
  assign new_n16802_ = new_n17947_ & new_n17946_ & new_n17945_;
  assign new_n16803_ = new_n17952_ & new_n17951_ & new_n17950_;
  assign new_n16804_ = new_n17405_ & new_n17965_ & new_n17966_;
  assign new_n16805_ = new_n17975_ & new_n17974_ & new_n17973_;
  assign new_n16806_ = new_n17980_ & new_n17979_ & new_n17978_;
  assign new_n16807_ = new_n17985_ & new_n17984_ & new_n17983_;
  assign new_n16808_ = new_n17990_ & new_n17989_ & new_n17988_;
  assign new_n16809_ = new_n17995_ & new_n17994_ & new_n17993_;
  assign new_n16810_ = new_n18000_ & new_n17999_ & new_n17998_;
  assign new_n16811_ = new_n18005_ & new_n18004_ & new_n18003_;
  assign new_n16812_ = new_n18010_ & new_n18009_ & new_n18008_;
  assign new_n16813_ = new_n17405_ & new_n18022_ & new_n18023_;
  assign new_n16814_ = new_n18032_ & new_n18031_ & new_n18030_;
  assign new_n16815_ = new_n18037_ & new_n18036_ & new_n18035_;
  assign new_n16816_ = new_n18042_ & new_n18041_ & new_n18040_;
  assign new_n16817_ = new_n18047_ & new_n18046_ & new_n18045_;
  assign new_n16818_ = new_n18052_ & new_n18051_ & new_n18050_;
  assign new_n16819_ = new_n18057_ & new_n18056_ & new_n18055_;
  assign new_n16820_ = new_n18062_ & new_n18061_ & new_n18060_;
  assign new_n16821_ = new_n18067_ & new_n18066_ & new_n18065_;
  assign new_n16822_ = new_n17405_ & new_n18080_ & new_n18081_;
  assign new_n16823_ = new_n18090_ & new_n18089_ & new_n18088_;
  assign new_n16824_ = new_n18095_ & new_n18094_ & new_n18093_;
  assign new_n16825_ = new_n18100_ & new_n18099_ & new_n18098_;
  assign new_n16826_ = new_n18105_ & new_n18104_ & new_n18103_;
  assign new_n16827_ = new_n18110_ & new_n18109_ & new_n18108_;
  assign new_n16828_ = new_n18115_ & new_n18114_ & new_n18113_;
  assign new_n16829_ = new_n18120_ & new_n18119_ & new_n18118_;
  assign new_n16830_ = new_n18125_ & new_n18124_ & new_n18123_;
  assign new_n16831_ = new_n17405_ & new_n18137_ & new_n18138_;
  assign new_n16832_ = new_n18147_ & new_n18146_ & new_n18145_;
  assign new_n16833_ = new_n18152_ & new_n18151_ & new_n18150_;
  assign new_n16834_ = new_n18157_ & new_n18156_ & new_n18155_;
  assign new_n16835_ = new_n18162_ & new_n18161_ & new_n18160_;
  assign new_n16836_ = new_n18167_ & new_n18166_ & new_n18165_;
  assign new_n16837_ = new_n18172_ & new_n18171_ & new_n18170_;
  assign new_n16838_ = new_n18177_ & new_n18176_ & new_n18175_;
  assign new_n16839_ = new_n18182_ & new_n18181_ & new_n18180_;
  assign new_n16840_ = new_n17405_ & new_n18193_ & new_n18194_;
  assign new_n16841_ = new_n18203_ & new_n18202_ & new_n18201_;
  assign new_n16842_ = new_n18208_ & new_n18207_ & new_n18206_;
  assign new_n16843_ = new_n18213_ & new_n18212_ & new_n18211_;
  assign new_n16844_ = new_n18218_ & new_n18217_ & new_n18216_;
  assign new_n16845_ = new_n18223_ & new_n18222_ & new_n18221_;
  assign new_n16846_ = new_n18228_ & new_n18227_ & new_n18226_;
  assign new_n16847_ = new_n18233_ & new_n18232_ & new_n18231_;
  assign new_n16848_ = new_n18238_ & new_n18237_ & new_n18236_;
  assign new_n16849_ = new_n17405_ & new_n18250_ & new_n18251_;
  assign new_n16850_ = new_n18260_ & new_n18259_ & new_n18258_;
  assign new_n16851_ = new_n18265_ & new_n18264_ & new_n18263_;
  assign new_n16852_ = new_n18270_ & new_n18269_ & new_n18268_;
  assign new_n16853_ = new_n18275_ & new_n18274_ & new_n18273_;
  assign new_n16854_ = new_n18280_ & new_n18279_ & new_n18278_;
  assign new_n16855_ = new_n18285_ & new_n18284_ & new_n18283_;
  assign new_n16856_ = new_n18290_ & new_n18289_ & new_n18288_;
  assign new_n16857_ = new_n18295_ & new_n18294_ & new_n18293_;
  assign new_n16858_ = new_n17405_ & new_n18308_ & new_n18309_;
  assign new_n16859_ = new_n18318_ & new_n18317_ & new_n18316_;
  assign new_n16860_ = new_n18323_ & new_n18322_ & new_n18321_;
  assign new_n16861_ = new_n18328_ & new_n18327_ & new_n18326_;
  assign new_n16862_ = new_n18333_ & new_n18332_ & new_n18331_;
  assign new_n16863_ = new_n18338_ & new_n18337_ & new_n18336_;
  assign new_n16864_ = new_n18343_ & new_n18342_ & new_n18341_;
  assign new_n16865_ = new_n18348_ & new_n18347_ & new_n18346_;
  assign new_n16866_ = new_n18353_ & new_n18352_ & new_n18351_;
  assign new_n16867_ = new_n17405_ & new_n18365_ & new_n18366_;
  assign new_n16868_ = new_n18375_ & new_n18374_ & new_n18373_;
  assign new_n16869_ = new_n18380_ & new_n18379_ & new_n18378_;
  assign new_n16870_ = new_n18385_ & new_n18384_ & new_n18383_;
  assign new_n16871_ = new_n18390_ & new_n18389_ & new_n18388_;
  assign new_n16872_ = new_n18395_ & new_n18394_ & new_n18393_;
  assign new_n16873_ = new_n18400_ & new_n18399_ & new_n18398_;
  assign new_n16874_ = new_n18405_ & new_n18404_ & new_n18403_;
  assign new_n16875_ = new_n18410_ & new_n18409_ & new_n18408_;
  assign new_n16876_ = new_n17405_ & new_n18423_ & new_n18424_;
  assign new_n16877_ = new_n18433_ & new_n18432_ & new_n18431_;
  assign new_n16878_ = new_n18438_ & new_n18437_ & new_n18436_;
  assign new_n16879_ = new_n18443_ & new_n18442_ & new_n18441_;
  assign new_n16880_ = new_n18448_ & new_n18447_ & new_n18446_;
  assign new_n16881_ = new_n18453_ & new_n18452_ & new_n18451_;
  assign new_n16882_ = new_n18458_ & new_n18457_ & new_n18456_;
  assign new_n16883_ = new_n18463_ & new_n18462_ & new_n18461_;
  assign new_n16884_ = new_n18468_ & new_n18467_ & new_n18466_;
  assign new_n16885_ = new_n17405_ & new_n18480_ & new_n18481_;
  assign new_n16886_ = new_n18490_ & new_n18489_ & new_n18488_;
  assign new_n16887_ = new_n18495_ & new_n18494_ & new_n18493_;
  assign new_n16888_ = new_n18500_ & new_n18499_ & new_n18498_;
  assign new_n16889_ = new_n18505_ & new_n18504_ & new_n18503_;
  assign new_n16890_ = new_n18510_ & new_n18509_ & new_n18508_;
  assign new_n16891_ = new_n18515_ & new_n18514_ & new_n18513_;
  assign new_n16892_ = new_n18520_ & new_n18519_ & new_n18518_;
  assign new_n16893_ = new_n18525_ & new_n18524_ & new_n18523_;
  assign new_n16894_ = new_n17405_ & new_n18538_ & new_n18539_;
  assign new_n16895_ = new_n18548_ & new_n18547_ & new_n18546_;
  assign new_n16896_ = new_n18553_ & new_n18552_ & new_n18551_;
  assign new_n16897_ = new_n18558_ & new_n18557_ & new_n18556_;
  assign new_n16898_ = new_n18563_ & new_n18562_ & new_n18561_;
  assign new_n16899_ = new_n18568_ & new_n18567_ & new_n18566_;
  assign new_n16900_ = new_n18573_ & new_n18572_ & new_n18571_;
  assign new_n16901_ = new_n18578_ & new_n18577_ & new_n18576_;
  assign new_n16902_ = new_n18583_ & new_n18582_ & new_n18581_;
  assign new_n16903_ = new_n17405_ & new_n18595_ & new_n18596_;
  assign new_n16904_ = new_n18605_ & new_n18604_ & new_n18603_;
  assign new_n16905_ = new_n18610_ & new_n18609_ & new_n18608_;
  assign new_n16906_ = new_n18615_ & new_n18614_ & new_n18613_;
  assign new_n16907_ = new_n18620_ & new_n18619_ & new_n18618_;
  assign new_n16908_ = new_n18624_ & new_n18623_ & new_n18622_;
  assign new_n16909_ = new_n18629_ & new_n18628_ & new_n18627_;
  assign new_n16910_ = new_n18634_ & new_n18633_ & new_n18632_;
  assign new_n16911_ = new_n18639_ & new_n18638_ & new_n18637_;
  assign new_n16912_ = pi1443 & pi1076;
  assign new_n16913_ = new_n17675_ & new_n17580_;
  assign new_n16914_ = new_n17678_ & new_n16438_;
  assign new_n16915_ = new_n17391_ & new_n16438_;
  assign new_n16916_ = new_n20677_ & new_n17398_;
  assign new_n16917_ = new_n18652_ & new_n18653_;
  assign new_n16918_ = new_n16917_ & new_n18651_;
  assign new_n16919_ = new_n16918_ & new_n15699_;
  assign new_n16920_ = new_n18656_ & new_n17423_;
  assign new_n16921_ = new_n18667_ & new_n18666_;
  assign new_n16922_ = new_n17630_ & new_n17581_;
  assign new_n16923_ = new_n18677_ & new_n16574_;
  assign new_n16924_ = new_n18679_ & new_n18678_;
  assign new_n16925_ = new_n20808_ & new_n16924_ & new_n16923_ & new_n18681_;
  assign new_n16926_ = new_n17444_ & new_n16578_;
  assign new_n16927_ = new_n16592_ & new_n16460_ & new_n15701_ & new_n16926_ & new_n16469_;
  assign new_n16928_ = new_n16929_ & new_n18683_;
  assign new_n16929_ = new_n18686_ & new_n18685_;
  assign new_n16930_ = new_n18694_ & new_n20898_ & new_n20897_;
  assign new_n16931_ = new_n18705_ & new_n18703_;
  assign new_n16932_ = new_n18724_ & new_n18725_;
  assign new_n16933_ = new_n18728_ & new_n18729_;
  assign new_n16934_ = new_n18733_ & new_n18734_;
  assign new_n16935_ = new_n18739_ & new_n16438_;
  assign new_n16936_ = new_n16465_ & new_n16588_;
  assign new_n16937_ = new_n18744_ & new_n18742_;
  assign new_n16938_ = new_n18748_ & new_n16579_ & new_n16580_;
  assign new_n16939_ = new_n16938_ & new_n15701_ & new_n18749_;
  assign new_n16940_ = new_n17367_ & new_n16465_;
  assign new_n16941_ = new_n16629_ & new_n16469_ & new_n17398_;
  assign new_n16942_ = new_n18747_ & new_n20688_;
  assign new_n16943_ = new_n20689_ & pi1074;
  assign new_n16944_ = new_n18752_ & new_n18751_;
  assign new_n16945_ = new_n18754_ & new_n18753_;
  assign new_n16946_ = new_n18756_ & new_n18757_;
  assign new_n16947_ = new_n16946_ & new_n18755_;
  assign new_n16948_ = new_n18759_ & new_n18758_;
  assign new_n16949_ = new_n18761_ & new_n18760_;
  assign new_n16950_ = new_n18763_ & new_n18764_;
  assign new_n16951_ = new_n16950_ & new_n18762_;
  assign new_n16952_ = new_n18766_ & new_n18765_;
  assign new_n16953_ = new_n18768_ & new_n18767_;
  assign new_n16954_ = new_n18770_ & new_n18771_;
  assign new_n16955_ = new_n16954_ & new_n18769_;
  assign new_n16956_ = new_n18775_ & new_n18773_ & new_n18772_;
  assign new_n16957_ = new_n18774_ & new_n16958_ & new_n18776_;
  assign new_n16958_ = new_n18777_ & new_n18778_;
  assign new_n16959_ = new_n18782_ & new_n18780_ & new_n18779_;
  assign new_n16960_ = new_n18784_ & new_n18785_;
  assign new_n16961_ = new_n16960_ & new_n18783_;
  assign new_n16962_ = new_n18789_ & new_n18787_ & new_n18786_;
  assign new_n16963_ = new_n18791_ & new_n18792_;
  assign new_n16964_ = new_n16963_ & new_n18790_;
  assign new_n16965_ = new_n18796_ & new_n18794_ & new_n18793_;
  assign new_n16966_ = new_n18798_ & new_n18799_;
  assign new_n16967_ = new_n16966_ & new_n18797_;
  assign new_n16968_ = new_n18803_ & new_n18801_ & new_n18800_;
  assign new_n16969_ = new_n18805_ & new_n18806_;
  assign new_n16970_ = new_n16969_ & new_n18804_;
  assign new_n16971_ = new_n18810_ & new_n18808_ & new_n18807_;
  assign new_n16972_ = new_n18812_ & new_n18813_;
  assign new_n16973_ = new_n16972_ & new_n18811_;
  assign new_n16974_ = new_n18817_ & new_n18815_ & new_n18814_;
  assign new_n16975_ = new_n18819_ & new_n18820_;
  assign new_n16976_ = new_n16975_ & new_n18818_;
  assign new_n16977_ = new_n18824_ & new_n18822_ & new_n18821_;
  assign new_n16978_ = new_n18826_ & new_n18827_;
  assign new_n16979_ = new_n16978_ & new_n18825_;
  assign new_n16980_ = new_n18831_ & new_n18829_ & new_n18828_;
  assign new_n16981_ = new_n18833_ & new_n18834_;
  assign new_n16982_ = new_n16981_ & new_n18832_;
  assign new_n16983_ = new_n18838_ & new_n18836_ & new_n18835_;
  assign new_n16984_ = new_n18840_ & new_n18841_;
  assign new_n16985_ = new_n16984_ & new_n18839_;
  assign new_n16986_ = new_n18843_ & new_n18845_;
  assign new_n16987_ = new_n18847_ & new_n18848_;
  assign new_n16988_ = new_n16987_ & new_n18846_;
  assign new_n16989_ = new_n18850_ & new_n18852_;
  assign new_n16990_ = new_n18854_ & new_n18855_;
  assign new_n16991_ = new_n16990_ & new_n18853_;
  assign new_n16992_ = new_n18857_ & new_n18859_;
  assign new_n16993_ = new_n18861_ & new_n18862_;
  assign new_n16994_ = new_n16993_ & new_n18860_;
  assign new_n16995_ = new_n18864_ & new_n18866_;
  assign new_n16996_ = new_n18868_ & new_n18869_;
  assign new_n16997_ = new_n16996_ & new_n18867_;
  assign new_n16998_ = new_n18871_ & new_n18873_;
  assign new_n16999_ = new_n18875_ & new_n18876_;
  assign new_n17000_ = new_n16999_ & new_n18874_;
  assign new_n17001_ = new_n18878_ & new_n18880_;
  assign new_n17002_ = new_n18882_ & new_n18883_;
  assign new_n17003_ = new_n17002_ & new_n18881_;
  assign new_n17004_ = new_n18885_ & new_n18887_;
  assign new_n17005_ = new_n18889_ & new_n18890_;
  assign new_n17006_ = new_n17005_ & new_n18888_;
  assign new_n17007_ = new_n18892_ & new_n18894_;
  assign new_n17008_ = new_n18896_ & new_n18897_;
  assign new_n17009_ = new_n17008_ & new_n18895_;
  assign new_n17010_ = new_n18899_ & new_n18901_;
  assign new_n17011_ = new_n18903_ & new_n18904_;
  assign new_n17012_ = new_n17011_ & new_n18902_;
  assign new_n17013_ = new_n18906_ & new_n18908_;
  assign new_n17014_ = new_n18910_ & new_n18911_;
  assign new_n17015_ = new_n17014_ & new_n18909_;
  assign new_n17016_ = new_n18913_ & new_n18915_;
  assign new_n17017_ = new_n18917_ & new_n18918_;
  assign new_n17018_ = new_n17017_ & new_n18916_;
  assign new_n17019_ = new_n18920_ & new_n18922_;
  assign new_n17020_ = new_n18924_ & new_n18925_;
  assign new_n17021_ = new_n17020_ & new_n18923_;
  assign new_n17022_ = new_n18927_ & new_n18929_;
  assign new_n17023_ = new_n18931_ & new_n18932_;
  assign new_n17024_ = new_n17023_ & new_n18930_;
  assign new_n17025_ = new_n18934_ & new_n18936_;
  assign new_n17026_ = new_n18938_ & new_n18939_;
  assign new_n17027_ = new_n17026_ & new_n18937_;
  assign new_n17028_ = new_n18941_ & new_n18943_;
  assign new_n17029_ = new_n18945_ & new_n18946_;
  assign new_n17030_ = new_n17029_ & new_n18944_;
  assign new_n17031_ = new_n18948_ & new_n18950_;
  assign new_n17032_ = new_n18952_ & new_n18953_;
  assign new_n17033_ = new_n17032_ & new_n18951_;
  assign new_n17034_ = new_n18955_ & new_n18957_;
  assign new_n17035_ = new_n18959_ & new_n18960_;
  assign new_n17036_ = new_n17035_ & new_n18958_;
  assign new_n17037_ = new_n18962_ & new_n18964_;
  assign new_n17038_ = new_n18966_ & new_n18967_;
  assign new_n17039_ = new_n17038_ & new_n18965_;
  assign new_n17040_ = new_n18969_ & new_n18971_;
  assign new_n17041_ = new_n18973_ & new_n18974_;
  assign new_n17042_ = new_n17041_ & new_n18972_;
  assign new_n17043_ = new_n20675_ & new_n16464_ & new_n16443_;
  assign new_n17044_ = new_n18975_ & new_n16589_;
  assign new_n17045_ = pi1075 & pi1445;
  assign new_n17046_ = new_n15549_ & new_n16465_;
  assign new_n17047_ = new_n15630_ & pi1076;
  assign new_n17048_ = new_n17389_ & new_n15549_;
  assign new_n17049_ = new_n19286_ & new_n19287_;
  assign new_n17050_ = new_n19289_ & new_n19290_;
  assign new_n17051_ = new_n19292_ & new_n19293_;
  assign new_n17052_ = new_n19295_ & new_n19296_;
  assign new_n17053_ = new_n19298_ & new_n19299_;
  assign new_n17054_ = new_n19301_ & new_n19302_;
  assign new_n17055_ = new_n19304_ & new_n19305_;
  assign new_n17056_ = new_n19307_ & new_n19308_;
  assign new_n17057_ = new_n19310_ & new_n19311_;
  assign new_n17058_ = new_n19313_ & new_n19314_;
  assign new_n17059_ = new_n19316_ & new_n19317_;
  assign new_n17060_ = new_n19319_ & new_n19320_;
  assign new_n17061_ = new_n19322_ & new_n19323_;
  assign new_n17062_ = new_n19325_ & new_n19326_;
  assign new_n17063_ = new_n19328_ & new_n19329_;
  assign new_n17064_ = new_n19332_ & new_n19331_;
  assign new_n17065_ = new_n15786_ & new_n16572_;
  assign new_n17066_ = new_n20675_ & pi1076 & new_n16452_;
  assign new_n17067_ = new_n17580_ & new_n17352_;
  assign new_n17068_ = new_n19543_ & new_n17422_ & new_n17425_;
  assign new_n17069_ = ~new_n2972_ & ~pi1445;
  assign new_n17070_ = new_n17675_ & new_n17367_;
  assign new_n17071_ = new_n19554_ & new_n19552_ & new_n19555_ & new_n19556_ & new_n19553_;
  assign new_n17072_ = new_n19562_ & new_n19560_ & new_n19563_ & new_n19564_ & new_n19561_;
  assign new_n17073_ = new_n19570_ & new_n19568_ & new_n19571_ & new_n19572_ & new_n19569_;
  assign new_n17074_ = new_n19578_ & new_n19576_ & new_n19579_ & new_n19580_ & new_n19577_;
  assign new_n17075_ = new_n19581_ & new_n17408_;
  assign new_n17076_ = new_n19585_ & new_n19587_ & new_n19588_ & new_n19586_;
  assign new_n17077_ = new_n19589_ & new_n17408_;
  assign new_n17078_ = new_n19594_ & new_n19592_ & new_n19595_ & new_n19596_ & new_n19593_;
  assign new_n17079_ = new_n19597_ & new_n17408_;
  assign new_n17080_ = new_n19602_ & new_n19603_ & new_n19600_;
  assign new_n17081_ = new_n19604_ & new_n17408_;
  assign new_n17082_ = new_n19609_ & new_n19610_ & new_n19607_;
  assign new_n17083_ = new_n19611_ & new_n17408_;
  assign new_n17084_ = new_n19616_ & new_n19617_ & new_n19614_;
  assign new_n17085_ = new_n19618_ & new_n17408_;
  assign new_n17086_ = new_n19623_ & new_n19624_ & new_n19621_;
  assign new_n17087_ = new_n19625_ & new_n17408_;
  assign new_n17088_ = new_n19630_ & new_n19631_ & new_n19628_;
  assign new_n17089_ = new_n19632_ & new_n17408_;
  assign new_n17090_ = new_n19637_ & new_n19638_ & new_n19635_;
  assign new_n17091_ = new_n19639_ & new_n17408_;
  assign new_n17092_ = new_n19644_ & new_n19645_ & new_n19642_;
  assign new_n17093_ = new_n19646_ & new_n17408_;
  assign new_n17094_ = new_n19651_ & new_n19652_ & new_n19649_;
  assign new_n17095_ = new_n19653_ & new_n17408_;
  assign new_n17096_ = new_n19658_ & new_n19659_ & new_n19656_;
  assign new_n17097_ = new_n19660_ & new_n17408_;
  assign new_n17098_ = new_n19665_ & new_n19666_ & new_n19663_;
  assign new_n17099_ = new_n19667_ & new_n17408_;
  assign new_n17100_ = new_n19672_ & new_n19673_ & new_n19670_;
  assign new_n17101_ = new_n17408_ & new_n19675_;
  assign new_n17102_ = new_n19679_ & new_n19680_ & new_n19677_;
  assign new_n17103_ = new_n17408_ & new_n19682_;
  assign new_n17104_ = new_n19686_ & new_n19687_ & new_n19684_;
  assign new_n17105_ = new_n17408_ & new_n19689_;
  assign new_n17106_ = new_n19693_ & new_n19694_ & new_n19691_;
  assign new_n17107_ = new_n19698_ & new_n19696_;
  assign new_n17108_ = new_n19700_ & new_n19701_;
  assign new_n17109_ = new_n19705_ & new_n19703_;
  assign new_n17110_ = new_n19707_ & new_n19708_;
  assign new_n17111_ = new_n19712_ & new_n19710_;
  assign new_n17112_ = new_n19714_ & new_n19715_;
  assign new_n17113_ = new_n19719_ & new_n19717_;
  assign new_n17114_ = new_n19721_ & new_n19722_;
  assign new_n17115_ = new_n19726_ & new_n19724_;
  assign new_n17116_ = new_n19728_ & new_n19729_;
  assign new_n17117_ = new_n19733_ & new_n19731_;
  assign new_n17118_ = new_n19735_ & new_n19736_;
  assign new_n17119_ = new_n19740_ & new_n19738_;
  assign new_n17120_ = new_n19742_ & new_n19743_;
  assign new_n17121_ = new_n19747_ & new_n19745_;
  assign new_n17122_ = new_n19749_ & new_n19750_;
  assign new_n17123_ = new_n19754_ & new_n19752_;
  assign new_n17124_ = new_n19756_ & new_n19757_;
  assign new_n17125_ = new_n19761_ & new_n19759_;
  assign new_n17126_ = new_n19763_ & new_n19764_;
  assign new_n17127_ = new_n19768_ & new_n19766_;
  assign new_n17128_ = new_n19770_ & new_n19771_;
  assign new_n17129_ = new_n19775_ & new_n19773_;
  assign new_n17130_ = new_n19777_ & new_n19778_;
  assign new_n17131_ = ~pi1044 & ~pi1043 & ~pi1046 & ~pi1045;
  assign new_n17132_ = ~pi1048 & ~pi1047 & ~pi1050 & ~pi1049;
  assign new_n17133_ = new_n17132_ & new_n17131_;
  assign new_n17134_ = ~pi1052 & ~pi1051 & ~pi1054 & ~pi1053;
  assign new_n17135_ = ~pi1056 & ~pi1055 & ~pi1058 & ~pi1057;
  assign new_n17136_ = new_n17135_ & new_n17134_;
  assign new_n17137_ = ~pi1060 & ~pi1059 & ~pi1062 & ~pi1061;
  assign new_n17138_ = ~pi1064 & ~pi1063 & ~pi1066 & ~pi1065;
  assign new_n17139_ = new_n17138_ & new_n17137_;
  assign new_n17140_ = ~pi1067 & ~pi1068;
  assign new_n17141_ = ~pi1069 & ~pi1070;
  assign new_n17142_ = ~pi1071 & ~pi1072;
  assign new_n17143_ = new_n19779_ & new_n17140_ & new_n17141_ & new_n17142_;
  assign new_n17144_ = ~pi1041 & ~pi1042 & ~pi1406;
  assign new_n17145_ = pi1074 & new_n16438_;
  assign new_n17146_ = new_n19789_ & new_n16479_;
  assign new_n17147_ = ~new_n2972_ & ~pi1076;
  assign new_n17148_ = new_n19783_ & new_n16488_ & new_n16589_;
  assign new_n17149_ = pi1074 & new_n16468_;
  assign new_n17150_ = new_n17416_ & new_n17387_;
  assign new_n17151_ = new_n19801_ & new_n19799_ & new_n19800_ & new_n19802_;
  assign new_n17152_ = new_n19805_ & new_n19803_ & new_n19804_ & new_n19806_;
  assign new_n17153_ = new_n19809_ & new_n19807_ & new_n19808_ & new_n19810_;
  assign new_n17154_ = new_n19813_ & new_n19811_ & new_n19812_ & new_n19814_;
  assign new_n17155_ = new_n19817_ & new_n19815_ & new_n19816_ & new_n19818_;
  assign new_n17156_ = new_n19821_ & new_n19819_ & new_n19820_ & new_n19822_;
  assign new_n17157_ = new_n19825_ & new_n19823_ & new_n19824_ & new_n19826_;
  assign new_n17158_ = new_n19829_ & new_n19827_ & new_n19828_ & new_n19830_;
  assign new_n17159_ = new_n19833_ & new_n19831_ & new_n19832_ & new_n19834_;
  assign new_n17160_ = new_n19837_ & new_n19835_ & new_n19836_ & new_n19838_;
  assign new_n17161_ = new_n19841_ & new_n19839_ & new_n19840_ & new_n19842_;
  assign new_n17162_ = new_n19845_ & new_n19843_ & new_n19844_ & new_n19846_;
  assign new_n17163_ = new_n19849_ & new_n19847_ & new_n19848_ & new_n19850_;
  assign new_n17164_ = new_n19853_ & new_n19851_ & new_n19852_ & new_n19854_;
  assign new_n17165_ = new_n19857_ & new_n19855_ & new_n19856_ & new_n19858_;
  assign new_n17166_ = new_n19861_ & new_n19859_ & new_n19860_ & new_n20794_;
  assign new_n17167_ = new_n19864_ & new_n19862_ & new_n19863_ & new_n19865_;
  assign new_n17168_ = new_n19868_ & new_n19866_ & new_n19867_ & new_n19869_;
  assign new_n17169_ = new_n19872_ & new_n19870_ & new_n19871_ & new_n19873_;
  assign new_n17170_ = new_n19876_ & new_n19874_ & new_n19875_ & new_n19877_;
  assign new_n17171_ = new_n19880_ & new_n19878_ & new_n19879_ & new_n19881_;
  assign new_n17172_ = new_n19884_ & new_n19882_ & new_n19883_ & new_n19885_;
  assign new_n17173_ = new_n19888_ & new_n19886_ & new_n19887_ & new_n19889_;
  assign new_n17174_ = new_n19892_ & new_n19890_ & new_n19891_ & new_n19893_;
  assign new_n17175_ = new_n19896_ & new_n19894_ & new_n19895_ & new_n19897_;
  assign new_n17176_ = new_n19900_ & new_n19898_ & new_n19899_ & new_n19901_;
  assign new_n17177_ = new_n19904_ & new_n19902_ & new_n19903_ & new_n19905_;
  assign new_n17178_ = new_n19908_ & new_n19906_ & new_n19907_ & new_n19909_;
  assign new_n17179_ = new_n19912_ & new_n19910_ & new_n19911_ & new_n19913_;
  assign new_n17180_ = new_n19916_ & new_n19914_ & new_n19915_ & new_n19917_;
  assign new_n17181_ = new_n19920_ & new_n19918_ & new_n19919_ & new_n19921_;
  assign new_n17182_ = new_n19924_ & new_n19922_ & new_n19923_ & new_n19925_;
  assign new_n17183_ = new_n19930_ & new_n19929_;
  assign new_n17184_ = new_n19933_ & new_n19932_;
  assign new_n17185_ = new_n19936_ & new_n19935_;
  assign new_n17186_ = new_n19939_ & new_n19938_;
  assign new_n17187_ = new_n19941_ & new_n17188_;
  assign new_n17188_ = new_n19943_ & new_n19942_;
  assign new_n17189_ = new_n19945_ & new_n19946_;
  assign new_n17190_ = new_n19955_ & new_n19953_ & new_n19954_;
  assign new_n17191_ = new_n19957_ & new_n19958_;
  assign new_n17192_ = new_n19964_ & new_n19962_ & new_n19963_;
  assign new_n17193_ = new_n19968_ & new_n19966_ & new_n19967_;
  assign new_n17194_ = new_n19972_ & new_n19970_ & new_n19971_;
  assign new_n17195_ = new_n19976_ & new_n19974_ & new_n19975_;
  assign new_n17196_ = new_n19980_ & new_n19978_ & new_n19979_;
  assign new_n17197_ = new_n19984_ & new_n19982_ & new_n19983_;
  assign new_n17198_ = new_n19988_ & new_n19986_ & new_n19987_;
  assign new_n17199_ = new_n19992_ & new_n19990_ & new_n19991_;
  assign new_n17200_ = new_n19996_ & new_n19994_ & new_n19995_;
  assign new_n17201_ = new_n20000_ & new_n19998_ & new_n19999_;
  assign new_n17202_ = new_n20002_ & new_n20003_;
  assign new_n17203_ = new_n20009_ & new_n20007_ & new_n20008_;
  assign new_n17204_ = new_n20013_ & new_n20011_ & new_n20012_;
  assign new_n17205_ = new_n20017_ & new_n20015_ & new_n20016_;
  assign new_n17206_ = new_n20021_ & new_n20019_ & new_n20020_;
  assign new_n17207_ = new_n20039_ & new_n20038_;
  assign new_n17208_ = new_n20041_ & new_n20042_;
  assign new_n17209_ = new_n16464_ & new_n20675_ & new_n20069_;
  assign new_n17210_ = new_n20075_ & new_n20073_ & new_n20074_ & new_n20076_;
  assign new_n17211_ = new_n20079_ & new_n20077_ & new_n20078_ & new_n20080_;
  assign new_n17212_ = new_n20083_ & new_n20081_ & new_n20082_ & new_n20084_;
  assign new_n17213_ = new_n20087_ & new_n20085_ & new_n20086_ & new_n20088_;
  assign new_n17214_ = new_n20093_ & new_n20091_ & new_n20092_ & new_n20094_;
  assign new_n17215_ = new_n20097_ & new_n20095_ & new_n20096_ & new_n20098_;
  assign new_n17216_ = new_n20101_ & new_n20099_ & new_n20100_ & new_n20102_;
  assign new_n17217_ = new_n20105_ & new_n20103_ & new_n20104_ & new_n20106_;
  assign new_n17218_ = new_n20124_ & new_n20122_ & new_n20123_ & new_n20125_;
  assign new_n17219_ = new_n20128_ & new_n20126_ & new_n20127_ & new_n20129_;
  assign new_n17220_ = new_n20132_ & new_n20130_ & new_n20131_ & new_n20133_;
  assign new_n17221_ = new_n20136_ & new_n20134_ & new_n20135_ & new_n20137_;
  assign new_n17222_ = new_n20141_ & new_n20139_ & new_n20140_ & new_n20142_;
  assign new_n17223_ = new_n20145_ & new_n20143_ & new_n20144_ & new_n20146_;
  assign new_n17224_ = new_n20149_ & new_n20147_ & new_n20148_ & new_n20150_;
  assign new_n17225_ = new_n20153_ & new_n20151_ & new_n20152_ & new_n20154_;
  assign new_n17226_ = new_n20158_ & new_n20156_ & new_n20157_ & new_n20159_;
  assign new_n17227_ = new_n20162_ & new_n20160_ & new_n20161_ & new_n20163_;
  assign new_n17228_ = new_n20166_ & new_n20164_ & new_n20165_ & new_n20167_;
  assign new_n17229_ = new_n20170_ & new_n20168_ & new_n20169_ & new_n20171_;
  assign new_n17230_ = new_n20175_ & new_n20173_ & new_n20174_ & new_n20176_;
  assign new_n17231_ = new_n20179_ & new_n20177_ & new_n20178_ & new_n20180_;
  assign new_n17232_ = new_n20183_ & new_n20181_ & new_n20182_ & new_n20184_;
  assign new_n17233_ = new_n20187_ & new_n20185_ & new_n20186_ & new_n20795_;
  assign new_n17234_ = new_n20190_ & new_n20188_ & new_n20189_ & new_n20191_;
  assign new_n17235_ = new_n20194_ & new_n20192_ & new_n20193_ & new_n20195_;
  assign new_n17236_ = new_n20198_ & new_n20196_ & new_n20197_ & new_n20199_;
  assign new_n17237_ = new_n20202_ & new_n20200_ & new_n20201_ & new_n20203_;
  assign new_n17238_ = new_n20207_ & new_n20205_ & new_n20206_ & new_n20208_;
  assign new_n17239_ = new_n20211_ & new_n20209_ & new_n20210_ & new_n20212_;
  assign new_n17240_ = new_n20215_ & new_n20213_ & new_n20214_ & new_n20216_;
  assign new_n17241_ = new_n20219_ & new_n20217_ & new_n20218_ & new_n20220_;
  assign new_n17242_ = new_n20240_ & new_n16624_;
  assign new_n17243_ = pi1076 & new_n20243_;
  assign new_n17244_ = new_n20249_ & new_n20247_ & new_n20248_ & new_n20250_;
  assign new_n17245_ = new_n20253_ & new_n20251_ & new_n20252_ & new_n20254_;
  assign new_n17246_ = new_n20257_ & new_n20255_ & new_n20256_ & new_n20258_;
  assign new_n17247_ = new_n20261_ & new_n20259_ & new_n20260_ & new_n20262_;
  assign new_n17248_ = new_n17437_ & pi1076;
  assign new_n17249_ = new_n17585_ & new_n17582_ & new_n17584_ & new_n17586_;
  assign new_n17250_ = new_n17589_ & new_n17588_ & new_n17587_;
  assign new_n17251_ = new_n17592_ & new_n17590_ & new_n17591_ & new_n17593_;
  assign new_n17252_ = new_n17595_ & new_n17594_;
  assign new_n17253_ = new_n17581_ & new_n16572_;
  assign new_n17254_ = pi1076 & new_n16465_;
  assign new_n17255_ = new_n20271_ & new_n20270_;
  assign new_n17256_ = new_n20654_ & new_n20653_ & new_n16615_;
  assign new_n17257_ = new_n20655_ & new_n20656_ & new_n20657_;
  assign new_n17258_ = new_n17257_ & new_n15787_ & new_n20658_;
  assign new_n17259_ = new_n20278_ & new_n20276_;
  assign new_n17260_ = new_n20281_ & new_n20279_ & new_n20280_ & new_n20282_;
  assign new_n17261_ = new_n20285_ & new_n20283_ & new_n20284_ & new_n20286_;
  assign new_n17262_ = new_n20289_ & new_n20287_ & new_n20288_ & new_n20290_;
  assign new_n17263_ = new_n20293_ & new_n20291_ & new_n20292_ & new_n20294_;
  assign new_n17264_ = new_n20298_ & new_n20296_ & new_n20297_ & new_n20299_;
  assign new_n17265_ = new_n20302_ & new_n20300_ & new_n20301_ & new_n20303_;
  assign new_n17266_ = new_n20306_ & new_n20304_ & new_n20305_ & new_n20307_;
  assign new_n17267_ = new_n20310_ & new_n20308_ & new_n20309_ & new_n20311_;
  assign new_n17268_ = new_n20315_ & new_n20313_ & new_n20314_ & new_n20316_;
  assign new_n17269_ = new_n20319_ & new_n20317_ & new_n20318_ & new_n20320_;
  assign new_n17270_ = new_n20323_ & new_n20321_ & new_n20322_ & new_n20324_;
  assign new_n17271_ = new_n20326_ & new_n20325_;
  assign new_n17272_ = new_n17271_ & new_n20798_ & new_n20327_;
  assign new_n17273_ = new_n20330_ & new_n20328_ & new_n20329_ & new_n20331_;
  assign new_n17274_ = new_n20334_ & new_n20332_ & new_n20333_ & new_n20335_;
  assign new_n17275_ = new_n20338_ & new_n20336_ & new_n20337_ & new_n20339_;
  assign new_n17276_ = new_n20342_ & new_n20340_ & new_n20341_ & new_n20343_;
  assign new_n17277_ = new_n20347_ & new_n20345_ & new_n20346_ & new_n20348_;
  assign new_n17278_ = new_n20351_ & new_n20349_ & new_n20350_ & new_n20352_;
  assign new_n17279_ = new_n20355_ & new_n20353_ & new_n20354_ & new_n20356_;
  assign new_n17280_ = new_n20359_ & new_n20357_ & new_n20358_ & new_n20360_;
  assign new_n17281_ = new_n20364_ & new_n20362_ & new_n20363_ & new_n20365_;
  assign new_n17282_ = new_n20368_ & new_n20366_ & new_n20367_ & new_n20369_;
  assign new_n17283_ = new_n20372_ & new_n20370_ & new_n20371_ & new_n20373_;
  assign new_n17284_ = new_n20376_ & new_n20374_ & new_n20375_ & new_n20377_;
  assign new_n17285_ = new_n20381_ & new_n20379_ & new_n20380_ & new_n20382_;
  assign new_n17286_ = new_n20385_ & new_n20383_ & new_n20384_ & new_n20386_;
  assign new_n17287_ = new_n20389_ & new_n20387_ & new_n20388_ & new_n20390_;
  assign new_n17288_ = new_n20393_ & new_n20391_ & new_n20392_ & new_n20394_;
  assign new_n17289_ = new_n20396_ & new_n16445_;
  assign new_n17290_ = new_n20397_ & new_n20396_;
  assign new_n17291_ = new_n20398_ & new_n16446_;
  assign new_n17292_ = new_n20270_ & new_n16608_;
  assign new_n17293_ = new_n20399_ & new_n20398_;
  assign new_n17294_ = new_n20654_ & new_n17293_ & new_n20653_;
  assign new_n17295_ = new_n16615_ & new_n17294_ & new_n17292_ & new_n20271_;
  assign new_n17296_ = new_n20661_ & new_n20655_ & new_n20657_ & new_n20667_;
  assign new_n17297_ = new_n20670_ & new_n20668_ & new_n20669_ & new_n20686_;
  assign new_n17298_ = new_n20271_ & new_n20270_;
  assign new_n17299_ = new_n20654_ & new_n20653_ & new_n16615_;
  assign new_n17300_ = new_n20655_ & new_n20656_ & new_n20657_;
  assign new_n17301_ = new_n20658_ & new_n17300_ & new_n15787_ & new_n15789_;
  assign new_n17302_ = new_n20403_ & new_n20401_ & new_n20402_ & new_n20404_;
  assign new_n17303_ = new_n20407_ & new_n20405_ & new_n20406_ & new_n20408_;
  assign new_n17304_ = new_n20411_ & new_n20409_ & new_n20410_ & new_n20412_;
  assign new_n17305_ = new_n20415_ & new_n20413_ & new_n20414_ & new_n20416_;
  assign new_n17306_ = new_n20420_ & new_n20418_ & new_n20419_ & new_n20421_;
  assign new_n17307_ = new_n20424_ & new_n20422_ & new_n20423_ & new_n20425_;
  assign new_n17308_ = new_n20428_ & new_n20426_ & new_n20427_ & new_n20429_;
  assign new_n17309_ = new_n20432_ & new_n20430_ & new_n20431_ & new_n20433_;
  assign new_n17310_ = new_n20437_ & new_n20435_ & new_n20436_ & new_n20438_;
  assign new_n17311_ = new_n20441_ & new_n20439_ & new_n20440_ & new_n20442_;
  assign new_n17312_ = new_n20445_ & new_n20443_ & new_n20444_ & new_n20446_;
  assign new_n17313_ = new_n20449_ & new_n20447_ & new_n20448_ & new_n20450_;
  assign new_n17314_ = new_n20454_ & new_n20452_ & new_n20453_ & new_n20455_;
  assign new_n17315_ = new_n20458_ & new_n20456_ & new_n20457_ & new_n20459_;
  assign new_n17316_ = new_n20462_ & new_n20460_ & new_n20461_ & new_n20463_;
  assign new_n17317_ = new_n20466_ & new_n20464_ & new_n20465_ & new_n20800_;
  assign new_n17318_ = new_n20469_ & new_n20467_ & new_n20468_ & new_n20470_;
  assign new_n17319_ = new_n20473_ & new_n20471_ & new_n20472_ & new_n20474_;
  assign new_n17320_ = new_n20477_ & new_n20475_ & new_n20476_ & new_n20478_;
  assign new_n17321_ = new_n20481_ & new_n20479_ & new_n20480_ & new_n20482_;
  assign new_n17322_ = new_n20486_ & new_n20484_ & new_n20485_ & new_n20487_;
  assign new_n17323_ = new_n20490_ & new_n20488_ & new_n20489_ & new_n20491_;
  assign new_n17324_ = new_n20494_ & new_n20492_ & new_n20493_ & new_n20495_;
  assign new_n17325_ = new_n20498_ & new_n20496_ & new_n20497_ & new_n20499_;
  assign new_n17326_ = new_n20503_ & new_n20501_ & new_n20502_ & new_n20504_;
  assign new_n17327_ = new_n20507_ & new_n20505_ & new_n20506_ & new_n20508_;
  assign new_n17328_ = new_n20511_ & new_n20509_ & new_n20510_ & new_n20512_;
  assign new_n17329_ = new_n20515_ & new_n20513_ & new_n20514_ & new_n20516_;
  assign new_n17330_ = new_n20520_ & new_n20518_ & new_n20519_ & new_n20521_;
  assign new_n17331_ = new_n20524_ & new_n20522_ & new_n20523_ & new_n20525_;
  assign new_n17332_ = new_n20528_ & new_n20526_ & new_n20527_ & new_n20529_;
  assign new_n17333_ = new_n20532_ & new_n20530_ & new_n20531_ & new_n20533_;
  assign new_n17334_ = new_n16465_ & new_n16600_;
  assign new_n17335_ = new_n16464_ & new_n16572_;
  assign new_n17336_ = new_n17444_ & new_n20538_ & new_n20539_;
  assign new_n17337_ = new_n17336_ & new_n20540_;
  assign new_n17338_ = pi1076 & new_n15608_;
  assign new_n17339_ = new_n17338_ & new_n20541_;
  assign new_n17340_ = new_n16452_ & new_n17354_;
  assign new_n17341_ = pi1076 & new_n17354_;
  assign new_n17342_ = new_n20550_ & pi1076;
  assign new_n17343_ = new_n20552_ & new_n15784_;
  assign new_n17344_ = new_n20554_ & pi1076;
  assign new_n17345_ = new_n20556_ & new_n15784_;
  assign new_n17346_ = new_n20563_ & new_n20564_;
  assign new_n17347_ = new_n16634_ & new_n20565_;
  assign new_n17348_ = new_n20568_ & new_n20570_ & new_n20569_;
  assign new_n17349_ = new_n20643_ & new_n20642_;
  assign new_n17350_ = new_n20646_ & new_n20645_;
  assign new_n17351_ = new_n20855_ & new_n20854_;
  assign new_n17352_ = ~new_n16752_ | ~new_n16750_ | ~new_n16751_ | ~new_n16753_;
  assign new_n17353_ = ~new_n16920_ | ~new_n18655_;
  assign new_n17354_ = ~new_n16757_ | ~new_n16754_ | ~new_n16755_ | ~new_n16756_ | ~new_n15788_;
  assign new_n17355_ = ~pi1246;
  assign new_n17356_ = new_n20907_ & new_n20906_;
  assign new_n17357_ = new_n20926_ & new_n20925_;
  assign new_n17358_ = ~new_n15549_ | ~new_n16466_;
  assign new_n17359_ = ~new_n17689_ | ~new_n16572_;
  assign new_n17360_ = ~pi0035;
  assign new_n17361_ = ~new_n17148_ | ~new_n17409_;
  assign new_n17362_ = ~new_n17409_ | ~new_n16613_;
  assign new_n17363_ = ~new_n16919_ | ~new_n20879_ | ~new_n20878_;
  assign new_n17364_ = ~pi1207 | ~new_n16450_;
  assign new_n17365_ = ~new_n16633_;
  assign new_n17366_ = ~pi0033 | ~new_n16438_;
  assign new_n17367_ = ~new_n16593_;
  assign new_n17368_ = ~new_n16621_;
  assign new_n17369_ = ~new_n16620_;
  assign new_n17370_ = ~new_n16574_;
  assign new_n17371_ = ~new_n16471_;
  assign new_n17372_ = ~new_n16630_;
  assign new_n17373_ = ~new_n16586_;
  assign new_n17374_ = ~new_n16615_;
  assign new_n17375_ = ~new_n16601_;
  assign new_n17376_ = ~new_n17446_ | ~new_n16452_;
  assign new_n17377_ = ~new_n17641_ | ~new_n15786_;
  assign new_n17378_ = ~new_n16577_;
  assign new_n17379_ = ~new_n16606_;
  assign new_n17380_ = ~new_n16470_;
  assign new_n17381_ = ~new_n16602_;
  assign new_n17382_ = ~new_n16603_;
  assign new_n17383_ = ~new_n16609_;
  assign new_n17384_ = ~new_n16589_;
  assign new_n17385_ = ~new_n16608_;
  assign new_n17386_ = ~new_n17378_ | ~new_n17066_ | ~new_n17370_;
  assign new_n17387_ = ~new_n16599_;
  assign new_n17388_ = ~new_n16624_;
  assign new_n17389_ = ~new_n16463_;
  assign new_n17390_ = ~new_n16488_;
  assign new_n17391_ = ~new_n16571_;
  assign new_n17392_ = ~new_n16627_;
  assign new_n17393_ = ~new_n16628_;
  assign new_n17394_ = ~new_n16629_;
  assign new_n17395_ = ~new_n16581_;
  assign new_n17396_ = ~new_n16469_;
  assign new_n17397_ = ~new_n16473_;
  assign new_n17398_ = ~new_n16759_ | ~new_n15612_;
  assign new_n17399_ = ~new_n16580_;
  assign new_n17400_ = ~new_n17630_ | ~new_n16452_;
  assign new_n17401_ = ~new_n16614_;
  assign new_n17402_ = ~new_n16430_;
  assign new_n17403_ = ~new_n16607_;
  assign new_n17404_ = ~new_n16605_;
  assign new_n17405_ = ~new_n16481_;
  assign new_n17406_ = ~new_n33286_;
  assign new_n17407_ = ~new_n16501_;
  assign new_n17408_ = ~new_n17436_ | ~new_n16612_;
  assign new_n17409_ = ~new_n17416_ | ~new_n20681_;
  assign new_n17410_ = ~new_n15543_ | ~new_n16453_;
  assign new_n17411_ = ~new_n15544_ | ~new_n17558_;
  assign new_n17412_ = ~new_n16588_;
  assign new_n17413_ = ~new_n16433_;
  assign new_n17414_ = ~new_n16431_;
  assign new_n17415_ = ~new_n16576_;
  assign new_n17416_ = ~new_n16478_;
  assign new_n17417_ = ~new_n16579_;
  assign new_n17418_ = ~new_n17359_;
  assign new_n17419_ = ~new_n16538_;
  assign new_n17420_ = ~new_n17658_ | ~new_n20562_;
  assign new_n17421_ = ~new_n17144_ | ~new_n17401_;
  assign new_n17422_ = ~new_n16765_ | ~new_n17442_;
  assign new_n17423_ = ~new_n16912_ | ~new_n15609_;
  assign new_n17424_ = ~new_n17545_ | ~new_n16439_;
  assign new_n17425_ = ~new_n15533_ | ~pi1075 | ~new_n16475_;
  assign new_n17426_ = ~new_n15609_ | ~new_n16584_;
  assign new_n17427_ = ~new_n2972_ | ~pi1076 | ~new_n16444_;
  assign new_n17428_ = ~new_n16575_;
  assign new_n17429_ = ~new_n15534_ | ~new_n15629_ | ~new_n17043_ | ~new_n15632_;
  assign new_n17430_ = ~new_n16468_;
  assign new_n17431_ = ~new_n16578_;
  assign new_n17432_ = ~new_n16596_;
  assign new_n17433_ = ~new_n16480_;
  assign new_n17434_ = ~new_n16590_;
  assign new_n17435_ = ~new_n16600_;
  assign new_n17436_ = ~new_n16613_;
  assign new_n17437_ = ~new_n16472_;
  assign new_n17438_ = ~new_n16570_;
  assign new_n17439_ = ~new_n16435_;
  assign new_n17440_ = ~new_n16462_;
  assign new_n17441_ = ~new_n16587_;
  assign new_n17442_ = ~new_n16479_;
  assign new_n17443_ = ~new_n16467_;
  assign new_n17444_ = ~new_n17417_ | ~new_n17580_;
  assign new_n17445_ = ~new_n16592_;
  assign new_n17446_ = ~new_n16634_;
  assign new_n17447_ = ~new_n16591_;
  assign new_n17448_ = ~pi1437 | ~new_n17414_;
  assign new_n17449_ = ~pi1436 | ~new_n17413_;
  assign new_n17450_ = ~pi1008 | ~new_n16430_;
  assign new_n17451_ = ~pi1436 | ~new_n17414_;
  assign new_n17452_ = ~pi1435 | ~new_n17413_;
  assign new_n17453_ = ~pi1009 | ~new_n16430_;
  assign new_n17454_ = ~pi1435 | ~new_n17414_;
  assign new_n17455_ = ~pi1434 | ~new_n17413_;
  assign new_n17456_ = ~pi1010 | ~new_n16430_;
  assign new_n17457_ = ~pi1434 | ~new_n17414_;
  assign new_n17458_ = ~pi1433 | ~new_n17413_;
  assign new_n17459_ = ~pi1011 | ~new_n16430_;
  assign new_n17460_ = ~pi1433 | ~new_n17414_;
  assign new_n17461_ = ~pi1432 | ~new_n17413_;
  assign new_n17462_ = ~pi1012 | ~new_n16430_;
  assign new_n17463_ = ~pi1432 | ~new_n17414_;
  assign new_n17464_ = ~pi1431 | ~new_n17413_;
  assign new_n17465_ = ~pi1013 | ~new_n16430_;
  assign new_n17466_ = ~pi1431 | ~new_n17414_;
  assign new_n17467_ = ~pi1430 | ~new_n17413_;
  assign new_n17468_ = ~pi1014 | ~new_n16430_;
  assign new_n17469_ = ~pi1430 | ~new_n17414_;
  assign new_n17470_ = ~pi1429 | ~new_n17413_;
  assign new_n17471_ = ~pi1015 | ~new_n16430_;
  assign new_n17472_ = ~pi1429 | ~new_n17414_;
  assign new_n17473_ = ~pi1428 | ~new_n17413_;
  assign new_n17474_ = ~pi1016 | ~new_n16430_;
  assign new_n17475_ = ~pi1428 | ~new_n17414_;
  assign new_n17476_ = ~pi1427 | ~new_n17413_;
  assign new_n17477_ = ~pi1017 | ~new_n16430_;
  assign new_n17478_ = ~pi1427 | ~new_n17414_;
  assign new_n17479_ = ~pi1426 | ~new_n17413_;
  assign new_n17480_ = ~pi1018 | ~new_n16430_;
  assign new_n17481_ = ~pi1426 | ~new_n17414_;
  assign new_n17482_ = ~pi1425 | ~new_n17413_;
  assign new_n17483_ = ~pi1019 | ~new_n16430_;
  assign new_n17484_ = ~pi1425 | ~new_n17414_;
  assign new_n17485_ = ~pi1424 | ~new_n17413_;
  assign new_n17486_ = ~pi1020 | ~new_n16430_;
  assign new_n17487_ = ~pi1424 | ~new_n17414_;
  assign new_n17488_ = ~pi1423 | ~new_n17413_;
  assign new_n17489_ = ~pi1021 | ~new_n16430_;
  assign new_n17490_ = ~pi1423 | ~new_n17414_;
  assign new_n17491_ = ~pi1422 | ~new_n17413_;
  assign new_n17492_ = ~pi1022 | ~new_n16430_;
  assign new_n17493_ = ~pi1422 | ~new_n17414_;
  assign new_n17494_ = ~pi1421 | ~new_n17413_;
  assign new_n17495_ = ~pi1023 | ~new_n16430_;
  assign new_n17496_ = ~pi1421 | ~new_n17414_;
  assign new_n17497_ = ~pi1420 | ~new_n17413_;
  assign new_n17498_ = ~pi1024 | ~new_n16430_;
  assign new_n17499_ = ~pi1420 | ~new_n17414_;
  assign new_n17500_ = ~pi1419 | ~new_n17413_;
  assign new_n17501_ = ~pi1025 | ~new_n16430_;
  assign new_n17502_ = ~pi1419 | ~new_n17414_;
  assign new_n17503_ = ~pi1418 | ~new_n17413_;
  assign new_n17504_ = ~pi1026 | ~new_n16430_;
  assign new_n17505_ = ~pi1418 | ~new_n17414_;
  assign new_n17506_ = ~pi1417 | ~new_n17413_;
  assign new_n17507_ = ~pi1027 | ~new_n16430_;
  assign new_n17508_ = ~pi1417 | ~new_n17414_;
  assign new_n17509_ = ~pi1416 | ~new_n17413_;
  assign new_n17510_ = ~pi1028 | ~new_n16430_;
  assign new_n17511_ = ~pi1416 | ~new_n17414_;
  assign new_n17512_ = ~pi1415 | ~new_n17413_;
  assign new_n17513_ = ~pi1029 | ~new_n16430_;
  assign new_n17514_ = ~pi1415 | ~new_n17414_;
  assign new_n17515_ = ~pi1414 | ~new_n17413_;
  assign new_n17516_ = ~pi1030 | ~new_n16430_;
  assign new_n17517_ = ~pi1414 | ~new_n17414_;
  assign new_n17518_ = ~pi1413 | ~new_n17413_;
  assign new_n17519_ = ~pi1031 | ~new_n16430_;
  assign new_n17520_ = ~pi1413 | ~new_n17414_;
  assign new_n17521_ = ~pi1412 | ~new_n17413_;
  assign new_n17522_ = ~pi1032 | ~new_n16430_;
  assign new_n17523_ = ~pi1412 | ~new_n17414_;
  assign new_n17524_ = ~pi1411 | ~new_n17413_;
  assign new_n17525_ = ~pi1033 | ~new_n16430_;
  assign new_n17526_ = ~pi1411 | ~new_n17414_;
  assign new_n17527_ = ~pi1410 | ~new_n17413_;
  assign new_n17528_ = ~pi1034 | ~new_n16430_;
  assign new_n17529_ = ~pi1410 | ~new_n17414_;
  assign new_n17530_ = ~pi1409 | ~new_n17413_;
  assign new_n17531_ = ~pi1035 | ~new_n16430_;
  assign new_n17532_ = ~pi1409 | ~new_n17414_;
  assign new_n17533_ = ~pi1408 | ~new_n17413_;
  assign new_n17534_ = ~pi1036 | ~new_n16430_;
  assign new_n17535_ = ~pi1408 | ~new_n17414_;
  assign new_n17536_ = ~pi1407 | ~new_n17413_;
  assign new_n17537_ = ~pi1037 | ~new_n16430_;
  assign new_n17538_ = ~new_n16441_;
  assign new_n17539_ = ~new_n17538_ | ~new_n16438_;
  assign new_n17540_ = ~pi0034 | ~new_n17439_;
  assign new_n17541_ = ~new_n16442_;
  assign new_n17542_ = ~new_n17541_ | ~new_n16438_;
  assign new_n17543_ = pi1040 | pi0034;
  assign new_n17544_ = ~new_n20804_ | ~new_n20803_ | ~new_n17543_;
  assign new_n17545_ = ~new_n16436_;
  assign new_n17546_ = ~new_n17545_ | ~pi0033 | ~new_n16428_;
  assign new_n17547_ = ~new_n2972_ | ~pi1039 | ~new_n16442_;
  assign new_n17548_ = ~new_n17547_ | ~new_n17546_;
  assign new_n17549_ = ~new_n17548_ | ~pi1040 | ~new_n17540_;
  assign new_n17550_ = ~pi1038 | ~new_n17544_;
  assign new_n17551_ = ~new_n2972_ | ~new_n17402_;
  assign new_n17552_ = ~new_n16677_ | ~new_n20806_;
  assign new_n17553_ = ~pi1038 | ~new_n16441_;
  assign new_n17554_ = ~pi0034 | ~new_n16439_;
  assign new_n17555_ = ~new_n17554_ | ~new_n17553_;
  assign new_n17556_ = ~new_n17555_ | ~new_n16429_;
  assign new_n17557_ = ~new_n17360_ | ~new_n16436_;
  assign new_n17558_ = ~new_n16461_;
  assign new_n17559_ = ~new_n16450_;
  assign new_n17560_ = ~new_n16625_;
  assign new_n17561_ = ~new_n16449_;
  assign new_n17562_ = ~new_n16455_;
  assign new_n17563_ = ~new_n16448_;
  assign new_n17564_ = ~pi1145 | ~new_n17563_;
  assign new_n17565_ = ~pi1201 | ~new_n15653_;
  assign new_n17566_ = ~pi1193 | ~new_n15652_;
  assign new_n17567_ = ~pi1185 | ~new_n15651_;
  assign new_n17568_ = ~pi1177 | ~new_n15649_;
  assign new_n17569_ = ~pi1169 | ~new_n15648_;
  assign new_n17570_ = ~pi1161 | ~new_n15647_;
  assign new_n17571_ = ~pi1153 | ~new_n15646_;
  assign new_n17572_ = ~pi1137 | ~new_n15645_;
  assign new_n17573_ = ~pi1129 | ~new_n15644_;
  assign new_n17574_ = ~pi1121 | ~new_n15642_;
  assign new_n17575_ = ~pi1113 | ~new_n15640_;
  assign new_n17576_ = ~pi1105 | ~new_n15639_;
  assign new_n17577_ = ~pi1097 | ~new_n15638_;
  assign new_n17578_ = ~pi1089 | ~new_n15636_;
  assign new_n17579_ = ~pi1081 | ~new_n15634_;
  assign new_n17580_ = ~new_n16464_;
  assign new_n17581_ = ~new_n16459_;
  assign new_n17582_ = ~pi1207 | ~pi1209 | ~pi1143 | ~pi1208 | ~new_n16451_;
  assign new_n17583_ = ~new_n17561_ | ~pi1199 | ~new_n16451_;
  assign new_n17584_ = ~new_n15650_ | ~new_n16446_ | ~pi1209 | ~pi1191;
  assign new_n17585_ = ~new_n15650_ | ~new_n16447_ | ~pi1208 | ~pi1183;
  assign new_n17586_ = ~new_n17559_ | ~new_n16451_ | ~pi1207 | ~pi1167;
  assign new_n17587_ = ~new_n16702_ | ~new_n16701_ | ~pi1207;
  assign new_n17588_ = ~new_n16704_ | ~new_n16703_ | ~pi1207;
  assign new_n17589_ = ~new_n16705_ | ~new_n17561_;
  assign new_n17590_ = ~new_n16707_ | ~new_n16706_ | ~pi1208;
  assign new_n17591_ = ~pi1208 | ~pi1206 | ~pi1111 | ~pi1209 | ~new_n16445_;
  assign new_n17592_ = ~new_n16708_ | ~new_n17559_ | ~pi1207;
  assign new_n17593_ = ~pi1207 | ~pi1206 | ~pi1095 | ~pi1209 | ~new_n16446_;
  assign new_n17594_ = ~pi1207 | ~pi1206 | ~pi1087 | ~pi1208 | ~new_n16447_;
  assign new_n17595_ = ~pi1208 | ~pi1206 | ~pi1079 | ~pi1209 | ~pi1207;
  assign new_n17596_ = ~new_n17354_;
  assign new_n17597_ = ~pi1146 | ~new_n17563_;
  assign new_n17598_ = ~pi1202 | ~new_n15653_;
  assign new_n17599_ = ~pi1194 | ~new_n15652_;
  assign new_n17600_ = ~pi1186 | ~new_n15651_;
  assign new_n17601_ = ~pi1178 | ~new_n15649_;
  assign new_n17602_ = ~pi1170 | ~new_n15648_;
  assign new_n17603_ = ~pi1162 | ~new_n15647_;
  assign new_n17604_ = ~pi1154 | ~new_n15646_;
  assign new_n17605_ = ~pi1138 | ~new_n15645_;
  assign new_n17606_ = ~pi1130 | ~new_n15644_;
  assign new_n17607_ = ~pi1122 | ~new_n15642_;
  assign new_n17608_ = ~pi1114 | ~new_n15640_;
  assign new_n17609_ = ~pi1106 | ~new_n15639_;
  assign new_n17610_ = ~pi1098 | ~new_n15638_;
  assign new_n17611_ = ~pi1090 | ~new_n15636_;
  assign new_n17612_ = ~pi1082 | ~new_n15634_;
  assign new_n17613_ = ~new_n17352_;
  assign new_n17614_ = ~pi1141 | ~new_n17563_;
  assign new_n17615_ = ~pi1197 | ~new_n15653_;
  assign new_n17616_ = ~pi1189 | ~new_n15652_;
  assign new_n17617_ = ~pi1181 | ~new_n15651_;
  assign new_n17618_ = ~pi1173 | ~new_n15649_;
  assign new_n17619_ = ~pi1165 | ~new_n15648_;
  assign new_n17620_ = ~pi1157 | ~new_n15647_;
  assign new_n17621_ = ~pi1149 | ~new_n15646_;
  assign new_n17622_ = ~pi1133 | ~new_n15645_;
  assign new_n17623_ = ~pi1125 | ~new_n15644_;
  assign new_n17624_ = ~pi1117 | ~new_n15642_;
  assign new_n17625_ = ~pi1109 | ~new_n15640_;
  assign new_n17626_ = ~pi1101 | ~new_n15639_;
  assign new_n17627_ = ~pi1093 | ~new_n15638_;
  assign new_n17628_ = ~pi1085 | ~new_n15636_;
  assign new_n17629_ = ~pi1077 | ~new_n15634_;
  assign new_n17630_ = ~new_n16572_;
  assign new_n17631_ = ~pi1142 | ~new_n16679_ | ~new_n17562_;
  assign new_n17632_ = ~new_n15637_ | ~pi1190 | ~new_n15650_;
  assign new_n17633_ = ~new_n15635_ | ~pi1182 | ~new_n15650_;
  assign new_n17634_ = ~new_n17562_ | ~pi1166 | ~new_n17559_;
  assign new_n17635_ = ~pi1158 | ~new_n15637_ | ~new_n17562_;
  assign new_n17636_ = ~pi1150 | ~new_n15635_ | ~new_n17562_;
  assign new_n17637_ = ~new_n16688_ | ~pi1102 | ~new_n17559_;
  assign new_n17638_ = ~pi1094 | ~new_n16688_ | ~new_n15637_;
  assign new_n17639_ = ~pi1086 | ~new_n16688_ | ~new_n15635_;
  assign new_n17640_ = ~pi1078 | ~new_n16688_ | ~new_n16679_;
  assign new_n17641_ = ~new_n16458_;
  assign new_n17642_ = ~pi1147 | ~new_n17563_;
  assign new_n17643_ = ~pi1203 | ~new_n15653_;
  assign new_n17644_ = ~pi1195 | ~new_n15652_;
  assign new_n17645_ = ~pi1187 | ~new_n15651_;
  assign new_n17646_ = ~pi1179 | ~new_n15649_;
  assign new_n17647_ = ~pi1171 | ~new_n15648_;
  assign new_n17648_ = ~pi1163 | ~new_n15647_;
  assign new_n17649_ = ~pi1155 | ~new_n15646_;
  assign new_n17650_ = ~pi1139 | ~new_n15645_;
  assign new_n17651_ = ~pi1131 | ~new_n15644_;
  assign new_n17652_ = ~pi1123 | ~new_n15642_;
  assign new_n17653_ = ~pi1115 | ~new_n15640_;
  assign new_n17654_ = ~pi1107 | ~new_n15639_;
  assign new_n17655_ = ~pi1099 | ~new_n15638_;
  assign new_n17656_ = ~pi1091 | ~new_n15636_;
  assign new_n17657_ = ~pi1083 | ~new_n15634_;
  assign new_n17658_ = ~new_n16452_;
  assign new_n17659_ = ~pi1148 | ~new_n17563_;
  assign new_n17660_ = ~pi1204 | ~new_n15653_;
  assign new_n17661_ = ~pi1196 | ~new_n15652_;
  assign new_n17662_ = ~pi1188 | ~new_n15651_;
  assign new_n17663_ = ~pi1180 | ~new_n15649_;
  assign new_n17664_ = ~pi1172 | ~new_n15648_;
  assign new_n17665_ = ~pi1164 | ~new_n15647_;
  assign new_n17666_ = ~pi1156 | ~new_n15646_;
  assign new_n17667_ = ~pi1140 | ~new_n15645_;
  assign new_n17668_ = ~pi1132 | ~new_n15644_;
  assign new_n17669_ = ~pi1124 | ~new_n15642_;
  assign new_n17670_ = ~pi1116 | ~new_n15640_;
  assign new_n17671_ = ~pi1108 | ~new_n15639_;
  assign new_n17672_ = ~pi1100 | ~new_n15638_;
  assign new_n17673_ = ~pi1092 | ~new_n15636_;
  assign new_n17674_ = ~pi1084 | ~new_n15634_;
  assign new_n17675_ = ~new_n16465_;
  assign new_n17676_ = ~pi1038 | ~new_n16429_;
  assign new_n17677_ = ~new_n16435_ | ~new_n17676_;
  assign new_n17678_ = ~new_n16453_;
  assign new_n17679_ = ~new_n17658_ | ~new_n16569_;
  assign new_n17680_ = ~new_n16618_;
  assign new_n17681_ = ~new_n16468_ | ~new_n16453_ | ~new_n16571_;
  assign new_n17682_ = ~new_n17681_ | ~new_n16438_;
  assign new_n17683_ = ~new_n16466_;
  assign new_n17684_ = ~new_n17641_ | ~new_n17354_;
  assign new_n17685_ = ~new_n17377_ | ~new_n16467_;
  assign new_n17686_ = ~new_n17685_ | ~new_n16760_;
  assign new_n17687_ = ~new_n16761_ | ~new_n17686_;
  assign new_n17688_ = ~new_n17396_ | ~new_n16569_;
  assign new_n17689_ = ~new_n17688_ | ~new_n20863_ | ~new_n20862_;
  assign new_n17690_ = ~new_n15629_ | ~new_n17443_;
  assign new_n17691_ = pi1444 | pi1443;
  assign new_n17692_ = ~new_n16474_;
  assign new_n17693_ = ~new_n17692_ | ~new_n16443_;
  assign new_n17694_ = ~pi1075 | ~new_n2972_;
  assign new_n17695_ = ~new_n16476_;
  assign new_n17696_ = ~pi1075 | ~new_n20869_ | ~new_n20868_;
  assign new_n17697_ = ~pi1074 | ~new_n16476_;
  assign new_n17698_ = ~new_n20785_ | ~new_n17427_;
  assign new_n17699_ = ~new_n16764_ | ~new_n17695_;
  assign new_n17700_ = ~pi1075 | ~new_n17698_;
  assign new_n17701_ = ~new_n15549_ | ~new_n20785_;
  assign new_n17702_ = ~new_n17433_ | ~new_n17442_;
  assign new_n17703_ = ~new_n20785_ | ~new_n17426_;
  assign new_n17704_ = ~new_n15549_ | ~new_n16474_;
  assign new_n17705_ = ~new_n16506_;
  assign new_n17706_ = ~new_n16512_;
  assign new_n17707_ = ~new_n16513_;
  assign new_n17708_ = ~new_n16495_;
  assign new_n17709_ = ~new_n16494_;
  assign new_n17710_ = ~new_n16523_;
  assign new_n17711_ = ~new_n31235_ | ~new_n16494_;
  assign new_n17712_ = ~new_n16539_;
  assign new_n17713_ = ~new_n16496_;
  assign new_n17714_ = ~new_n16486_;
  assign new_n17715_ = ~new_n16487_;
  assign new_n17716_ = ~new_n15619_ | ~new_n15623_;
  assign new_n17717_ = ~new_n16502_;
  assign new_n17718_ = ~new_n16537_;
  assign new_n17719_ = ~new_n16521_;
  assign new_n17720_ = ~pi1211 | ~new_n16486_;
  assign new_n17721_ = ~new_n16541_;
  assign new_n17722_ = ~new_n16510_;
  assign new_n17723_ = ~new_n16504_;
  assign new_n17724_ = ~new_n16416_;
  assign new_n17725_ = ~new_n15613_ | ~new_n15617_;
  assign new_n17726_ = ~new_n16503_;
  assign new_n17727_ = ~pi1075 | ~new_n16444_;
  assign new_n17728_ = ~new_n16480_ | ~new_n17727_ | ~new_n16478_;
  assign new_n17729_ = ~new_n17709_ | ~new_n15657_;
  assign new_n17730_ = ~new_n15661_ | ~new_n15539_;
  assign new_n17731_ = ~new_n16501_ | ~new_n17730_;
  assign new_n17732_ = ~new_n17717_ | ~new_n17731_;
  assign new_n17733_ = ~pi1073 | ~new_n16487_;
  assign new_n17734_ = ~new_n17726_ | ~pi1074;
  assign new_n17735_ = ~new_n17732_ | ~new_n16768_;
  assign new_n17736_ = ~new_n15661_ | ~new_n15569_;
  assign new_n17737_ = ~new_n16501_ | ~new_n17736_;
  assign new_n17738_ = ~new_n17737_ | ~new_n16502_;
  assign new_n17739_ = ~pi1074 | ~new_n16503_;
  assign new_n17740_ = ~new_n17739_ | ~new_n17738_;
  assign new_n17741_ = ~new_n15596_ | ~new_n17715_;
  assign new_n17742_ = ~new_n15594_ | ~new_n15658_;
  assign new_n17743_ = ~new_n15593_ | ~new_n17713_;
  assign new_n17744_ = ~new_n15578_ | ~new_n17740_;
  assign new_n17745_ = ~pi1077 | ~new_n17735_;
  assign new_n17746_ = ~new_n15597_ | ~new_n17715_;
  assign new_n17747_ = ~new_n15592_ | ~new_n15658_;
  assign new_n17748_ = ~new_n15591_ | ~new_n17713_;
  assign new_n17749_ = ~new_n15577_ | ~new_n17740_;
  assign new_n17750_ = ~pi1078 | ~new_n17735_;
  assign new_n17751_ = ~new_n15601_ | ~new_n17715_;
  assign new_n17752_ = ~new_n15590_ | ~new_n15658_;
  assign new_n17753_ = ~new_n15589_ | ~new_n17713_;
  assign new_n17754_ = ~new_n15576_ | ~new_n17740_;
  assign new_n17755_ = ~pi1079 | ~new_n17735_;
  assign new_n17756_ = ~new_n15600_ | ~new_n17715_;
  assign new_n17757_ = ~new_n15588_ | ~new_n15658_;
  assign new_n17758_ = ~new_n15587_ | ~new_n17713_;
  assign new_n17759_ = ~new_n15575_ | ~new_n17740_;
  assign new_n17760_ = ~pi1080 | ~new_n17735_;
  assign new_n17761_ = ~new_n15599_ | ~new_n17715_;
  assign new_n17762_ = ~new_n15586_ | ~new_n15658_;
  assign new_n17763_ = ~new_n15585_ | ~new_n17713_;
  assign new_n17764_ = ~new_n15574_ | ~new_n17740_;
  assign new_n17765_ = ~pi1081 | ~new_n17735_;
  assign new_n17766_ = ~new_n15602_ | ~new_n17715_;
  assign new_n17767_ = ~new_n15584_ | ~new_n15658_;
  assign new_n17768_ = ~new_n15583_ | ~new_n17713_;
  assign new_n17769_ = ~new_n15573_ | ~new_n17740_;
  assign new_n17770_ = ~pi1082 | ~new_n17735_;
  assign new_n17771_ = ~new_n15595_ | ~new_n17715_;
  assign new_n17772_ = ~new_n15582_ | ~new_n15658_;
  assign new_n17773_ = ~new_n15581_ | ~new_n17713_;
  assign new_n17774_ = ~new_n15572_ | ~new_n17740_;
  assign new_n17775_ = ~pi1083 | ~new_n17735_;
  assign new_n17776_ = ~new_n15598_ | ~new_n17715_;
  assign new_n17777_ = ~new_n15580_ | ~new_n15658_;
  assign new_n17778_ = ~new_n15579_ | ~new_n17713_;
  assign new_n17779_ = ~new_n15571_ | ~new_n17740_;
  assign new_n17780_ = ~pi1084 | ~new_n17735_;
  assign new_n17781_ = ~new_n16507_;
  assign new_n17782_ = ~new_n16508_;
  assign new_n17783_ = ~new_n16505_;
  assign new_n17784_ = ~new_n15624_ | ~new_n15619_;
  assign new_n17785_ = ~new_n16509_;
  assign new_n17786_ = ~new_n16417_;
  assign new_n17787_ = ~new_n17705_ | ~new_n15657_;
  assign new_n17788_ = ~new_n15663_ | ~new_n15539_;
  assign new_n17789_ = ~new_n16501_ | ~new_n17788_;
  assign new_n17790_ = ~new_n17785_ | ~new_n17789_;
  assign new_n17791_ = ~pi1073 | ~new_n16505_;
  assign new_n17792_ = ~pi1074 | ~new_n16417_;
  assign new_n17793_ = ~new_n17790_ | ~new_n16777_;
  assign new_n17794_ = ~new_n15663_ | ~new_n15569_;
  assign new_n17795_ = ~new_n16501_ | ~new_n17794_;
  assign new_n17796_ = ~new_n17795_ | ~new_n16509_;
  assign new_n17797_ = ~pi1074 | ~new_n17786_;
  assign new_n17798_ = ~new_n17797_ | ~new_n17796_;
  assign new_n17799_ = ~new_n17783_ | ~new_n15596_;
  assign new_n17800_ = ~new_n15662_ | ~new_n15594_;
  assign new_n17801_ = ~new_n17782_ | ~new_n15593_;
  assign new_n17802_ = ~new_n15578_ | ~new_n17798_;
  assign new_n17803_ = ~pi1085 | ~new_n17793_;
  assign new_n17804_ = ~new_n17783_ | ~new_n15597_;
  assign new_n17805_ = ~new_n15662_ | ~new_n15592_;
  assign new_n17806_ = ~new_n17782_ | ~new_n15591_;
  assign new_n17807_ = ~new_n15577_ | ~new_n17798_;
  assign new_n17808_ = ~pi1086 | ~new_n17793_;
  assign new_n17809_ = ~new_n17783_ | ~new_n15601_;
  assign new_n17810_ = ~new_n15662_ | ~new_n15590_;
  assign new_n17811_ = ~new_n17782_ | ~new_n15589_;
  assign new_n17812_ = ~new_n15576_ | ~new_n17798_;
  assign new_n17813_ = ~pi1087 | ~new_n17793_;
  assign new_n17814_ = ~new_n17783_ | ~new_n15600_;
  assign new_n17815_ = ~new_n15662_ | ~new_n15588_;
  assign new_n17816_ = ~new_n17782_ | ~new_n15587_;
  assign new_n17817_ = ~new_n15575_ | ~new_n17798_;
  assign new_n17818_ = ~pi1088 | ~new_n17793_;
  assign new_n17819_ = ~new_n17783_ | ~new_n15599_;
  assign new_n17820_ = ~new_n15662_ | ~new_n15586_;
  assign new_n17821_ = ~new_n17782_ | ~new_n15585_;
  assign new_n17822_ = ~new_n15574_ | ~new_n17798_;
  assign new_n17823_ = ~pi1089 | ~new_n17793_;
  assign new_n17824_ = ~new_n17783_ | ~new_n15602_;
  assign new_n17825_ = ~new_n15662_ | ~new_n15584_;
  assign new_n17826_ = ~new_n17782_ | ~new_n15583_;
  assign new_n17827_ = ~new_n15573_ | ~new_n17798_;
  assign new_n17828_ = ~pi1090 | ~new_n17793_;
  assign new_n17829_ = ~new_n17783_ | ~new_n15595_;
  assign new_n17830_ = ~new_n15662_ | ~new_n15582_;
  assign new_n17831_ = ~new_n17782_ | ~new_n15581_;
  assign new_n17832_ = ~new_n15572_ | ~new_n17798_;
  assign new_n17833_ = ~pi1091 | ~new_n17793_;
  assign new_n17834_ = ~new_n17783_ | ~new_n15598_;
  assign new_n17835_ = ~new_n15662_ | ~new_n15580_;
  assign new_n17836_ = ~new_n17782_ | ~new_n15579_;
  assign new_n17837_ = ~new_n15571_ | ~new_n17798_;
  assign new_n17838_ = ~pi1092 | ~new_n17793_;
  assign new_n17839_ = ~new_n16514_;
  assign new_n17840_ = ~new_n16515_;
  assign new_n17841_ = ~new_n16511_;
  assign new_n17842_ = ~new_n15625_ | ~new_n15619_;
  assign new_n17843_ = ~new_n16516_;
  assign new_n17844_ = ~new_n15618_ | ~new_n15613_;
  assign new_n17845_ = ~new_n16517_;
  assign new_n17846_ = ~new_n17706_ | ~new_n15657_;
  assign new_n17847_ = ~new_n15665_ | ~new_n15539_;
  assign new_n17848_ = ~new_n16501_ | ~new_n17847_;
  assign new_n17849_ = ~new_n17843_ | ~new_n17848_;
  assign new_n17850_ = ~pi1073 | ~new_n16511_;
  assign new_n17851_ = ~new_n17845_ | ~pi1074;
  assign new_n17852_ = ~new_n17849_ | ~new_n16786_;
  assign new_n17853_ = ~new_n15665_ | ~new_n15569_;
  assign new_n17854_ = ~new_n16501_ | ~new_n17853_;
  assign new_n17855_ = ~new_n17854_ | ~new_n16516_;
  assign new_n17856_ = ~pi1074 | ~new_n16517_;
  assign new_n17857_ = ~new_n17856_ | ~new_n17855_;
  assign new_n17858_ = ~new_n17841_ | ~new_n15596_;
  assign new_n17859_ = ~new_n15664_ | ~new_n15594_;
  assign new_n17860_ = ~new_n17840_ | ~new_n15593_;
  assign new_n17861_ = ~new_n15578_ | ~new_n17857_;
  assign new_n17862_ = ~pi1093 | ~new_n17852_;
  assign new_n17863_ = ~new_n17841_ | ~new_n15597_;
  assign new_n17864_ = ~new_n15664_ | ~new_n15592_;
  assign new_n17865_ = ~new_n17840_ | ~new_n15591_;
  assign new_n17866_ = ~new_n15577_ | ~new_n17857_;
  assign new_n17867_ = ~pi1094 | ~new_n17852_;
  assign new_n17868_ = ~new_n17841_ | ~new_n15601_;
  assign new_n17869_ = ~new_n15664_ | ~new_n15590_;
  assign new_n17870_ = ~new_n17840_ | ~new_n15589_;
  assign new_n17871_ = ~new_n15576_ | ~new_n17857_;
  assign new_n17872_ = ~pi1095 | ~new_n17852_;
  assign new_n17873_ = ~new_n17841_ | ~new_n15600_;
  assign new_n17874_ = ~new_n15664_ | ~new_n15588_;
  assign new_n17875_ = ~new_n17840_ | ~new_n15587_;
  assign new_n17876_ = ~new_n15575_ | ~new_n17857_;
  assign new_n17877_ = ~pi1096 | ~new_n17852_;
  assign new_n17878_ = ~new_n17841_ | ~new_n15599_;
  assign new_n17879_ = ~new_n15664_ | ~new_n15586_;
  assign new_n17880_ = ~new_n17840_ | ~new_n15585_;
  assign new_n17881_ = ~new_n15574_ | ~new_n17857_;
  assign new_n17882_ = ~pi1097 | ~new_n17852_;
  assign new_n17883_ = ~new_n17841_ | ~new_n15602_;
  assign new_n17884_ = ~new_n15664_ | ~new_n15584_;
  assign new_n17885_ = ~new_n17840_ | ~new_n15583_;
  assign new_n17886_ = ~new_n15573_ | ~new_n17857_;
  assign new_n17887_ = ~pi1098 | ~new_n17852_;
  assign new_n17888_ = ~new_n17841_ | ~new_n15595_;
  assign new_n17889_ = ~new_n15664_ | ~new_n15582_;
  assign new_n17890_ = ~new_n17840_ | ~new_n15581_;
  assign new_n17891_ = ~new_n15572_ | ~new_n17857_;
  assign new_n17892_ = ~pi1099 | ~new_n17852_;
  assign new_n17893_ = ~new_n17841_ | ~new_n15598_;
  assign new_n17894_ = ~new_n15664_ | ~new_n15580_;
  assign new_n17895_ = ~new_n17840_ | ~new_n15579_;
  assign new_n17896_ = ~new_n15571_ | ~new_n17857_;
  assign new_n17897_ = ~pi1100 | ~new_n17852_;
  assign new_n17898_ = ~new_n16519_;
  assign new_n17899_ = ~new_n16518_;
  assign new_n17900_ = ~new_n15626_ | ~new_n15619_;
  assign new_n17901_ = ~new_n16520_;
  assign new_n17902_ = ~new_n16418_;
  assign new_n17903_ = ~new_n15667_ | ~new_n15657_;
  assign new_n17904_ = ~new_n15670_ | ~new_n15539_;
  assign new_n17905_ = ~new_n16501_ | ~new_n17904_;
  assign new_n17906_ = ~new_n17901_ | ~new_n17905_;
  assign new_n17907_ = ~pi1073 | ~new_n16518_;
  assign new_n17908_ = ~pi1074 | ~new_n16418_;
  assign new_n17909_ = ~new_n17906_ | ~new_n16795_;
  assign new_n17910_ = ~new_n15670_ | ~new_n15569_;
  assign new_n17911_ = ~new_n16501_ | ~new_n17910_;
  assign new_n17912_ = ~new_n17911_ | ~new_n16520_;
  assign new_n17913_ = ~pi1074 | ~new_n17902_;
  assign new_n17914_ = ~new_n17913_ | ~new_n17912_;
  assign new_n17915_ = ~new_n17899_ | ~new_n15596_;
  assign new_n17916_ = ~new_n15668_ | ~new_n15594_;
  assign new_n17917_ = ~new_n17898_ | ~new_n15593_;
  assign new_n17918_ = ~new_n15578_ | ~new_n17914_;
  assign new_n17919_ = ~pi1101 | ~new_n17909_;
  assign new_n17920_ = ~new_n17899_ | ~new_n15597_;
  assign new_n17921_ = ~new_n15668_ | ~new_n15592_;
  assign new_n17922_ = ~new_n17898_ | ~new_n15591_;
  assign new_n17923_ = ~new_n15577_ | ~new_n17914_;
  assign new_n17924_ = ~pi1102 | ~new_n17909_;
  assign new_n17925_ = ~new_n17899_ | ~new_n15601_;
  assign new_n17926_ = ~new_n15668_ | ~new_n15590_;
  assign new_n17927_ = ~new_n17898_ | ~new_n15589_;
  assign new_n17928_ = ~new_n15576_ | ~new_n17914_;
  assign new_n17929_ = ~pi1103 | ~new_n17909_;
  assign new_n17930_ = ~new_n17899_ | ~new_n15600_;
  assign new_n17931_ = ~new_n15668_ | ~new_n15588_;
  assign new_n17932_ = ~new_n17898_ | ~new_n15587_;
  assign new_n17933_ = ~new_n15575_ | ~new_n17914_;
  assign new_n17934_ = ~pi1104 | ~new_n17909_;
  assign new_n17935_ = ~new_n17899_ | ~new_n15599_;
  assign new_n17936_ = ~new_n15668_ | ~new_n15586_;
  assign new_n17937_ = ~new_n17898_ | ~new_n15585_;
  assign new_n17938_ = ~new_n15574_ | ~new_n17914_;
  assign new_n17939_ = ~pi1105 | ~new_n17909_;
  assign new_n17940_ = ~new_n17899_ | ~new_n15602_;
  assign new_n17941_ = ~new_n15668_ | ~new_n15584_;
  assign new_n17942_ = ~new_n17898_ | ~new_n15583_;
  assign new_n17943_ = ~new_n15573_ | ~new_n17914_;
  assign new_n17944_ = ~pi1106 | ~new_n17909_;
  assign new_n17945_ = ~new_n17899_ | ~new_n15595_;
  assign new_n17946_ = ~new_n15668_ | ~new_n15582_;
  assign new_n17947_ = ~new_n17898_ | ~new_n15581_;
  assign new_n17948_ = ~new_n15572_ | ~new_n17914_;
  assign new_n17949_ = ~pi1107 | ~new_n17909_;
  assign new_n17950_ = ~new_n17899_ | ~new_n15598_;
  assign new_n17951_ = ~new_n15668_ | ~new_n15580_;
  assign new_n17952_ = ~new_n17898_ | ~new_n15579_;
  assign new_n17953_ = ~new_n15571_ | ~new_n17914_;
  assign new_n17954_ = ~pi1108 | ~new_n17909_;
  assign new_n17955_ = ~new_n16524_;
  assign new_n17956_ = ~new_n16522_;
  assign new_n17957_ = ~new_n15621_ | ~new_n15623_;
  assign new_n17958_ = ~new_n16525_;
  assign new_n17959_ = ~new_n15615_ | ~new_n15617_;
  assign new_n17960_ = ~new_n16526_;
  assign new_n17961_ = ~new_n17710_ | ~new_n17709_;
  assign new_n17962_ = ~new_n15673_ | ~new_n15539_;
  assign new_n17963_ = ~new_n16501_ | ~new_n17962_;
  assign new_n17964_ = ~new_n17958_ | ~new_n17963_;
  assign new_n17965_ = ~pi1073 | ~new_n16522_;
  assign new_n17966_ = ~new_n17960_ | ~pi1074;
  assign new_n17967_ = ~new_n17964_ | ~new_n16804_;
  assign new_n17968_ = ~new_n15673_ | ~new_n15569_;
  assign new_n17969_ = ~new_n16501_ | ~new_n17968_;
  assign new_n17970_ = ~new_n17969_ | ~new_n16525_;
  assign new_n17971_ = ~pi1074 | ~new_n16526_;
  assign new_n17972_ = ~new_n17971_ | ~new_n17970_;
  assign new_n17973_ = ~new_n17956_ | ~new_n15596_;
  assign new_n17974_ = ~new_n15672_ | ~new_n15594_;
  assign new_n17975_ = ~new_n17955_ | ~new_n15593_;
  assign new_n17976_ = ~new_n15578_ | ~new_n17972_;
  assign new_n17977_ = ~pi1109 | ~new_n17967_;
  assign new_n17978_ = ~new_n17956_ | ~new_n15597_;
  assign new_n17979_ = ~new_n15672_ | ~new_n15592_;
  assign new_n17980_ = ~new_n17955_ | ~new_n15591_;
  assign new_n17981_ = ~new_n15577_ | ~new_n17972_;
  assign new_n17982_ = ~pi1110 | ~new_n17967_;
  assign new_n17983_ = ~new_n17956_ | ~new_n15601_;
  assign new_n17984_ = ~new_n15672_ | ~new_n15590_;
  assign new_n17985_ = ~new_n17955_ | ~new_n15589_;
  assign new_n17986_ = ~new_n15576_ | ~new_n17972_;
  assign new_n17987_ = ~pi1111 | ~new_n17967_;
  assign new_n17988_ = ~new_n17956_ | ~new_n15600_;
  assign new_n17989_ = ~new_n15672_ | ~new_n15588_;
  assign new_n17990_ = ~new_n17955_ | ~new_n15587_;
  assign new_n17991_ = ~new_n15575_ | ~new_n17972_;
  assign new_n17992_ = ~pi1112 | ~new_n17967_;
  assign new_n17993_ = ~new_n17956_ | ~new_n15599_;
  assign new_n17994_ = ~new_n15672_ | ~new_n15586_;
  assign new_n17995_ = ~new_n17955_ | ~new_n15585_;
  assign new_n17996_ = ~new_n15574_ | ~new_n17972_;
  assign new_n17997_ = ~pi1113 | ~new_n17967_;
  assign new_n17998_ = ~new_n17956_ | ~new_n15602_;
  assign new_n17999_ = ~new_n15672_ | ~new_n15584_;
  assign new_n18000_ = ~new_n17955_ | ~new_n15583_;
  assign new_n18001_ = ~new_n15573_ | ~new_n17972_;
  assign new_n18002_ = ~pi1114 | ~new_n17967_;
  assign new_n18003_ = ~new_n17956_ | ~new_n15595_;
  assign new_n18004_ = ~new_n15672_ | ~new_n15582_;
  assign new_n18005_ = ~new_n17955_ | ~new_n15581_;
  assign new_n18006_ = ~new_n15572_ | ~new_n17972_;
  assign new_n18007_ = ~pi1115 | ~new_n17967_;
  assign new_n18008_ = ~new_n17956_ | ~new_n15598_;
  assign new_n18009_ = ~new_n15672_ | ~new_n15580_;
  assign new_n18010_ = ~new_n17955_ | ~new_n15579_;
  assign new_n18011_ = ~new_n15571_ | ~new_n17972_;
  assign new_n18012_ = ~pi1116 | ~new_n17967_;
  assign new_n18013_ = ~new_n16528_;
  assign new_n18014_ = ~new_n16527_;
  assign new_n18015_ = ~new_n15621_ | ~new_n15624_;
  assign new_n18016_ = ~new_n16529_;
  assign new_n18017_ = ~new_n16419_;
  assign new_n18018_ = ~new_n17710_ | ~new_n17705_;
  assign new_n18019_ = ~new_n15675_ | ~new_n15539_;
  assign new_n18020_ = ~new_n16501_ | ~new_n18019_;
  assign new_n18021_ = ~new_n18016_ | ~new_n18020_;
  assign new_n18022_ = ~pi1073 | ~new_n16527_;
  assign new_n18023_ = ~pi1074 | ~new_n16419_;
  assign new_n18024_ = ~new_n18021_ | ~new_n16813_;
  assign new_n18025_ = ~new_n15675_ | ~new_n15569_;
  assign new_n18026_ = ~new_n16501_ | ~new_n18025_;
  assign new_n18027_ = ~new_n18026_ | ~new_n16529_;
  assign new_n18028_ = ~pi1074 | ~new_n18017_;
  assign new_n18029_ = ~new_n18028_ | ~new_n18027_;
  assign new_n18030_ = ~new_n18014_ | ~new_n15596_;
  assign new_n18031_ = ~new_n15674_ | ~new_n15594_;
  assign new_n18032_ = ~new_n18013_ | ~new_n15593_;
  assign new_n18033_ = ~new_n15578_ | ~new_n18029_;
  assign new_n18034_ = ~pi1117 | ~new_n18024_;
  assign new_n18035_ = ~new_n18014_ | ~new_n15597_;
  assign new_n18036_ = ~new_n15674_ | ~new_n15592_;
  assign new_n18037_ = ~new_n18013_ | ~new_n15591_;
  assign new_n18038_ = ~new_n15577_ | ~new_n18029_;
  assign new_n18039_ = ~pi1118 | ~new_n18024_;
  assign new_n18040_ = ~new_n18014_ | ~new_n15601_;
  assign new_n18041_ = ~new_n15674_ | ~new_n15590_;
  assign new_n18042_ = ~new_n18013_ | ~new_n15589_;
  assign new_n18043_ = ~new_n15576_ | ~new_n18029_;
  assign new_n18044_ = ~pi1119 | ~new_n18024_;
  assign new_n18045_ = ~new_n18014_ | ~new_n15600_;
  assign new_n18046_ = ~new_n15674_ | ~new_n15588_;
  assign new_n18047_ = ~new_n18013_ | ~new_n15587_;
  assign new_n18048_ = ~new_n15575_ | ~new_n18029_;
  assign new_n18049_ = ~pi1120 | ~new_n18024_;
  assign new_n18050_ = ~new_n18014_ | ~new_n15599_;
  assign new_n18051_ = ~new_n15674_ | ~new_n15586_;
  assign new_n18052_ = ~new_n18013_ | ~new_n15585_;
  assign new_n18053_ = ~new_n15574_ | ~new_n18029_;
  assign new_n18054_ = ~pi1121 | ~new_n18024_;
  assign new_n18055_ = ~new_n18014_ | ~new_n15602_;
  assign new_n18056_ = ~new_n15674_ | ~new_n15584_;
  assign new_n18057_ = ~new_n18013_ | ~new_n15583_;
  assign new_n18058_ = ~new_n15573_ | ~new_n18029_;
  assign new_n18059_ = ~pi1122 | ~new_n18024_;
  assign new_n18060_ = ~new_n18014_ | ~new_n15595_;
  assign new_n18061_ = ~new_n15674_ | ~new_n15582_;
  assign new_n18062_ = ~new_n18013_ | ~new_n15581_;
  assign new_n18063_ = ~new_n15572_ | ~new_n18029_;
  assign new_n18064_ = ~pi1123 | ~new_n18024_;
  assign new_n18065_ = ~new_n18014_ | ~new_n15598_;
  assign new_n18066_ = ~new_n15674_ | ~new_n15580_;
  assign new_n18067_ = ~new_n18013_ | ~new_n15579_;
  assign new_n18068_ = ~new_n15571_ | ~new_n18029_;
  assign new_n18069_ = ~pi1124 | ~new_n18024_;
  assign new_n18070_ = ~new_n16531_;
  assign new_n18071_ = ~new_n16530_;
  assign new_n18072_ = ~new_n15621_ | ~new_n15625_;
  assign new_n18073_ = ~new_n16532_;
  assign new_n18074_ = ~new_n15615_ | ~new_n15618_;
  assign new_n18075_ = ~new_n16533_;
  assign new_n18076_ = ~new_n17710_ | ~new_n17706_;
  assign new_n18077_ = ~new_n15677_ | ~new_n15539_;
  assign new_n18078_ = ~new_n16501_ | ~new_n18077_;
  assign new_n18079_ = ~new_n18073_ | ~new_n18078_;
  assign new_n18080_ = ~pi1073 | ~new_n16530_;
  assign new_n18081_ = ~new_n18075_ | ~pi1074;
  assign new_n18082_ = ~new_n18079_ | ~new_n16822_;
  assign new_n18083_ = ~new_n15677_ | ~new_n15569_;
  assign new_n18084_ = ~new_n16501_ | ~new_n18083_;
  assign new_n18085_ = ~new_n18084_ | ~new_n16532_;
  assign new_n18086_ = ~pi1074 | ~new_n16533_;
  assign new_n18087_ = ~new_n18086_ | ~new_n18085_;
  assign new_n18088_ = ~new_n18071_ | ~new_n15596_;
  assign new_n18089_ = ~new_n15676_ | ~new_n15594_;
  assign new_n18090_ = ~new_n18070_ | ~new_n15593_;
  assign new_n18091_ = ~new_n15578_ | ~new_n18087_;
  assign new_n18092_ = ~pi1125 | ~new_n18082_;
  assign new_n18093_ = ~new_n18071_ | ~new_n15597_;
  assign new_n18094_ = ~new_n15676_ | ~new_n15592_;
  assign new_n18095_ = ~new_n18070_ | ~new_n15591_;
  assign new_n18096_ = ~new_n15577_ | ~new_n18087_;
  assign new_n18097_ = ~pi1126 | ~new_n18082_;
  assign new_n18098_ = ~new_n18071_ | ~new_n15601_;
  assign new_n18099_ = ~new_n15676_ | ~new_n15590_;
  assign new_n18100_ = ~new_n18070_ | ~new_n15589_;
  assign new_n18101_ = ~new_n15576_ | ~new_n18087_;
  assign new_n18102_ = ~pi1127 | ~new_n18082_;
  assign new_n18103_ = ~new_n18071_ | ~new_n15600_;
  assign new_n18104_ = ~new_n15676_ | ~new_n15588_;
  assign new_n18105_ = ~new_n18070_ | ~new_n15587_;
  assign new_n18106_ = ~new_n15575_ | ~new_n18087_;
  assign new_n18107_ = ~pi1128 | ~new_n18082_;
  assign new_n18108_ = ~new_n18071_ | ~new_n15599_;
  assign new_n18109_ = ~new_n15676_ | ~new_n15586_;
  assign new_n18110_ = ~new_n18070_ | ~new_n15585_;
  assign new_n18111_ = ~new_n15574_ | ~new_n18087_;
  assign new_n18112_ = ~pi1129 | ~new_n18082_;
  assign new_n18113_ = ~new_n18071_ | ~new_n15602_;
  assign new_n18114_ = ~new_n15676_ | ~new_n15584_;
  assign new_n18115_ = ~new_n18070_ | ~new_n15583_;
  assign new_n18116_ = ~new_n15573_ | ~new_n18087_;
  assign new_n18117_ = ~pi1130 | ~new_n18082_;
  assign new_n18118_ = ~new_n18071_ | ~new_n15595_;
  assign new_n18119_ = ~new_n15676_ | ~new_n15582_;
  assign new_n18120_ = ~new_n18070_ | ~new_n15581_;
  assign new_n18121_ = ~new_n15572_ | ~new_n18087_;
  assign new_n18122_ = ~pi1131 | ~new_n18082_;
  assign new_n18123_ = ~new_n18071_ | ~new_n15598_;
  assign new_n18124_ = ~new_n15676_ | ~new_n15580_;
  assign new_n18125_ = ~new_n18070_ | ~new_n15579_;
  assign new_n18126_ = ~new_n15571_ | ~new_n18087_;
  assign new_n18127_ = ~pi1132 | ~new_n18082_;
  assign new_n18128_ = ~new_n16535_;
  assign new_n18129_ = ~new_n16534_;
  assign new_n18130_ = ~new_n15621_ | ~new_n15626_;
  assign new_n18131_ = ~new_n16536_;
  assign new_n18132_ = ~new_n16420_;
  assign new_n18133_ = ~new_n17710_ | ~new_n15667_;
  assign new_n18134_ = ~new_n15679_ | ~new_n15539_;
  assign new_n18135_ = ~new_n16501_ | ~new_n18134_;
  assign new_n18136_ = ~new_n18131_ | ~new_n18135_;
  assign new_n18137_ = ~pi1073 | ~new_n16534_;
  assign new_n18138_ = ~pi1074 | ~new_n16420_;
  assign new_n18139_ = ~new_n18136_ | ~new_n16831_;
  assign new_n18140_ = ~new_n15679_ | ~new_n15569_;
  assign new_n18141_ = ~new_n16501_ | ~new_n18140_;
  assign new_n18142_ = ~new_n18141_ | ~new_n16536_;
  assign new_n18143_ = ~pi1074 | ~new_n18132_;
  assign new_n18144_ = ~new_n18143_ | ~new_n18142_;
  assign new_n18145_ = ~new_n18129_ | ~new_n15596_;
  assign new_n18146_ = ~new_n15678_ | ~new_n15594_;
  assign new_n18147_ = ~new_n18128_ | ~new_n15593_;
  assign new_n18148_ = ~new_n15578_ | ~new_n18144_;
  assign new_n18149_ = ~pi1133 | ~new_n18139_;
  assign new_n18150_ = ~new_n18129_ | ~new_n15597_;
  assign new_n18151_ = ~new_n15678_ | ~new_n15592_;
  assign new_n18152_ = ~new_n18128_ | ~new_n15591_;
  assign new_n18153_ = ~new_n15577_ | ~new_n18144_;
  assign new_n18154_ = ~pi1134 | ~new_n18139_;
  assign new_n18155_ = ~new_n18129_ | ~new_n15601_;
  assign new_n18156_ = ~new_n15678_ | ~new_n15590_;
  assign new_n18157_ = ~new_n18128_ | ~new_n15589_;
  assign new_n18158_ = ~new_n15576_ | ~new_n18144_;
  assign new_n18159_ = ~pi1135 | ~new_n18139_;
  assign new_n18160_ = ~new_n18129_ | ~new_n15600_;
  assign new_n18161_ = ~new_n15678_ | ~new_n15588_;
  assign new_n18162_ = ~new_n18128_ | ~new_n15587_;
  assign new_n18163_ = ~new_n15575_ | ~new_n18144_;
  assign new_n18164_ = ~pi1136 | ~new_n18139_;
  assign new_n18165_ = ~new_n18129_ | ~new_n15599_;
  assign new_n18166_ = ~new_n15678_ | ~new_n15586_;
  assign new_n18167_ = ~new_n18128_ | ~new_n15585_;
  assign new_n18168_ = ~new_n15574_ | ~new_n18144_;
  assign new_n18169_ = ~pi1137 | ~new_n18139_;
  assign new_n18170_ = ~new_n18129_ | ~new_n15602_;
  assign new_n18171_ = ~new_n15678_ | ~new_n15584_;
  assign new_n18172_ = ~new_n18128_ | ~new_n15583_;
  assign new_n18173_ = ~new_n15573_ | ~new_n18144_;
  assign new_n18174_ = ~pi1138 | ~new_n18139_;
  assign new_n18175_ = ~new_n18129_ | ~new_n15595_;
  assign new_n18176_ = ~new_n15678_ | ~new_n15582_;
  assign new_n18177_ = ~new_n18128_ | ~new_n15581_;
  assign new_n18178_ = ~new_n15572_ | ~new_n18144_;
  assign new_n18179_ = ~pi1139 | ~new_n18139_;
  assign new_n18180_ = ~new_n18129_ | ~new_n15598_;
  assign new_n18181_ = ~new_n15678_ | ~new_n15580_;
  assign new_n18182_ = ~new_n18128_ | ~new_n15579_;
  assign new_n18183_ = ~new_n15571_ | ~new_n18144_;
  assign new_n18184_ = ~pi1140 | ~new_n18139_;
  assign new_n18185_ = ~new_n16540_;
  assign new_n18186_ = ~new_n15620_ | ~new_n15623_;
  assign new_n18187_ = ~new_n16542_;
  assign new_n18188_ = ~new_n15614_ | ~new_n15617_;
  assign new_n18189_ = ~new_n16543_;
  assign new_n18190_ = ~new_n15681_ | ~new_n15539_;
  assign new_n18191_ = ~new_n16501_ | ~new_n18190_;
  assign new_n18192_ = ~new_n18187_ | ~new_n18191_;
  assign new_n18193_ = ~pi1073 | ~new_n16537_;
  assign new_n18194_ = ~new_n18189_ | ~pi1074;
  assign new_n18195_ = ~new_n18192_ | ~new_n16840_;
  assign new_n18196_ = ~new_n15681_ | ~new_n15569_;
  assign new_n18197_ = ~new_n16501_ | ~new_n18196_;
  assign new_n18198_ = ~new_n18197_ | ~new_n16542_;
  assign new_n18199_ = ~pi1074 | ~new_n16543_;
  assign new_n18200_ = ~new_n18199_ | ~new_n18198_;
  assign new_n18201_ = ~new_n17718_ | ~new_n15596_;
  assign new_n18202_ = ~new_n17419_ | ~new_n15594_;
  assign new_n18203_ = ~new_n18185_ | ~new_n15593_;
  assign new_n18204_ = ~new_n15578_ | ~new_n18200_;
  assign new_n18205_ = ~pi1141 | ~new_n18195_;
  assign new_n18206_ = ~new_n17718_ | ~new_n15597_;
  assign new_n18207_ = ~new_n17419_ | ~new_n15592_;
  assign new_n18208_ = ~new_n18185_ | ~new_n15591_;
  assign new_n18209_ = ~new_n15577_ | ~new_n18200_;
  assign new_n18210_ = ~pi1142 | ~new_n18195_;
  assign new_n18211_ = ~new_n17718_ | ~new_n15601_;
  assign new_n18212_ = ~new_n17419_ | ~new_n15590_;
  assign new_n18213_ = ~new_n18185_ | ~new_n15589_;
  assign new_n18214_ = ~new_n15576_ | ~new_n18200_;
  assign new_n18215_ = ~pi1143 | ~new_n18195_;
  assign new_n18216_ = ~new_n17718_ | ~new_n15600_;
  assign new_n18217_ = ~new_n17419_ | ~new_n15588_;
  assign new_n18218_ = ~new_n18185_ | ~new_n15587_;
  assign new_n18219_ = ~new_n15575_ | ~new_n18200_;
  assign new_n18220_ = ~pi1144 | ~new_n18195_;
  assign new_n18221_ = ~new_n17718_ | ~new_n15599_;
  assign new_n18222_ = ~new_n17419_ | ~new_n15586_;
  assign new_n18223_ = ~new_n18185_ | ~new_n15585_;
  assign new_n18224_ = ~new_n15574_ | ~new_n18200_;
  assign new_n18225_ = ~pi1145 | ~new_n18195_;
  assign new_n18226_ = ~new_n17718_ | ~new_n15602_;
  assign new_n18227_ = ~new_n17419_ | ~new_n15584_;
  assign new_n18228_ = ~new_n18185_ | ~new_n15583_;
  assign new_n18229_ = ~new_n15573_ | ~new_n18200_;
  assign new_n18230_ = ~pi1146 | ~new_n18195_;
  assign new_n18231_ = ~new_n17718_ | ~new_n15595_;
  assign new_n18232_ = ~new_n17419_ | ~new_n15582_;
  assign new_n18233_ = ~new_n18185_ | ~new_n15581_;
  assign new_n18234_ = ~new_n15572_ | ~new_n18200_;
  assign new_n18235_ = ~pi1147 | ~new_n18195_;
  assign new_n18236_ = ~new_n17718_ | ~new_n15598_;
  assign new_n18237_ = ~new_n17419_ | ~new_n15580_;
  assign new_n18238_ = ~new_n18185_ | ~new_n15579_;
  assign new_n18239_ = ~new_n15571_ | ~new_n18200_;
  assign new_n18240_ = ~pi1148 | ~new_n18195_;
  assign new_n18241_ = ~new_n16545_;
  assign new_n18242_ = ~new_n16544_;
  assign new_n18243_ = ~new_n15620_ | ~new_n15624_;
  assign new_n18244_ = ~new_n16546_;
  assign new_n18245_ = ~new_n16421_;
  assign new_n18246_ = ~new_n17705_ | ~new_n15655_;
  assign new_n18247_ = ~new_n15683_ | ~new_n15539_;
  assign new_n18248_ = ~new_n16501_ | ~new_n18247_;
  assign new_n18249_ = ~new_n18244_ | ~new_n18248_;
  assign new_n18250_ = ~pi1073 | ~new_n16544_;
  assign new_n18251_ = ~pi1074 | ~new_n16421_;
  assign new_n18252_ = ~new_n18249_ | ~new_n16849_;
  assign new_n18253_ = ~new_n15683_ | ~new_n15569_;
  assign new_n18254_ = ~new_n16501_ | ~new_n18253_;
  assign new_n18255_ = ~new_n18254_ | ~new_n16546_;
  assign new_n18256_ = ~pi1074 | ~new_n18245_;
  assign new_n18257_ = ~new_n18256_ | ~new_n18255_;
  assign new_n18258_ = ~new_n18242_ | ~new_n15596_;
  assign new_n18259_ = ~new_n15682_ | ~new_n15594_;
  assign new_n18260_ = ~new_n18241_ | ~new_n15593_;
  assign new_n18261_ = ~new_n15578_ | ~new_n18257_;
  assign new_n18262_ = ~pi1149 | ~new_n18252_;
  assign new_n18263_ = ~new_n18242_ | ~new_n15597_;
  assign new_n18264_ = ~new_n15682_ | ~new_n15592_;
  assign new_n18265_ = ~new_n18241_ | ~new_n15591_;
  assign new_n18266_ = ~new_n15577_ | ~new_n18257_;
  assign new_n18267_ = ~pi1150 | ~new_n18252_;
  assign new_n18268_ = ~new_n18242_ | ~new_n15601_;
  assign new_n18269_ = ~new_n15682_ | ~new_n15590_;
  assign new_n18270_ = ~new_n18241_ | ~new_n15589_;
  assign new_n18271_ = ~new_n15576_ | ~new_n18257_;
  assign new_n18272_ = ~pi1151 | ~new_n18252_;
  assign new_n18273_ = ~new_n18242_ | ~new_n15600_;
  assign new_n18274_ = ~new_n15682_ | ~new_n15588_;
  assign new_n18275_ = ~new_n18241_ | ~new_n15587_;
  assign new_n18276_ = ~new_n15575_ | ~new_n18257_;
  assign new_n18277_ = ~pi1152 | ~new_n18252_;
  assign new_n18278_ = ~new_n18242_ | ~new_n15599_;
  assign new_n18279_ = ~new_n15682_ | ~new_n15586_;
  assign new_n18280_ = ~new_n18241_ | ~new_n15585_;
  assign new_n18281_ = ~new_n15574_ | ~new_n18257_;
  assign new_n18282_ = ~pi1153 | ~new_n18252_;
  assign new_n18283_ = ~new_n18242_ | ~new_n15602_;
  assign new_n18284_ = ~new_n15682_ | ~new_n15584_;
  assign new_n18285_ = ~new_n18241_ | ~new_n15583_;
  assign new_n18286_ = ~new_n15573_ | ~new_n18257_;
  assign new_n18287_ = ~pi1154 | ~new_n18252_;
  assign new_n18288_ = ~new_n18242_ | ~new_n15595_;
  assign new_n18289_ = ~new_n15682_ | ~new_n15582_;
  assign new_n18290_ = ~new_n18241_ | ~new_n15581_;
  assign new_n18291_ = ~new_n15572_ | ~new_n18257_;
  assign new_n18292_ = ~pi1155 | ~new_n18252_;
  assign new_n18293_ = ~new_n18242_ | ~new_n15598_;
  assign new_n18294_ = ~new_n15682_ | ~new_n15580_;
  assign new_n18295_ = ~new_n18241_ | ~new_n15579_;
  assign new_n18296_ = ~new_n15571_ | ~new_n18257_;
  assign new_n18297_ = ~pi1156 | ~new_n18252_;
  assign new_n18298_ = ~new_n16548_;
  assign new_n18299_ = ~new_n16547_;
  assign new_n18300_ = ~new_n15620_ | ~new_n15625_;
  assign new_n18301_ = ~new_n16549_;
  assign new_n18302_ = ~new_n15614_ | ~new_n15618_;
  assign new_n18303_ = ~new_n16550_;
  assign new_n18304_ = ~new_n17706_ | ~new_n15655_;
  assign new_n18305_ = ~new_n15685_ | ~new_n15539_;
  assign new_n18306_ = ~new_n16501_ | ~new_n18305_;
  assign new_n18307_ = ~new_n18301_ | ~new_n18306_;
  assign new_n18308_ = ~pi1073 | ~new_n16547_;
  assign new_n18309_ = ~new_n18303_ | ~pi1074;
  assign new_n18310_ = ~new_n18307_ | ~new_n16858_;
  assign new_n18311_ = ~new_n15685_ | ~new_n15569_;
  assign new_n18312_ = ~new_n16501_ | ~new_n18311_;
  assign new_n18313_ = ~new_n18312_ | ~new_n16549_;
  assign new_n18314_ = ~pi1074 | ~new_n16550_;
  assign new_n18315_ = ~new_n18314_ | ~new_n18313_;
  assign new_n18316_ = ~new_n18299_ | ~new_n15596_;
  assign new_n18317_ = ~new_n15684_ | ~new_n15594_;
  assign new_n18318_ = ~new_n18298_ | ~new_n15593_;
  assign new_n18319_ = ~new_n15578_ | ~new_n18315_;
  assign new_n18320_ = ~pi1157 | ~new_n18310_;
  assign new_n18321_ = ~new_n18299_ | ~new_n15597_;
  assign new_n18322_ = ~new_n15684_ | ~new_n15592_;
  assign new_n18323_ = ~new_n18298_ | ~new_n15591_;
  assign new_n18324_ = ~new_n15577_ | ~new_n18315_;
  assign new_n18325_ = ~pi1158 | ~new_n18310_;
  assign new_n18326_ = ~new_n18299_ | ~new_n15601_;
  assign new_n18327_ = ~new_n15684_ | ~new_n15590_;
  assign new_n18328_ = ~new_n18298_ | ~new_n15589_;
  assign new_n18329_ = ~new_n15576_ | ~new_n18315_;
  assign new_n18330_ = ~pi1159 | ~new_n18310_;
  assign new_n18331_ = ~new_n18299_ | ~new_n15600_;
  assign new_n18332_ = ~new_n15684_ | ~new_n15588_;
  assign new_n18333_ = ~new_n18298_ | ~new_n15587_;
  assign new_n18334_ = ~new_n15575_ | ~new_n18315_;
  assign new_n18335_ = ~pi1160 | ~new_n18310_;
  assign new_n18336_ = ~new_n18299_ | ~new_n15599_;
  assign new_n18337_ = ~new_n15684_ | ~new_n15586_;
  assign new_n18338_ = ~new_n18298_ | ~new_n15585_;
  assign new_n18339_ = ~new_n15574_ | ~new_n18315_;
  assign new_n18340_ = ~pi1161 | ~new_n18310_;
  assign new_n18341_ = ~new_n18299_ | ~new_n15602_;
  assign new_n18342_ = ~new_n15684_ | ~new_n15584_;
  assign new_n18343_ = ~new_n18298_ | ~new_n15583_;
  assign new_n18344_ = ~new_n15573_ | ~new_n18315_;
  assign new_n18345_ = ~pi1162 | ~new_n18310_;
  assign new_n18346_ = ~new_n18299_ | ~new_n15595_;
  assign new_n18347_ = ~new_n15684_ | ~new_n15582_;
  assign new_n18348_ = ~new_n18298_ | ~new_n15581_;
  assign new_n18349_ = ~new_n15572_ | ~new_n18315_;
  assign new_n18350_ = ~pi1163 | ~new_n18310_;
  assign new_n18351_ = ~new_n18299_ | ~new_n15598_;
  assign new_n18352_ = ~new_n15684_ | ~new_n15580_;
  assign new_n18353_ = ~new_n18298_ | ~new_n15579_;
  assign new_n18354_ = ~new_n15571_ | ~new_n18315_;
  assign new_n18355_ = ~pi1164 | ~new_n18310_;
  assign new_n18356_ = ~new_n16552_;
  assign new_n18357_ = ~new_n16551_;
  assign new_n18358_ = ~new_n15620_ | ~new_n15626_;
  assign new_n18359_ = ~new_n16553_;
  assign new_n18360_ = ~new_n16422_;
  assign new_n18361_ = ~new_n15667_ | ~new_n15655_;
  assign new_n18362_ = ~new_n15687_ | ~new_n15539_;
  assign new_n18363_ = ~new_n16501_ | ~new_n18362_;
  assign new_n18364_ = ~new_n18359_ | ~new_n18363_;
  assign new_n18365_ = ~pi1073 | ~new_n16551_;
  assign new_n18366_ = ~pi1074 | ~new_n16422_;
  assign new_n18367_ = ~new_n18364_ | ~new_n16867_;
  assign new_n18368_ = ~new_n15687_ | ~new_n15569_;
  assign new_n18369_ = ~new_n16501_ | ~new_n18368_;
  assign new_n18370_ = ~new_n18369_ | ~new_n16553_;
  assign new_n18371_ = ~pi1074 | ~new_n18360_;
  assign new_n18372_ = ~new_n18371_ | ~new_n18370_;
  assign new_n18373_ = ~new_n18357_ | ~new_n15596_;
  assign new_n18374_ = ~new_n15686_ | ~new_n15594_;
  assign new_n18375_ = ~new_n18356_ | ~new_n15593_;
  assign new_n18376_ = ~new_n15578_ | ~new_n18372_;
  assign new_n18377_ = ~pi1165 | ~new_n18367_;
  assign new_n18378_ = ~new_n18357_ | ~new_n15597_;
  assign new_n18379_ = ~new_n15686_ | ~new_n15592_;
  assign new_n18380_ = ~new_n18356_ | ~new_n15591_;
  assign new_n18381_ = ~new_n15577_ | ~new_n18372_;
  assign new_n18382_ = ~pi1166 | ~new_n18367_;
  assign new_n18383_ = ~new_n18357_ | ~new_n15601_;
  assign new_n18384_ = ~new_n15686_ | ~new_n15590_;
  assign new_n18385_ = ~new_n18356_ | ~new_n15589_;
  assign new_n18386_ = ~new_n15576_ | ~new_n18372_;
  assign new_n18387_ = ~pi1167 | ~new_n18367_;
  assign new_n18388_ = ~new_n18357_ | ~new_n15600_;
  assign new_n18389_ = ~new_n15686_ | ~new_n15588_;
  assign new_n18390_ = ~new_n18356_ | ~new_n15587_;
  assign new_n18391_ = ~new_n15575_ | ~new_n18372_;
  assign new_n18392_ = ~pi1168 | ~new_n18367_;
  assign new_n18393_ = ~new_n18357_ | ~new_n15599_;
  assign new_n18394_ = ~new_n15686_ | ~new_n15586_;
  assign new_n18395_ = ~new_n18356_ | ~new_n15585_;
  assign new_n18396_ = ~new_n15574_ | ~new_n18372_;
  assign new_n18397_ = ~pi1169 | ~new_n18367_;
  assign new_n18398_ = ~new_n18357_ | ~new_n15602_;
  assign new_n18399_ = ~new_n15686_ | ~new_n15584_;
  assign new_n18400_ = ~new_n18356_ | ~new_n15583_;
  assign new_n18401_ = ~new_n15573_ | ~new_n18372_;
  assign new_n18402_ = ~pi1170 | ~new_n18367_;
  assign new_n18403_ = ~new_n18357_ | ~new_n15595_;
  assign new_n18404_ = ~new_n15686_ | ~new_n15582_;
  assign new_n18405_ = ~new_n18356_ | ~new_n15581_;
  assign new_n18406_ = ~new_n15572_ | ~new_n18372_;
  assign new_n18407_ = ~pi1171 | ~new_n18367_;
  assign new_n18408_ = ~new_n18357_ | ~new_n15598_;
  assign new_n18409_ = ~new_n15686_ | ~new_n15580_;
  assign new_n18410_ = ~new_n18356_ | ~new_n15579_;
  assign new_n18411_ = ~new_n15571_ | ~new_n18372_;
  assign new_n18412_ = ~pi1172 | ~new_n18367_;
  assign new_n18413_ = ~new_n16555_;
  assign new_n18414_ = ~new_n16554_;
  assign new_n18415_ = ~new_n15622_ | ~new_n15623_;
  assign new_n18416_ = ~new_n16556_;
  assign new_n18417_ = ~new_n15616_ | ~new_n15617_;
  assign new_n18418_ = ~new_n16557_;
  assign new_n18419_ = ~new_n15689_ | ~new_n17709_;
  assign new_n18420_ = ~new_n15692_ | ~new_n15539_;
  assign new_n18421_ = ~new_n16501_ | ~new_n18420_;
  assign new_n18422_ = ~new_n18416_ | ~new_n18421_;
  assign new_n18423_ = ~pi1073 | ~new_n16554_;
  assign new_n18424_ = ~new_n18418_ | ~pi1074;
  assign new_n18425_ = ~new_n18422_ | ~new_n16876_;
  assign new_n18426_ = ~new_n15692_ | ~new_n15569_;
  assign new_n18427_ = ~new_n16501_ | ~new_n18426_;
  assign new_n18428_ = ~new_n18427_ | ~new_n16556_;
  assign new_n18429_ = ~pi1074 | ~new_n16557_;
  assign new_n18430_ = ~new_n18429_ | ~new_n18428_;
  assign new_n18431_ = ~new_n18414_ | ~new_n15596_;
  assign new_n18432_ = ~new_n15690_ | ~new_n15594_;
  assign new_n18433_ = ~new_n18413_ | ~new_n15593_;
  assign new_n18434_ = ~new_n15578_ | ~new_n18430_;
  assign new_n18435_ = ~pi1173 | ~new_n18425_;
  assign new_n18436_ = ~new_n18414_ | ~new_n15597_;
  assign new_n18437_ = ~new_n15690_ | ~new_n15592_;
  assign new_n18438_ = ~new_n18413_ | ~new_n15591_;
  assign new_n18439_ = ~new_n15577_ | ~new_n18430_;
  assign new_n18440_ = ~pi1174 | ~new_n18425_;
  assign new_n18441_ = ~new_n18414_ | ~new_n15601_;
  assign new_n18442_ = ~new_n15690_ | ~new_n15590_;
  assign new_n18443_ = ~new_n18413_ | ~new_n15589_;
  assign new_n18444_ = ~new_n15576_ | ~new_n18430_;
  assign new_n18445_ = ~pi1175 | ~new_n18425_;
  assign new_n18446_ = ~new_n18414_ | ~new_n15600_;
  assign new_n18447_ = ~new_n15690_ | ~new_n15588_;
  assign new_n18448_ = ~new_n18413_ | ~new_n15587_;
  assign new_n18449_ = ~new_n15575_ | ~new_n18430_;
  assign new_n18450_ = ~pi1176 | ~new_n18425_;
  assign new_n18451_ = ~new_n18414_ | ~new_n15599_;
  assign new_n18452_ = ~new_n15690_ | ~new_n15586_;
  assign new_n18453_ = ~new_n18413_ | ~new_n15585_;
  assign new_n18454_ = ~new_n15574_ | ~new_n18430_;
  assign new_n18455_ = ~pi1177 | ~new_n18425_;
  assign new_n18456_ = ~new_n18414_ | ~new_n15602_;
  assign new_n18457_ = ~new_n15690_ | ~new_n15584_;
  assign new_n18458_ = ~new_n18413_ | ~new_n15583_;
  assign new_n18459_ = ~new_n15573_ | ~new_n18430_;
  assign new_n18460_ = ~pi1178 | ~new_n18425_;
  assign new_n18461_ = ~new_n18414_ | ~new_n15595_;
  assign new_n18462_ = ~new_n15690_ | ~new_n15582_;
  assign new_n18463_ = ~new_n18413_ | ~new_n15581_;
  assign new_n18464_ = ~new_n15572_ | ~new_n18430_;
  assign new_n18465_ = ~pi1179 | ~new_n18425_;
  assign new_n18466_ = ~new_n18414_ | ~new_n15598_;
  assign new_n18467_ = ~new_n15690_ | ~new_n15580_;
  assign new_n18468_ = ~new_n18413_ | ~new_n15579_;
  assign new_n18469_ = ~new_n15571_ | ~new_n18430_;
  assign new_n18470_ = ~pi1180 | ~new_n18425_;
  assign new_n18471_ = ~new_n16559_;
  assign new_n18472_ = ~new_n16558_;
  assign new_n18473_ = ~new_n15622_ | ~new_n15624_;
  assign new_n18474_ = ~new_n16560_;
  assign new_n18475_ = ~new_n16423_;
  assign new_n18476_ = ~new_n15689_ | ~new_n17705_;
  assign new_n18477_ = ~new_n15694_ | ~new_n15539_;
  assign new_n18478_ = ~new_n16501_ | ~new_n18477_;
  assign new_n18479_ = ~new_n18474_ | ~new_n18478_;
  assign new_n18480_ = ~pi1073 | ~new_n16558_;
  assign new_n18481_ = ~pi1074 | ~new_n16423_;
  assign new_n18482_ = ~new_n18479_ | ~new_n16885_;
  assign new_n18483_ = ~new_n15694_ | ~new_n15569_;
  assign new_n18484_ = ~new_n16501_ | ~new_n18483_;
  assign new_n18485_ = ~new_n18484_ | ~new_n16560_;
  assign new_n18486_ = ~pi1074 | ~new_n18475_;
  assign new_n18487_ = ~new_n18486_ | ~new_n18485_;
  assign new_n18488_ = ~new_n18472_ | ~new_n15596_;
  assign new_n18489_ = ~new_n15693_ | ~new_n15594_;
  assign new_n18490_ = ~new_n18471_ | ~new_n15593_;
  assign new_n18491_ = ~new_n15578_ | ~new_n18487_;
  assign new_n18492_ = ~pi1181 | ~new_n18482_;
  assign new_n18493_ = ~new_n18472_ | ~new_n15597_;
  assign new_n18494_ = ~new_n15693_ | ~new_n15592_;
  assign new_n18495_ = ~new_n18471_ | ~new_n15591_;
  assign new_n18496_ = ~new_n15577_ | ~new_n18487_;
  assign new_n18497_ = ~pi1182 | ~new_n18482_;
  assign new_n18498_ = ~new_n18472_ | ~new_n15601_;
  assign new_n18499_ = ~new_n15693_ | ~new_n15590_;
  assign new_n18500_ = ~new_n18471_ | ~new_n15589_;
  assign new_n18501_ = ~new_n15576_ | ~new_n18487_;
  assign new_n18502_ = ~pi1183 | ~new_n18482_;
  assign new_n18503_ = ~new_n18472_ | ~new_n15600_;
  assign new_n18504_ = ~new_n15693_ | ~new_n15588_;
  assign new_n18505_ = ~new_n18471_ | ~new_n15587_;
  assign new_n18506_ = ~new_n15575_ | ~new_n18487_;
  assign new_n18507_ = ~pi1184 | ~new_n18482_;
  assign new_n18508_ = ~new_n18472_ | ~new_n15599_;
  assign new_n18509_ = ~new_n15693_ | ~new_n15586_;
  assign new_n18510_ = ~new_n18471_ | ~new_n15585_;
  assign new_n18511_ = ~new_n15574_ | ~new_n18487_;
  assign new_n18512_ = ~pi1185 | ~new_n18482_;
  assign new_n18513_ = ~new_n18472_ | ~new_n15602_;
  assign new_n18514_ = ~new_n15693_ | ~new_n15584_;
  assign new_n18515_ = ~new_n18471_ | ~new_n15583_;
  assign new_n18516_ = ~new_n15573_ | ~new_n18487_;
  assign new_n18517_ = ~pi1186 | ~new_n18482_;
  assign new_n18518_ = ~new_n18472_ | ~new_n15595_;
  assign new_n18519_ = ~new_n15693_ | ~new_n15582_;
  assign new_n18520_ = ~new_n18471_ | ~new_n15581_;
  assign new_n18521_ = ~new_n15572_ | ~new_n18487_;
  assign new_n18522_ = ~pi1187 | ~new_n18482_;
  assign new_n18523_ = ~new_n18472_ | ~new_n15598_;
  assign new_n18524_ = ~new_n15693_ | ~new_n15580_;
  assign new_n18525_ = ~new_n18471_ | ~new_n15579_;
  assign new_n18526_ = ~new_n15571_ | ~new_n18487_;
  assign new_n18527_ = ~pi1188 | ~new_n18482_;
  assign new_n18528_ = ~new_n16562_;
  assign new_n18529_ = ~new_n16561_;
  assign new_n18530_ = ~new_n15622_ | ~new_n15625_;
  assign new_n18531_ = ~new_n16563_;
  assign new_n18532_ = ~new_n15616_ | ~new_n15618_;
  assign new_n18533_ = ~new_n16564_;
  assign new_n18534_ = ~new_n15689_ | ~new_n17706_;
  assign new_n18535_ = ~new_n15696_ | ~new_n15539_;
  assign new_n18536_ = ~new_n16501_ | ~new_n18535_;
  assign new_n18537_ = ~new_n18531_ | ~new_n18536_;
  assign new_n18538_ = ~pi1073 | ~new_n16561_;
  assign new_n18539_ = ~new_n18533_ | ~pi1074;
  assign new_n18540_ = ~new_n18537_ | ~new_n16894_;
  assign new_n18541_ = ~new_n15696_ | ~new_n15569_;
  assign new_n18542_ = ~new_n16501_ | ~new_n18541_;
  assign new_n18543_ = ~new_n18542_ | ~new_n16563_;
  assign new_n18544_ = ~pi1074 | ~new_n16564_;
  assign new_n18545_ = ~new_n18544_ | ~new_n18543_;
  assign new_n18546_ = ~new_n18529_ | ~new_n15596_;
  assign new_n18547_ = ~new_n15695_ | ~new_n15594_;
  assign new_n18548_ = ~new_n18528_ | ~new_n15593_;
  assign new_n18549_ = ~new_n15578_ | ~new_n18545_;
  assign new_n18550_ = ~pi1189 | ~new_n18540_;
  assign new_n18551_ = ~new_n18529_ | ~new_n15597_;
  assign new_n18552_ = ~new_n15695_ | ~new_n15592_;
  assign new_n18553_ = ~new_n18528_ | ~new_n15591_;
  assign new_n18554_ = ~new_n15577_ | ~new_n18545_;
  assign new_n18555_ = ~pi1190 | ~new_n18540_;
  assign new_n18556_ = ~new_n18529_ | ~new_n15601_;
  assign new_n18557_ = ~new_n15695_ | ~new_n15590_;
  assign new_n18558_ = ~new_n18528_ | ~new_n15589_;
  assign new_n18559_ = ~new_n15576_ | ~new_n18545_;
  assign new_n18560_ = ~pi1191 | ~new_n18540_;
  assign new_n18561_ = ~new_n18529_ | ~new_n15600_;
  assign new_n18562_ = ~new_n15695_ | ~new_n15588_;
  assign new_n18563_ = ~new_n18528_ | ~new_n15587_;
  assign new_n18564_ = ~new_n15575_ | ~new_n18545_;
  assign new_n18565_ = ~pi1192 | ~new_n18540_;
  assign new_n18566_ = ~new_n18529_ | ~new_n15599_;
  assign new_n18567_ = ~new_n15695_ | ~new_n15586_;
  assign new_n18568_ = ~new_n18528_ | ~new_n15585_;
  assign new_n18569_ = ~new_n15574_ | ~new_n18545_;
  assign new_n18570_ = ~pi1193 | ~new_n18540_;
  assign new_n18571_ = ~new_n18529_ | ~new_n15602_;
  assign new_n18572_ = ~new_n15695_ | ~new_n15584_;
  assign new_n18573_ = ~new_n18528_ | ~new_n15583_;
  assign new_n18574_ = ~new_n15573_ | ~new_n18545_;
  assign new_n18575_ = ~pi1194 | ~new_n18540_;
  assign new_n18576_ = ~new_n18529_ | ~new_n15595_;
  assign new_n18577_ = ~new_n15695_ | ~new_n15582_;
  assign new_n18578_ = ~new_n18528_ | ~new_n15581_;
  assign new_n18579_ = ~new_n15572_ | ~new_n18545_;
  assign new_n18580_ = ~pi1195 | ~new_n18540_;
  assign new_n18581_ = ~new_n18529_ | ~new_n15598_;
  assign new_n18582_ = ~new_n15695_ | ~new_n15580_;
  assign new_n18583_ = ~new_n18528_ | ~new_n15579_;
  assign new_n18584_ = ~new_n15571_ | ~new_n18545_;
  assign new_n18585_ = ~pi1196 | ~new_n18540_;
  assign new_n18586_ = ~new_n16566_;
  assign new_n18587_ = ~new_n16565_;
  assign new_n18588_ = ~new_n15622_ | ~new_n15626_;
  assign new_n18589_ = ~new_n16567_;
  assign new_n18590_ = ~new_n16424_;
  assign new_n18591_ = ~new_n15689_ | ~new_n15667_;
  assign new_n18592_ = ~new_n15698_ | ~new_n15539_;
  assign new_n18593_ = ~new_n16501_ | ~new_n18592_;
  assign new_n18594_ = ~new_n18589_ | ~new_n18593_;
  assign new_n18595_ = ~pi1073 | ~new_n16565_;
  assign new_n18596_ = ~pi1074 | ~new_n16424_;
  assign new_n18597_ = ~new_n18594_ | ~new_n16903_;
  assign new_n18598_ = ~new_n15698_ | ~new_n15569_;
  assign new_n18599_ = ~new_n16501_ | ~new_n18598_;
  assign new_n18600_ = ~new_n18599_ | ~new_n16567_;
  assign new_n18601_ = ~pi1074 | ~new_n18590_;
  assign new_n18602_ = ~new_n18601_ | ~new_n18600_;
  assign new_n18603_ = ~new_n18587_ | ~new_n15596_;
  assign new_n18604_ = ~new_n15697_ | ~new_n15594_;
  assign new_n18605_ = ~new_n18586_ | ~new_n15593_;
  assign new_n18606_ = ~new_n15578_ | ~new_n18602_;
  assign new_n18607_ = ~pi1197 | ~new_n18597_;
  assign new_n18608_ = ~new_n18587_ | ~new_n15597_;
  assign new_n18609_ = ~new_n15697_ | ~new_n15592_;
  assign new_n18610_ = ~new_n18586_ | ~new_n15591_;
  assign new_n18611_ = ~new_n15577_ | ~new_n18602_;
  assign new_n18612_ = ~pi1198 | ~new_n18597_;
  assign new_n18613_ = ~new_n18587_ | ~new_n15601_;
  assign new_n18614_ = ~new_n15697_ | ~new_n15590_;
  assign new_n18615_ = ~new_n18586_ | ~new_n15589_;
  assign new_n18616_ = ~new_n15576_ | ~new_n18602_;
  assign new_n18617_ = ~pi1199 | ~new_n18597_;
  assign new_n18618_ = ~new_n18587_ | ~new_n15600_;
  assign new_n18619_ = ~new_n15697_ | ~new_n15588_;
  assign new_n18620_ = ~new_n18586_ | ~new_n15587_;
  assign new_n18621_ = ~new_n15575_ | ~new_n18602_;
  assign new_n18622_ = ~new_n18587_ | ~new_n15599_;
  assign new_n18623_ = ~new_n15697_ | ~new_n15586_;
  assign new_n18624_ = ~new_n18586_ | ~new_n15585_;
  assign new_n18625_ = ~new_n15574_ | ~new_n18602_;
  assign new_n18626_ = ~pi1201 | ~new_n18597_;
  assign new_n18627_ = ~new_n18587_ | ~new_n15602_;
  assign new_n18628_ = ~new_n15697_ | ~new_n15584_;
  assign new_n18629_ = ~new_n18586_ | ~new_n15583_;
  assign new_n18630_ = ~new_n15573_ | ~new_n18602_;
  assign new_n18631_ = ~pi1202 | ~new_n18597_;
  assign new_n18632_ = ~new_n18587_ | ~new_n15595_;
  assign new_n18633_ = ~new_n15697_ | ~new_n15582_;
  assign new_n18634_ = ~new_n18586_ | ~new_n15581_;
  assign new_n18635_ = ~new_n15572_ | ~new_n18602_;
  assign new_n18636_ = ~pi1203 | ~new_n18597_;
  assign new_n18637_ = ~new_n18587_ | ~new_n15598_;
  assign new_n18638_ = ~new_n15697_ | ~new_n15580_;
  assign new_n18639_ = ~new_n18586_ | ~new_n15579_;
  assign new_n18640_ = ~new_n15571_ | ~new_n18602_;
  assign new_n18641_ = ~pi1204 | ~new_n18597_;
  assign new_n18642_ = ~new_n16604_;
  assign new_n18643_ = ~new_n17684_ | ~new_n16572_ | ~new_n16575_;
  assign new_n18644_ = ~new_n17641_ | ~new_n17581_ | ~new_n17354_;
  assign new_n18645_ = ~new_n16425_;
  assign new_n18646_ = ~new_n17675_ | ~new_n16470_;
  assign new_n18647_ = ~new_n18645_ | ~new_n18646_ | ~new_n16464_;
  assign new_n18648_ = ~new_n16913_ | ~new_n15633_;
  assign new_n18649_ = ~new_n17389_ | ~new_n18643_;
  assign new_n18650_ = ~new_n16914_ | ~new_n20790_;
  assign new_n18651_ = ~new_n9378_ | ~new_n17396_ | ~new_n16438_;
  assign new_n18652_ = ~new_n15630_ | ~new_n20675_;
  assign new_n18653_ = ~new_n17438_ | ~new_n17684_;
  assign new_n18654_ = ~new_n17363_;
  assign new_n18655_ = ~new_n15549_ | ~new_n17363_;
  assign new_n18656_ = ~pi1073 | ~new_n16475_;
  assign new_n18657_ = ~new_n17353_;
  assign new_n18658_ = ~pi1208 | ~pi1207;
  assign new_n18659_ = ~pi1206 | ~new_n18658_;
  assign new_n18660_ = ~new_n17562_ | ~pi1208;
  assign new_n18661_ = ~new_n16623_;
  assign new_n18662_ = ~new_n16679_ | ~pi1207;
  assign new_n18663_ = ~pi1206 | ~new_n18662_;
  assign new_n18664_ = ~new_n16619_;
  assign new_n18665_ = ~new_n16456_ | ~new_n16445_;
  assign new_n18666_ = ~pi1206 | ~new_n18665_;
  assign new_n18667_ = ~new_n15650_ | ~new_n16456_;
  assign new_n18668_ = ~new_n17675_ | ~new_n16471_;
  assign new_n18669_ = ~new_n17581_ | ~new_n15786_;
  assign new_n18670_ = ~new_n20675_ | ~new_n20885_ | ~new_n20884_;
  assign new_n18671_ = ~new_n17630_ | ~new_n18669_;
  assign new_n18672_ = ~new_n16590_ | ~new_n17581_ | ~new_n16575_;
  assign new_n18673_ = ~new_n18672_ | ~new_n17352_;
  assign new_n18674_ = ~new_n20810_ | ~new_n18673_;
  assign new_n18675_ = ~new_n17641_ | ~new_n17352_;
  assign new_n18676_ = ~new_n16576_ | ~new_n18675_;
  assign new_n18677_ = ~new_n17389_ | ~new_n18643_;
  assign new_n18678_ = ~new_n17438_ | ~new_n17684_;
  assign new_n18679_ = ~new_n18676_ | ~new_n16452_;
  assign new_n18680_ = ~new_n17675_ | ~new_n20888_;
  assign new_n18681_ = ~new_n17371_ | ~new_n16425_;
  assign new_n18682_ = ~new_n16473_ | ~new_n17398_;
  assign new_n18683_ = ~new_n16921_ | ~new_n18682_;
  assign new_n18684_ = ~new_n31170_ | ~new_n20690_;
  assign new_n18685_ = ~new_n17399_ | ~new_n16619_;
  assign new_n18686_ = ~new_n17395_ | ~new_n16623_;
  assign new_n18687_ = ~new_n18684_ | ~new_n16928_;
  assign new_n18688_ = ~new_n17433_ | ~new_n16619_;
  assign new_n18689_ = ~new_n15608_ | ~new_n18687_;
  assign new_n18690_ = ~new_n18689_ | ~new_n18688_;
  assign new_n18691_ = ~pi1207 | ~new_n16456_;
  assign new_n18692_ = ~new_n16582_;
  assign new_n18693_ = ~new_n31187_ | ~new_n20690_;
  assign new_n18694_ = ~new_n17395_ | ~new_n16637_;
  assign new_n18695_ = ~new_n16930_ | ~new_n18693_;
  assign new_n18696_ = ~new_n15627_ | ~new_n16651_;
  assign new_n18697_ = ~new_n17433_ | ~new_n16582_;
  assign new_n18698_ = ~new_n15608_ | ~new_n18695_;
  assign new_n18699_ = ~new_n18697_ | ~new_n18698_ | ~new_n18696_;
  assign new_n18700_ = ~new_n16583_;
  assign new_n18701_ = ~new_n15612_ | ~new_n17430_;
  assign new_n18702_ = ~new_n16473_ | ~new_n18701_;
  assign new_n18703_ = ~new_n18700_ | ~new_n18702_;
  assign new_n18704_ = ~new_n31178_ | ~new_n20690_;
  assign new_n18705_ = ~new_n17395_ | ~new_n16446_;
  assign new_n18706_ = ~new_n16931_ | ~new_n18704_;
  assign new_n18707_ = ~new_n20893_ | ~new_n15627_;
  assign new_n18708_ = ~new_n18700_ | ~new_n17433_;
  assign new_n18709_ = ~new_n15608_ | ~new_n18706_;
  assign new_n18710_ = ~new_n18708_ | ~new_n18709_ | ~new_n18707_;
  assign new_n18711_ = ~new_n31179_ | ~new_n20690_;
  assign new_n18712_ = ~new_n17356_ | ~new_n18711_;
  assign new_n18713_ = ~new_n17433_ | ~new_n16447_;
  assign new_n18714_ = ~new_n15608_ | ~new_n18712_;
  assign new_n18715_ = ~new_n20896_ | ~pi1075;
  assign new_n18716_ = ~new_n18713_ | ~new_n18714_ | ~new_n18715_;
  assign new_n18717_ = ~new_n32701_ | ~new_n15609_ | ~pi1076;
  assign new_n18718_ = ~new_n16585_;
  assign new_n18719_ = ~pi1075 | ~new_n16477_;
  assign new_n18720_ = ~new_n17708_ | ~new_n16635_;
  assign new_n18721_ = ~new_n16539_ | ~new_n18720_;
  assign new_n18722_ = ~new_n16540_ | ~new_n18721_;
  assign new_n18723_ = ~new_n15569_ | ~new_n18722_;
  assign new_n18724_ = ~new_n31170_ | ~new_n18719_;
  assign new_n18725_ = ~new_n17407_ | ~new_n31235_;
  assign new_n18726_ = ~new_n16932_ | ~new_n18723_;
  assign new_n18727_ = ~new_n15569_ | ~new_n20914_;
  assign new_n18728_ = ~new_n31187_ | ~new_n18719_;
  assign new_n18729_ = ~new_n17407_ | ~new_n31276_;
  assign new_n18730_ = ~new_n16933_ | ~new_n18727_;
  assign new_n18731_ = ~new_n16507_ | ~new_n16514_;
  assign new_n18732_ = ~new_n15569_ | ~new_n18731_;
  assign new_n18733_ = ~new_n31178_ | ~new_n18719_;
  assign new_n18734_ = ~new_n17407_ | ~new_n31277_;
  assign new_n18735_ = ~new_n16934_ | ~new_n18732_;
  assign new_n18736_ = ~new_n31179_ | ~new_n18719_;
  assign new_n18737_ = ~new_n31270_ | ~new_n17390_;
  assign new_n18738_ = ~new_n17426_ | ~new_n18736_ | ~new_n18737_;
  assign new_n18739_ = ~new_n17658_ | ~new_n16453_;
  assign new_n18740_ = ~new_n17441_ | ~new_n15612_;
  assign new_n18741_ = ~new_n18740_ | ~new_n20923_ | ~new_n20924_ | ~new_n15699_;
  assign new_n18742_ = ~new_n17373_ | ~new_n17416_ | ~new_n17684_;
  assign new_n18743_ = ~new_n15549_ | ~new_n18741_;
  assign new_n18744_ = ~new_n17384_ | ~new_n16444_;
  assign new_n18745_ = ~new_n16595_;
  assign new_n18746_ = ~new_n17443_ | ~new_n17389_;
  assign new_n18747_ = ~new_n17437_ | ~new_n15570_;
  assign new_n18748_ = ~new_n17447_ | ~new_n17431_;
  assign new_n18749_ = ~new_n17445_ | ~new_n17675_;
  assign new_n18750_ = ~new_n16939_ | ~new_n15700_;
  assign new_n18751_ = ~new_n32790_ | ~new_n15561_;
  assign new_n18752_ = ~new_n30952_ | ~new_n15559_;
  assign new_n18753_ = ~new_n31582_ | ~new_n15558_;
  assign new_n18754_ = ~new_n33660_ | ~new_n15556_;
  assign new_n18755_ = ~pi1215 | ~new_n15555_;
  assign new_n18756_ = ~pi1406 | ~new_n15551_;
  assign new_n18757_ = ~new_n18745_ | ~pi1215;
  assign new_n18758_ = ~new_n32791_ | ~new_n15561_;
  assign new_n18759_ = ~new_n31018_ | ~new_n15559_;
  assign new_n18760_ = ~new_n31502_ | ~new_n15558_;
  assign new_n18761_ = ~new_n33741_ | ~new_n15556_;
  assign new_n18762_ = ~new_n9376_ | ~new_n15555_;
  assign new_n18763_ = ~new_n15551_ | ~pi1407;
  assign new_n18764_ = ~new_n18745_ | ~pi1216;
  assign new_n18765_ = ~new_n32842_ | ~new_n15561_;
  assign new_n18766_ = ~new_n31007_ | ~new_n15559_;
  assign new_n18767_ = ~new_n31590_ | ~new_n15558_;
  assign new_n18768_ = ~new_n33661_ | ~new_n15556_;
  assign new_n18769_ = ~new_n9313_ | ~new_n15555_;
  assign new_n18770_ = ~new_n15551_ | ~pi1408;
  assign new_n18771_ = ~pi1217 | ~new_n18745_;
  assign new_n18772_ = ~new_n32746_ | ~new_n15561_;
  assign new_n18773_ = ~new_n31004_ | ~new_n15559_;
  assign new_n18774_ = ~new_n31588_ | ~new_n15558_;
  assign new_n18775_ = ~new_n20994_ | ~new_n15556_;
  assign new_n18776_ = ~new_n9295_ | ~new_n15555_;
  assign new_n18777_ = ~new_n15551_ | ~pi1409;
  assign new_n18778_ = ~pi1218 | ~new_n18745_;
  assign new_n18779_ = ~new_n32745_ | ~new_n15561_;
  assign new_n18780_ = ~new_n31003_ | ~new_n15559_;
  assign new_n18781_ = ~new_n31587_ | ~new_n15558_;
  assign new_n18782_ = ~new_n33732_ | ~new_n15556_;
  assign new_n18783_ = ~new_n9304_ | ~new_n15555_;
  assign new_n18784_ = ~new_n15551_ | ~pi1410;
  assign new_n18785_ = ~pi1219 | ~new_n18745_;
  assign new_n18786_ = ~new_n32744_ | ~new_n15561_;
  assign new_n18787_ = ~new_n31002_ | ~new_n15559_;
  assign new_n18788_ = ~new_n31500_ | ~new_n15558_;
  assign new_n18789_ = ~new_n33735_ | ~new_n15556_;
  assign new_n18790_ = ~new_n9301_ | ~new_n15555_;
  assign new_n18791_ = ~new_n15551_ | ~pi1411;
  assign new_n18792_ = ~pi1220 | ~new_n18745_;
  assign new_n18793_ = ~new_n32743_ | ~new_n15561_;
  assign new_n18794_ = ~new_n31001_ | ~new_n15559_;
  assign new_n18795_ = ~new_n31586_ | ~new_n15558_;
  assign new_n18796_ = ~new_n33719_ | ~new_n15556_;
  assign new_n18797_ = ~new_n9318_ | ~new_n15555_;
  assign new_n18798_ = ~new_n15551_ | ~pi1412;
  assign new_n18799_ = ~pi1221 | ~new_n18745_;
  assign new_n18800_ = ~new_n32742_ | ~new_n15561_;
  assign new_n18801_ = ~new_n31000_ | ~new_n15559_;
  assign new_n18802_ = ~new_n31501_ | ~new_n15558_;
  assign new_n18803_ = ~new_n21000_ | ~new_n15556_;
  assign new_n18804_ = ~new_n9291_ | ~new_n15555_;
  assign new_n18805_ = ~new_n15551_ | ~pi1413;
  assign new_n18806_ = ~pi1222 | ~new_n18745_;
  assign new_n18807_ = ~new_n32741_ | ~new_n15561_;
  assign new_n18808_ = ~new_n30999_ | ~new_n15559_;
  assign new_n18809_ = ~new_n31585_ | ~new_n15558_;
  assign new_n18810_ = ~new_n33736_ | ~new_n15556_;
  assign new_n18811_ = ~new_n9300_ | ~new_n15555_;
  assign new_n18812_ = ~new_n15551_ | ~pi1414;
  assign new_n18813_ = ~pi1223 | ~new_n18745_;
  assign new_n18814_ = ~new_n32740_ | ~new_n15561_;
  assign new_n18815_ = ~new_n30998_ | ~new_n15559_;
  assign new_n18816_ = ~new_n31584_ | ~new_n15558_;
  assign new_n18817_ = ~new_n33726_ | ~new_n15556_;
  assign new_n18818_ = ~new_n9310_ | ~new_n15555_;
  assign new_n18819_ = ~new_n15551_ | ~pi1415;
  assign new_n18820_ = ~pi1224 | ~new_n18745_;
  assign new_n18821_ = ~new_n32789_ | ~new_n15561_;
  assign new_n18822_ = ~new_n31028_ | ~new_n15559_;
  assign new_n18823_ = ~new_n31609_ | ~new_n15558_;
  assign new_n18824_ = ~new_n33739_ | ~new_n15556_;
  assign new_n18825_ = ~new_n9297_ | ~new_n15555_;
  assign new_n18826_ = ~new_n15551_ | ~pi1416;
  assign new_n18827_ = ~pi1225 | ~new_n18745_;
  assign new_n18828_ = ~new_n32788_ | ~new_n15561_;
  assign new_n18829_ = ~new_n31027_ | ~new_n15559_;
  assign new_n18830_ = ~new_n31498_ | ~new_n15558_;
  assign new_n18831_ = ~new_n33729_ | ~new_n15556_;
  assign new_n18832_ = ~new_n9307_ | ~new_n15555_;
  assign new_n18833_ = ~new_n15551_ | ~pi1417;
  assign new_n18834_ = ~pi1226 | ~new_n18745_;
  assign new_n18835_ = ~new_n32787_ | ~new_n15561_;
  assign new_n18836_ = ~new_n31026_ | ~new_n15559_;
  assign new_n18837_ = ~new_n31608_ | ~new_n15558_;
  assign new_n18838_ = ~new_n21001_ | ~new_n15556_;
  assign new_n18839_ = ~new_n9292_ | ~new_n15555_;
  assign new_n18840_ = ~new_n15551_ | ~pi1418;
  assign new_n18841_ = ~pi1227 | ~new_n18745_;
  assign new_n18842_ = ~new_n32786_ | ~new_n15561_;
  assign new_n18843_ = ~new_n31025_ | ~new_n15559_;
  assign new_n18844_ = ~new_n31606_ | ~new_n15558_;
  assign new_n18845_ = ~new_n33725_ | ~new_n15556_;
  assign new_n18846_ = ~new_n9311_ | ~new_n15555_;
  assign new_n18847_ = ~new_n15551_ | ~pi1419;
  assign new_n18848_ = ~pi1228 | ~new_n18745_;
  assign new_n18849_ = ~new_n32785_ | ~new_n15561_;
  assign new_n18850_ = ~new_n31024_ | ~new_n15559_;
  assign new_n18851_ = ~new_n31605_ | ~new_n15558_;
  assign new_n18852_ = ~new_n33734_ | ~new_n15556_;
  assign new_n18853_ = ~new_n9302_ | ~new_n15555_;
  assign new_n18854_ = ~new_n15551_ | ~pi1420;
  assign new_n18855_ = ~pi1229 | ~new_n18745_;
  assign new_n18856_ = ~new_n32784_ | ~new_n15561_;
  assign new_n18857_ = ~new_n31023_ | ~new_n15559_;
  assign new_n18858_ = ~new_n31503_ | ~new_n15558_;
  assign new_n18859_ = ~new_n33731_ | ~new_n15556_;
  assign new_n18860_ = ~new_n9305_ | ~new_n15555_;
  assign new_n18861_ = ~new_n15551_ | ~pi1421;
  assign new_n18862_ = ~pi1230 | ~new_n18745_;
  assign new_n18863_ = ~new_n32783_ | ~new_n15561_;
  assign new_n18864_ = ~new_n31022_ | ~new_n15559_;
  assign new_n18865_ = ~new_n31604_ | ~new_n15558_;
  assign new_n18866_ = ~new_n20998_ | ~new_n15556_;
  assign new_n18867_ = ~new_n9289_ | ~new_n15555_;
  assign new_n18868_ = ~new_n15551_ | ~pi1422;
  assign new_n18869_ = ~pi1231 | ~new_n18745_;
  assign new_n18870_ = ~new_n32782_ | ~new_n15561_;
  assign new_n18871_ = ~new_n31021_ | ~new_n15559_;
  assign new_n18872_ = ~new_n31603_ | ~new_n15558_;
  assign new_n18873_ = ~new_n33723_ | ~new_n15556_;
  assign new_n18874_ = ~new_n9314_ | ~new_n15555_;
  assign new_n18875_ = ~new_n15551_ | ~pi1423;
  assign new_n18876_ = ~pi1232 | ~new_n18745_;
  assign new_n18877_ = ~new_n32781_ | ~new_n15561_;
  assign new_n18878_ = ~new_n31020_ | ~new_n15559_;
  assign new_n18879_ = ~new_n31602_ | ~new_n15558_;
  assign new_n18880_ = ~new_n33728_ | ~new_n15556_;
  assign new_n18881_ = ~new_n9308_ | ~new_n15555_;
  assign new_n18882_ = ~new_n15551_ | ~pi1424;
  assign new_n18883_ = ~pi1233 | ~new_n18745_;
  assign new_n18884_ = ~new_n32780_ | ~new_n15561_;
  assign new_n18885_ = ~new_n31019_ | ~new_n15559_;
  assign new_n18886_ = ~new_n31601_ | ~new_n15558_;
  assign new_n18887_ = ~new_n33738_ | ~new_n15556_;
  assign new_n18888_ = ~new_n9298_ | ~new_n15555_;
  assign new_n18889_ = ~new_n15551_ | ~pi1425;
  assign new_n18890_ = ~pi1234 | ~new_n18745_;
  assign new_n18891_ = ~new_n32779_ | ~new_n15561_;
  assign new_n18892_ = ~new_n31017_ | ~new_n15559_;
  assign new_n18893_ = ~new_n31600_ | ~new_n15558_;
  assign new_n18894_ = ~new_n33724_ | ~new_n15556_;
  assign new_n18895_ = ~new_n9312_ | ~new_n15555_;
  assign new_n18896_ = ~new_n15551_ | ~pi1426;
  assign new_n18897_ = ~pi1235 | ~new_n18745_;
  assign new_n18898_ = ~new_n32778_ | ~new_n15561_;
  assign new_n18899_ = ~new_n31016_ | ~new_n15559_;
  assign new_n18900_ = ~new_n31599_ | ~new_n15558_;
  assign new_n18901_ = ~new_n21002_ | ~new_n15556_;
  assign new_n18902_ = ~new_n9293_ | ~new_n15555_;
  assign new_n18903_ = ~new_n15551_ | ~pi1427;
  assign new_n18904_ = ~pi1236 | ~new_n18745_;
  assign new_n18905_ = ~new_n32777_ | ~new_n15561_;
  assign new_n18906_ = ~new_n31015_ | ~new_n15559_;
  assign new_n18907_ = ~new_n31598_ | ~new_n15558_;
  assign new_n18908_ = ~new_n33727_ | ~new_n15556_;
  assign new_n18909_ = ~new_n9309_ | ~new_n15555_;
  assign new_n18910_ = ~new_n15551_ | ~pi1428;
  assign new_n18911_ = ~pi1237 | ~new_n18745_;
  assign new_n18912_ = ~new_n32776_ | ~new_n15561_;
  assign new_n18913_ = ~new_n31014_ | ~new_n15559_;
  assign new_n18914_ = ~new_n31597_ | ~new_n15558_;
  assign new_n18915_ = ~new_n33737_ | ~new_n15556_;
  assign new_n18916_ = ~new_n9299_ | ~new_n15555_;
  assign new_n18917_ = ~new_n15551_ | ~pi1429;
  assign new_n18918_ = ~pi1238 | ~new_n18745_;
  assign new_n18919_ = ~new_n32775_ | ~new_n15561_;
  assign new_n18920_ = ~new_n31013_ | ~new_n15559_;
  assign new_n18921_ = ~new_n31596_ | ~new_n15558_;
  assign new_n18922_ = ~new_n33722_ | ~new_n15556_;
  assign new_n18923_ = ~new_n9315_ | ~new_n15555_;
  assign new_n18924_ = ~new_n15551_ | ~pi1430;
  assign new_n18925_ = ~pi1239 | ~new_n18745_;
  assign new_n18926_ = ~new_n32774_ | ~new_n15561_;
  assign new_n18927_ = ~new_n31012_ | ~new_n15559_;
  assign new_n18928_ = ~new_n31595_ | ~new_n15558_;
  assign new_n18929_ = ~new_n20999_ | ~new_n15556_;
  assign new_n18930_ = ~new_n9290_ | ~new_n15555_;
  assign new_n18931_ = ~new_n15551_ | ~pi1431;
  assign new_n18932_ = ~pi1240 | ~new_n18745_;
  assign new_n18933_ = ~new_n32773_ | ~new_n15561_;
  assign new_n18934_ = ~new_n31011_ | ~new_n15559_;
  assign new_n18935_ = ~new_n31594_ | ~new_n15558_;
  assign new_n18936_ = ~new_n33730_ | ~new_n15556_;
  assign new_n18937_ = ~new_n9306_ | ~new_n15555_;
  assign new_n18938_ = ~new_n15551_ | ~pi1432;
  assign new_n18939_ = ~pi1241 | ~new_n18745_;
  assign new_n18940_ = ~new_n32772_ | ~new_n15561_;
  assign new_n18941_ = ~new_n31010_ | ~new_n15559_;
  assign new_n18942_ = ~new_n31593_ | ~new_n15558_;
  assign new_n18943_ = ~new_n33733_ | ~new_n15556_;
  assign new_n18944_ = ~new_n9303_ | ~new_n15555_;
  assign new_n18945_ = ~new_n15551_ | ~pi1433;
  assign new_n18946_ = ~pi1242 | ~new_n18745_;
  assign new_n18947_ = ~new_n32771_ | ~new_n15561_;
  assign new_n18948_ = ~new_n31009_ | ~new_n15559_;
  assign new_n18949_ = ~new_n31592_ | ~new_n15558_;
  assign new_n18950_ = ~new_n33742_ | ~new_n15556_;
  assign new_n18951_ = ~new_n9294_ | ~new_n15555_;
  assign new_n18952_ = ~new_n15551_ | ~pi1434;
  assign new_n18953_ = ~pi1243 | ~new_n18745_;
  assign new_n18954_ = ~new_n32770_ | ~new_n15561_;
  assign new_n18955_ = ~new_n31008_ | ~new_n15559_;
  assign new_n18956_ = ~new_n31591_ | ~new_n15558_;
  assign new_n18957_ = ~new_n33721_ | ~new_n15556_;
  assign new_n18958_ = ~new_n9316_ | ~new_n15555_;
  assign new_n18959_ = ~new_n15551_ | ~pi1435;
  assign new_n18960_ = ~pi1244 | ~new_n18745_;
  assign new_n18961_ = ~new_n32769_ | ~new_n15561_;
  assign new_n18962_ = ~new_n31006_ | ~new_n15559_;
  assign new_n18963_ = ~new_n31589_ | ~new_n15558_;
  assign new_n18964_ = ~new_n33720_ | ~new_n15556_;
  assign new_n18965_ = ~new_n9317_ | ~new_n15555_;
  assign new_n18966_ = ~new_n15551_ | ~pi1436;
  assign new_n18967_ = ~pi1245 | ~new_n18745_;
  assign new_n18968_ = ~new_n32768_ | ~new_n15561_;
  assign new_n18969_ = ~new_n31005_ | ~new_n15559_;
  assign new_n18970_ = ~new_n31499_ | ~new_n15558_;
  assign new_n18971_ = ~new_n33740_ | ~new_n15556_;
  assign new_n18972_ = ~new_n9296_ | ~new_n15555_;
  assign new_n18973_ = ~new_n15551_ | ~pi1437;
  assign new_n18974_ = ~pi1246 | ~new_n18745_;
  assign new_n18975_ = ~new_n17390_ | ~new_n16475_;
  assign new_n18976_ = ~new_n16597_;
  assign new_n18977_ = ~pi1074 | ~new_n16475_;
  assign new_n18978_ = ~pi1075 | ~new_n16489_;
  assign new_n18979_ = ~new_n18978_ | ~new_n18977_;
  assign new_n18980_ = ~pi1247 | ~new_n15557_;
  assign new_n18981_ = ~new_n15553_ | ~new_n31582_;
  assign new_n18982_ = ~new_n15546_ | ~pi1406;
  assign new_n18983_ = ~new_n32165_ | ~new_n15545_;
  assign new_n18984_ = ~pi1247 | ~new_n18976_;
  assign new_n18985_ = ~new_n33099_ | ~new_n15557_;
  assign new_n18986_ = ~new_n15553_ | ~new_n31502_;
  assign new_n18987_ = ~new_n15546_ | ~pi1407;
  assign new_n18988_ = ~new_n32196_ | ~new_n15545_;
  assign new_n18989_ = ~pi1248 | ~new_n18976_;
  assign new_n18990_ = ~new_n33166_ | ~new_n15557_;
  assign new_n18991_ = ~new_n15553_ | ~new_n31590_;
  assign new_n18992_ = ~new_n15546_ | ~pi1408;
  assign new_n18993_ = ~new_n32107_ | ~new_n15545_;
  assign new_n18994_ = ~pi1249 | ~new_n18976_;
  assign new_n18995_ = ~new_n33163_ | ~new_n15557_;
  assign new_n18996_ = ~new_n15553_ | ~new_n31588_;
  assign new_n18997_ = ~new_n15546_ | ~pi1409;
  assign new_n18998_ = ~new_n32108_ | ~new_n15545_;
  assign new_n18999_ = ~pi1250 | ~new_n18976_;
  assign new_n19000_ = ~new_n33162_ | ~new_n15557_;
  assign new_n19001_ = ~new_n15553_ | ~new_n31587_;
  assign new_n19002_ = ~new_n15546_ | ~pi1410;
  assign new_n19003_ = ~new_n32173_ | ~new_n15545_;
  assign new_n19004_ = ~pi1251 | ~new_n18976_;
  assign new_n19005_ = ~new_n33161_ | ~new_n15557_;
  assign new_n19006_ = ~new_n15553_ | ~new_n31500_;
  assign new_n19007_ = ~new_n15546_ | ~pi1411;
  assign new_n19008_ = ~new_n32171_ | ~new_n15545_;
  assign new_n19009_ = ~pi1252 | ~new_n18976_;
  assign new_n19010_ = ~new_n33160_ | ~new_n15557_;
  assign new_n19011_ = ~new_n15553_ | ~new_n31586_;
  assign new_n19012_ = ~new_n15546_ | ~pi1412;
  assign new_n19013_ = ~new_n32109_ | ~new_n15545_;
  assign new_n19014_ = ~pi1253 | ~new_n18976_;
  assign new_n19015_ = ~new_n33159_ | ~new_n15557_;
  assign new_n19016_ = ~new_n15553_ | ~new_n31501_;
  assign new_n19017_ = ~new_n15546_ | ~pi1413;
  assign new_n19018_ = ~new_n32110_ | ~new_n15545_;
  assign new_n19019_ = ~pi1254 | ~new_n18976_;
  assign new_n19020_ = ~new_n33158_ | ~new_n15557_;
  assign new_n19021_ = ~new_n15553_ | ~new_n31585_;
  assign new_n19022_ = ~new_n15546_ | ~pi1414;
  assign new_n19023_ = ~new_n32169_ | ~new_n15545_;
  assign new_n19024_ = ~pi1255 | ~new_n18976_;
  assign new_n19025_ = ~new_n33157_ | ~new_n15557_;
  assign new_n19026_ = ~new_n15553_ | ~new_n31584_;
  assign new_n19027_ = ~new_n15546_ | ~pi1415;
  assign new_n19028_ = ~new_n32167_ | ~new_n15545_;
  assign new_n19029_ = ~pi1256 | ~new_n18976_;
  assign new_n19030_ = ~new_n33186_ | ~new_n15557_;
  assign new_n19031_ = ~new_n15553_ | ~new_n31609_;
  assign new_n19032_ = ~new_n15546_ | ~pi1416;
  assign new_n19033_ = ~new_n32103_ | ~new_n15545_;
  assign new_n19034_ = ~pi1257 | ~new_n18976_;
  assign new_n19035_ = ~new_n33185_ | ~new_n15557_;
  assign new_n19036_ = ~new_n15553_ | ~new_n31498_;
  assign new_n19037_ = ~new_n15546_ | ~pi1417;
  assign new_n19038_ = ~new_n32104_ | ~new_n15545_;
  assign new_n19039_ = ~pi1258 | ~new_n18976_;
  assign new_n19040_ = ~new_n33184_ | ~new_n15557_;
  assign new_n19041_ = ~new_n15553_ | ~new_n31608_;
  assign new_n19042_ = ~new_n15546_ | ~pi1418;
  assign new_n19043_ = ~new_n32208_ | ~new_n15545_;
  assign new_n19044_ = ~pi1259 | ~new_n18976_;
  assign new_n19045_ = ~new_n33183_ | ~new_n15557_;
  assign new_n19046_ = ~new_n15553_ | ~new_n31606_;
  assign new_n19047_ = ~new_n15546_ | ~pi1419;
  assign new_n19048_ = ~new_n32206_ | ~new_n15545_;
  assign new_n19049_ = ~pi1260 | ~new_n18976_;
  assign new_n19050_ = ~new_n33182_ | ~new_n15557_;
  assign new_n19051_ = ~new_n15553_ | ~new_n31605_;
  assign new_n19052_ = ~new_n15546_ | ~pi1420;
  assign new_n19053_ = ~new_n32105_ | ~new_n15545_;
  assign new_n19054_ = ~pi1261 | ~new_n18976_;
  assign new_n19055_ = ~new_n33181_ | ~new_n15557_;
  assign new_n19056_ = ~new_n15553_ | ~new_n31503_;
  assign new_n19057_ = ~new_n15546_ | ~pi1421;
  assign new_n19058_ = ~new_n32106_ | ~new_n15545_;
  assign new_n19059_ = ~pi1262 | ~new_n18976_;
  assign new_n19060_ = ~new_n33180_ | ~new_n15557_;
  assign new_n19061_ = ~new_n15553_ | ~new_n31604_;
  assign new_n19062_ = ~new_n15546_ | ~pi1422;
  assign new_n19063_ = ~new_n32204_ | ~new_n15545_;
  assign new_n19064_ = ~pi1263 | ~new_n18976_;
  assign new_n19065_ = ~new_n33179_ | ~new_n15557_;
  assign new_n19066_ = ~new_n15553_ | ~new_n31603_;
  assign new_n19067_ = ~new_n15546_ | ~pi1423;
  assign new_n19068_ = ~new_n32202_ | ~new_n15545_;
  assign new_n19069_ = ~pi1264 | ~new_n18976_;
  assign new_n19070_ = ~new_n33178_ | ~new_n15557_;
  assign new_n19071_ = ~new_n15553_ | ~new_n31602_;
  assign new_n19072_ = ~new_n15546_ | ~pi1424;
  assign new_n19073_ = ~new_n32200_ | ~new_n15545_;
  assign new_n19074_ = ~pi1265 | ~new_n18976_;
  assign new_n19075_ = ~new_n33177_ | ~new_n15557_;
  assign new_n19076_ = ~new_n15553_ | ~new_n31601_;
  assign new_n19077_ = ~new_n15546_ | ~pi1425;
  assign new_n19078_ = ~new_n32198_ | ~new_n15545_;
  assign new_n19079_ = ~pi1266 | ~new_n18976_;
  assign new_n19080_ = ~new_n33176_ | ~new_n15557_;
  assign new_n19081_ = ~new_n15553_ | ~new_n31600_;
  assign new_n19082_ = ~new_n15546_ | ~pi1426;
  assign new_n19083_ = ~new_n32194_ | ~new_n15545_;
  assign new_n19084_ = ~pi1267 | ~new_n18976_;
  assign new_n19085_ = ~new_n33175_ | ~new_n15557_;
  assign new_n19086_ = ~new_n15553_ | ~new_n31599_;
  assign new_n19087_ = ~new_n15546_ | ~pi1427;
  assign new_n19088_ = ~new_n32192_ | ~new_n15545_;
  assign new_n19089_ = ~pi1268 | ~new_n18976_;
  assign new_n19090_ = ~new_n33174_ | ~new_n15557_;
  assign new_n19091_ = ~new_n15553_ | ~new_n31598_;
  assign new_n19092_ = ~new_n15546_ | ~pi1428;
  assign new_n19093_ = ~new_n32190_ | ~new_n15545_;
  assign new_n19094_ = ~pi1269 | ~new_n18976_;
  assign new_n19095_ = ~new_n33173_ | ~new_n15557_;
  assign new_n19096_ = ~new_n15553_ | ~new_n31597_;
  assign new_n19097_ = ~new_n15546_ | ~pi1429;
  assign new_n19098_ = ~new_n32188_ | ~new_n15545_;
  assign new_n19099_ = ~pi1270 | ~new_n18976_;
  assign new_n19100_ = ~new_n33172_ | ~new_n15557_;
  assign new_n19101_ = ~new_n15553_ | ~new_n31596_;
  assign new_n19102_ = ~new_n15546_ | ~pi1430;
  assign new_n19103_ = ~new_n32186_ | ~new_n15545_;
  assign new_n19104_ = ~pi1271 | ~new_n18976_;
  assign new_n19105_ = ~new_n33171_ | ~new_n15557_;
  assign new_n19106_ = ~new_n15553_ | ~new_n31595_;
  assign new_n19107_ = ~new_n15546_ | ~pi1431;
  assign new_n19108_ = ~new_n32184_ | ~new_n15545_;
  assign new_n19109_ = ~pi1272 | ~new_n18976_;
  assign new_n19110_ = ~new_n33170_ | ~new_n15557_;
  assign new_n19111_ = ~new_n15553_ | ~new_n31594_;
  assign new_n19112_ = ~new_n15546_ | ~pi1432;
  assign new_n19113_ = ~new_n32182_ | ~new_n15545_;
  assign new_n19114_ = ~pi1273 | ~new_n18976_;
  assign new_n19115_ = ~new_n33169_ | ~new_n15557_;
  assign new_n19116_ = ~new_n15553_ | ~new_n31593_;
  assign new_n19117_ = ~new_n15546_ | ~pi1433;
  assign new_n19118_ = ~new_n32180_ | ~new_n15545_;
  assign new_n19119_ = ~pi1274 | ~new_n18976_;
  assign new_n19120_ = ~new_n33168_ | ~new_n15557_;
  assign new_n19121_ = ~new_n15553_ | ~new_n31592_;
  assign new_n19122_ = ~new_n15546_ | ~pi1434;
  assign new_n19123_ = ~new_n32178_ | ~new_n15545_;
  assign new_n19124_ = ~pi1275 | ~new_n18976_;
  assign new_n19125_ = ~new_n33167_ | ~new_n15557_;
  assign new_n19126_ = ~new_n15553_ | ~new_n31591_;
  assign new_n19127_ = ~new_n15546_ | ~pi1435;
  assign new_n19128_ = ~new_n32176_ | ~new_n15545_;
  assign new_n19129_ = ~pi1276 | ~new_n18976_;
  assign new_n19130_ = ~new_n33165_ | ~new_n15557_;
  assign new_n19131_ = ~new_n15553_ | ~new_n31589_;
  assign new_n19132_ = ~new_n15546_ | ~pi1436;
  assign new_n19133_ = ~new_n32174_ | ~new_n15545_;
  assign new_n19134_ = ~pi1277 | ~new_n18976_;
  assign new_n19135_ = ~new_n33164_ | ~new_n15557_;
  assign new_n19136_ = ~new_n15553_ | ~new_n31499_;
  assign new_n19137_ = ~new_n15546_ | ~pi1437;
  assign new_n19138_ = ~new_n32111_ | ~new_n15545_;
  assign new_n19139_ = ~pi1278 | ~new_n18976_;
  assign new_n19140_ = ~new_n2972_ | ~new_n16463_;
  assign new_n19141_ = ~pi1357 | ~new_n15563_;
  assign new_n19142_ = ~new_n3102_ | ~new_n15562_;
  assign new_n19143_ = ~new_n19142_ | ~new_n19141_;
  assign new_n19144_ = ~pi1356 | ~new_n15563_;
  assign new_n19145_ = ~new_n3103_ | ~new_n15562_;
  assign new_n19146_ = ~new_n19145_ | ~new_n19144_;
  assign new_n19147_ = ~pi1355 | ~new_n15563_;
  assign new_n19148_ = ~new_n3104_ | ~new_n15562_;
  assign new_n19149_ = ~new_n19148_ | ~new_n19147_;
  assign new_n19150_ = ~pi1354 | ~new_n15563_;
  assign new_n19151_ = ~new_n3105_ | ~new_n15562_;
  assign new_n19152_ = ~new_n19151_ | ~new_n19150_;
  assign new_n19153_ = ~pi1353 | ~new_n15563_;
  assign new_n19154_ = ~new_n3106_ | ~new_n15562_;
  assign new_n19155_ = ~new_n19154_ | ~new_n19153_;
  assign new_n19156_ = ~pi1352 | ~new_n15563_;
  assign new_n19157_ = ~new_n3107_ | ~new_n15562_;
  assign new_n19158_ = ~new_n19157_ | ~new_n19156_;
  assign new_n19159_ = ~pi1351 | ~new_n15563_;
  assign new_n19160_ = ~new_n3077_ | ~new_n15562_;
  assign new_n19161_ = ~new_n19160_ | ~new_n19159_;
  assign new_n19162_ = ~pi1350 | ~new_n15563_;
  assign new_n19163_ = ~new_n3078_ | ~new_n15562_;
  assign new_n19164_ = ~new_n19163_ | ~new_n19162_;
  assign new_n19165_ = ~pi1349 | ~new_n15563_;
  assign new_n19166_ = ~new_n15562_ | ~new_n3079_;
  assign new_n19167_ = ~new_n19166_ | ~new_n19165_;
  assign new_n19168_ = ~pi1348 | ~new_n15563_;
  assign new_n19169_ = ~new_n15562_ | ~new_n3080_;
  assign new_n19170_ = ~new_n19169_ | ~new_n19168_;
  assign new_n19171_ = ~pi1347 | ~new_n15563_;
  assign new_n19172_ = ~new_n15562_ | ~new_n3081_;
  assign new_n19173_ = ~new_n19172_ | ~new_n19171_;
  assign new_n19174_ = ~pi1346 | ~new_n15563_;
  assign new_n19175_ = ~new_n15562_ | ~new_n3082_;
  assign new_n19176_ = ~new_n19175_ | ~new_n19174_;
  assign new_n19177_ = ~pi1345 | ~new_n15563_;
  assign new_n19178_ = ~new_n15562_ | ~new_n3083_;
  assign new_n19179_ = ~new_n19178_ | ~new_n19177_;
  assign new_n19180_ = ~pi1344 | ~new_n15563_;
  assign new_n19181_ = ~new_n15562_ | ~new_n3086_;
  assign new_n19182_ = ~new_n19181_ | ~new_n19180_;
  assign new_n19183_ = ~pi1343 | ~new_n15563_;
  assign new_n19184_ = ~new_n15562_ | ~new_n3097_;
  assign new_n19185_ = ~new_n19184_ | ~new_n19183_;
  assign new_n19186_ = ~pi1342 | ~new_n15563_;
  assign new_n19187_ = ~new_n15562_ | ~new_n3108_;
  assign new_n19188_ = ~new_n19187_ | ~new_n19186_;
  assign new_n19189_ = ~pi1372 | ~new_n15563_;
  assign new_n19190_ = ~new_n3103_ | ~new_n15562_;
  assign new_n19191_ = ~new_n19190_ | ~new_n19189_;
  assign new_n19192_ = ~pi1371 | ~new_n15563_;
  assign new_n19193_ = ~new_n3104_ | ~new_n15562_;
  assign new_n19194_ = ~new_n19193_ | ~new_n19192_;
  assign new_n19195_ = ~pi1370 | ~new_n15563_;
  assign new_n19196_ = ~new_n3105_ | ~new_n15562_;
  assign new_n19197_ = ~new_n19196_ | ~new_n19195_;
  assign new_n19198_ = ~pi1369 | ~new_n15563_;
  assign new_n19199_ = ~new_n3106_ | ~new_n15562_;
  assign new_n19200_ = ~new_n19199_ | ~new_n19198_;
  assign new_n19201_ = ~pi1368 | ~new_n15563_;
  assign new_n19202_ = ~new_n3107_ | ~new_n15562_;
  assign new_n19203_ = ~new_n19202_ | ~new_n19201_;
  assign new_n19204_ = ~pi1367 | ~new_n15563_;
  assign new_n19205_ = ~new_n3077_ | ~new_n15562_;
  assign new_n19206_ = ~new_n19205_ | ~new_n19204_;
  assign new_n19207_ = ~pi1366 | ~new_n15563_;
  assign new_n19208_ = ~new_n3078_ | ~new_n15562_;
  assign new_n19209_ = ~new_n19208_ | ~new_n19207_;
  assign new_n19210_ = ~pi1365 | ~new_n15563_;
  assign new_n19211_ = ~new_n15562_ | ~new_n3079_;
  assign new_n19212_ = ~new_n19211_ | ~new_n19210_;
  assign new_n19213_ = ~pi1364 | ~new_n15563_;
  assign new_n19214_ = ~new_n15562_ | ~new_n3080_;
  assign new_n19215_ = ~new_n19214_ | ~new_n19213_;
  assign new_n19216_ = ~pi1363 | ~new_n15563_;
  assign new_n19217_ = ~new_n15562_ | ~new_n3081_;
  assign new_n19218_ = ~new_n19217_ | ~new_n19216_;
  assign new_n19219_ = ~pi1362 | ~new_n15563_;
  assign new_n19220_ = ~new_n15562_ | ~new_n3082_;
  assign new_n19221_ = ~new_n19220_ | ~new_n19219_;
  assign new_n19222_ = ~pi1361 | ~new_n15563_;
  assign new_n19223_ = ~new_n15562_ | ~new_n3083_;
  assign new_n19224_ = ~new_n19223_ | ~new_n19222_;
  assign new_n19225_ = ~pi1360 | ~new_n15563_;
  assign new_n19226_ = ~new_n15562_ | ~new_n3086_;
  assign new_n19227_ = ~new_n19226_ | ~new_n19225_;
  assign new_n19228_ = ~pi1359 | ~new_n15563_;
  assign new_n19229_ = ~new_n15562_ | ~new_n3097_;
  assign new_n19230_ = ~new_n19229_ | ~new_n19228_;
  assign new_n19231_ = ~pi1358 | ~new_n15563_;
  assign new_n19232_ = ~new_n15562_ | ~new_n3108_;
  assign new_n19233_ = ~new_n19232_ | ~new_n19231_;
  assign new_n19234_ = ~new_n17440_ | ~new_n17416_ | ~new_n20787_;
  assign new_n19235_ = ~new_n15609_ | ~new_n16475_;
  assign new_n19236_ = ~new_n16598_;
  assign new_n19237_ = ~new_n15566_ | ~pi1294;
  assign new_n19238_ = ~new_n15565_ | ~pi1342;
  assign new_n19239_ = ~pi1310 | ~new_n19236_;
  assign new_n19240_ = ~new_n15566_ | ~pi1293;
  assign new_n19241_ = ~new_n15565_ | ~pi1343;
  assign new_n19242_ = ~pi1311 | ~new_n19236_;
  assign new_n19243_ = ~new_n15566_ | ~pi1292;
  assign new_n19244_ = ~new_n15565_ | ~pi1344;
  assign new_n19245_ = ~pi1312 | ~new_n19236_;
  assign new_n19246_ = ~new_n15566_ | ~pi1291;
  assign new_n19247_ = ~new_n15565_ | ~pi1345;
  assign new_n19248_ = ~pi1313 | ~new_n19236_;
  assign new_n19249_ = ~new_n15566_ | ~pi1290;
  assign new_n19250_ = ~new_n15565_ | ~pi1346;
  assign new_n19251_ = ~pi1314 | ~new_n19236_;
  assign new_n19252_ = ~new_n15566_ | ~pi1289;
  assign new_n19253_ = ~new_n15565_ | ~pi1347;
  assign new_n19254_ = ~pi1315 | ~new_n19236_;
  assign new_n19255_ = ~new_n15566_ | ~pi1288;
  assign new_n19256_ = ~new_n15565_ | ~pi1348;
  assign new_n19257_ = ~pi1316 | ~new_n19236_;
  assign new_n19258_ = ~new_n15566_ | ~pi1287;
  assign new_n19259_ = ~new_n15565_ | ~pi1349;
  assign new_n19260_ = ~pi1317 | ~new_n19236_;
  assign new_n19261_ = ~new_n15566_ | ~pi1286;
  assign new_n19262_ = ~new_n15565_ | ~pi1350;
  assign new_n19263_ = ~pi1318 | ~new_n19236_;
  assign new_n19264_ = ~new_n15566_ | ~pi1285;
  assign new_n19265_ = ~new_n15565_ | ~pi1351;
  assign new_n19266_ = ~pi1319 | ~new_n19236_;
  assign new_n19267_ = ~new_n15566_ | ~pi1284;
  assign new_n19268_ = ~new_n15565_ | ~pi1352;
  assign new_n19269_ = ~pi1320 | ~new_n19236_;
  assign new_n19270_ = ~new_n15566_ | ~pi1283;
  assign new_n19271_ = ~new_n15565_ | ~pi1353;
  assign new_n19272_ = ~pi1321 | ~new_n19236_;
  assign new_n19273_ = ~new_n15566_ | ~pi1282;
  assign new_n19274_ = ~new_n15565_ | ~pi1354;
  assign new_n19275_ = ~pi1322 | ~new_n19236_;
  assign new_n19276_ = ~new_n15566_ | ~pi1281;
  assign new_n19277_ = ~new_n15565_ | ~pi1355;
  assign new_n19278_ = ~pi1323 | ~new_n19236_;
  assign new_n19279_ = ~new_n15566_ | ~pi1280;
  assign new_n19280_ = ~new_n15565_ | ~pi1356;
  assign new_n19281_ = ~pi1324 | ~new_n19236_;
  assign new_n19282_ = ~new_n15566_ | ~pi1279;
  assign new_n19283_ = ~new_n15565_ | ~pi1357;
  assign new_n19284_ = ~pi1325 | ~new_n19236_;
  assign new_n19285_ = ~new_n15605_ | ~pi1358;
  assign new_n19286_ = ~new_n15566_ | ~pi1309;
  assign new_n19287_ = ~pi1326 | ~new_n19236_;
  assign new_n19288_ = ~new_n15605_ | ~pi1359;
  assign new_n19289_ = ~new_n15566_ | ~pi1308;
  assign new_n19290_ = ~pi1327 | ~new_n19236_;
  assign new_n19291_ = ~new_n15605_ | ~pi1360;
  assign new_n19292_ = ~new_n15566_ | ~pi1307;
  assign new_n19293_ = ~pi1328 | ~new_n19236_;
  assign new_n19294_ = ~new_n15605_ | ~pi1361;
  assign new_n19295_ = ~new_n15566_ | ~pi1306;
  assign new_n19296_ = ~pi1329 | ~new_n19236_;
  assign new_n19297_ = ~new_n15605_ | ~pi1362;
  assign new_n19298_ = ~new_n15566_ | ~pi1305;
  assign new_n19299_ = ~pi1330 | ~new_n19236_;
  assign new_n19300_ = ~new_n15605_ | ~pi1363;
  assign new_n19301_ = ~new_n15566_ | ~pi1304;
  assign new_n19302_ = ~pi1331 | ~new_n19236_;
  assign new_n19303_ = ~new_n15605_ | ~pi1364;
  assign new_n19304_ = ~new_n15566_ | ~pi1303;
  assign new_n19305_ = ~pi1332 | ~new_n19236_;
  assign new_n19306_ = ~new_n15605_ | ~pi1365;
  assign new_n19307_ = ~new_n15566_ | ~pi1302;
  assign new_n19308_ = ~pi1333 | ~new_n19236_;
  assign new_n19309_ = ~new_n15605_ | ~pi1366;
  assign new_n19310_ = ~new_n15566_ | ~pi1301;
  assign new_n19311_ = ~pi1334 | ~new_n19236_;
  assign new_n19312_ = ~new_n15605_ | ~pi1367;
  assign new_n19313_ = ~new_n15566_ | ~pi1300;
  assign new_n19314_ = ~pi1335 | ~new_n19236_;
  assign new_n19315_ = ~new_n15605_ | ~pi1368;
  assign new_n19316_ = ~new_n15566_ | ~pi1299;
  assign new_n19317_ = ~pi1336 | ~new_n19236_;
  assign new_n19318_ = ~new_n15605_ | ~pi1369;
  assign new_n19319_ = ~new_n15566_ | ~pi1298;
  assign new_n19320_ = ~pi1337 | ~new_n19236_;
  assign new_n19321_ = ~new_n15605_ | ~pi1370;
  assign new_n19322_ = ~new_n15566_ | ~pi1297;
  assign new_n19323_ = ~pi1338 | ~new_n19236_;
  assign new_n19324_ = ~new_n15605_ | ~pi1371;
  assign new_n19325_ = ~new_n15566_ | ~pi1296;
  assign new_n19326_ = ~pi1339 | ~new_n19236_;
  assign new_n19327_ = ~new_n15605_ | ~pi1372;
  assign new_n19328_ = ~new_n15566_ | ~pi1295;
  assign new_n19329_ = ~pi1340 | ~new_n19236_;
  assign new_n19330_ = ~new_n9378_ | ~new_n17375_ | ~new_n15628_;
  assign new_n19331_ = ~new_n17375_ | ~new_n17435_ | ~new_n17378_;
  assign new_n19332_ = ~new_n33065_ | ~new_n17381_ | ~new_n16464_;
  assign new_n19333_ = ~new_n20684_ | ~new_n16438_;
  assign new_n19334_ = ~new_n17064_ | ~new_n19333_;
  assign new_n19335_ = ~new_n15603_ | ~new_n3108_;
  assign new_n19336_ = ~new_n15567_ | ~new_n32165_;
  assign new_n19337_ = ~pi1342 | ~new_n16605_;
  assign new_n19338_ = ~new_n15603_ | ~new_n3097_;
  assign new_n19339_ = ~new_n15567_ | ~new_n32196_;
  assign new_n19340_ = ~pi1343 | ~new_n16605_;
  assign new_n19341_ = ~new_n15603_ | ~new_n3086_;
  assign new_n19342_ = ~new_n15567_ | ~new_n32107_;
  assign new_n19343_ = ~pi1344 | ~new_n16605_;
  assign new_n19344_ = ~new_n15603_ | ~new_n3083_;
  assign new_n19345_ = ~new_n15567_ | ~new_n32108_;
  assign new_n19346_ = ~pi1345 | ~new_n16605_;
  assign new_n19347_ = ~new_n15603_ | ~new_n3082_;
  assign new_n19348_ = ~new_n15567_ | ~new_n32173_;
  assign new_n19349_ = ~pi1346 | ~new_n16605_;
  assign new_n19350_ = ~new_n15603_ | ~new_n3081_;
  assign new_n19351_ = ~new_n15567_ | ~new_n32171_;
  assign new_n19352_ = ~pi1347 | ~new_n16605_;
  assign new_n19353_ = ~new_n15603_ | ~new_n3080_;
  assign new_n19354_ = ~new_n15567_ | ~new_n32109_;
  assign new_n19355_ = ~pi1348 | ~new_n16605_;
  assign new_n19356_ = ~new_n15603_ | ~new_n3079_;
  assign new_n19357_ = ~new_n15567_ | ~new_n32110_;
  assign new_n19358_ = ~pi1349 | ~new_n16605_;
  assign new_n19359_ = ~new_n15603_ | ~new_n3078_;
  assign new_n19360_ = ~new_n15567_ | ~new_n32169_;
  assign new_n19361_ = ~pi1350 | ~new_n16605_;
  assign new_n19362_ = ~new_n15603_ | ~new_n3077_;
  assign new_n19363_ = ~new_n15567_ | ~new_n32167_;
  assign new_n19364_ = ~pi1351 | ~new_n16605_;
  assign new_n19365_ = ~new_n15603_ | ~new_n3107_;
  assign new_n19366_ = ~new_n15567_ | ~new_n32103_;
  assign new_n19367_ = ~pi1352 | ~new_n16605_;
  assign new_n19368_ = ~new_n15603_ | ~new_n3106_;
  assign new_n19369_ = ~new_n15567_ | ~new_n32104_;
  assign new_n19370_ = ~pi1353 | ~new_n16605_;
  assign new_n19371_ = ~new_n15603_ | ~new_n3105_;
  assign new_n19372_ = ~new_n15567_ | ~new_n32208_;
  assign new_n19373_ = ~pi1354 | ~new_n16605_;
  assign new_n19374_ = ~new_n15603_ | ~new_n3104_;
  assign new_n19375_ = ~new_n15567_ | ~new_n32206_;
  assign new_n19376_ = ~pi1355 | ~new_n16605_;
  assign new_n19377_ = ~new_n15603_ | ~new_n3103_;
  assign new_n19378_ = ~new_n15567_ | ~new_n32105_;
  assign new_n19379_ = ~pi1356 | ~new_n16605_;
  assign new_n19380_ = ~new_n15603_ | ~new_n3102_;
  assign new_n19381_ = ~new_n15567_ | ~new_n32106_;
  assign new_n19382_ = ~pi1357 | ~new_n16605_;
  assign new_n19383_ = ~new_n15604_ | ~new_n3101_;
  assign new_n19384_ = ~new_n15568_ | ~new_n3108_;
  assign new_n19385_ = ~new_n15567_ | ~new_n32204_;
  assign new_n19386_ = ~pi1358 | ~new_n16605_;
  assign new_n19387_ = ~new_n15604_ | ~new_n3100_;
  assign new_n19388_ = ~new_n15568_ | ~new_n3097_;
  assign new_n19389_ = ~new_n15567_ | ~new_n32202_;
  assign new_n19390_ = ~pi1359 | ~new_n16605_;
  assign new_n19391_ = ~new_n15604_ | ~new_n3099_;
  assign new_n19392_ = ~new_n15568_ | ~new_n3086_;
  assign new_n19393_ = ~new_n15567_ | ~new_n32200_;
  assign new_n19394_ = ~pi1360 | ~new_n16605_;
  assign new_n19395_ = ~new_n15604_ | ~new_n3098_;
  assign new_n19396_ = ~new_n15568_ | ~new_n3083_;
  assign new_n19397_ = ~new_n15567_ | ~new_n32198_;
  assign new_n19398_ = ~pi1361 | ~new_n16605_;
  assign new_n19399_ = ~new_n15604_ | ~new_n3096_;
  assign new_n19400_ = ~new_n15568_ | ~new_n3082_;
  assign new_n19401_ = ~new_n15567_ | ~new_n32194_;
  assign new_n19402_ = ~pi1362 | ~new_n16605_;
  assign new_n19403_ = ~new_n15604_ | ~new_n3095_;
  assign new_n19404_ = ~new_n15568_ | ~new_n3081_;
  assign new_n19405_ = ~new_n15567_ | ~new_n32192_;
  assign new_n19406_ = ~pi1363 | ~new_n16605_;
  assign new_n19407_ = ~new_n15604_ | ~new_n3094_;
  assign new_n19408_ = ~new_n15568_ | ~new_n3080_;
  assign new_n19409_ = ~new_n15567_ | ~new_n32190_;
  assign new_n19410_ = ~pi1364 | ~new_n16605_;
  assign new_n19411_ = ~new_n15604_ | ~new_n3093_;
  assign new_n19412_ = ~new_n15568_ | ~new_n3079_;
  assign new_n19413_ = ~new_n15567_ | ~new_n32188_;
  assign new_n19414_ = ~pi1365 | ~new_n16605_;
  assign new_n19415_ = ~new_n15604_ | ~new_n3092_;
  assign new_n19416_ = ~new_n15568_ | ~new_n3078_;
  assign new_n19417_ = ~new_n15567_ | ~new_n32186_;
  assign new_n19418_ = ~pi1366 | ~new_n16605_;
  assign new_n19419_ = ~new_n15604_ | ~new_n3091_;
  assign new_n19420_ = ~new_n15568_ | ~new_n3077_;
  assign new_n19421_ = ~new_n15567_ | ~new_n32184_;
  assign new_n19422_ = ~pi1367 | ~new_n16605_;
  assign new_n19423_ = ~new_n15604_ | ~new_n3090_;
  assign new_n19424_ = ~new_n15568_ | ~new_n3107_;
  assign new_n19425_ = ~new_n15567_ | ~new_n32182_;
  assign new_n19426_ = ~pi1368 | ~new_n16605_;
  assign new_n19427_ = ~new_n15604_ | ~new_n3089_;
  assign new_n19428_ = ~new_n15568_ | ~new_n3106_;
  assign new_n19429_ = ~new_n15567_ | ~new_n32180_;
  assign new_n19430_ = ~pi1369 | ~new_n16605_;
  assign new_n19431_ = ~new_n15604_ | ~new_n3088_;
  assign new_n19432_ = ~new_n15568_ | ~new_n3105_;
  assign new_n19433_ = ~new_n15567_ | ~new_n32178_;
  assign new_n19434_ = ~pi1370 | ~new_n16605_;
  assign new_n19435_ = ~new_n15604_ | ~new_n3087_;
  assign new_n19436_ = ~new_n15568_ | ~new_n3104_;
  assign new_n19437_ = ~new_n15567_ | ~new_n32176_;
  assign new_n19438_ = ~pi1371 | ~new_n16605_;
  assign new_n19439_ = ~new_n15604_ | ~new_n3085_;
  assign new_n19440_ = ~new_n15568_ | ~new_n3103_;
  assign new_n19441_ = ~new_n15567_ | ~new_n32174_;
  assign new_n19442_ = ~pi1372 | ~new_n16605_;
  assign new_n19443_ = ~new_n15604_ | ~new_n3084_;
  assign new_n19444_ = ~new_n17379_ | ~new_n16454_;
  assign new_n19445_ = ~new_n17386_ | ~new_n19444_;
  assign new_n19446_ = ~new_n15564_ | ~new_n32165_;
  assign new_n19447_ = ~new_n15552_ | ~new_n32790_;
  assign new_n19448_ = ~pi1374 | ~new_n16607_;
  assign new_n19449_ = ~new_n15564_ | ~new_n32196_;
  assign new_n19450_ = ~new_n15552_ | ~new_n32791_;
  assign new_n19451_ = ~pi1375 | ~new_n16607_;
  assign new_n19452_ = ~new_n15564_ | ~new_n32107_;
  assign new_n19453_ = ~new_n15552_ | ~new_n32842_;
  assign new_n19454_ = ~pi1376 | ~new_n16607_;
  assign new_n19455_ = ~new_n15564_ | ~new_n32108_;
  assign new_n19456_ = ~new_n15552_ | ~new_n32746_;
  assign new_n19457_ = ~pi1377 | ~new_n16607_;
  assign new_n19458_ = ~new_n15564_ | ~new_n32173_;
  assign new_n19459_ = ~new_n15552_ | ~new_n32745_;
  assign new_n19460_ = ~pi1378 | ~new_n16607_;
  assign new_n19461_ = ~new_n15564_ | ~new_n32171_;
  assign new_n19462_ = ~new_n15552_ | ~new_n32744_;
  assign new_n19463_ = ~pi1379 | ~new_n16607_;
  assign new_n19464_ = ~new_n15564_ | ~new_n32109_;
  assign new_n19465_ = ~new_n15552_ | ~new_n32743_;
  assign new_n19466_ = ~pi1380 | ~new_n16607_;
  assign new_n19467_ = ~new_n15564_ | ~new_n32110_;
  assign new_n19468_ = ~new_n15552_ | ~new_n32742_;
  assign new_n19469_ = ~pi1381 | ~new_n16607_;
  assign new_n19470_ = ~new_n15564_ | ~new_n32169_;
  assign new_n19471_ = ~new_n15552_ | ~new_n32741_;
  assign new_n19472_ = ~pi1382 | ~new_n16607_;
  assign new_n19473_ = ~new_n15564_ | ~new_n32167_;
  assign new_n19474_ = ~new_n15552_ | ~new_n32740_;
  assign new_n19475_ = ~pi1383 | ~new_n16607_;
  assign new_n19476_ = ~new_n15564_ | ~new_n32103_;
  assign new_n19477_ = ~new_n15552_ | ~new_n32789_;
  assign new_n19478_ = ~pi1384 | ~new_n16607_;
  assign new_n19479_ = ~new_n15564_ | ~new_n32104_;
  assign new_n19480_ = ~new_n15552_ | ~new_n32788_;
  assign new_n19481_ = ~pi1385 | ~new_n16607_;
  assign new_n19482_ = ~new_n15564_ | ~new_n32208_;
  assign new_n19483_ = ~new_n15552_ | ~new_n32787_;
  assign new_n19484_ = ~pi1386 | ~new_n16607_;
  assign new_n19485_ = ~new_n15564_ | ~new_n32206_;
  assign new_n19486_ = ~new_n15552_ | ~new_n32786_;
  assign new_n19487_ = ~pi1387 | ~new_n16607_;
  assign new_n19488_ = ~new_n15564_ | ~new_n32105_;
  assign new_n19489_ = ~new_n15552_ | ~new_n32785_;
  assign new_n19490_ = ~pi1388 | ~new_n16607_;
  assign new_n19491_ = ~new_n15564_ | ~new_n32106_;
  assign new_n19492_ = ~new_n15552_ | ~new_n32784_;
  assign new_n19493_ = ~pi1389 | ~new_n16607_;
  assign new_n19494_ = ~new_n15564_ | ~new_n32204_;
  assign new_n19495_ = ~new_n15552_ | ~new_n32783_;
  assign new_n19496_ = ~pi1390 | ~new_n16607_;
  assign new_n19497_ = ~new_n15564_ | ~new_n32202_;
  assign new_n19498_ = ~new_n15552_ | ~new_n32782_;
  assign new_n19499_ = ~pi1391 | ~new_n16607_;
  assign new_n19500_ = ~new_n15564_ | ~new_n32200_;
  assign new_n19501_ = ~new_n15552_ | ~new_n32781_;
  assign new_n19502_ = ~pi1392 | ~new_n16607_;
  assign new_n19503_ = ~new_n15564_ | ~new_n32198_;
  assign new_n19504_ = ~new_n15552_ | ~new_n32780_;
  assign new_n19505_ = ~pi1393 | ~new_n16607_;
  assign new_n19506_ = ~new_n15564_ | ~new_n32194_;
  assign new_n19507_ = ~new_n15552_ | ~new_n32779_;
  assign new_n19508_ = ~pi1394 | ~new_n16607_;
  assign new_n19509_ = ~new_n15564_ | ~new_n32192_;
  assign new_n19510_ = ~new_n15552_ | ~new_n32778_;
  assign new_n19511_ = ~pi1395 | ~new_n16607_;
  assign new_n19512_ = ~new_n15564_ | ~new_n32190_;
  assign new_n19513_ = ~new_n15552_ | ~new_n32777_;
  assign new_n19514_ = ~pi1396 | ~new_n16607_;
  assign new_n19515_ = ~new_n15564_ | ~new_n32188_;
  assign new_n19516_ = ~new_n15552_ | ~new_n32776_;
  assign new_n19517_ = ~pi1397 | ~new_n16607_;
  assign new_n19518_ = ~new_n15564_ | ~new_n32186_;
  assign new_n19519_ = ~new_n15552_ | ~new_n32775_;
  assign new_n19520_ = ~pi1398 | ~new_n16607_;
  assign new_n19521_ = ~new_n15564_ | ~new_n32184_;
  assign new_n19522_ = ~new_n15552_ | ~new_n32774_;
  assign new_n19523_ = ~pi1399 | ~new_n16607_;
  assign new_n19524_ = ~new_n15564_ | ~new_n32182_;
  assign new_n19525_ = ~new_n15552_ | ~new_n32773_;
  assign new_n19526_ = ~pi1400 | ~new_n16607_;
  assign new_n19527_ = ~new_n15564_ | ~new_n32180_;
  assign new_n19528_ = ~new_n15552_ | ~new_n32772_;
  assign new_n19529_ = ~pi1401 | ~new_n16607_;
  assign new_n19530_ = ~new_n15564_ | ~new_n32178_;
  assign new_n19531_ = ~new_n15552_ | ~new_n32771_;
  assign new_n19532_ = ~pi1402 | ~new_n16607_;
  assign new_n19533_ = ~new_n15564_ | ~new_n32176_;
  assign new_n19534_ = ~new_n15552_ | ~new_n32770_;
  assign new_n19535_ = ~pi1403 | ~new_n16607_;
  assign new_n19536_ = ~new_n15564_ | ~new_n32174_;
  assign new_n19537_ = ~new_n15552_ | ~new_n32769_;
  assign new_n19538_ = ~pi1404 | ~new_n16607_;
  assign new_n19539_ = ~new_n15552_ | ~new_n32768_;
  assign new_n19540_ = ~pi1405 | ~new_n16607_;
  assign new_n19541_ = ~new_n17385_ | ~new_n9378_;
  assign new_n19542_ = ~new_n17383_ | ~new_n33065_;
  assign new_n19543_ = ~new_n17384_ | ~new_n16444_;
  assign new_n19544_ = ~new_n16612_;
  assign new_n19545_ = ~new_n17430_ | ~pi1074;
  assign new_n19546_ = ~new_n33164_ | ~pi1075;
  assign new_n19547_ = ~new_n19546_ | ~new_n19545_;
  assign new_n19548_ = pi1445 | new_n2972_;
  assign new_n19549_ = ~new_n15785_ | ~new_n32790_;
  assign new_n19550_ = ~pi1406 | ~new_n20666_;
  assign new_n19551_ = ~pi1374 | ~new_n20665_;
  assign new_n19552_ = ~new_n15610_ | ~new_n32165_;
  assign new_n19553_ = ~new_n15607_ | ~new_n31179_;
  assign new_n19554_ = ~new_n15554_ | ~pi1247;
  assign new_n19555_ = ~new_n15547_ | ~pi1247;
  assign new_n19556_ = ~new_n19544_ | ~pi1406;
  assign new_n19557_ = ~new_n15785_ | ~new_n32791_;
  assign new_n19558_ = ~new_n33295_ | ~new_n20666_;
  assign new_n19559_ = ~pi1375 | ~new_n20665_;
  assign new_n19560_ = ~new_n15610_ | ~new_n32196_;
  assign new_n19561_ = ~new_n15607_ | ~new_n31178_;
  assign new_n19562_ = ~new_n15554_ | ~pi1248;
  assign new_n19563_ = ~new_n15547_ | ~new_n33099_;
  assign new_n19564_ = ~new_n19544_ | ~pi1407;
  assign new_n19565_ = ~new_n15785_ | ~new_n32842_;
  assign new_n19566_ = ~new_n33362_ | ~new_n20666_;
  assign new_n19567_ = ~pi1376 | ~new_n20665_;
  assign new_n19568_ = ~new_n15610_ | ~new_n32107_;
  assign new_n19569_ = ~new_n15607_ | ~new_n31187_;
  assign new_n19570_ = ~new_n15554_ | ~pi1249;
  assign new_n19571_ = ~new_n15547_ | ~new_n33166_;
  assign new_n19572_ = ~new_n19544_ | ~pi1408;
  assign new_n19573_ = ~new_n15785_ | ~new_n32746_;
  assign new_n19574_ = ~new_n33359_ | ~new_n20666_;
  assign new_n19575_ = ~pi1377 | ~new_n20665_;
  assign new_n19576_ = ~new_n15610_ | ~new_n32108_;
  assign new_n19577_ = ~new_n15607_ | ~new_n31170_;
  assign new_n19578_ = ~new_n15554_ | ~pi1250;
  assign new_n19579_ = ~new_n15547_ | ~new_n33163_;
  assign new_n19580_ = ~new_n19544_ | ~pi1409;
  assign new_n19581_ = ~new_n15785_ | ~new_n32745_;
  assign new_n19582_ = ~new_n33358_ | ~new_n20666_;
  assign new_n19583_ = ~pi1378 | ~new_n20665_;
  assign new_n19584_ = ~new_n15610_ | ~new_n32173_;
  assign new_n19585_ = ~new_n15607_ | ~new_n31169_;
  assign new_n19586_ = ~new_n15554_ | ~pi1251;
  assign new_n19587_ = ~new_n15547_ | ~new_n33162_;
  assign new_n19588_ = ~new_n19544_ | ~pi1410;
  assign new_n19589_ = ~new_n15785_ | ~new_n32744_;
  assign new_n19590_ = ~new_n33357_ | ~new_n20666_;
  assign new_n19591_ = ~pi1379 | ~new_n20665_;
  assign new_n19592_ = ~new_n15610_ | ~new_n32171_;
  assign new_n19593_ = ~new_n31150_ | ~new_n15607_;
  assign new_n19594_ = ~new_n15554_ | ~pi1252;
  assign new_n19595_ = ~new_n15547_ | ~new_n33161_;
  assign new_n19596_ = ~new_n19544_ | ~pi1411;
  assign new_n19597_ = ~new_n15785_ | ~new_n32743_;
  assign new_n19598_ = ~new_n33356_ | ~new_n20666_;
  assign new_n19599_ = ~pi1380 | ~new_n20665_;
  assign new_n19600_ = ~new_n15554_ | ~pi1253;
  assign new_n19601_ = ~new_n15548_ | ~new_n32109_;
  assign new_n19602_ = ~new_n15547_ | ~new_n33160_;
  assign new_n19603_ = ~new_n19544_ | ~pi1412;
  assign new_n19604_ = ~new_n15785_ | ~new_n32742_;
  assign new_n19605_ = ~new_n33355_ | ~new_n20666_;
  assign new_n19606_ = ~pi1381 | ~new_n20665_;
  assign new_n19607_ = ~new_n15554_ | ~pi1254;
  assign new_n19608_ = ~new_n15548_ | ~new_n32110_;
  assign new_n19609_ = ~new_n15547_ | ~new_n33159_;
  assign new_n19610_ = ~new_n19544_ | ~pi1413;
  assign new_n19611_ = ~new_n15785_ | ~new_n32741_;
  assign new_n19612_ = ~new_n33354_ | ~new_n20666_;
  assign new_n19613_ = ~pi1382 | ~new_n20665_;
  assign new_n19614_ = ~new_n15554_ | ~pi1255;
  assign new_n19615_ = ~new_n15548_ | ~new_n32169_;
  assign new_n19616_ = ~new_n15547_ | ~new_n33158_;
  assign new_n19617_ = ~new_n19544_ | ~pi1414;
  assign new_n19618_ = ~new_n15785_ | ~new_n32740_;
  assign new_n19619_ = ~new_n33353_ | ~new_n20666_;
  assign new_n19620_ = ~pi1383 | ~new_n20665_;
  assign new_n19621_ = ~new_n15554_ | ~pi1256;
  assign new_n19622_ = ~new_n15548_ | ~new_n32167_;
  assign new_n19623_ = ~new_n15547_ | ~new_n33157_;
  assign new_n19624_ = ~new_n19544_ | ~pi1415;
  assign new_n19625_ = ~new_n15785_ | ~new_n32789_;
  assign new_n19626_ = ~new_n33382_ | ~new_n20666_;
  assign new_n19627_ = ~pi1384 | ~new_n20665_;
  assign new_n19628_ = ~new_n15554_ | ~pi1257;
  assign new_n19629_ = ~new_n15548_ | ~new_n32103_;
  assign new_n19630_ = ~new_n15547_ | ~new_n33186_;
  assign new_n19631_ = ~new_n19544_ | ~pi1416;
  assign new_n19632_ = ~new_n15785_ | ~new_n32788_;
  assign new_n19633_ = ~new_n33381_ | ~new_n20666_;
  assign new_n19634_ = ~pi1385 | ~new_n20665_;
  assign new_n19635_ = ~new_n15554_ | ~pi1258;
  assign new_n19636_ = ~new_n15548_ | ~new_n32104_;
  assign new_n19637_ = ~new_n15547_ | ~new_n33185_;
  assign new_n19638_ = ~new_n19544_ | ~pi1417;
  assign new_n19639_ = ~new_n15785_ | ~new_n32787_;
  assign new_n19640_ = ~new_n33380_ | ~new_n20666_;
  assign new_n19641_ = ~pi1386 | ~new_n20665_;
  assign new_n19642_ = ~new_n15554_ | ~pi1259;
  assign new_n19643_ = ~new_n15548_ | ~new_n32208_;
  assign new_n19644_ = ~new_n15547_ | ~new_n33184_;
  assign new_n19645_ = ~new_n19544_ | ~pi1418;
  assign new_n19646_ = ~new_n15785_ | ~new_n32786_;
  assign new_n19647_ = ~new_n33379_ | ~new_n20666_;
  assign new_n19648_ = ~pi1387 | ~new_n20665_;
  assign new_n19649_ = ~new_n15554_ | ~pi1260;
  assign new_n19650_ = ~new_n15548_ | ~new_n32206_;
  assign new_n19651_ = ~new_n15547_ | ~new_n33183_;
  assign new_n19652_ = ~new_n19544_ | ~pi1419;
  assign new_n19653_ = ~new_n15785_ | ~new_n32785_;
  assign new_n19654_ = ~new_n33378_ | ~new_n20666_;
  assign new_n19655_ = ~pi1388 | ~new_n20665_;
  assign new_n19656_ = ~new_n15554_ | ~pi1261;
  assign new_n19657_ = ~new_n15548_ | ~new_n32105_;
  assign new_n19658_ = ~new_n15547_ | ~new_n33182_;
  assign new_n19659_ = ~new_n19544_ | ~pi1420;
  assign new_n19660_ = ~new_n15785_ | ~new_n32784_;
  assign new_n19661_ = ~new_n33377_ | ~new_n20666_;
  assign new_n19662_ = ~pi1389 | ~new_n20665_;
  assign new_n19663_ = ~new_n15554_ | ~pi1262;
  assign new_n19664_ = ~new_n15548_ | ~new_n32106_;
  assign new_n19665_ = ~new_n15547_ | ~new_n33181_;
  assign new_n19666_ = ~new_n19544_ | ~pi1421;
  assign new_n19667_ = ~new_n15785_ | ~new_n32783_;
  assign new_n19668_ = ~new_n33376_ | ~new_n20666_;
  assign new_n19669_ = ~pi1390 | ~new_n20665_;
  assign new_n19670_ = ~new_n15554_ | ~pi1263;
  assign new_n19671_ = ~new_n15548_ | ~new_n32204_;
  assign new_n19672_ = ~new_n15547_ | ~new_n33180_;
  assign new_n19673_ = ~new_n19544_ | ~pi1422;
  assign new_n19674_ = ~new_n15785_ | ~new_n32782_;
  assign new_n19675_ = ~new_n33375_ | ~new_n20666_;
  assign new_n19676_ = ~pi1391 | ~new_n20665_;
  assign new_n19677_ = ~new_n15554_ | ~pi1264;
  assign new_n19678_ = ~new_n15548_ | ~new_n32202_;
  assign new_n19679_ = ~new_n15547_ | ~new_n33179_;
  assign new_n19680_ = ~new_n19544_ | ~pi1423;
  assign new_n19681_ = ~new_n15785_ | ~new_n32781_;
  assign new_n19682_ = ~new_n33374_ | ~new_n20666_;
  assign new_n19683_ = ~pi1392 | ~new_n20665_;
  assign new_n19684_ = ~new_n15554_ | ~pi1265;
  assign new_n19685_ = ~new_n15548_ | ~new_n32200_;
  assign new_n19686_ = ~new_n15547_ | ~new_n33178_;
  assign new_n19687_ = ~new_n19544_ | ~pi1424;
  assign new_n19688_ = ~new_n15785_ | ~new_n32780_;
  assign new_n19689_ = ~new_n33373_ | ~new_n20666_;
  assign new_n19690_ = ~pi1393 | ~new_n20665_;
  assign new_n19691_ = ~new_n15554_ | ~pi1266;
  assign new_n19692_ = ~new_n15548_ | ~new_n32198_;
  assign new_n19693_ = ~new_n15547_ | ~new_n33177_;
  assign new_n19694_ = ~new_n19544_ | ~pi1425;
  assign new_n19695_ = ~new_n15785_ | ~new_n32779_;
  assign new_n19696_ = ~new_n33372_ | ~new_n20666_;
  assign new_n19697_ = ~pi1394 | ~new_n20665_;
  assign new_n19698_ = ~new_n15554_ | ~pi1267;
  assign new_n19699_ = ~new_n15548_ | ~new_n32194_;
  assign new_n19700_ = ~new_n15547_ | ~new_n33176_;
  assign new_n19701_ = ~new_n19544_ | ~pi1426;
  assign new_n19702_ = ~new_n15785_ | ~new_n32778_;
  assign new_n19703_ = ~new_n33371_ | ~new_n20666_;
  assign new_n19704_ = ~pi1395 | ~new_n20665_;
  assign new_n19705_ = ~new_n15554_ | ~pi1268;
  assign new_n19706_ = ~new_n15548_ | ~new_n32192_;
  assign new_n19707_ = ~new_n15547_ | ~new_n33175_;
  assign new_n19708_ = ~new_n19544_ | ~pi1427;
  assign new_n19709_ = ~new_n15785_ | ~new_n32777_;
  assign new_n19710_ = ~new_n33370_ | ~new_n20666_;
  assign new_n19711_ = ~pi1396 | ~new_n20665_;
  assign new_n19712_ = ~new_n15554_ | ~pi1269;
  assign new_n19713_ = ~new_n15548_ | ~new_n32190_;
  assign new_n19714_ = ~new_n15547_ | ~new_n33174_;
  assign new_n19715_ = ~new_n19544_ | ~pi1428;
  assign new_n19716_ = ~new_n15785_ | ~new_n32776_;
  assign new_n19717_ = ~new_n33369_ | ~new_n20666_;
  assign new_n19718_ = ~pi1397 | ~new_n20665_;
  assign new_n19719_ = ~new_n15554_ | ~pi1270;
  assign new_n19720_ = ~new_n15548_ | ~new_n32188_;
  assign new_n19721_ = ~new_n15547_ | ~new_n33173_;
  assign new_n19722_ = ~new_n19544_ | ~pi1429;
  assign new_n19723_ = ~new_n15785_ | ~new_n32775_;
  assign new_n19724_ = ~new_n33368_ | ~new_n20666_;
  assign new_n19725_ = ~pi1398 | ~new_n20665_;
  assign new_n19726_ = ~new_n15554_ | ~pi1271;
  assign new_n19727_ = ~new_n15548_ | ~new_n32186_;
  assign new_n19728_ = ~new_n15547_ | ~new_n33172_;
  assign new_n19729_ = ~new_n19544_ | ~pi1430;
  assign new_n19730_ = ~new_n15785_ | ~new_n32774_;
  assign new_n19731_ = ~new_n33367_ | ~new_n20666_;
  assign new_n19732_ = ~pi1399 | ~new_n20665_;
  assign new_n19733_ = ~new_n15554_ | ~pi1272;
  assign new_n19734_ = ~new_n15548_ | ~new_n32184_;
  assign new_n19735_ = ~new_n15547_ | ~new_n33171_;
  assign new_n19736_ = ~new_n19544_ | ~pi1431;
  assign new_n19737_ = ~new_n15785_ | ~new_n32773_;
  assign new_n19738_ = ~new_n33366_ | ~new_n20666_;
  assign new_n19739_ = ~pi1400 | ~new_n20665_;
  assign new_n19740_ = ~new_n15554_ | ~pi1273;
  assign new_n19741_ = ~new_n15548_ | ~new_n32182_;
  assign new_n19742_ = ~new_n15547_ | ~new_n33170_;
  assign new_n19743_ = ~new_n19544_ | ~pi1432;
  assign new_n19744_ = ~new_n15785_ | ~new_n32772_;
  assign new_n19745_ = ~new_n33365_ | ~new_n20666_;
  assign new_n19746_ = ~pi1401 | ~new_n20665_;
  assign new_n19747_ = ~new_n15554_ | ~pi1274;
  assign new_n19748_ = ~new_n15548_ | ~new_n32180_;
  assign new_n19749_ = ~new_n15547_ | ~new_n33169_;
  assign new_n19750_ = ~new_n19544_ | ~pi1433;
  assign new_n19751_ = ~new_n15785_ | ~new_n32771_;
  assign new_n19752_ = ~new_n33364_ | ~new_n20666_;
  assign new_n19753_ = ~pi1402 | ~new_n20665_;
  assign new_n19754_ = ~new_n15554_ | ~pi1275;
  assign new_n19755_ = ~new_n15548_ | ~new_n32178_;
  assign new_n19756_ = ~new_n15547_ | ~new_n33168_;
  assign new_n19757_ = ~new_n19544_ | ~pi1434;
  assign new_n19758_ = ~new_n15785_ | ~new_n32770_;
  assign new_n19759_ = ~new_n33363_ | ~new_n20666_;
  assign new_n19760_ = ~pi1403 | ~new_n20665_;
  assign new_n19761_ = ~new_n15554_ | ~pi1276;
  assign new_n19762_ = ~new_n15548_ | ~new_n32176_;
  assign new_n19763_ = ~new_n15547_ | ~new_n33167_;
  assign new_n19764_ = ~new_n19544_ | ~pi1435;
  assign new_n19765_ = ~new_n15785_ | ~new_n32769_;
  assign new_n19766_ = ~new_n33361_ | ~new_n20666_;
  assign new_n19767_ = ~pi1404 | ~new_n20665_;
  assign new_n19768_ = ~new_n15554_ | ~pi1277;
  assign new_n19769_ = ~new_n15548_ | ~new_n32174_;
  assign new_n19770_ = ~new_n15547_ | ~new_n33165_;
  assign new_n19771_ = ~new_n19544_ | ~pi1436;
  assign new_n19772_ = ~new_n15785_ | ~new_n32768_;
  assign new_n19773_ = ~new_n33360_ | ~new_n20666_;
  assign new_n19774_ = ~pi1405 | ~new_n20665_;
  assign new_n19775_ = ~new_n15554_ | ~pi1278;
  assign new_n19776_ = ~new_n15548_ | ~new_n32111_;
  assign new_n19777_ = ~new_n15547_ | ~new_n33164_;
  assign new_n19778_ = ~new_n19544_ | ~pi1437;
  assign new_n19779_ = ~pi1042 | ~pi1041;
  assign new_n19780_ = pi1407 | pi1406;
  assign new_n19781_ = ~new_n17358_;
  assign new_n19782_ = ~pi1443 | ~new_n17358_;
  assign new_n19783_ = ~new_n17147_ | ~new_n15609_;
  assign new_n19784_ = ~new_n17361_;
  assign new_n19785_ = ~pi1445 | ~new_n17678_;
  assign new_n19786_ = ~new_n17389_ | ~new_n19785_;
  assign new_n19787_ = ~new_n17145_ | ~new_n19786_;
  assign new_n19788_ = ~pi1076 | ~new_n19787_;
  assign new_n19789_ = ~new_n17374_ | ~new_n16453_;
  assign new_n19790_ = ~new_n17146_ | ~new_n19788_;
  assign new_n19791_ = ~new_n15549_ | ~new_n15654_;
  assign new_n19792_ = ~pi1449 | ~new_n19791_;
  assign new_n19793_ = ~new_n17436_ | ~pi1076;
  assign new_n19794_ = ~pi1450 | ~pi1040;
  assign new_n19795_ = ~new_n17362_;
  assign new_n19796_ = ~new_n17149_ | ~new_n16472_;
  assign new_n19797_ = ~new_n16587_ | ~new_n17680_ | ~new_n17150_;
  assign new_n19798_ = ~pi1452 | ~new_n19797_;
  assign new_n19799_ = ~new_n15725_ | ~pi1077;
  assign new_n19800_ = ~new_n15724_ | ~pi1085;
  assign new_n19801_ = ~new_n15723_ | ~pi1093;
  assign new_n19802_ = ~new_n15722_ | ~pi1101;
  assign new_n19803_ = ~new_n15720_ | ~pi1109;
  assign new_n19804_ = ~new_n15719_ | ~pi1117;
  assign new_n19805_ = ~new_n15718_ | ~pi1125;
  assign new_n19806_ = ~new_n15717_ | ~pi1133;
  assign new_n19807_ = ~new_n15715_ | ~pi1141;
  assign new_n19808_ = ~new_n15714_ | ~pi1149;
  assign new_n19809_ = ~new_n15713_ | ~pi1157;
  assign new_n19810_ = ~new_n15712_ | ~pi1165;
  assign new_n19811_ = ~new_n15710_ | ~pi1173;
  assign new_n19812_ = ~new_n15708_ | ~pi1181;
  assign new_n19813_ = ~new_n15706_ | ~pi1189;
  assign new_n19814_ = ~new_n15704_ | ~pi1197;
  assign new_n19815_ = ~new_n15725_ | ~pi1078;
  assign new_n19816_ = ~new_n15724_ | ~pi1086;
  assign new_n19817_ = ~new_n15723_ | ~pi1094;
  assign new_n19818_ = ~new_n15722_ | ~pi1102;
  assign new_n19819_ = ~new_n15720_ | ~pi1110;
  assign new_n19820_ = ~new_n15719_ | ~pi1118;
  assign new_n19821_ = ~new_n15718_ | ~pi1126;
  assign new_n19822_ = ~new_n15717_ | ~pi1134;
  assign new_n19823_ = ~new_n15715_ | ~pi1142;
  assign new_n19824_ = ~new_n15714_ | ~pi1150;
  assign new_n19825_ = ~new_n15713_ | ~pi1158;
  assign new_n19826_ = ~new_n15712_ | ~pi1166;
  assign new_n19827_ = ~new_n15710_ | ~pi1174;
  assign new_n19828_ = ~new_n15708_ | ~pi1182;
  assign new_n19829_ = ~new_n15706_ | ~pi1190;
  assign new_n19830_ = ~new_n15704_ | ~pi1198;
  assign new_n19831_ = ~new_n15725_ | ~pi1079;
  assign new_n19832_ = ~new_n15724_ | ~pi1087;
  assign new_n19833_ = ~new_n15723_ | ~pi1095;
  assign new_n19834_ = ~new_n15722_ | ~pi1103;
  assign new_n19835_ = ~new_n15720_ | ~pi1111;
  assign new_n19836_ = ~new_n15719_ | ~pi1119;
  assign new_n19837_ = ~new_n15718_ | ~pi1127;
  assign new_n19838_ = ~new_n15717_ | ~pi1135;
  assign new_n19839_ = ~new_n15715_ | ~pi1143;
  assign new_n19840_ = ~new_n15714_ | ~pi1151;
  assign new_n19841_ = ~new_n15713_ | ~pi1159;
  assign new_n19842_ = ~new_n15712_ | ~pi1167;
  assign new_n19843_ = ~new_n15710_ | ~pi1175;
  assign new_n19844_ = ~new_n15708_ | ~pi1183;
  assign new_n19845_ = ~new_n15706_ | ~pi1191;
  assign new_n19846_ = ~new_n15704_ | ~pi1199;
  assign new_n19847_ = ~new_n15725_ | ~pi1080;
  assign new_n19848_ = ~new_n15724_ | ~pi1088;
  assign new_n19849_ = ~new_n15723_ | ~pi1096;
  assign new_n19850_ = ~new_n15722_ | ~pi1104;
  assign new_n19851_ = ~new_n15720_ | ~pi1112;
  assign new_n19852_ = ~new_n15719_ | ~pi1120;
  assign new_n19853_ = ~new_n15718_ | ~pi1128;
  assign new_n19854_ = ~new_n15717_ | ~pi1136;
  assign new_n19855_ = ~new_n15715_ | ~pi1144;
  assign new_n19856_ = ~new_n15714_ | ~pi1152;
  assign new_n19857_ = ~new_n15713_ | ~pi1160;
  assign new_n19858_ = ~new_n15712_ | ~pi1168;
  assign new_n19859_ = ~new_n15710_ | ~pi1176;
  assign new_n19860_ = ~new_n15708_ | ~pi1184;
  assign new_n19861_ = ~new_n15706_ | ~pi1192;
  assign new_n19862_ = ~new_n15725_ | ~pi1081;
  assign new_n19863_ = ~new_n15724_ | ~pi1089;
  assign new_n19864_ = ~new_n15723_ | ~pi1097;
  assign new_n19865_ = ~new_n15722_ | ~pi1105;
  assign new_n19866_ = ~new_n15720_ | ~pi1113;
  assign new_n19867_ = ~new_n15719_ | ~pi1121;
  assign new_n19868_ = ~new_n15718_ | ~pi1129;
  assign new_n19869_ = ~new_n15717_ | ~pi1137;
  assign new_n19870_ = ~new_n15715_ | ~pi1145;
  assign new_n19871_ = ~new_n15714_ | ~pi1153;
  assign new_n19872_ = ~new_n15713_ | ~pi1161;
  assign new_n19873_ = ~new_n15712_ | ~pi1169;
  assign new_n19874_ = ~new_n15710_ | ~pi1177;
  assign new_n19875_ = ~new_n15708_ | ~pi1185;
  assign new_n19876_ = ~new_n15706_ | ~pi1193;
  assign new_n19877_ = ~new_n15704_ | ~pi1201;
  assign new_n19878_ = ~new_n15725_ | ~pi1082;
  assign new_n19879_ = ~new_n15724_ | ~pi1090;
  assign new_n19880_ = ~new_n15723_ | ~pi1098;
  assign new_n19881_ = ~new_n15722_ | ~pi1106;
  assign new_n19882_ = ~new_n15720_ | ~pi1114;
  assign new_n19883_ = ~new_n15719_ | ~pi1122;
  assign new_n19884_ = ~new_n15718_ | ~pi1130;
  assign new_n19885_ = ~new_n15717_ | ~pi1138;
  assign new_n19886_ = ~new_n15715_ | ~pi1146;
  assign new_n19887_ = ~new_n15714_ | ~pi1154;
  assign new_n19888_ = ~new_n15713_ | ~pi1162;
  assign new_n19889_ = ~new_n15712_ | ~pi1170;
  assign new_n19890_ = ~new_n15710_ | ~pi1178;
  assign new_n19891_ = ~new_n15708_ | ~pi1186;
  assign new_n19892_ = ~new_n15706_ | ~pi1194;
  assign new_n19893_ = ~new_n15704_ | ~pi1202;
  assign new_n19894_ = ~new_n15725_ | ~pi1083;
  assign new_n19895_ = ~new_n15724_ | ~pi1091;
  assign new_n19896_ = ~new_n15723_ | ~pi1099;
  assign new_n19897_ = ~new_n15722_ | ~pi1107;
  assign new_n19898_ = ~new_n15720_ | ~pi1115;
  assign new_n19899_ = ~new_n15719_ | ~pi1123;
  assign new_n19900_ = ~new_n15718_ | ~pi1131;
  assign new_n19901_ = ~new_n15717_ | ~pi1139;
  assign new_n19902_ = ~new_n15715_ | ~pi1147;
  assign new_n19903_ = ~new_n15714_ | ~pi1155;
  assign new_n19904_ = ~new_n15713_ | ~pi1163;
  assign new_n19905_ = ~new_n15712_ | ~pi1171;
  assign new_n19906_ = ~new_n15710_ | ~pi1179;
  assign new_n19907_ = ~new_n15708_ | ~pi1187;
  assign new_n19908_ = ~new_n15706_ | ~pi1195;
  assign new_n19909_ = ~new_n15704_ | ~pi1203;
  assign new_n19910_ = ~new_n15725_ | ~pi1084;
  assign new_n19911_ = ~new_n15724_ | ~pi1092;
  assign new_n19912_ = ~new_n15723_ | ~pi1100;
  assign new_n19913_ = ~new_n15722_ | ~pi1108;
  assign new_n19914_ = ~new_n15720_ | ~pi1116;
  assign new_n19915_ = ~new_n15719_ | ~pi1124;
  assign new_n19916_ = ~new_n15718_ | ~pi1132;
  assign new_n19917_ = ~new_n15717_ | ~pi1140;
  assign new_n19918_ = ~new_n15715_ | ~pi1148;
  assign new_n19919_ = ~new_n15714_ | ~pi1156;
  assign new_n19920_ = ~new_n15713_ | ~pi1164;
  assign new_n19921_ = ~new_n15712_ | ~pi1172;
  assign new_n19922_ = ~new_n15710_ | ~pi1180;
  assign new_n19923_ = ~new_n15708_ | ~pi1188;
  assign new_n19924_ = ~new_n15706_ | ~pi1196;
  assign new_n19925_ = ~new_n15704_ | ~pi1204;
  assign new_n19926_ = ~new_n17641_ | ~pi1074;
  assign new_n19927_ = ~new_n16593_ | ~new_n19926_;
  assign new_n19928_ = ~new_n17369_ | ~pi1351;
  assign new_n19929_ = ~new_n17368_ | ~pi1256;
  assign new_n19930_ = ~new_n33157_ | ~new_n15533_;
  assign new_n19931_ = ~new_n17369_ | ~pi1350;
  assign new_n19932_ = ~new_n17368_ | ~pi1255;
  assign new_n19933_ = ~new_n33158_ | ~new_n15533_;
  assign new_n19934_ = ~new_n17369_ | ~pi1349;
  assign new_n19935_ = ~new_n17368_ | ~pi1254;
  assign new_n19936_ = ~new_n33159_ | ~new_n15533_;
  assign new_n19937_ = ~new_n17369_ | ~pi1348;
  assign new_n19938_ = ~new_n17368_ | ~pi1253;
  assign new_n19939_ = ~new_n33160_ | ~new_n15533_;
  assign new_n19940_ = ~new_n31150_ | ~new_n19927_;
  assign new_n19941_ = ~new_n17369_ | ~pi1347;
  assign new_n19942_ = ~new_n17368_ | ~pi1252;
  assign new_n19943_ = ~new_n33161_ | ~new_n15533_;
  assign new_n19944_ = ~new_n31169_ | ~new_n19927_;
  assign new_n19945_ = ~new_n17369_ | ~pi1346;
  assign new_n19946_ = ~new_n17368_ | ~pi1251;
  assign new_n19947_ = ~new_n33162_ | ~new_n15533_;
  assign new_n19948_ = ~new_n15534_ | ~pi1205;
  assign new_n19949_ = ~new_n17369_ | ~pi1373;
  assign new_n19950_ = ~new_n17368_ | ~pi1278;
  assign new_n19951_ = ~new_n33164_ | ~new_n15533_;
  assign new_n19952_ = ~new_n31171_ | ~new_n19927_;
  assign new_n19953_ = ~new_n17369_ | ~pi1372;
  assign new_n19954_ = ~new_n17368_ | ~pi1277;
  assign new_n19955_ = ~new_n33165_ | ~new_n15533_;
  assign new_n19956_ = ~new_n31170_ | ~new_n19927_;
  assign new_n19957_ = ~new_n17369_ | ~pi1345;
  assign new_n19958_ = ~new_n17368_ | ~pi1250;
  assign new_n19959_ = ~new_n33163_ | ~new_n15533_;
  assign new_n19960_ = ~new_n15534_ | ~pi1206;
  assign new_n19961_ = ~new_n31172_ | ~new_n19927_;
  assign new_n19962_ = ~new_n17369_ | ~pi1371;
  assign new_n19963_ = ~new_n17368_ | ~pi1276;
  assign new_n19964_ = ~new_n33167_ | ~new_n15533_;
  assign new_n19965_ = ~new_n31173_ | ~new_n19927_;
  assign new_n19966_ = ~new_n17369_ | ~pi1370;
  assign new_n19967_ = ~new_n17368_ | ~pi1275;
  assign new_n19968_ = ~new_n33168_ | ~new_n15533_;
  assign new_n19969_ = ~new_n31174_ | ~new_n19927_;
  assign new_n19970_ = ~new_n17369_ | ~pi1369;
  assign new_n19971_ = ~new_n17368_ | ~pi1274;
  assign new_n19972_ = ~new_n33169_ | ~new_n15533_;
  assign new_n19973_ = ~new_n31175_ | ~new_n19927_;
  assign new_n19974_ = ~new_n17369_ | ~pi1368;
  assign new_n19975_ = ~new_n17368_ | ~pi1273;
  assign new_n19976_ = ~new_n33170_ | ~new_n15533_;
  assign new_n19977_ = ~new_n31176_ | ~new_n19927_;
  assign new_n19978_ = ~new_n17369_ | ~pi1367;
  assign new_n19979_ = ~new_n17368_ | ~pi1272;
  assign new_n19980_ = ~new_n33171_ | ~new_n15533_;
  assign new_n19981_ = ~new_n31177_ | ~new_n19927_;
  assign new_n19982_ = ~new_n17369_ | ~pi1366;
  assign new_n19983_ = ~new_n17368_ | ~pi1271;
  assign new_n19984_ = ~new_n33172_ | ~new_n15533_;
  assign new_n19985_ = ~new_n31151_ | ~new_n19927_;
  assign new_n19986_ = ~new_n17369_ | ~pi1365;
  assign new_n19987_ = ~new_n17368_ | ~pi1270;
  assign new_n19988_ = ~new_n33173_ | ~new_n15533_;
  assign new_n19989_ = ~new_n15905_ | ~new_n19927_;
  assign new_n19990_ = ~new_n17369_ | ~pi1364;
  assign new_n19991_ = ~new_n17368_ | ~pi1269;
  assign new_n19992_ = ~new_n33174_ | ~new_n15533_;
  assign new_n19993_ = ~new_n15906_ | ~new_n19927_;
  assign new_n19994_ = ~new_n17369_ | ~pi1363;
  assign new_n19995_ = ~new_n17368_ | ~pi1268;
  assign new_n19996_ = ~new_n33175_ | ~new_n15533_;
  assign new_n19997_ = ~new_n15907_ | ~new_n19927_;
  assign new_n19998_ = ~new_n17369_ | ~pi1362;
  assign new_n19999_ = ~new_n17368_ | ~pi1267;
  assign new_n20000_ = ~new_n33176_ | ~new_n15533_;
  assign new_n20001_ = ~new_n31187_ | ~new_n19927_;
  assign new_n20002_ = ~new_n17369_ | ~pi1344;
  assign new_n20003_ = ~new_n17368_ | ~pi1249;
  assign new_n20004_ = ~new_n33166_ | ~new_n15533_;
  assign new_n20005_ = ~new_n15534_ | ~pi1207;
  assign new_n20006_ = ~new_n15908_ | ~new_n19927_;
  assign new_n20007_ = ~new_n17369_ | ~pi1361;
  assign new_n20008_ = ~new_n17368_ | ~pi1266;
  assign new_n20009_ = ~new_n33177_ | ~new_n15533_;
  assign new_n20010_ = ~new_n15909_ | ~new_n19927_;
  assign new_n20011_ = ~new_n17369_ | ~pi1360;
  assign new_n20012_ = ~new_n17368_ | ~pi1265;
  assign new_n20013_ = ~new_n33178_ | ~new_n15533_;
  assign new_n20014_ = ~new_n15910_ | ~new_n19927_;
  assign new_n20015_ = ~new_n17369_ | ~pi1359;
  assign new_n20016_ = ~new_n17368_ | ~pi1264;
  assign new_n20017_ = ~new_n33179_ | ~new_n15533_;
  assign new_n20018_ = ~new_n15911_ | ~new_n19927_;
  assign new_n20019_ = ~new_n17369_ | ~pi1358;
  assign new_n20020_ = ~new_n17368_ | ~pi1263;
  assign new_n20021_ = ~new_n33180_ | ~new_n15533_;
  assign new_n20022_ = ~new_n17369_ | ~pi1357;
  assign new_n20023_ = ~new_n17368_ | ~pi1262;
  assign new_n20024_ = ~new_n33181_ | ~new_n15533_;
  assign new_n20025_ = ~new_n17369_ | ~pi1356;
  assign new_n20026_ = ~new_n17368_ | ~pi1261;
  assign new_n20027_ = ~new_n33182_ | ~new_n15533_;
  assign new_n20028_ = ~new_n17369_ | ~pi1355;
  assign new_n20029_ = ~new_n17368_ | ~pi1260;
  assign new_n20030_ = ~new_n33183_ | ~new_n15533_;
  assign new_n20031_ = ~new_n17369_ | ~pi1354;
  assign new_n20032_ = ~new_n17368_ | ~pi1259;
  assign new_n20033_ = ~new_n33184_ | ~new_n15533_;
  assign new_n20034_ = ~new_n17369_ | ~pi1353;
  assign new_n20035_ = ~new_n17368_ | ~pi1258;
  assign new_n20036_ = ~new_n33185_ | ~new_n15533_;
  assign new_n20037_ = ~new_n17369_ | ~pi1352;
  assign new_n20038_ = ~new_n17368_ | ~pi1257;
  assign new_n20039_ = ~new_n33186_ | ~new_n15533_;
  assign new_n20040_ = ~new_n31178_ | ~new_n19927_;
  assign new_n20041_ = ~new_n17369_ | ~pi1343;
  assign new_n20042_ = ~new_n17368_ | ~pi1248;
  assign new_n20043_ = ~new_n33099_ | ~new_n15533_;
  assign new_n20044_ = ~new_n15534_ | ~pi1208;
  assign new_n20045_ = ~new_n31179_ | ~new_n19927_;
  assign new_n20046_ = ~new_n17369_ | ~pi1342;
  assign new_n20047_ = ~new_n17368_ | ~pi1247;
  assign new_n20048_ = ~pi1247 | ~new_n15533_;
  assign new_n20049_ = ~new_n15534_ | ~pi1209;
  assign new_n20050_ = ~new_n31276_ | ~new_n19927_;
  assign new_n20051_ = ~new_n16490_ | ~new_n16620_ | ~new_n17641_;
  assign new_n20052_ = ~new_n17340_ | ~new_n31307_;
  assign new_n20053_ = ~new_n33621_ | ~new_n17389_;
  assign new_n20054_ = ~new_n17340_ | ~new_n31237_;
  assign new_n20055_ = ~new_n33636_ | ~new_n17389_;
  assign new_n20056_ = ~new_n17340_ | ~new_n31236_;
  assign new_n20057_ = ~new_n33632_ | ~new_n17389_;
  assign new_n20058_ = ~new_n17340_ | ~new_n31272_;
  assign new_n20059_ = ~new_n33634_ | ~new_n17389_;
  assign new_n20060_ = ~new_n17340_ | ~new_n31274_;
  assign new_n20061_ = ~new_n33633_ | ~new_n17389_;
  assign new_n20062_ = ~new_n17340_ | ~new_n31235_;
  assign new_n20063_ = ~new_n33639_ | ~new_n17389_;
  assign new_n20064_ = ~new_n17340_ | ~new_n31276_;
  assign new_n20065_ = ~new_n33620_ | ~new_n17389_;
  assign new_n20066_ = ~new_n17675_ | ~new_n16464_;
  assign new_n20067_ = ~new_n17340_ | ~new_n31277_;
  assign new_n20068_ = ~new_n33635_ | ~new_n17389_;
  assign new_n20069_ = ~new_n15786_ | ~new_n16465_;
  assign new_n20070_ = ~new_n17340_ | ~new_n31270_;
  assign new_n20071_ = ~new_n33619_ | ~new_n17389_;
  assign new_n20072_ = ~new_n17675_ | ~new_n16464_;
  assign new_n20073_ = ~new_n15745_ | ~pi1083;
  assign new_n20074_ = ~new_n15744_ | ~pi1091;
  assign new_n20075_ = ~new_n15743_ | ~pi1099;
  assign new_n20076_ = ~new_n15742_ | ~pi1107;
  assign new_n20077_ = ~new_n15740_ | ~pi1115;
  assign new_n20078_ = ~new_n15739_ | ~pi1123;
  assign new_n20079_ = ~new_n15738_ | ~pi1131;
  assign new_n20080_ = ~new_n15737_ | ~pi1139;
  assign new_n20081_ = ~new_n15735_ | ~pi1147;
  assign new_n20082_ = ~new_n15734_ | ~pi1155;
  assign new_n20083_ = ~new_n15733_ | ~pi1163;
  assign new_n20084_ = ~new_n15732_ | ~pi1171;
  assign new_n20085_ = ~new_n15730_ | ~pi1179;
  assign new_n20086_ = ~new_n15729_ | ~pi1187;
  assign new_n20087_ = ~new_n15728_ | ~pi1195;
  assign new_n20088_ = ~new_n15727_ | ~pi1203;
  assign new_n20089_ = ~new_n17212_ | ~new_n17210_ | ~new_n17211_ | ~new_n17213_;
  assign new_n20090_ = ~new_n16586_ | ~new_n16599_;
  assign new_n20091_ = ~new_n15745_ | ~pi1084;
  assign new_n20092_ = ~new_n15744_ | ~pi1092;
  assign new_n20093_ = ~new_n15743_ | ~pi1100;
  assign new_n20094_ = ~new_n15742_ | ~pi1108;
  assign new_n20095_ = ~new_n15740_ | ~pi1116;
  assign new_n20096_ = ~new_n15739_ | ~pi1124;
  assign new_n20097_ = ~new_n15738_ | ~pi1132;
  assign new_n20098_ = ~new_n15737_ | ~pi1140;
  assign new_n20099_ = ~new_n15735_ | ~pi1148;
  assign new_n20100_ = ~new_n15734_ | ~pi1156;
  assign new_n20101_ = ~new_n15733_ | ~pi1164;
  assign new_n20102_ = ~new_n15732_ | ~pi1172;
  assign new_n20103_ = ~new_n15730_ | ~pi1180;
  assign new_n20104_ = ~new_n15729_ | ~pi1188;
  assign new_n20105_ = ~new_n15728_ | ~pi1196;
  assign new_n20106_ = ~new_n15727_ | ~pi1204;
  assign new_n20107_ = ~new_n17216_ | ~new_n17214_ | ~new_n17215_ | ~new_n17217_;
  assign new_n20108_ = ~new_n17388_ | ~new_n16415_;
  assign new_n20109_ = ~new_n15536_ | ~new_n33280_;
  assign new_n20110_ = ~new_n17388_ | ~new_n16414_;
  assign new_n20111_ = ~new_n33278_ | ~new_n15536_;
  assign new_n20112_ = ~new_n17388_ | ~new_n16413_;
  assign new_n20113_ = ~new_n33281_ | ~new_n15536_;
  assign new_n20114_ = ~new_n17388_ | ~new_n16412_;
  assign new_n20115_ = ~new_n33285_ | ~new_n15536_;
  assign new_n20116_ = ~new_n17388_ | ~new_n16411_;
  assign new_n20117_ = ~new_n33283_ | ~new_n15536_;
  assign new_n20118_ = ~new_n31170_ | ~new_n16475_;
  assign new_n20119_ = ~new_n17388_ | ~new_n16410_;
  assign new_n20120_ = ~new_n33284_ | ~new_n15536_;
  assign new_n20121_ = ~new_n31187_ | ~new_n16475_;
  assign new_n20122_ = ~new_n15745_ | ~pi1077;
  assign new_n20123_ = ~new_n15744_ | ~pi1085;
  assign new_n20124_ = ~new_n15743_ | ~pi1093;
  assign new_n20125_ = ~new_n15742_ | ~pi1101;
  assign new_n20126_ = ~new_n15740_ | ~pi1109;
  assign new_n20127_ = ~new_n15739_ | ~pi1117;
  assign new_n20128_ = ~new_n15738_ | ~pi1125;
  assign new_n20129_ = ~new_n15737_ | ~pi1133;
  assign new_n20130_ = ~new_n15735_ | ~pi1141;
  assign new_n20131_ = ~new_n15734_ | ~pi1149;
  assign new_n20132_ = ~new_n15733_ | ~pi1157;
  assign new_n20133_ = ~new_n15732_ | ~pi1165;
  assign new_n20134_ = ~new_n15730_ | ~pi1173;
  assign new_n20135_ = ~new_n15729_ | ~pi1181;
  assign new_n20136_ = ~new_n15728_ | ~pi1189;
  assign new_n20137_ = ~new_n15727_ | ~pi1197;
  assign new_n20138_ = ~new_n17220_ | ~new_n17218_ | ~new_n17219_ | ~new_n17221_;
  assign new_n20139_ = ~new_n15745_ | ~pi1078;
  assign new_n20140_ = ~new_n15744_ | ~pi1086;
  assign new_n20141_ = ~new_n15743_ | ~pi1094;
  assign new_n20142_ = ~new_n15742_ | ~pi1102;
  assign new_n20143_ = ~new_n15740_ | ~pi1110;
  assign new_n20144_ = ~new_n15739_ | ~pi1118;
  assign new_n20145_ = ~new_n15738_ | ~pi1126;
  assign new_n20146_ = ~new_n15737_ | ~pi1134;
  assign new_n20147_ = ~new_n15735_ | ~pi1142;
  assign new_n20148_ = ~new_n15734_ | ~pi1150;
  assign new_n20149_ = ~new_n15733_ | ~pi1158;
  assign new_n20150_ = ~new_n15732_ | ~pi1166;
  assign new_n20151_ = ~new_n15730_ | ~pi1174;
  assign new_n20152_ = ~new_n15729_ | ~pi1182;
  assign new_n20153_ = ~new_n15728_ | ~pi1190;
  assign new_n20154_ = ~new_n15727_ | ~pi1198;
  assign new_n20155_ = ~new_n17224_ | ~new_n17222_ | ~new_n17223_ | ~new_n17225_;
  assign new_n20156_ = ~new_n15745_ | ~pi1079;
  assign new_n20157_ = ~new_n15744_ | ~pi1087;
  assign new_n20158_ = ~new_n15743_ | ~pi1095;
  assign new_n20159_ = ~new_n15742_ | ~pi1103;
  assign new_n20160_ = ~new_n15740_ | ~pi1111;
  assign new_n20161_ = ~new_n15739_ | ~pi1119;
  assign new_n20162_ = ~new_n15738_ | ~pi1127;
  assign new_n20163_ = ~new_n15737_ | ~pi1135;
  assign new_n20164_ = ~new_n15735_ | ~pi1143;
  assign new_n20165_ = ~new_n15734_ | ~pi1151;
  assign new_n20166_ = ~new_n15733_ | ~pi1159;
  assign new_n20167_ = ~new_n15732_ | ~pi1167;
  assign new_n20168_ = ~new_n15730_ | ~pi1175;
  assign new_n20169_ = ~new_n15729_ | ~pi1183;
  assign new_n20170_ = ~new_n15728_ | ~pi1191;
  assign new_n20171_ = ~new_n15727_ | ~pi1199;
  assign new_n20172_ = ~new_n17228_ | ~new_n17226_ | ~new_n17227_ | ~new_n17229_;
  assign new_n20173_ = ~new_n15745_ | ~pi1080;
  assign new_n20174_ = ~new_n15744_ | ~pi1088;
  assign new_n20175_ = ~new_n15743_ | ~pi1096;
  assign new_n20176_ = ~new_n15742_ | ~pi1104;
  assign new_n20177_ = ~new_n15740_ | ~pi1112;
  assign new_n20178_ = ~new_n15739_ | ~pi1120;
  assign new_n20179_ = ~new_n15738_ | ~pi1128;
  assign new_n20180_ = ~new_n15737_ | ~pi1136;
  assign new_n20181_ = ~new_n15735_ | ~pi1144;
  assign new_n20182_ = ~new_n15734_ | ~pi1152;
  assign new_n20183_ = ~new_n15733_ | ~pi1160;
  assign new_n20184_ = ~new_n15732_ | ~pi1168;
  assign new_n20185_ = ~new_n15730_ | ~pi1176;
  assign new_n20186_ = ~new_n15729_ | ~pi1184;
  assign new_n20187_ = ~new_n15728_ | ~pi1192;
  assign new_n20188_ = ~new_n15745_ | ~pi1081;
  assign new_n20189_ = ~new_n15744_ | ~pi1089;
  assign new_n20190_ = ~new_n15743_ | ~pi1097;
  assign new_n20191_ = ~new_n15742_ | ~pi1105;
  assign new_n20192_ = ~new_n15740_ | ~pi1113;
  assign new_n20193_ = ~new_n15739_ | ~pi1121;
  assign new_n20194_ = ~new_n15738_ | ~pi1129;
  assign new_n20195_ = ~new_n15737_ | ~pi1137;
  assign new_n20196_ = ~new_n15735_ | ~pi1145;
  assign new_n20197_ = ~new_n15734_ | ~pi1153;
  assign new_n20198_ = ~new_n15733_ | ~pi1161;
  assign new_n20199_ = ~new_n15732_ | ~pi1169;
  assign new_n20200_ = ~new_n15730_ | ~pi1177;
  assign new_n20201_ = ~new_n15729_ | ~pi1185;
  assign new_n20202_ = ~new_n15728_ | ~pi1193;
  assign new_n20203_ = ~new_n15727_ | ~pi1201;
  assign new_n20204_ = ~new_n17236_ | ~new_n17234_ | ~new_n17235_ | ~new_n17237_;
  assign new_n20205_ = ~new_n15745_ | ~pi1082;
  assign new_n20206_ = ~new_n15744_ | ~pi1090;
  assign new_n20207_ = ~new_n15743_ | ~pi1098;
  assign new_n20208_ = ~new_n15742_ | ~pi1106;
  assign new_n20209_ = ~new_n15740_ | ~pi1114;
  assign new_n20210_ = ~new_n15739_ | ~pi1122;
  assign new_n20211_ = ~new_n15738_ | ~pi1130;
  assign new_n20212_ = ~new_n15737_ | ~pi1138;
  assign new_n20213_ = ~new_n15735_ | ~pi1146;
  assign new_n20214_ = ~new_n15734_ | ~pi1154;
  assign new_n20215_ = ~new_n15733_ | ~pi1162;
  assign new_n20216_ = ~new_n15732_ | ~pi1170;
  assign new_n20217_ = ~new_n15730_ | ~pi1178;
  assign new_n20218_ = ~new_n15729_ | ~pi1186;
  assign new_n20219_ = ~new_n15728_ | ~pi1194;
  assign new_n20220_ = ~new_n15727_ | ~pi1202;
  assign new_n20221_ = ~new_n17240_ | ~new_n17238_ | ~new_n17239_ | ~new_n17241_;
  assign new_n20222_ = ~new_n17388_ | ~new_n16409_;
  assign new_n20223_ = ~new_n33279_ | ~new_n15536_;
  assign new_n20224_ = ~new_n31178_ | ~new_n16475_;
  assign new_n20225_ = ~new_n17388_ | ~new_n16408_;
  assign new_n20226_ = ~new_n33282_ | ~new_n15536_;
  assign new_n20227_ = ~new_n31179_ | ~new_n16475_;
  assign new_n20228_ = ~new_n17387_ | ~new_n16415_;
  assign new_n20229_ = ~new_n17373_ | ~pi1197;
  assign new_n20230_ = ~new_n17387_ | ~new_n16414_;
  assign new_n20231_ = ~new_n17373_ | ~pi1198;
  assign new_n20232_ = ~new_n17387_ | ~new_n16413_;
  assign new_n20233_ = ~new_n17373_ | ~pi1199;
  assign new_n20234_ = ~new_n17387_ | ~new_n16412_;
  assign new_n20235_ = ~new_n17387_ | ~new_n16411_;
  assign new_n20236_ = ~new_n17373_ | ~pi1201;
  assign new_n20237_ = ~new_n17387_ | ~new_n16410_;
  assign new_n20238_ = ~new_n17373_ | ~pi1202;
  assign new_n20239_ = ~new_n17387_ | ~new_n16409_;
  assign new_n20240_ = ~new_n17373_ | ~pi1203;
  assign new_n20241_ = ~new_n17387_ | ~new_n16408_;
  assign new_n20242_ = ~new_n16415_ | ~new_n17581_;
  assign new_n20243_ = ~new_n17373_ | ~pi1204;
  assign new_n20244_ = ~new_n16609_ | ~new_n16608_;
  assign new_n20245_ = ~pi1206 | ~new_n16445_;
  assign new_n20246_ = ~new_n16626_;
  assign new_n20247_ = ~new_n15763_ | ~pi1133;
  assign new_n20248_ = ~new_n15762_ | ~pi1125;
  assign new_n20249_ = ~new_n15761_ | ~pi1117;
  assign new_n20250_ = ~new_n15760_ | ~pi1109;
  assign new_n20251_ = ~new_n15758_ | ~pi1101;
  assign new_n20252_ = ~new_n15757_ | ~pi1093;
  assign new_n20253_ = ~new_n15756_ | ~pi1085;
  assign new_n20254_ = ~new_n15755_ | ~pi1077;
  assign new_n20255_ = ~new_n15754_ | ~pi1197;
  assign new_n20256_ = ~new_n15753_ | ~pi1189;
  assign new_n20257_ = ~new_n15752_ | ~pi1181;
  assign new_n20258_ = ~new_n15751_ | ~pi1173;
  assign new_n20259_ = ~new_n15749_ | ~pi1165;
  assign new_n20260_ = ~new_n15748_ | ~pi1157;
  assign new_n20261_ = ~new_n15747_ | ~pi1149;
  assign new_n20262_ = ~new_n15746_ | ~pi1141;
  assign new_n20263_ = ~new_n17246_ | ~new_n17244_ | ~new_n17245_ | ~new_n17247_;
  assign new_n20264_ = ~new_n16606_ | ~new_n16602_;
  assign new_n20265_ = ~new_n17254_ | ~new_n17372_;
  assign new_n20266_ = ~new_n20265_ | ~new_n16603_;
  assign new_n20267_ = ~new_n17684_ | ~new_n16459_;
  assign new_n20268_ = ~new_n16426_;
  assign new_n20269_ = ~new_n17684_ | ~new_n16575_ | ~new_n17335_ | ~new_n17581_;
  assign new_n20270_ = ~new_n17370_ | ~pi1076;
  assign new_n20271_ = ~new_n17248_ | ~new_n16426_;
  assign new_n20272_ = ~new_n16632_;
  assign new_n20273_ = ~new_n20810_ | ~new_n16632_ | ~new_n18673_;
  assign new_n20274_ = ~new_n17375_ | ~new_n20273_;
  assign new_n20275_ = ~new_n16631_;
  assign new_n20276_ = ~pi1211 | ~new_n16478_;
  assign new_n20277_ = ~pi1206 | ~new_n16631_;
  assign new_n20278_ = ~new_n17384_ | ~new_n16541_;
  assign new_n20279_ = ~new_n15763_ | ~pi1134;
  assign new_n20280_ = ~new_n15762_ | ~pi1126;
  assign new_n20281_ = ~new_n15761_ | ~pi1118;
  assign new_n20282_ = ~new_n15760_ | ~pi1110;
  assign new_n20283_ = ~new_n15758_ | ~pi1102;
  assign new_n20284_ = ~new_n15757_ | ~pi1094;
  assign new_n20285_ = ~new_n15756_ | ~pi1086;
  assign new_n20286_ = ~new_n15755_ | ~pi1078;
  assign new_n20287_ = ~new_n15754_ | ~pi1198;
  assign new_n20288_ = ~new_n15753_ | ~pi1190;
  assign new_n20289_ = ~new_n15752_ | ~pi1182;
  assign new_n20290_ = ~new_n15751_ | ~pi1174;
  assign new_n20291_ = ~new_n15749_ | ~pi1166;
  assign new_n20292_ = ~new_n15748_ | ~pi1158;
  assign new_n20293_ = ~new_n15747_ | ~pi1150;
  assign new_n20294_ = ~new_n15746_ | ~pi1142;
  assign new_n20295_ = ~new_n17262_ | ~new_n17260_ | ~new_n17261_ | ~new_n17263_;
  assign new_n20296_ = ~new_n15763_ | ~pi1135;
  assign new_n20297_ = ~new_n15762_ | ~pi1127;
  assign new_n20298_ = ~new_n15761_ | ~pi1119;
  assign new_n20299_ = ~new_n15760_ | ~pi1111;
  assign new_n20300_ = ~new_n15758_ | ~pi1103;
  assign new_n20301_ = ~new_n15757_ | ~pi1095;
  assign new_n20302_ = ~new_n15756_ | ~pi1087;
  assign new_n20303_ = ~new_n15755_ | ~pi1079;
  assign new_n20304_ = ~new_n15754_ | ~pi1199;
  assign new_n20305_ = ~new_n15753_ | ~pi1191;
  assign new_n20306_ = ~new_n15752_ | ~pi1183;
  assign new_n20307_ = ~new_n15751_ | ~pi1175;
  assign new_n20308_ = ~new_n15749_ | ~pi1167;
  assign new_n20309_ = ~new_n15748_ | ~pi1159;
  assign new_n20310_ = ~new_n15747_ | ~pi1151;
  assign new_n20311_ = ~new_n15746_ | ~pi1143;
  assign new_n20312_ = ~new_n17266_ | ~new_n17264_ | ~new_n17265_ | ~new_n17267_;
  assign new_n20313_ = ~new_n15763_ | ~pi1136;
  assign new_n20314_ = ~new_n15762_ | ~pi1128;
  assign new_n20315_ = ~new_n15761_ | ~pi1120;
  assign new_n20316_ = ~new_n15760_ | ~pi1112;
  assign new_n20317_ = ~new_n15758_ | ~pi1104;
  assign new_n20318_ = ~new_n15757_ | ~pi1096;
  assign new_n20319_ = ~new_n15756_ | ~pi1088;
  assign new_n20320_ = ~new_n15755_ | ~pi1080;
  assign new_n20321_ = ~new_n15753_ | ~pi1192;
  assign new_n20322_ = ~new_n15752_ | ~pi1184;
  assign new_n20323_ = ~new_n15751_ | ~pi1176;
  assign new_n20324_ = ~new_n15749_ | ~pi1168;
  assign new_n20325_ = ~new_n15748_ | ~pi1160;
  assign new_n20326_ = ~new_n15747_ | ~pi1152;
  assign new_n20327_ = ~new_n15746_ | ~pi1144;
  assign new_n20328_ = ~new_n15763_ | ~pi1137;
  assign new_n20329_ = ~new_n15762_ | ~pi1129;
  assign new_n20330_ = ~new_n15761_ | ~pi1121;
  assign new_n20331_ = ~new_n15760_ | ~pi1113;
  assign new_n20332_ = ~new_n15758_ | ~pi1105;
  assign new_n20333_ = ~new_n15757_ | ~pi1097;
  assign new_n20334_ = ~new_n15756_ | ~pi1089;
  assign new_n20335_ = ~new_n15755_ | ~pi1081;
  assign new_n20336_ = ~new_n15754_ | ~pi1201;
  assign new_n20337_ = ~new_n15753_ | ~pi1193;
  assign new_n20338_ = ~new_n15752_ | ~pi1185;
  assign new_n20339_ = ~new_n15751_ | ~pi1177;
  assign new_n20340_ = ~new_n15749_ | ~pi1169;
  assign new_n20341_ = ~new_n15748_ | ~pi1161;
  assign new_n20342_ = ~new_n15747_ | ~pi1153;
  assign new_n20343_ = ~new_n15746_ | ~pi1145;
  assign new_n20344_ = ~new_n17275_ | ~new_n17273_ | ~new_n17274_ | ~new_n17276_;
  assign new_n20345_ = ~new_n15763_ | ~pi1138;
  assign new_n20346_ = ~new_n15762_ | ~pi1130;
  assign new_n20347_ = ~new_n15761_ | ~pi1122;
  assign new_n20348_ = ~new_n15760_ | ~pi1114;
  assign new_n20349_ = ~new_n15758_ | ~pi1106;
  assign new_n20350_ = ~new_n15757_ | ~pi1098;
  assign new_n20351_ = ~new_n15756_ | ~pi1090;
  assign new_n20352_ = ~new_n15755_ | ~pi1082;
  assign new_n20353_ = ~new_n15754_ | ~pi1202;
  assign new_n20354_ = ~new_n15753_ | ~pi1194;
  assign new_n20355_ = ~new_n15752_ | ~pi1186;
  assign new_n20356_ = ~new_n15751_ | ~pi1178;
  assign new_n20357_ = ~new_n15749_ | ~pi1170;
  assign new_n20358_ = ~new_n15748_ | ~pi1162;
  assign new_n20359_ = ~new_n15747_ | ~pi1154;
  assign new_n20360_ = ~new_n15746_ | ~pi1146;
  assign new_n20361_ = ~new_n17279_ | ~new_n17277_ | ~new_n17278_ | ~new_n17280_;
  assign new_n20362_ = ~new_n15763_ | ~pi1139;
  assign new_n20363_ = ~new_n15762_ | ~pi1131;
  assign new_n20364_ = ~new_n15761_ | ~pi1123;
  assign new_n20365_ = ~new_n15760_ | ~pi1115;
  assign new_n20366_ = ~new_n15758_ | ~pi1107;
  assign new_n20367_ = ~new_n15757_ | ~pi1099;
  assign new_n20368_ = ~new_n15756_ | ~pi1091;
  assign new_n20369_ = ~new_n15755_ | ~pi1083;
  assign new_n20370_ = ~new_n15754_ | ~pi1203;
  assign new_n20371_ = ~new_n15753_ | ~pi1195;
  assign new_n20372_ = ~new_n15752_ | ~pi1187;
  assign new_n20373_ = ~new_n15751_ | ~pi1179;
  assign new_n20374_ = ~new_n15749_ | ~pi1171;
  assign new_n20375_ = ~new_n15748_ | ~pi1163;
  assign new_n20376_ = ~new_n15747_ | ~pi1155;
  assign new_n20377_ = ~new_n15746_ | ~pi1147;
  assign new_n20378_ = ~new_n17283_ | ~new_n17281_ | ~new_n17282_ | ~new_n17284_;
  assign new_n20379_ = ~new_n15763_ | ~pi1140;
  assign new_n20380_ = ~new_n15762_ | ~pi1132;
  assign new_n20381_ = ~new_n15761_ | ~pi1124;
  assign new_n20382_ = ~new_n15760_ | ~pi1116;
  assign new_n20383_ = ~new_n15758_ | ~pi1108;
  assign new_n20384_ = ~new_n15757_ | ~pi1100;
  assign new_n20385_ = ~new_n15756_ | ~pi1092;
  assign new_n20386_ = ~new_n15755_ | ~pi1084;
  assign new_n20387_ = ~new_n15754_ | ~pi1204;
  assign new_n20388_ = ~new_n15753_ | ~pi1196;
  assign new_n20389_ = ~new_n15752_ | ~pi1188;
  assign new_n20390_ = ~new_n15751_ | ~pi1180;
  assign new_n20391_ = ~new_n15749_ | ~pi1172;
  assign new_n20392_ = ~new_n15748_ | ~pi1164;
  assign new_n20393_ = ~new_n15747_ | ~pi1156;
  assign new_n20394_ = ~new_n15746_ | ~pi1148;
  assign new_n20395_ = ~new_n17287_ | ~new_n17285_ | ~new_n17286_ | ~new_n17288_;
  assign new_n20396_ = ~pi1212 | ~new_n16478_;
  assign new_n20397_ = ~new_n17384_ | ~new_n16636_;
  assign new_n20398_ = ~pi1213 | ~new_n16478_;
  assign new_n20399_ = ~new_n17384_ | ~new_n16416_;
  assign new_n20400_ = ~new_n17364_;
  assign new_n20401_ = ~new_n15783_ | ~pi1133;
  assign new_n20402_ = ~new_n15782_ | ~pi1125;
  assign new_n20403_ = ~new_n15781_ | ~pi1117;
  assign new_n20404_ = ~new_n15780_ | ~pi1109;
  assign new_n20405_ = ~new_n15778_ | ~pi1101;
  assign new_n20406_ = ~new_n15777_ | ~pi1093;
  assign new_n20407_ = ~new_n15776_ | ~pi1085;
  assign new_n20408_ = ~new_n15775_ | ~pi1077;
  assign new_n20409_ = ~new_n15773_ | ~pi1197;
  assign new_n20410_ = ~new_n15772_ | ~pi1189;
  assign new_n20411_ = ~new_n15771_ | ~pi1181;
  assign new_n20412_ = ~new_n15770_ | ~pi1173;
  assign new_n20413_ = ~new_n15768_ | ~pi1165;
  assign new_n20414_ = ~new_n15767_ | ~pi1157;
  assign new_n20415_ = ~new_n15766_ | ~pi1149;
  assign new_n20416_ = ~new_n15765_ | ~pi1141;
  assign new_n20417_ = ~new_n17304_ | ~new_n17302_ | ~new_n17303_ | ~new_n17305_;
  assign new_n20418_ = ~new_n15783_ | ~pi1134;
  assign new_n20419_ = ~new_n15782_ | ~pi1126;
  assign new_n20420_ = ~new_n15781_ | ~pi1118;
  assign new_n20421_ = ~new_n15780_ | ~pi1110;
  assign new_n20422_ = ~new_n15778_ | ~pi1102;
  assign new_n20423_ = ~new_n15777_ | ~pi1094;
  assign new_n20424_ = ~new_n15776_ | ~pi1086;
  assign new_n20425_ = ~new_n15775_ | ~pi1078;
  assign new_n20426_ = ~new_n15773_ | ~pi1198;
  assign new_n20427_ = ~new_n15772_ | ~pi1190;
  assign new_n20428_ = ~new_n15771_ | ~pi1182;
  assign new_n20429_ = ~new_n15770_ | ~pi1174;
  assign new_n20430_ = ~new_n15768_ | ~pi1166;
  assign new_n20431_ = ~new_n15767_ | ~pi1158;
  assign new_n20432_ = ~new_n15766_ | ~pi1150;
  assign new_n20433_ = ~new_n15765_ | ~pi1142;
  assign new_n20434_ = ~new_n17308_ | ~new_n17306_ | ~new_n17307_ | ~new_n17309_;
  assign new_n20435_ = ~new_n15783_ | ~pi1135;
  assign new_n20436_ = ~new_n15782_ | ~pi1127;
  assign new_n20437_ = ~new_n15781_ | ~pi1119;
  assign new_n20438_ = ~new_n15780_ | ~pi1111;
  assign new_n20439_ = ~new_n15778_ | ~pi1103;
  assign new_n20440_ = ~new_n15777_ | ~pi1095;
  assign new_n20441_ = ~new_n15776_ | ~pi1087;
  assign new_n20442_ = ~new_n15775_ | ~pi1079;
  assign new_n20443_ = ~new_n15773_ | ~pi1199;
  assign new_n20444_ = ~new_n15772_ | ~pi1191;
  assign new_n20445_ = ~new_n15771_ | ~pi1183;
  assign new_n20446_ = ~new_n15770_ | ~pi1175;
  assign new_n20447_ = ~new_n15768_ | ~pi1167;
  assign new_n20448_ = ~new_n15767_ | ~pi1159;
  assign new_n20449_ = ~new_n15766_ | ~pi1151;
  assign new_n20450_ = ~new_n15765_ | ~pi1143;
  assign new_n20451_ = ~new_n17312_ | ~new_n17310_ | ~new_n17311_ | ~new_n17313_;
  assign new_n20452_ = ~new_n15783_ | ~pi1136;
  assign new_n20453_ = ~new_n15782_ | ~pi1128;
  assign new_n20454_ = ~new_n15781_ | ~pi1120;
  assign new_n20455_ = ~new_n15780_ | ~pi1112;
  assign new_n20456_ = ~new_n15778_ | ~pi1104;
  assign new_n20457_ = ~new_n15777_ | ~pi1096;
  assign new_n20458_ = ~new_n15776_ | ~pi1088;
  assign new_n20459_ = ~new_n15775_ | ~pi1080;
  assign new_n20460_ = ~new_n15772_ | ~pi1192;
  assign new_n20461_ = ~new_n15771_ | ~pi1184;
  assign new_n20462_ = ~new_n15770_ | ~pi1176;
  assign new_n20463_ = ~new_n15768_ | ~pi1168;
  assign new_n20464_ = ~new_n15767_ | ~pi1160;
  assign new_n20465_ = ~new_n15766_ | ~pi1152;
  assign new_n20466_ = ~new_n15765_ | ~pi1144;
  assign new_n20467_ = ~new_n15783_ | ~pi1137;
  assign new_n20468_ = ~new_n15782_ | ~pi1129;
  assign new_n20469_ = ~new_n15781_ | ~pi1121;
  assign new_n20470_ = ~new_n15780_ | ~pi1113;
  assign new_n20471_ = ~new_n15778_ | ~pi1105;
  assign new_n20472_ = ~new_n15777_ | ~pi1097;
  assign new_n20473_ = ~new_n15776_ | ~pi1089;
  assign new_n20474_ = ~new_n15775_ | ~pi1081;
  assign new_n20475_ = ~new_n15773_ | ~pi1201;
  assign new_n20476_ = ~new_n15772_ | ~pi1193;
  assign new_n20477_ = ~new_n15771_ | ~pi1185;
  assign new_n20478_ = ~new_n15770_ | ~pi1177;
  assign new_n20479_ = ~new_n15768_ | ~pi1169;
  assign new_n20480_ = ~new_n15767_ | ~pi1161;
  assign new_n20481_ = ~new_n15766_ | ~pi1153;
  assign new_n20482_ = ~new_n15765_ | ~pi1145;
  assign new_n20483_ = ~new_n17320_ | ~new_n17318_ | ~new_n17319_ | ~new_n17321_;
  assign new_n20484_ = ~new_n15783_ | ~pi1138;
  assign new_n20485_ = ~new_n15782_ | ~pi1130;
  assign new_n20486_ = ~new_n15781_ | ~pi1122;
  assign new_n20487_ = ~new_n15780_ | ~pi1114;
  assign new_n20488_ = ~new_n15778_ | ~pi1106;
  assign new_n20489_ = ~new_n15777_ | ~pi1098;
  assign new_n20490_ = ~new_n15776_ | ~pi1090;
  assign new_n20491_ = ~new_n15775_ | ~pi1082;
  assign new_n20492_ = ~new_n15773_ | ~pi1202;
  assign new_n20493_ = ~new_n15772_ | ~pi1194;
  assign new_n20494_ = ~new_n15771_ | ~pi1186;
  assign new_n20495_ = ~new_n15770_ | ~pi1178;
  assign new_n20496_ = ~new_n15768_ | ~pi1170;
  assign new_n20497_ = ~new_n15767_ | ~pi1162;
  assign new_n20498_ = ~new_n15766_ | ~pi1154;
  assign new_n20499_ = ~new_n15765_ | ~pi1146;
  assign new_n20500_ = ~new_n17324_ | ~new_n17322_ | ~new_n17323_ | ~new_n17325_;
  assign new_n20501_ = ~new_n15783_ | ~pi1139;
  assign new_n20502_ = ~new_n15782_ | ~pi1131;
  assign new_n20503_ = ~new_n15781_ | ~pi1123;
  assign new_n20504_ = ~new_n15780_ | ~pi1115;
  assign new_n20505_ = ~new_n15778_ | ~pi1107;
  assign new_n20506_ = ~new_n15777_ | ~pi1099;
  assign new_n20507_ = ~new_n15776_ | ~pi1091;
  assign new_n20508_ = ~new_n15775_ | ~pi1083;
  assign new_n20509_ = ~new_n15773_ | ~pi1203;
  assign new_n20510_ = ~new_n15772_ | ~pi1195;
  assign new_n20511_ = ~new_n15771_ | ~pi1187;
  assign new_n20512_ = ~new_n15770_ | ~pi1179;
  assign new_n20513_ = ~new_n15768_ | ~pi1171;
  assign new_n20514_ = ~new_n15767_ | ~pi1163;
  assign new_n20515_ = ~new_n15766_ | ~pi1155;
  assign new_n20516_ = ~new_n15765_ | ~pi1147;
  assign new_n20517_ = ~new_n17328_ | ~new_n17326_ | ~new_n17327_ | ~new_n17329_;
  assign new_n20518_ = ~new_n15783_ | ~pi1140;
  assign new_n20519_ = ~new_n15782_ | ~pi1132;
  assign new_n20520_ = ~new_n15781_ | ~pi1124;
  assign new_n20521_ = ~new_n15780_ | ~pi1116;
  assign new_n20522_ = ~new_n15778_ | ~pi1108;
  assign new_n20523_ = ~new_n15777_ | ~pi1100;
  assign new_n20524_ = ~new_n15776_ | ~pi1092;
  assign new_n20525_ = ~new_n15775_ | ~pi1084;
  assign new_n20526_ = ~new_n15773_ | ~pi1204;
  assign new_n20527_ = ~new_n15772_ | ~pi1196;
  assign new_n20528_ = ~new_n15771_ | ~pi1188;
  assign new_n20529_ = ~new_n15770_ | ~pi1180;
  assign new_n20530_ = ~new_n15768_ | ~pi1172;
  assign new_n20531_ = ~new_n15767_ | ~pi1164;
  assign new_n20532_ = ~new_n15766_ | ~pi1156;
  assign new_n20533_ = ~new_n15765_ | ~pi1148;
  assign new_n20534_ = ~new_n17332_ | ~new_n17330_ | ~new_n17331_ | ~new_n17333_;
  assign new_n20535_ = ~new_n17415_ | ~new_n17412_ | ~new_n15535_;
  assign new_n20536_ = ~new_n17334_ | ~new_n20268_;
  assign new_n20537_ = ~new_n16577_ | ~new_n16591_;
  assign new_n20538_ = ~new_n17415_ | ~new_n20537_;
  assign new_n20539_ = ~new_n17371_ | ~new_n15633_;
  assign new_n20540_ = ~new_n20536_ | ~new_n16452_;
  assign new_n20541_ = ~new_n17389_ | ~new_n20269_;
  assign new_n20542_ = ~new_n17341_ | ~new_n17389_;
  assign new_n20543_ = ~new_n15632_ | ~new_n17391_;
  assign new_n20544_ = ~new_n16601_ | ~new_n20542_ | ~new_n20543_ | ~new_n17376_ | ~new_n16615_;
  assign new_n20545_ = ~new_n33497_ | ~new_n20544_;
  assign new_n20546_ = ~new_n33558_ | ~new_n15535_;
  assign new_n20547_ = ~new_n33510_ | ~new_n20544_;
  assign new_n20548_ = ~new_n33571_ | ~new_n15535_;
  assign new_n20549_ = ~new_n33511_ | ~new_n20544_;
  assign new_n20550_ = ~new_n33572_ | ~new_n15535_;
  assign new_n20551_ = ~new_n33512_ | ~new_n20544_;
  assign new_n20552_ = ~new_n33573_ | ~new_n15535_;
  assign new_n20553_ = ~new_n33513_ | ~new_n20544_;
  assign new_n20554_ = ~new_n33574_ | ~new_n15535_;
  assign new_n20555_ = ~new_n33498_ | ~new_n20544_;
  assign new_n20556_ = ~new_n33559_ | ~new_n15535_;
  assign new_n20557_ = ~new_n33510_ | ~new_n17373_;
  assign new_n20558_ = ~pi1205 | ~new_n16475_;
  assign new_n20559_ = ~new_n33511_ | ~new_n17373_;
  assign new_n20560_ = ~pi1206 | ~new_n16475_;
  assign new_n20561_ = ~pi1076 | ~new_n17354_;
  assign new_n20562_ = ~new_n16601_ | ~new_n20561_;
  assign new_n20563_ = ~new_n33512_ | ~new_n17373_;
  assign new_n20564_ = ~pi1207 | ~new_n16475_;
  assign new_n20565_ = ~new_n15631_ | ~new_n16452_;
  assign new_n20566_ = ~new_n33513_ | ~new_n17373_;
  assign new_n20567_ = ~pi1208 | ~new_n16475_;
  assign new_n20568_ = ~new_n15632_ | ~new_n16465_;
  assign new_n20569_ = ~new_n33498_ | ~new_n17373_;
  assign new_n20570_ = ~pi1209 | ~new_n16475_;
  assign new_n20571_ = ~new_n16574_ | ~new_n16471_;
  assign new_n20572_ = ~new_n16465_ | ~new_n16630_;
  assign new_n20573_ = ~pi1224 | ~new_n20572_;
  assign new_n20574_ = ~pi1383 | ~new_n20571_;
  assign new_n20575_ = ~pi1223 | ~new_n20572_;
  assign new_n20576_ = ~pi1382 | ~new_n20571_;
  assign new_n20577_ = ~pi1222 | ~new_n20572_;
  assign new_n20578_ = ~pi1381 | ~new_n20571_;
  assign new_n20579_ = ~pi1221 | ~new_n20572_;
  assign new_n20580_ = ~pi1380 | ~new_n20571_;
  assign new_n20581_ = ~pi1220 | ~new_n20572_;
  assign new_n20582_ = ~pi1379 | ~new_n20571_;
  assign new_n20583_ = ~pi1219 | ~new_n20572_;
  assign new_n20584_ = ~pi1378 | ~new_n20571_;
  assign new_n20585_ = ~pi1246 | ~new_n20572_;
  assign new_n20586_ = ~pi1405 | ~new_n20571_;
  assign new_n20587_ = ~pi1245 | ~new_n20572_;
  assign new_n20588_ = ~pi1404 | ~new_n20571_;
  assign new_n20589_ = ~pi1218 | ~new_n20572_;
  assign new_n20590_ = ~pi1377 | ~new_n20571_;
  assign new_n20591_ = ~pi1244 | ~new_n20572_;
  assign new_n20592_ = ~pi1403 | ~new_n20571_;
  assign new_n20593_ = ~pi1243 | ~new_n20572_;
  assign new_n20594_ = ~pi1402 | ~new_n20571_;
  assign new_n20595_ = ~pi1242 | ~new_n20572_;
  assign new_n20596_ = ~pi1401 | ~new_n20571_;
  assign new_n20597_ = ~pi1241 | ~new_n20572_;
  assign new_n20598_ = ~pi1400 | ~new_n20571_;
  assign new_n20599_ = ~pi1240 | ~new_n20572_;
  assign new_n20600_ = ~pi1399 | ~new_n20571_;
  assign new_n20601_ = ~pi1239 | ~new_n20572_;
  assign new_n20602_ = ~pi1398 | ~new_n20571_;
  assign new_n20603_ = ~pi1238 | ~new_n20572_;
  assign new_n20604_ = ~pi1397 | ~new_n20571_;
  assign new_n20605_ = ~pi1237 | ~new_n20572_;
  assign new_n20606_ = ~pi1396 | ~new_n20571_;
  assign new_n20607_ = ~pi1236 | ~new_n20572_;
  assign new_n20608_ = ~pi1395 | ~new_n20571_;
  assign new_n20609_ = ~pi1235 | ~new_n20572_;
  assign new_n20610_ = ~pi1394 | ~new_n20571_;
  assign new_n20611_ = ~pi1217 | ~new_n20572_;
  assign new_n20612_ = ~pi1376 | ~new_n20571_;
  assign new_n20613_ = ~pi1234 | ~new_n20572_;
  assign new_n20614_ = ~pi1393 | ~new_n20571_;
  assign new_n20615_ = ~pi1233 | ~new_n20572_;
  assign new_n20616_ = ~pi1392 | ~new_n20571_;
  assign new_n20617_ = ~pi1232 | ~new_n20572_;
  assign new_n20618_ = ~pi1391 | ~new_n20571_;
  assign new_n20619_ = ~pi1231 | ~new_n20572_;
  assign new_n20620_ = ~pi1390 | ~new_n20571_;
  assign new_n20621_ = ~pi1230 | ~new_n20572_;
  assign new_n20622_ = ~pi1389 | ~new_n20571_;
  assign new_n20623_ = ~pi1229 | ~new_n20572_;
  assign new_n20624_ = ~pi1388 | ~new_n20571_;
  assign new_n20625_ = ~pi1228 | ~new_n20572_;
  assign new_n20626_ = ~pi1387 | ~new_n20571_;
  assign new_n20627_ = ~pi1227 | ~new_n20572_;
  assign new_n20628_ = ~pi1386 | ~new_n20571_;
  assign new_n20629_ = ~pi1226 | ~new_n20572_;
  assign new_n20630_ = ~pi1385 | ~new_n20571_;
  assign new_n20631_ = ~pi1225 | ~new_n20572_;
  assign new_n20632_ = ~pi1384 | ~new_n20571_;
  assign new_n20633_ = ~pi1216 | ~new_n20572_;
  assign new_n20634_ = ~pi1375 | ~new_n20571_;
  assign new_n20635_ = ~pi1215 | ~new_n20572_;
  assign new_n20636_ = ~pi1374 | ~new_n20571_;
  assign new_n20637_ = ~new_n17658_ | ~new_n17677_;
  assign new_n20638_ = ~new_n15611_ | ~pi1205;
  assign new_n20639_ = ~new_n16670_ | ~new_n16443_;
  assign new_n20640_ = ~new_n15611_ | ~pi1206;
  assign new_n20641_ = ~new_n16671_ | ~new_n16443_;
  assign new_n20642_ = ~new_n16651_ | ~pi1443 | ~new_n15627_;
  assign new_n20643_ = ~new_n15611_ | ~pi1207;
  assign new_n20644_ = ~new_n16672_ | ~new_n16443_;
  assign new_n20645_ = ~new_n20893_ | ~new_n15627_ | ~pi1443;
  assign new_n20646_ = ~new_n15611_ | ~pi1208;
  assign new_n20647_ = ~new_n16673_ | ~new_n16443_;
  assign new_n20648_ = ~new_n15611_ | ~pi1209;
  assign new_n20649_ = ~pi1040 | ~new_n17366_;
  assign new_n20650_ = new_n2972_ | pi1074;
  assign new_n20651_ = ~new_n17291_ | ~new_n20399_;
  assign new_n20652_ = ~new_n20265_ | ~new_n16603_;
  assign new_n20653_ = ~new_n17392_ | ~pi1076;
  assign new_n20654_ = ~new_n17393_ | ~pi1076;
  assign new_n20655_ = ~new_n17394_ | ~pi1076;
  assign new_n20656_ = ~new_n17417_ | ~pi1076;
  assign new_n20657_ = ~new_n17445_ | ~pi1076;
  assign new_n20658_ = ~pi1076 | ~new_n20813_;
  assign new_n20659_ = ~new_n15789_ | ~new_n16447_;
  assign new_n20660_ = ~new_n20274_ | ~new_n17301_ | ~new_n17299_ | ~new_n17298_;
  assign new_n20661_ = ~pi1076 | ~new_n20813_;
  assign new_n20662_ = ~new_n15560_ | ~new_n16610_;
  assign new_n20663_ = ~new_n15550_ | ~new_n19548_;
  assign new_n20664_ = ~new_n17069_ | ~new_n15550_;
  assign new_n20665_ = ~new_n20663_ | ~new_n20662_ | ~new_n17410_;
  assign new_n20666_ = ~new_n20664_ | ~new_n17411_;
  assign new_n20667_ = ~new_n17375_ | ~new_n18672_ | ~new_n17352_;
  assign new_n20668_ = ~new_n20272_ | ~new_n17375_;
  assign new_n20669_ = ~new_n17375_ | ~new_n16573_;
  assign new_n20670_ = ~new_n17417_ | ~pi1076;
  assign new_n20671_ = ~new_n17253_ | ~new_n20966_ | ~new_n20965_;
  assign new_n20672_ = ~new_n17289_ | ~new_n20397_;
  assign new_n20673_ = ~new_n17290_ | ~new_n20275_;
  assign new_n20674_ = ~new_n16460_;
  assign new_n20675_ = ~new_n16457_;
  assign new_n20676_ = ~new_n17252_ | ~new_n17249_ | ~new_n17250_ | ~new_n17251_ | ~new_n15788_;
  assign new_n20677_ = ~new_n16915_ | ~new_n20674_;
  assign new_n20678_ = ~new_n16916_ | ~new_n18650_;
  assign new_n20679_ = ~new_n15606_ | ~new_n20674_;
  assign new_n20680_ = ~new_n15606_ | ~new_n20674_;
  assign new_n20681_ = ~new_n20680_ | ~new_n19542_ | ~new_n19541_;
  assign new_n20682_ = ~new_n20674_ | ~new_n33065_;
  assign new_n20683_ = ~new_n33065_ | ~new_n20674_ | ~new_n17382_;
  assign new_n20684_ = ~new_n20683_ | ~new_n19330_;
  assign new_n20685_ = ~new_n20674_ | ~new_n20266_;
  assign new_n20686_ = ~new_n20674_ | ~new_n20652_;
  assign new_n20687_ = ~new_n17295_ | ~new_n17297_ | ~new_n17296_;
  assign new_n20688_ = ~new_n16940_ | ~new_n20674_;
  assign new_n20689_ = ~new_n16941_ | ~new_n16942_ | ~new_n18746_;
  assign new_n20690_ = ~new_n16927_ | ~new_n15700_;
  assign new_n20691_ = ~new_n20674_ | ~new_n19143_;
  assign new_n20692_ = ~new_n20674_ | ~new_n19146_;
  assign new_n20693_ = ~new_n20674_ | ~new_n19149_;
  assign new_n20694_ = ~new_n20674_ | ~new_n19152_;
  assign new_n20695_ = ~new_n20674_ | ~new_n19155_;
  assign new_n20696_ = ~new_n20674_ | ~new_n19158_;
  assign new_n20697_ = ~new_n20674_ | ~new_n19161_;
  assign new_n20698_ = ~new_n20674_ | ~new_n19164_;
  assign new_n20699_ = ~new_n20674_ | ~new_n19167_;
  assign new_n20700_ = ~new_n20674_ | ~new_n19170_;
  assign new_n20701_ = ~new_n20674_ | ~new_n19173_;
  assign new_n20702_ = ~new_n20674_ | ~new_n19176_;
  assign new_n20703_ = ~new_n20674_ | ~new_n19179_;
  assign new_n20704_ = ~new_n20674_ | ~new_n19182_;
  assign new_n20705_ = ~new_n20674_ | ~new_n19185_;
  assign new_n20706_ = ~new_n20674_ | ~new_n19188_;
  assign new_n20707_ = ~new_n20674_ | ~new_n19191_;
  assign new_n20708_ = ~new_n20674_ | ~new_n19194_;
  assign new_n20709_ = ~new_n20674_ | ~new_n19197_;
  assign new_n20710_ = ~new_n20674_ | ~new_n19200_;
  assign new_n20711_ = ~new_n20674_ | ~new_n19203_;
  assign new_n20712_ = ~new_n20674_ | ~new_n19206_;
  assign new_n20713_ = ~new_n20674_ | ~new_n19209_;
  assign new_n20714_ = ~new_n20674_ | ~new_n19212_;
  assign new_n20715_ = ~new_n20674_ | ~new_n19215_;
  assign new_n20716_ = ~new_n20674_ | ~new_n19218_;
  assign new_n20717_ = ~new_n20674_ | ~new_n19221_;
  assign new_n20718_ = ~new_n20674_ | ~new_n19224_;
  assign new_n20719_ = ~new_n20674_ | ~new_n19227_;
  assign new_n20720_ = ~new_n20674_ | ~new_n19230_;
  assign new_n20721_ = ~new_n20674_ | ~new_n19233_;
  assign new_n20722_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20723_ = ~pi1309 | ~new_n20722_;
  assign new_n20724_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20725_ = ~pi1308 | ~new_n20724_;
  assign new_n20726_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20727_ = ~pi1307 | ~new_n20726_;
  assign new_n20728_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20729_ = ~pi1306 | ~new_n20728_;
  assign new_n20730_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20731_ = ~pi1305 | ~new_n20730_;
  assign new_n20732_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20733_ = ~pi1304 | ~new_n20732_;
  assign new_n20734_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20735_ = ~pi1303 | ~new_n20734_;
  assign new_n20736_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20737_ = ~pi1302 | ~new_n20736_;
  assign new_n20738_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20739_ = ~pi1301 | ~new_n20738_;
  assign new_n20740_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20741_ = ~pi1300 | ~new_n20740_;
  assign new_n20742_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20743_ = ~pi1299 | ~new_n20742_;
  assign new_n20744_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20745_ = ~pi1298 | ~new_n20744_;
  assign new_n20746_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20747_ = ~pi1297 | ~new_n20746_;
  assign new_n20748_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20749_ = ~pi1296 | ~new_n20748_;
  assign new_n20750_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20751_ = ~pi1295 | ~new_n20750_;
  assign new_n20752_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20753_ = ~pi1294 | ~new_n20752_;
  assign new_n20754_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20755_ = ~pi1293 | ~new_n20754_;
  assign new_n20756_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20757_ = ~pi1292 | ~new_n20756_;
  assign new_n20758_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20759_ = ~pi1291 | ~new_n20758_;
  assign new_n20760_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20761_ = ~pi1290 | ~new_n20760_;
  assign new_n20762_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20763_ = ~pi1289 | ~new_n20762_;
  assign new_n20764_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20765_ = ~pi1288 | ~new_n20764_;
  assign new_n20766_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20767_ = ~pi1287 | ~new_n20766_;
  assign new_n20768_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20769_ = ~pi1286 | ~new_n20768_;
  assign new_n20770_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20771_ = ~pi1285 | ~new_n20770_;
  assign new_n20772_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20773_ = ~pi1284 | ~new_n20772_;
  assign new_n20774_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20775_ = ~pi1283 | ~new_n20774_;
  assign new_n20776_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20777_ = ~pi1282 | ~new_n20776_;
  assign new_n20778_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20779_ = ~pi1281 | ~new_n20778_;
  assign new_n20780_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20781_ = ~pi1280 | ~new_n20780_;
  assign new_n20782_ = ~new_n15538_ | ~new_n20674_;
  assign new_n20783_ = ~pi1279 | ~new_n20782_;
  assign new_n20784_ = ~new_n17440_ | ~new_n20674_ | ~new_n16749_;
  assign new_n20785_ = ~new_n16762_ | ~new_n20865_ | ~new_n20864_;
  assign new_n20786_ = ~new_n17048_ | ~new_n20674_;
  assign new_n20787_ = ~new_n20786_ | ~new_n16609_;
  assign new_n20788_ = ~new_n17389_ | ~new_n20674_;
  assign new_n20789_ = ~new_n20788_ | ~new_n16628_;
  assign new_n20790_ = ~new_n16460_ | ~new_n16581_;
  assign new_n20791_ = ~new_n16935_ | ~new_n20674_;
  assign new_n20792_ = ~new_n16936_ | ~new_n20791_;
  assign new_n20793_ = ~pi1200 | ~new_n18597_;
  assign new_n20794_ = ~new_n15704_ | ~pi1200;
  assign new_n20795_ = ~new_n15727_ | ~pi1200;
  assign new_n20796_ = ~new_n17232_ | ~new_n17230_ | ~new_n17231_ | ~new_n17233_;
  assign new_n20797_ = ~new_n17373_ | ~pi1200;
  assign new_n20798_ = ~new_n15754_ | ~pi1200;
  assign new_n20799_ = ~new_n17270_ | ~new_n17268_ | ~new_n17269_ | ~new_n17272_;
  assign new_n20800_ = ~new_n15773_ | ~pi1200;
  assign new_n20801_ = ~new_n17316_ | ~new_n17314_ | ~new_n17315_ | ~new_n17317_;
  assign new_n20802_ = ~new_n16440_;
  assign new_n20803_ = ~new_n20802_ | ~new_n16442_;
  assign new_n20804_ = ~new_n17539_ | ~new_n17542_ | ~pi1039;
  assign new_n20805_ = ~pi1038 | ~new_n20649_;
  assign new_n20806_ = ~pi1039 | ~new_n17539_;
  assign new_n20807_ = ~new_n17683_ | ~new_n17691_;
  assign new_n20808_ = ~new_n18668_ | ~new_n17352_;
  assign new_n20809_ = ~new_n16464_ | ~new_n16470_;
  assign new_n20810_ = ~new_n16573_;
  assign new_n20811_ = ~new_n17389_ | ~new_n20671_;
  assign new_n20812_ = ~new_n18668_ | ~new_n17352_;
  assign new_n20813_ = ~new_n20812_ | ~new_n20811_;
  assign new_n20814_ = ~pi1004 | ~new_n16430_;
  assign new_n20815_ = ~pi1438 | ~new_n17402_;
  assign new_n20816_ = ~pi1005 | ~new_n16430_;
  assign new_n20817_ = ~pi1439 | ~new_n17402_;
  assign new_n20818_ = ~pi1006 | ~new_n16430_;
  assign new_n20819_ = ~pi1440 | ~new_n17402_;
  assign new_n20820_ = ~pi1007 | ~new_n16430_;
  assign new_n20821_ = ~pi1441 | ~new_n17402_;
  assign new_n20822_ = ~new_n16432_ | ~pi1040 | ~pi1446;
  assign new_n20823_ = ~pi1038 | ~new_n16440_;
  assign new_n20824_ = ~new_n20823_ | ~new_n20822_;
  assign new_n20825_ = ~pi1039 | ~new_n20805_ | ~new_n17542_;
  assign new_n20826_ = ~new_n20824_ | ~new_n16429_;
  assign new_n20827_ = ~pi1038 | ~pi1040 | ~new_n16441_;
  assign new_n20828_ = ~new_n17552_ | ~new_n16432_;
  assign new_n20829_ = pi1040 | pi1039;
  assign new_n20830_ = ~pi1040 | ~new_n17439_;
  assign new_n20831_ = ~new_n16643_;
  assign new_n20832_ = ~new_n20831_ | ~pi1041;
  assign new_n20833_ = ~new_n16644_ | ~new_n16643_;
  assign new_n20834_ = ~new_n16643_ | ~new_n17557_;
  assign new_n20835_ = ~new_n20831_ | ~pi1042;
  assign new_n20836_ = ~new_n16446_ | ~new_n16722_ | ~new_n16721_;
  assign new_n20837_ = ~pi1144 | ~pi1208 | ~new_n16451_ | ~pi1207 | ~pi1209;
  assign new_n20838_ = ~pi1160 | ~new_n16446_ | ~new_n16451_ | ~pi1207 | ~pi1209;
  assign new_n20839_ = ~pi1184 | ~pi1208 | ~new_n16447_ | ~new_n16445_ | ~new_n16451_;
  assign new_n20840_ = ~new_n16451_ | ~new_n16724_ | ~new_n16723_;
  assign new_n20841_ = ~pi1206 | ~new_n16726_ | ~new_n16725_;
  assign new_n20842_ = ~new_n16446_ | ~new_n16728_ | ~new_n16727_;
  assign new_n20843_ = ~pi1208 | ~new_n16730_ | ~new_n16729_;
  assign new_n20844_ = ~new_n16447_ | ~new_n16732_ | ~new_n16731_;
  assign new_n20845_ = ~pi1080 | ~pi1209 | ~pi1207 | ~pi1208 | ~pi1206;
  assign new_n20846_ = ~pi1200 | ~new_n16451_ | ~new_n16447_ | ~new_n16446_ | ~new_n16445_;
  assign new_n20847_ = ~pi1136 | ~pi1206 | ~new_n16447_ | ~new_n16446_ | ~new_n16445_;
  assign new_n20848_ = ~pi1120 | ~new_n16447_ | ~new_n16445_ | ~pi1208 | ~pi1206;
  assign new_n20849_ = ~pi1209 | ~new_n16734_ | ~new_n16733_;
  assign new_n20850_ = ~pi1176 | ~new_n16451_ | ~new_n16445_ | ~pi1208 | ~pi1209;
  assign new_n20851_ = ~pi1112 | ~pi1206 | ~new_n16445_ | ~pi1208 | ~pi1209;
  assign new_n20852_ = ~pi1175 | ~new_n16451_ | ~new_n16445_ | ~pi1208 | ~pi1209;
  assign new_n20853_ = ~pi1206 | ~new_n16710_ | ~new_n16709_;
  assign new_n20854_ = ~pi1126 | ~new_n16446_ | ~new_n16445_ | ~pi1209 | ~pi1206;
  assign new_n20855_ = ~pi1208 | ~new_n16716_ | ~new_n16715_;
  assign new_n20856_ = ~pi1118 | ~new_n16447_ | ~new_n16445_ | ~pi1208 | ~pi1206;
  assign new_n20857_ = ~pi1110 | ~pi1209 | ~new_n16445_ | ~pi1208 | ~pi1206;
  assign new_n20858_ = ~pi1198 | ~new_n16451_ | ~new_n16447_ | ~new_n16446_ | ~new_n16445_;
  assign new_n20859_ = ~pi1134 | ~pi1206 | ~new_n16447_ | ~new_n16446_ | ~new_n16445_;
  assign new_n20860_ = ~new_n17675_ | ~new_n16618_;
  assign new_n20861_ = ~new_n20682_ | ~new_n16465_;
  assign new_n20862_ = ~new_n17397_ | ~new_n33065_;
  assign new_n20863_ = ~new_n17687_ | ~new_n16454_;
  assign new_n20864_ = ~pi1076 | ~new_n17693_;
  assign new_n20865_ = ~new_n17694_ | ~new_n16475_;
  assign new_n20866_ = ~pi1073 | ~new_n16476_;
  assign new_n20867_ = ~new_n15609_ | ~new_n17695_;
  assign new_n20868_ = pi1445 | pi1076;
  assign new_n20869_ = ~pi1076 | ~new_n20650_;
  assign new_n20870_ = ~pi1076 | ~new_n17703_;
  assign new_n20871_ = ~new_n16475_ | ~new_n20785_ | ~new_n17702_;
  assign new_n20872_ = ~new_n31276_ | ~new_n16494_;
  assign new_n20873_ = ~new_n17709_ | ~new_n16492_;
  assign new_n20874_ = ~new_n16635_;
  assign new_n20875_ = ~pi1212 | ~new_n16486_;
  assign new_n20876_ = ~new_n17714_ | ~new_n16485_;
  assign new_n20877_ = ~new_n16636_;
  assign new_n20878_ = ~new_n17397_ | ~new_n16454_;
  assign new_n20879_ = ~new_n33065_ | ~new_n20678_;
  assign new_n20880_ = ~new_n17613_ | ~new_n18647_;
  assign new_n20881_ = ~new_n18648_ | ~new_n17352_;
  assign new_n20882_ = ~new_n16648_ | ~new_n17353_;
  assign new_n20883_ = ~new_n18657_ | ~pi1205;
  assign new_n20884_ = ~new_n17641_ | ~new_n16459_;
  assign new_n20885_ = ~new_n17596_ | ~new_n16458_;
  assign new_n20886_ = ~new_n16452_ | ~new_n16596_;
  assign new_n20887_ = ~new_n17658_ | ~new_n18674_;
  assign new_n20888_ = ~new_n20887_ | ~new_n20886_;
  assign new_n20889_ = ~new_n18657_ | ~pi1206;
  assign new_n20890_ = ~new_n18690_ | ~new_n17353_;
  assign new_n20891_ = ~pi1216 | ~new_n17355_;
  assign new_n20892_ = ~new_n33290_ | ~pi1246;
  assign new_n20893_ = ~new_n16651_;
  assign new_n20894_ = ~pi1215 | ~new_n17355_;
  assign new_n20895_ = ~pi1215 | ~pi1246;
  assign new_n20896_ = ~new_n16652_;
  assign new_n20897_ = ~new_n18692_ | ~new_n18682_;
  assign new_n20898_ = ~new_n17399_ | ~new_n16582_;
  assign new_n20899_ = ~pi1208 | ~new_n16445_;
  assign new_n20900_ = ~pi1207 | ~new_n16446_;
  assign new_n20901_ = ~new_n16637_;
  assign new_n20902_ = ~new_n18657_ | ~pi1207;
  assign new_n20903_ = ~new_n18699_ | ~new_n17353_;
  assign new_n20904_ = ~new_n18657_ | ~pi1208;
  assign new_n20905_ = ~new_n18710_ | ~new_n17353_;
  assign new_n20906_ = ~new_n17395_ | ~pi1209;
  assign new_n20907_ = ~new_n18702_ | ~new_n16447_;
  assign new_n20908_ = ~new_n18657_ | ~pi1209;
  assign new_n20909_ = ~new_n18716_ | ~new_n17353_;
  assign new_n20910_ = ~new_n18718_ | ~pi1211;
  assign new_n20911_ = ~new_n18726_ | ~new_n16585_;
  assign new_n20912_ = ~new_n20874_ | ~new_n17708_;
  assign new_n20913_ = ~new_n16635_ | ~new_n16495_;
  assign new_n20914_ = ~new_n20913_ | ~new_n20912_;
  assign new_n20915_ = ~new_n18718_ | ~pi1212;
  assign new_n20916_ = ~new_n18730_ | ~new_n16585_;
  assign new_n20917_ = ~new_n18718_ | ~pi1213;
  assign new_n20918_ = ~new_n18735_ | ~new_n16585_;
  assign new_n20919_ = ~new_n18718_ | ~pi1214;
  assign new_n20920_ = ~new_n18738_ | ~new_n16585_;
  assign new_n20921_ = ~new_n17658_ | ~new_n16569_;
  assign new_n20922_ = ~new_n16452_ | ~new_n16462_;
  assign new_n20923_ = ~new_n20921_ | ~new_n17352_ | ~new_n16438_ | ~new_n20922_;
  assign new_n20924_ = ~new_n17613_ | ~new_n33065_ | ~new_n20792_;
  assign new_n20925_ = ~pi1373 | ~new_n16605_;
  assign new_n20926_ = ~new_n16660_ | ~new_n17404_;
  assign new_n20927_ = ~pi1438 | ~new_n16614_;
  assign new_n20928_ = ~new_n16661_ | ~new_n17401_;
  assign new_n20929_ = pi1041 | pi1042;
  assign new_n20930_ = ~pi1041 | ~new_n16594_;
  assign new_n20931_ = ~new_n20930_ | ~new_n20929_;
  assign new_n20932_ = ~new_n20931_ | ~new_n16434_;
  assign new_n20933_ = ~pi1406 | ~pi1407;
  assign new_n20934_ = ~new_n20933_ | ~new_n20932_;
  assign new_n20935_ = ~pi1439 | ~new_n16614_;
  assign new_n20936_ = ~new_n20934_ | ~new_n17401_;
  assign new_n20937_ = ~pi1440 | ~new_n16614_;
  assign new_n20938_ = ~new_n17401_ | ~pi1407;
  assign new_n20939_ = ~pi1441 | ~new_n16614_;
  assign new_n20940_ = ~new_n17401_ | ~new_n19780_;
  assign new_n20941_ = ~new_n17402_ | ~new_n16617_;
  assign new_n20942_ = ~pi1442 | ~new_n16430_;
  assign new_n20943_ = ~pi1444 | ~new_n17358_;
  assign new_n20944_ = ~new_n17418_ | ~new_n19781_;
  assign new_n20945_ = ~new_n20831_ | ~pi1445;
  assign new_n20946_ = ~pi0035 | ~new_n16643_;
  assign new_n20947_ = ~new_n19784_ | ~pi1446;
  assign new_n20948_ = ~new_n19790_ | ~new_n17361_;
  assign new_n20949_ = ~new_n17402_ | ~new_n16616_;
  assign new_n20950_ = ~pi1447 | ~new_n16430_;
  assign new_n20951_ = ~pi1448 | ~new_n16430_;
  assign new_n20952_ = ~pi1452 | ~new_n17402_;
  assign new_n20953_ = ~new_n19795_ | ~pi1451;
  assign new_n20954_ = ~new_n19796_ | ~new_n17362_;
  assign new_n20955_ = ~new_n16669_ | ~new_n17363_;
  assign new_n20956_ = ~new_n18654_ | ~pi1205;
  assign new_n20957_ = ~new_n18654_ | ~pi1206;
  assign new_n20958_ = ~new_n18687_ | ~new_n17363_;
  assign new_n20959_ = ~new_n18654_ | ~pi1207;
  assign new_n20960_ = ~new_n18695_ | ~new_n17363_;
  assign new_n20961_ = ~new_n18654_ | ~pi1208;
  assign new_n20962_ = ~new_n18706_ | ~new_n17363_;
  assign new_n20963_ = ~new_n18654_ | ~pi1209;
  assign new_n20964_ = ~new_n18712_ | ~new_n17363_;
  assign new_n20965_ = ~new_n15786_ | ~new_n16458_;
  assign new_n20966_ = ~new_n17641_ | ~new_n20676_;
  assign new_n20967_ = ~new_n17384_ | ~new_n16482_;
  assign new_n20968_ = ~pi1214 | ~new_n16478_;
  assign new_n20969_ = ~pi1206 | ~new_n17364_;
  assign new_n20970_ = ~new_n20400_ | ~new_n16451_;
  assign new_n20971_ = ~new_n16638_;
  assign new_n20972_ = ~new_n16457_ | ~new_n16465_;
  assign new_n20973_ = ~new_n20888_ | ~new_n17675_;
  assign new_n20974_ = ~new_n16674_ | ~new_n16443_;
  assign new_n20975_ = ~pi1075 | ~pi1443 | ~new_n20896_;
  assign new_n20976_ = ~new_n33694_;
  assign new_n20977_ = ~new_n33692_;
  assign new_n20978_ = ~new_n33690_;
  assign new_n20979_ = ~new_n33688_;
  assign new_n20980_ = ~new_n33686_;
  assign new_n20981_ = ~new_n33684_;
  assign new_n20982_ = ~new_n33682_;
  assign new_n20983_ = ~new_n33680_;
  assign new_n20984_ = ~new_n33678_;
  assign new_n20985_ = ~new_n33676_;
  assign new_n20986_ = ~new_n33674_;
  assign new_n20987_ = ~new_n33672_;
  assign new_n20988_ = ~new_n33670_;
  assign new_n20989_ = ~new_n33669_;
  assign new_n20990_ = ~new_n33666_;
  assign new_n20991_ = ~new_n33664_;
  assign new_n20992_ = ~new_n20995_;
  assign new_n20993_ = ~pi1216 | ~pi1215;
  assign new_n20994_ = new_n9738_ & new_n15476_;
  assign new_n20995_ = ~new_n33718_ | ~new_n20993_;
  assign new_n20996_ = ~new_n15523_ | ~pi1245;
  assign new_n20997_ = ~pi1246;
  assign new_n20998_ = ~new_n9379_ | ~new_n9380_;
  assign new_n20999_ = ~new_n9381_ | ~new_n9382_;
  assign new_n21000_ = ~new_n9383_ | ~new_n9384_;
  assign new_n21001_ = ~new_n9385_ | ~new_n9386_;
  assign new_n21002_ = ~new_n9387_ | ~new_n9388_;
  assign new_n21003_ = ~pi0442 | ~new_n21004_;
  assign new_n21004_ = ~pi0443;
  assign new_n21005_ = ~pi1340 | ~new_n21006_;
  assign new_n21006_ = ~pi1341;
  assign new_n21007_ = ~pi0559;
  assign new_n21008_ = pi0559 & new_n21017_;
  assign new_n21009_ = pi0579 | pi0571 | pi0566 | pi0581;
  assign new_n21010_ = ~pi0578 & ~new_n21009_ & ~pi0569 & ~pi0564 & ~pi0563;
  assign new_n21011_ = pi0588 | pi0572 | pi0580 | pi0570;
  assign new_n21012_ = ~pi0565 & ~new_n21011_ & ~pi0577 & ~pi0587;
  assign new_n21013_ = pi0567 | pi0562 | pi0582 | pi0560;
  assign new_n21014_ = ~pi0576 & ~new_n21013_ & ~pi0584 & ~pi0574;
  assign new_n21015_ = pi0568 | pi0575 | pi0561 | pi0585;
  assign new_n21016_ = ~pi0586 & ~new_n21015_ & ~pi0573 & ~pi0583;
  assign new_n21017_ = ~new_n21014_ | ~new_n21010_ | ~new_n21012_ | ~new_n21016_;
  assign new_n21018_ = pi1008 & new_n21027_;
  assign new_n21019_ = pi1028 | pi1020 | pi1015 | pi1030;
  assign new_n21020_ = ~pi1027 & ~new_n21019_ & ~pi1018 & ~pi1013 & ~pi1012;
  assign new_n21021_ = pi1037 | pi1021 | pi1029 | pi1019;
  assign new_n21022_ = ~pi1014 & ~new_n21021_ & ~pi1026 & ~pi1036;
  assign new_n21023_ = pi1016 | pi1011 | pi1031 | pi1009;
  assign new_n21024_ = ~pi1025 & ~new_n21023_ & ~pi1033 & ~pi1023;
  assign new_n21025_ = pi1017 | pi1024 | pi1010 | pi1034;
  assign new_n21026_ = ~pi1035 & ~new_n21025_ & ~pi1022 & ~pi1032;
  assign new_n21027_ = ~new_n21024_ | ~new_n21020_ | ~new_n21022_ | ~new_n21026_;
  assign new_n21028_ = ~pi0891 | ~new_n21029_;
  assign new_n21029_ = ~pi0892;
  assign new_n21030_ = ~pi0317;
  assign new_n21031_ = ~pi0319;
  assign new_n21032_ = ~pi0318;
  assign new_n21033_ = ~pi0321;
  assign new_n21034_ = ~pi0320;
  assign new_n21035_ = ~pi0318 | ~pi0319 | ~pi0317;
  assign new_n21036_ = ~pi0323;
  assign new_n21037_ = ~pi0322;
  assign new_n21038_ = ~new_n21107_ | ~new_n21136_;
  assign new_n21039_ = ~pi0325;
  assign new_n21040_ = ~pi0324;
  assign new_n21041_ = ~new_n21108_ | ~new_n21137_;
  assign new_n21042_ = ~new_n21109_ | ~new_n21143_;
  assign new_n21043_ = ~pi0326;
  assign new_n21044_ = ~pi0327;
  assign new_n21045_ = ~pi0329;
  assign new_n21046_ = ~pi0328;
  assign new_n21047_ = ~new_n21110_ | ~new_n21145_;
  assign new_n21048_ = ~pi0331;
  assign new_n21049_ = ~pi0330;
  assign new_n21050_ = ~new_n21111_ | ~new_n21138_;
  assign new_n21051_ = ~pi0332;
  assign new_n21052_ = ~new_n21112_ | ~new_n21144_;
  assign new_n21053_ = ~pi0333;
  assign new_n21054_ = ~pi0335;
  assign new_n21055_ = ~pi0334;
  assign new_n21056_ = ~new_n21113_ | ~new_n21149_;
  assign new_n21057_ = ~pi0337;
  assign new_n21058_ = ~pi0336;
  assign new_n21059_ = ~new_n21114_ | ~new_n21142_;
  assign new_n21060_ = ~pi0338;
  assign new_n21061_ = ~new_n21115_ | ~new_n21139_;
  assign new_n21062_ = ~pi0339;
  assign new_n21063_ = ~pi0341;
  assign new_n21064_ = ~pi0340;
  assign new_n21065_ = ~new_n21116_ | ~new_n21146_;
  assign new_n21066_ = ~pi0343;
  assign new_n21067_ = ~pi0342;
  assign new_n21068_ = ~new_n21117_ | ~new_n21140_;
  assign new_n21069_ = ~pi0344;
  assign new_n21070_ = ~pi0345;
  assign new_n21071_ = ~new_n21118_ | ~new_n21141_;
  assign new_n21072_ = ~pi0346;
  assign new_n21073_ = ~new_n21119_ | ~new_n21147_;
  assign new_n21074_ = ~new_n21148_ | ~pi0346;
  assign new_n21075_ = ~pi0347;
  assign new_n21076_ = ~new_n21167_ | ~new_n21166_;
  assign new_n21077_ = ~new_n21169_ | ~new_n21168_;
  assign new_n21078_ = ~new_n21171_ | ~new_n21170_;
  assign new_n21079_ = ~new_n21173_ | ~new_n21172_;
  assign new_n21080_ = ~new_n21175_ | ~new_n21174_;
  assign new_n21081_ = ~new_n21177_ | ~new_n21176_;
  assign new_n21082_ = ~new_n21179_ | ~new_n21178_;
  assign new_n21083_ = ~new_n21181_ | ~new_n21180_;
  assign new_n21084_ = ~new_n21183_ | ~new_n21182_;
  assign new_n21085_ = ~new_n21185_ | ~new_n21184_;
  assign new_n21086_ = ~new_n21187_ | ~new_n21186_;
  assign new_n21087_ = ~new_n21189_ | ~new_n21188_;
  assign new_n21088_ = ~new_n21191_ | ~new_n21190_;
  assign new_n21089_ = ~new_n21193_ | ~new_n21192_;
  assign new_n21090_ = ~new_n21195_ | ~new_n21194_;
  assign new_n21091_ = ~new_n21197_ | ~new_n21196_;
  assign new_n21092_ = ~new_n21199_ | ~new_n21198_;
  assign new_n21093_ = ~new_n21201_ | ~new_n21200_;
  assign new_n21094_ = ~new_n21203_ | ~new_n21202_;
  assign new_n21095_ = ~new_n21205_ | ~new_n21204_;
  assign new_n21096_ = ~new_n21207_ | ~new_n21206_;
  assign new_n21097_ = ~new_n21209_ | ~new_n21208_;
  assign new_n21098_ = ~new_n21211_ | ~new_n21210_;
  assign new_n21099_ = ~new_n21213_ | ~new_n21212_;
  assign new_n21100_ = ~new_n21215_ | ~new_n21214_;
  assign new_n21101_ = ~new_n21217_ | ~new_n21216_;
  assign new_n21102_ = ~new_n21219_ | ~new_n21218_;
  assign new_n21103_ = ~new_n21221_ | ~new_n21220_;
  assign new_n21104_ = ~new_n21223_ | ~new_n21222_;
  assign new_n21105_ = ~new_n21225_ | ~new_n21224_;
  assign new_n21106_ = ~new_n21227_ | ~new_n21226_;
  assign new_n21107_ = pi0320 & pi0321;
  assign new_n21108_ = pi0322 & pi0323;
  assign new_n21109_ = pi0324 & pi0325;
  assign new_n21110_ = pi0326 & pi0327;
  assign new_n21111_ = pi0328 & pi0329;
  assign new_n21112_ = pi0330 & pi0331;
  assign new_n21113_ = pi0333 & pi0332;
  assign new_n21114_ = pi0334 & pi0335;
  assign new_n21115_ = pi0336 & pi0337;
  assign new_n21116_ = pi0339 & pi0338;
  assign new_n21117_ = pi0340 & pi0341;
  assign new_n21118_ = pi0342 & pi0343;
  assign new_n21119_ = pi0345 & pi0344;
  assign new_n21120_ = ~new_n21143_ | ~pi0324;
  assign new_n21121_ = ~new_n21137_ | ~pi0322;
  assign new_n21122_ = ~new_n21136_ | ~pi0320;
  assign new_n21123_ = ~pi0348;
  assign new_n21124_ = ~pi0347 | ~new_n21153_;
  assign new_n21125_ = ~pi0318 | ~pi0317;
  assign new_n21126_ = ~new_n21147_ | ~pi0344;
  assign new_n21127_ = ~new_n21141_ | ~pi0342;
  assign new_n21128_ = ~new_n21140_ | ~pi0340;
  assign new_n21129_ = ~new_n21146_ | ~pi0338;
  assign new_n21130_ = ~new_n21139_ | ~pi0336;
  assign new_n21131_ = ~new_n21142_ | ~pi0334;
  assign new_n21132_ = ~new_n21149_ | ~pi0332;
  assign new_n21133_ = ~new_n21144_ | ~pi0330;
  assign new_n21134_ = ~new_n21138_ | ~pi0328;
  assign new_n21135_ = ~pi0326 | ~new_n21145_;
  assign new_n21136_ = ~new_n21035_;
  assign new_n21137_ = ~new_n21038_;
  assign new_n21138_ = ~new_n21047_;
  assign new_n21139_ = ~new_n21059_;
  assign new_n21140_ = ~new_n21065_;
  assign new_n21141_ = ~new_n21068_;
  assign new_n21142_ = ~new_n21056_;
  assign new_n21143_ = ~new_n21041_;
  assign new_n21144_ = ~new_n21050_;
  assign new_n21145_ = ~new_n21042_;
  assign new_n21146_ = ~new_n21061_;
  assign new_n21147_ = ~new_n21071_;
  assign new_n21148_ = ~new_n21073_;
  assign new_n21149_ = ~new_n21052_;
  assign new_n21150_ = ~new_n21120_;
  assign new_n21151_ = ~new_n21121_;
  assign new_n21152_ = ~new_n21122_;
  assign new_n21153_ = ~new_n21074_;
  assign new_n21154_ = ~new_n21124_;
  assign new_n21155_ = ~new_n21125_;
  assign new_n21156_ = ~new_n21126_;
  assign new_n21157_ = ~new_n21127_;
  assign new_n21158_ = ~new_n21128_;
  assign new_n21159_ = ~new_n21129_;
  assign new_n21160_ = ~new_n21130_;
  assign new_n21161_ = ~new_n21131_;
  assign new_n21162_ = ~new_n21132_;
  assign new_n21163_ = ~new_n21133_;
  assign new_n21164_ = ~new_n21134_;
  assign new_n21165_ = ~new_n21135_;
  assign new_n21166_ = ~new_n21145_ | ~new_n21043_;
  assign new_n21167_ = ~pi0326 | ~new_n21042_;
  assign new_n21168_ = ~pi0325 | ~new_n21120_;
  assign new_n21169_ = ~new_n21150_ | ~new_n21039_;
  assign new_n21170_ = ~new_n21143_ | ~new_n21040_;
  assign new_n21171_ = ~pi0324 | ~new_n21041_;
  assign new_n21172_ = ~pi0323 | ~new_n21121_;
  assign new_n21173_ = ~new_n21151_ | ~new_n21036_;
  assign new_n21174_ = ~new_n21137_ | ~new_n21037_;
  assign new_n21175_ = ~pi0322 | ~new_n21038_;
  assign new_n21176_ = ~pi0321 | ~new_n21122_;
  assign new_n21177_ = ~new_n21152_ | ~new_n21033_;
  assign new_n21178_ = ~new_n21136_ | ~new_n21034_;
  assign new_n21179_ = ~pi0320 | ~new_n21035_;
  assign new_n21180_ = ~pi0348 | ~new_n21124_;
  assign new_n21181_ = ~new_n21154_ | ~new_n21123_;
  assign new_n21182_ = ~pi0347 | ~new_n21074_;
  assign new_n21183_ = ~new_n21153_ | ~new_n21075_;
  assign new_n21184_ = ~pi0319 | ~new_n21125_;
  assign new_n21185_ = ~new_n21155_ | ~new_n21031_;
  assign new_n21186_ = ~new_n21148_ | ~new_n21072_;
  assign new_n21187_ = ~pi0346 | ~new_n21073_;
  assign new_n21188_ = ~pi0345 | ~new_n21126_;
  assign new_n21189_ = ~new_n21156_ | ~new_n21070_;
  assign new_n21190_ = ~new_n21147_ | ~new_n21069_;
  assign new_n21191_ = ~pi0344 | ~new_n21071_;
  assign new_n21192_ = ~pi0343 | ~new_n21127_;
  assign new_n21193_ = ~new_n21157_ | ~new_n21066_;
  assign new_n21194_ = ~new_n21141_ | ~new_n21067_;
  assign new_n21195_ = ~pi0342 | ~new_n21068_;
  assign new_n21196_ = ~pi0341 | ~new_n21128_;
  assign new_n21197_ = ~new_n21158_ | ~new_n21063_;
  assign new_n21198_ = ~new_n21140_ | ~new_n21064_;
  assign new_n21199_ = ~pi0340 | ~new_n21065_;
  assign new_n21200_ = ~pi0339 | ~new_n21129_;
  assign new_n21201_ = ~new_n21159_ | ~new_n21062_;
  assign new_n21202_ = ~new_n21146_ | ~new_n21060_;
  assign new_n21203_ = ~pi0338 | ~new_n21061_;
  assign new_n21204_ = ~pi0337 | ~new_n21130_;
  assign new_n21205_ = ~new_n21160_ | ~new_n21057_;
  assign new_n21206_ = ~pi0317 | ~new_n21032_;
  assign new_n21207_ = ~pi0318 | ~new_n21030_;
  assign new_n21208_ = ~new_n21139_ | ~new_n21058_;
  assign new_n21209_ = ~pi0336 | ~new_n21059_;
  assign new_n21210_ = ~pi0335 | ~new_n21131_;
  assign new_n21211_ = ~new_n21161_ | ~new_n21054_;
  assign new_n21212_ = ~new_n21142_ | ~new_n21055_;
  assign new_n21213_ = ~pi0334 | ~new_n21056_;
  assign new_n21214_ = ~pi0333 | ~new_n21132_;
  assign new_n21215_ = ~new_n21162_ | ~new_n21053_;
  assign new_n21216_ = ~new_n21149_ | ~new_n21051_;
  assign new_n21217_ = ~pi0332 | ~new_n21052_;
  assign new_n21218_ = ~pi0331 | ~new_n21133_;
  assign new_n21219_ = ~new_n21163_ | ~new_n21048_;
  assign new_n21220_ = ~new_n21144_ | ~new_n21049_;
  assign new_n21221_ = ~pi0330 | ~new_n21050_;
  assign new_n21222_ = ~pi0329 | ~new_n21134_;
  assign new_n21223_ = ~new_n21164_ | ~new_n21045_;
  assign new_n21224_ = ~new_n21138_ | ~new_n21046_;
  assign new_n21225_ = ~pi0328 | ~new_n21047_;
  assign new_n21226_ = ~pi0327 | ~new_n21135_;
  assign new_n21227_ = ~new_n21165_ | ~new_n21044_;
  assign new_n21228_ = ~pi0476;
  assign new_n21229_ = ~pi0478;
  assign new_n21230_ = ~pi0477;
  assign new_n21231_ = ~pi0480;
  assign new_n21232_ = ~pi0479;
  assign new_n21233_ = ~pi0477 | ~pi0478 | ~pi0476;
  assign new_n21234_ = ~pi0482;
  assign new_n21235_ = ~pi0481;
  assign new_n21236_ = ~new_n21305_ | ~new_n21334_;
  assign new_n21237_ = ~pi0484;
  assign new_n21238_ = ~pi0483;
  assign new_n21239_ = ~new_n21306_ | ~new_n21335_;
  assign new_n21240_ = ~new_n21307_ | ~new_n21341_;
  assign new_n21241_ = ~pi0485;
  assign new_n21242_ = ~pi0486;
  assign new_n21243_ = ~pi0488;
  assign new_n21244_ = ~pi0487;
  assign new_n21245_ = ~new_n21308_ | ~new_n21343_;
  assign new_n21246_ = ~pi0490;
  assign new_n21247_ = ~pi0489;
  assign new_n21248_ = ~new_n21309_ | ~new_n21336_;
  assign new_n21249_ = ~pi0491;
  assign new_n21250_ = ~new_n21310_ | ~new_n21342_;
  assign new_n21251_ = ~pi0492;
  assign new_n21252_ = ~pi0494;
  assign new_n21253_ = ~pi0493;
  assign new_n21254_ = ~new_n21311_ | ~new_n21347_;
  assign new_n21255_ = ~pi0496;
  assign new_n21256_ = ~pi0495;
  assign new_n21257_ = ~new_n21312_ | ~new_n21340_;
  assign new_n21258_ = ~pi0497;
  assign new_n21259_ = ~new_n21313_ | ~new_n21337_;
  assign new_n21260_ = ~pi0498;
  assign new_n21261_ = ~pi0500;
  assign new_n21262_ = ~pi0499;
  assign new_n21263_ = ~new_n21314_ | ~new_n21344_;
  assign new_n21264_ = ~pi0502;
  assign new_n21265_ = ~pi0501;
  assign new_n21266_ = ~new_n21315_ | ~new_n21338_;
  assign new_n21267_ = ~pi0503;
  assign new_n21268_ = ~pi0504;
  assign new_n21269_ = ~new_n21316_ | ~new_n21339_;
  assign new_n21270_ = ~pi0505;
  assign new_n21271_ = ~new_n21317_ | ~new_n21345_;
  assign new_n21272_ = ~new_n21346_ | ~pi0505;
  assign new_n21273_ = ~pi0506;
  assign new_n21274_ = ~new_n21365_ | ~new_n21364_;
  assign new_n21275_ = ~new_n21367_ | ~new_n21366_;
  assign new_n21276_ = ~new_n21369_ | ~new_n21368_;
  assign new_n21277_ = ~new_n21371_ | ~new_n21370_;
  assign new_n21278_ = ~new_n21373_ | ~new_n21372_;
  assign new_n21279_ = ~new_n21375_ | ~new_n21374_;
  assign new_n21280_ = ~new_n21377_ | ~new_n21376_;
  assign new_n21281_ = ~new_n21379_ | ~new_n21378_;
  assign new_n21282_ = ~new_n21381_ | ~new_n21380_;
  assign new_n21283_ = ~new_n21383_ | ~new_n21382_;
  assign new_n21284_ = ~new_n21385_ | ~new_n21384_;
  assign new_n21285_ = ~new_n21387_ | ~new_n21386_;
  assign new_n21286_ = ~new_n21389_ | ~new_n21388_;
  assign new_n21287_ = ~new_n21391_ | ~new_n21390_;
  assign new_n21288_ = ~new_n21393_ | ~new_n21392_;
  assign new_n21289_ = ~new_n21395_ | ~new_n21394_;
  assign new_n21290_ = ~new_n21397_ | ~new_n21396_;
  assign new_n21291_ = ~new_n21399_ | ~new_n21398_;
  assign new_n21292_ = ~new_n21401_ | ~new_n21400_;
  assign new_n21293_ = ~new_n21403_ | ~new_n21402_;
  assign new_n21294_ = ~new_n21405_ | ~new_n21404_;
  assign new_n21295_ = ~new_n21407_ | ~new_n21406_;
  assign new_n21296_ = ~new_n21409_ | ~new_n21408_;
  assign new_n21297_ = ~new_n21411_ | ~new_n21410_;
  assign new_n21298_ = ~new_n21413_ | ~new_n21412_;
  assign new_n21299_ = ~new_n21415_ | ~new_n21414_;
  assign new_n21300_ = ~new_n21417_ | ~new_n21416_;
  assign new_n21301_ = ~new_n21419_ | ~new_n21418_;
  assign new_n21302_ = ~new_n21421_ | ~new_n21420_;
  assign new_n21303_ = ~new_n21423_ | ~new_n21422_;
  assign new_n21304_ = ~new_n21425_ | ~new_n21424_;
  assign new_n21305_ = pi0479 & pi0480;
  assign new_n21306_ = pi0481 & pi0482;
  assign new_n21307_ = pi0483 & pi0484;
  assign new_n21308_ = pi0485 & pi0486;
  assign new_n21309_ = pi0487 & pi0488;
  assign new_n21310_ = pi0489 & pi0490;
  assign new_n21311_ = pi0492 & pi0491;
  assign new_n21312_ = pi0493 & pi0494;
  assign new_n21313_ = pi0495 & pi0496;
  assign new_n21314_ = pi0498 & pi0497;
  assign new_n21315_ = pi0499 & pi0500;
  assign new_n21316_ = pi0501 & pi0502;
  assign new_n21317_ = pi0504 & pi0503;
  assign new_n21318_ = ~new_n21341_ | ~pi0483;
  assign new_n21319_ = ~new_n21335_ | ~pi0481;
  assign new_n21320_ = ~new_n21334_ | ~pi0479;
  assign new_n21321_ = ~pi0507;
  assign new_n21322_ = ~pi0506 | ~new_n21351_;
  assign new_n21323_ = ~pi0477 | ~pi0476;
  assign new_n21324_ = ~new_n21345_ | ~pi0503;
  assign new_n21325_ = ~new_n21339_ | ~pi0501;
  assign new_n21326_ = ~new_n21338_ | ~pi0499;
  assign new_n21327_ = ~new_n21344_ | ~pi0497;
  assign new_n21328_ = ~new_n21337_ | ~pi0495;
  assign new_n21329_ = ~new_n21340_ | ~pi0493;
  assign new_n21330_ = ~new_n21347_ | ~pi0491;
  assign new_n21331_ = ~new_n21342_ | ~pi0489;
  assign new_n21332_ = ~new_n21336_ | ~pi0487;
  assign new_n21333_ = ~pi0485 | ~new_n21343_;
  assign new_n21334_ = ~new_n21233_;
  assign new_n21335_ = ~new_n21236_;
  assign new_n21336_ = ~new_n21245_;
  assign new_n21337_ = ~new_n21257_;
  assign new_n21338_ = ~new_n21263_;
  assign new_n21339_ = ~new_n21266_;
  assign new_n21340_ = ~new_n21254_;
  assign new_n21341_ = ~new_n21239_;
  assign new_n21342_ = ~new_n21248_;
  assign new_n21343_ = ~new_n21240_;
  assign new_n21344_ = ~new_n21259_;
  assign new_n21345_ = ~new_n21269_;
  assign new_n21346_ = ~new_n21271_;
  assign new_n21347_ = ~new_n21250_;
  assign new_n21348_ = ~new_n21318_;
  assign new_n21349_ = ~new_n21319_;
  assign new_n21350_ = ~new_n21320_;
  assign new_n21351_ = ~new_n21272_;
  assign new_n21352_ = ~new_n21322_;
  assign new_n21353_ = ~new_n21323_;
  assign new_n21354_ = ~new_n21324_;
  assign new_n21355_ = ~new_n21325_;
  assign new_n21356_ = ~new_n21326_;
  assign new_n21357_ = ~new_n21327_;
  assign new_n21358_ = ~new_n21328_;
  assign new_n21359_ = ~new_n21329_;
  assign new_n21360_ = ~new_n21330_;
  assign new_n21361_ = ~new_n21331_;
  assign new_n21362_ = ~new_n21332_;
  assign new_n21363_ = ~new_n21333_;
  assign new_n21364_ = ~new_n21343_ | ~new_n21241_;
  assign new_n21365_ = ~pi0485 | ~new_n21240_;
  assign new_n21366_ = ~pi0484 | ~new_n21318_;
  assign new_n21367_ = ~new_n21348_ | ~new_n21237_;
  assign new_n21368_ = ~new_n21341_ | ~new_n21238_;
  assign new_n21369_ = ~pi0483 | ~new_n21239_;
  assign new_n21370_ = ~pi0482 | ~new_n21319_;
  assign new_n21371_ = ~new_n21349_ | ~new_n21234_;
  assign new_n21372_ = ~new_n21335_ | ~new_n21235_;
  assign new_n21373_ = ~pi0481 | ~new_n21236_;
  assign new_n21374_ = ~pi0480 | ~new_n21320_;
  assign new_n21375_ = ~new_n21350_ | ~new_n21231_;
  assign new_n21376_ = ~new_n21334_ | ~new_n21232_;
  assign new_n21377_ = ~pi0479 | ~new_n21233_;
  assign new_n21378_ = ~pi0507 | ~new_n21322_;
  assign new_n21379_ = ~new_n21352_ | ~new_n21321_;
  assign new_n21380_ = ~pi0506 | ~new_n21272_;
  assign new_n21381_ = ~new_n21351_ | ~new_n21273_;
  assign new_n21382_ = ~pi0478 | ~new_n21323_;
  assign new_n21383_ = ~new_n21353_ | ~new_n21229_;
  assign new_n21384_ = ~new_n21346_ | ~new_n21270_;
  assign new_n21385_ = ~pi0505 | ~new_n21271_;
  assign new_n21386_ = ~pi0504 | ~new_n21324_;
  assign new_n21387_ = ~new_n21354_ | ~new_n21268_;
  assign new_n21388_ = ~new_n21345_ | ~new_n21267_;
  assign new_n21389_ = ~pi0503 | ~new_n21269_;
  assign new_n21390_ = ~pi0502 | ~new_n21325_;
  assign new_n21391_ = ~new_n21355_ | ~new_n21264_;
  assign new_n21392_ = ~new_n21339_ | ~new_n21265_;
  assign new_n21393_ = ~pi0501 | ~new_n21266_;
  assign new_n21394_ = ~pi0500 | ~new_n21326_;
  assign new_n21395_ = ~new_n21356_ | ~new_n21261_;
  assign new_n21396_ = ~new_n21338_ | ~new_n21262_;
  assign new_n21397_ = ~pi0499 | ~new_n21263_;
  assign new_n21398_ = ~pi0498 | ~new_n21327_;
  assign new_n21399_ = ~new_n21357_ | ~new_n21260_;
  assign new_n21400_ = ~new_n21344_ | ~new_n21258_;
  assign new_n21401_ = ~pi0497 | ~new_n21259_;
  assign new_n21402_ = ~pi0496 | ~new_n21328_;
  assign new_n21403_ = ~new_n21358_ | ~new_n21255_;
  assign new_n21404_ = ~pi0476 | ~new_n21230_;
  assign new_n21405_ = ~pi0477 | ~new_n21228_;
  assign new_n21406_ = ~new_n21337_ | ~new_n21256_;
  assign new_n21407_ = ~pi0495 | ~new_n21257_;
  assign new_n21408_ = ~pi0494 | ~new_n21329_;
  assign new_n21409_ = ~new_n21359_ | ~new_n21252_;
  assign new_n21410_ = ~new_n21340_ | ~new_n21253_;
  assign new_n21411_ = ~pi0493 | ~new_n21254_;
  assign new_n21412_ = ~pi0492 | ~new_n21330_;
  assign new_n21413_ = ~new_n21360_ | ~new_n21251_;
  assign new_n21414_ = ~new_n21347_ | ~new_n21249_;
  assign new_n21415_ = ~pi0491 | ~new_n21250_;
  assign new_n21416_ = ~pi0490 | ~new_n21331_;
  assign new_n21417_ = ~new_n21361_ | ~new_n21246_;
  assign new_n21418_ = ~new_n21342_ | ~new_n21247_;
  assign new_n21419_ = ~pi0489 | ~new_n21248_;
  assign new_n21420_ = ~pi0488 | ~new_n21332_;
  assign new_n21421_ = ~new_n21362_ | ~new_n21243_;
  assign new_n21422_ = ~new_n21336_ | ~new_n21244_;
  assign new_n21423_ = ~pi0487 | ~new_n21245_;
  assign new_n21424_ = ~pi0486 | ~new_n21333_;
  assign new_n21425_ = ~new_n21363_ | ~new_n21242_;
  assign new_n21426_ = ~pi0444;
  assign new_n21427_ = ~pi0446;
  assign new_n21428_ = ~pi0445;
  assign new_n21429_ = ~pi0448;
  assign new_n21430_ = ~pi0447;
  assign new_n21431_ = ~pi0445 | ~pi0446 | ~pi0444;
  assign new_n21432_ = ~pi0450;
  assign new_n21433_ = ~pi0449;
  assign new_n21434_ = ~new_n21503_ | ~new_n21532_;
  assign new_n21435_ = ~pi0452;
  assign new_n21436_ = ~pi0451;
  assign new_n21437_ = ~new_n21504_ | ~new_n21533_;
  assign new_n21438_ = ~new_n21505_ | ~new_n21539_;
  assign new_n21439_ = ~pi0453;
  assign new_n21440_ = ~pi0454;
  assign new_n21441_ = ~pi0456;
  assign new_n21442_ = ~pi0455;
  assign new_n21443_ = ~new_n21506_ | ~new_n21541_;
  assign new_n21444_ = ~pi0458;
  assign new_n21445_ = ~pi0457;
  assign new_n21446_ = ~new_n21507_ | ~new_n21534_;
  assign new_n21447_ = ~pi0459;
  assign new_n21448_ = ~new_n21508_ | ~new_n21540_;
  assign new_n21449_ = ~pi0460;
  assign new_n21450_ = ~pi0462;
  assign new_n21451_ = ~pi0461;
  assign new_n21452_ = ~new_n21509_ | ~new_n21545_;
  assign new_n21453_ = ~pi0464;
  assign new_n21454_ = ~pi0463;
  assign new_n21455_ = ~new_n21510_ | ~new_n21538_;
  assign new_n21456_ = ~pi0465;
  assign new_n21457_ = ~new_n21511_ | ~new_n21535_;
  assign new_n21458_ = ~pi0466;
  assign new_n21459_ = ~pi0468;
  assign new_n21460_ = ~pi0467;
  assign new_n21461_ = ~new_n21512_ | ~new_n21542_;
  assign new_n21462_ = ~pi0470;
  assign new_n21463_ = ~pi0469;
  assign new_n21464_ = ~new_n21513_ | ~new_n21536_;
  assign new_n21465_ = ~pi0471;
  assign new_n21466_ = ~pi0472;
  assign new_n21467_ = ~new_n21514_ | ~new_n21537_;
  assign new_n21468_ = ~pi0473;
  assign new_n21469_ = ~new_n21515_ | ~new_n21543_;
  assign new_n21470_ = ~new_n21544_ | ~pi0473;
  assign new_n21471_ = ~pi0474;
  assign new_n21472_ = ~new_n21563_ | ~new_n21562_;
  assign new_n21473_ = ~new_n21565_ | ~new_n21564_;
  assign new_n21474_ = ~new_n21567_ | ~new_n21566_;
  assign new_n21475_ = ~new_n21569_ | ~new_n21568_;
  assign new_n21476_ = ~new_n21571_ | ~new_n21570_;
  assign new_n21477_ = ~new_n21573_ | ~new_n21572_;
  assign new_n21478_ = ~new_n21575_ | ~new_n21574_;
  assign new_n21479_ = ~new_n21577_ | ~new_n21576_;
  assign new_n21480_ = ~new_n21579_ | ~new_n21578_;
  assign new_n21481_ = ~new_n21581_ | ~new_n21580_;
  assign new_n21482_ = ~new_n21583_ | ~new_n21582_;
  assign new_n21483_ = ~new_n21585_ | ~new_n21584_;
  assign new_n21484_ = ~new_n21587_ | ~new_n21586_;
  assign new_n21485_ = ~new_n21589_ | ~new_n21588_;
  assign new_n21486_ = ~new_n21591_ | ~new_n21590_;
  assign new_n21487_ = ~new_n21593_ | ~new_n21592_;
  assign new_n21488_ = ~new_n21595_ | ~new_n21594_;
  assign new_n21489_ = ~new_n21597_ | ~new_n21596_;
  assign new_n21490_ = ~new_n21599_ | ~new_n21598_;
  assign new_n21491_ = ~new_n21601_ | ~new_n21600_;
  assign new_n21492_ = ~new_n21603_ | ~new_n21602_;
  assign new_n21493_ = ~new_n21605_ | ~new_n21604_;
  assign new_n21494_ = ~new_n21607_ | ~new_n21606_;
  assign new_n21495_ = ~new_n21609_ | ~new_n21608_;
  assign new_n21496_ = ~new_n21611_ | ~new_n21610_;
  assign new_n21497_ = ~new_n21613_ | ~new_n21612_;
  assign new_n21498_ = ~new_n21615_ | ~new_n21614_;
  assign new_n21499_ = ~new_n21617_ | ~new_n21616_;
  assign new_n21500_ = ~new_n21619_ | ~new_n21618_;
  assign new_n21501_ = ~new_n21621_ | ~new_n21620_;
  assign new_n21502_ = ~new_n21623_ | ~new_n21622_;
  assign new_n21503_ = pi0447 & pi0448;
  assign new_n21504_ = pi0449 & pi0450;
  assign new_n21505_ = pi0451 & pi0452;
  assign new_n21506_ = pi0453 & pi0454;
  assign new_n21507_ = pi0455 & pi0456;
  assign new_n21508_ = pi0457 & pi0458;
  assign new_n21509_ = pi0460 & pi0459;
  assign new_n21510_ = pi0461 & pi0462;
  assign new_n21511_ = pi0463 & pi0464;
  assign new_n21512_ = pi0466 & pi0465;
  assign new_n21513_ = pi0467 & pi0468;
  assign new_n21514_ = pi0469 & pi0470;
  assign new_n21515_ = pi0472 & pi0471;
  assign new_n21516_ = ~new_n21539_ | ~pi0451;
  assign new_n21517_ = ~new_n21533_ | ~pi0449;
  assign new_n21518_ = ~new_n21532_ | ~pi0447;
  assign new_n21519_ = ~pi0475;
  assign new_n21520_ = ~pi0474 | ~new_n21549_;
  assign new_n21521_ = ~pi0445 | ~pi0444;
  assign new_n21522_ = ~new_n21543_ | ~pi0471;
  assign new_n21523_ = ~new_n21537_ | ~pi0469;
  assign new_n21524_ = ~new_n21536_ | ~pi0467;
  assign new_n21525_ = ~new_n21542_ | ~pi0465;
  assign new_n21526_ = ~new_n21535_ | ~pi0463;
  assign new_n21527_ = ~new_n21538_ | ~pi0461;
  assign new_n21528_ = ~new_n21545_ | ~pi0459;
  assign new_n21529_ = ~new_n21540_ | ~pi0457;
  assign new_n21530_ = ~new_n21534_ | ~pi0455;
  assign new_n21531_ = ~pi0453 | ~new_n21541_;
  assign new_n21532_ = ~new_n21431_;
  assign new_n21533_ = ~new_n21434_;
  assign new_n21534_ = ~new_n21443_;
  assign new_n21535_ = ~new_n21455_;
  assign new_n21536_ = ~new_n21461_;
  assign new_n21537_ = ~new_n21464_;
  assign new_n21538_ = ~new_n21452_;
  assign new_n21539_ = ~new_n21437_;
  assign new_n21540_ = ~new_n21446_;
  assign new_n21541_ = ~new_n21438_;
  assign new_n21542_ = ~new_n21457_;
  assign new_n21543_ = ~new_n21467_;
  assign new_n21544_ = ~new_n21469_;
  assign new_n21545_ = ~new_n21448_;
  assign new_n21546_ = ~new_n21516_;
  assign new_n21547_ = ~new_n21517_;
  assign new_n21548_ = ~new_n21518_;
  assign new_n21549_ = ~new_n21470_;
  assign new_n21550_ = ~new_n21520_;
  assign new_n21551_ = ~new_n21521_;
  assign new_n21552_ = ~new_n21522_;
  assign new_n21553_ = ~new_n21523_;
  assign new_n21554_ = ~new_n21524_;
  assign new_n21555_ = ~new_n21525_;
  assign new_n21556_ = ~new_n21526_;
  assign new_n21557_ = ~new_n21527_;
  assign new_n21558_ = ~new_n21528_;
  assign new_n21559_ = ~new_n21529_;
  assign new_n21560_ = ~new_n21530_;
  assign new_n21561_ = ~new_n21531_;
  assign new_n21562_ = ~new_n21541_ | ~new_n21439_;
  assign new_n21563_ = ~pi0453 | ~new_n21438_;
  assign new_n21564_ = ~pi0452 | ~new_n21516_;
  assign new_n21565_ = ~new_n21546_ | ~new_n21435_;
  assign new_n21566_ = ~new_n21539_ | ~new_n21436_;
  assign new_n21567_ = ~pi0451 | ~new_n21437_;
  assign new_n21568_ = ~pi0450 | ~new_n21517_;
  assign new_n21569_ = ~new_n21547_ | ~new_n21432_;
  assign new_n21570_ = ~new_n21533_ | ~new_n21433_;
  assign new_n21571_ = ~pi0449 | ~new_n21434_;
  assign new_n21572_ = ~pi0448 | ~new_n21518_;
  assign new_n21573_ = ~new_n21548_ | ~new_n21429_;
  assign new_n21574_ = ~new_n21532_ | ~new_n21430_;
  assign new_n21575_ = ~pi0447 | ~new_n21431_;
  assign new_n21576_ = ~pi0475 | ~new_n21520_;
  assign new_n21577_ = ~new_n21550_ | ~new_n21519_;
  assign new_n21578_ = ~pi0474 | ~new_n21470_;
  assign new_n21579_ = ~new_n21549_ | ~new_n21471_;
  assign new_n21580_ = ~pi0446 | ~new_n21521_;
  assign new_n21581_ = ~new_n21551_ | ~new_n21427_;
  assign new_n21582_ = ~new_n21544_ | ~new_n21468_;
  assign new_n21583_ = ~pi0473 | ~new_n21469_;
  assign new_n21584_ = ~pi0472 | ~new_n21522_;
  assign new_n21585_ = ~new_n21552_ | ~new_n21466_;
  assign new_n21586_ = ~new_n21543_ | ~new_n21465_;
  assign new_n21587_ = ~pi0471 | ~new_n21467_;
  assign new_n21588_ = ~pi0470 | ~new_n21523_;
  assign new_n21589_ = ~new_n21553_ | ~new_n21462_;
  assign new_n21590_ = ~new_n21537_ | ~new_n21463_;
  assign new_n21591_ = ~pi0469 | ~new_n21464_;
  assign new_n21592_ = ~pi0468 | ~new_n21524_;
  assign new_n21593_ = ~new_n21554_ | ~new_n21459_;
  assign new_n21594_ = ~new_n21536_ | ~new_n21460_;
  assign new_n21595_ = ~pi0467 | ~new_n21461_;
  assign new_n21596_ = ~pi0466 | ~new_n21525_;
  assign new_n21597_ = ~new_n21555_ | ~new_n21458_;
  assign new_n21598_ = ~new_n21542_ | ~new_n21456_;
  assign new_n21599_ = ~pi0465 | ~new_n21457_;
  assign new_n21600_ = ~pi0464 | ~new_n21526_;
  assign new_n21601_ = ~new_n21556_ | ~new_n21453_;
  assign new_n21602_ = ~pi0444 | ~new_n21428_;
  assign new_n21603_ = ~pi0445 | ~new_n21426_;
  assign new_n21604_ = ~new_n21535_ | ~new_n21454_;
  assign new_n21605_ = ~pi0463 | ~new_n21455_;
  assign new_n21606_ = ~pi0462 | ~new_n21527_;
  assign new_n21607_ = ~new_n21557_ | ~new_n21450_;
  assign new_n21608_ = ~new_n21538_ | ~new_n21451_;
  assign new_n21609_ = ~pi0461 | ~new_n21452_;
  assign new_n21610_ = ~pi0460 | ~new_n21528_;
  assign new_n21611_ = ~new_n21558_ | ~new_n21449_;
  assign new_n21612_ = ~new_n21545_ | ~new_n21447_;
  assign new_n21613_ = ~pi0459 | ~new_n21448_;
  assign new_n21614_ = ~pi0458 | ~new_n21529_;
  assign new_n21615_ = ~new_n21559_ | ~new_n21444_;
  assign new_n21616_ = ~new_n21540_ | ~new_n21445_;
  assign new_n21617_ = ~pi0457 | ~new_n21446_;
  assign new_n21618_ = ~pi0456 | ~new_n21530_;
  assign new_n21619_ = ~new_n21560_ | ~new_n21441_;
  assign new_n21620_ = ~new_n21534_ | ~new_n21442_;
  assign new_n21621_ = ~pi0455 | ~new_n21443_;
  assign new_n21622_ = ~pi0454 | ~new_n21531_;
  assign new_n21623_ = ~new_n21561_ | ~new_n21440_;
  assign new_n21624_ = ~new_n26956_ & ~new_n21626_;
  assign new_n21625_ = new_n26971_ & new_n21627_;
  assign new_n21626_ = ~new_n26970_ & ~new_n21625_ & ~new_n26969_;
  assign new_n21627_ = new_n26957_ | new_n26972_;
  assign new_n21628_ = ~new_n3769_;
  assign new_n21629_ = ~new_n4225_;
  assign new_n21630_ = ~new_n4225_ | ~new_n3769_;
  assign new_n21631_ = ~new_n3770_;
  assign new_n21632_ = ~new_n3770_ | ~new_n21652_;
  assign new_n21633_ = ~new_n3771_;
  assign new_n21634_ = ~new_n3771_ | ~new_n21653_;
  assign new_n21635_ = ~new_n3772_;
  assign new_n21636_ = ~new_n3772_ | ~new_n21654_;
  assign new_n21637_ = ~new_n3773_;
  assign new_n21638_ = ~new_n3773_ | ~new_n21655_;
  assign new_n21639_ = ~new_n3774_;
  assign new_n21640_ = ~new_n3774_ | ~new_n21656_;
  assign new_n21641_ = ~new_n3775_;
  assign new_n21642_ = ~new_n21660_ | ~new_n21659_;
  assign new_n21643_ = ~new_n21662_ | ~new_n21661_;
  assign new_n21644_ = ~new_n21664_ | ~new_n21663_;
  assign new_n21645_ = ~new_n21666_ | ~new_n21665_;
  assign new_n21646_ = ~new_n21668_ | ~new_n21667_;
  assign new_n21647_ = ~new_n21670_ | ~new_n21669_;
  assign new_n21648_ = ~new_n21672_ | ~new_n21671_;
  assign new_n21649_ = ~new_n21674_ | ~new_n21673_;
  assign new_n21650_ = ~new_n3776_;
  assign new_n21651_ = ~new_n3775_ | ~new_n21657_;
  assign new_n21652_ = ~new_n21630_;
  assign new_n21653_ = ~new_n21632_;
  assign new_n21654_ = ~new_n21634_;
  assign new_n21655_ = ~new_n21636_;
  assign new_n21656_ = ~new_n21638_;
  assign new_n21657_ = ~new_n21640_;
  assign new_n21658_ = ~new_n21651_;
  assign new_n21659_ = ~new_n3776_ | ~new_n21651_;
  assign new_n21660_ = ~new_n21658_ | ~new_n21650_;
  assign new_n21661_ = ~new_n3775_ | ~new_n21640_;
  assign new_n21662_ = ~new_n21657_ | ~new_n21641_;
  assign new_n21663_ = ~new_n3774_ | ~new_n21638_;
  assign new_n21664_ = ~new_n21656_ | ~new_n21639_;
  assign new_n21665_ = ~new_n3773_ | ~new_n21636_;
  assign new_n21666_ = ~new_n21655_ | ~new_n21637_;
  assign new_n21667_ = ~new_n3772_ | ~new_n21634_;
  assign new_n21668_ = ~new_n21654_ | ~new_n21635_;
  assign new_n21669_ = ~new_n3771_ | ~new_n21632_;
  assign new_n21670_ = ~new_n21653_ | ~new_n21633_;
  assign new_n21671_ = ~new_n3770_ | ~new_n21630_;
  assign new_n21672_ = ~new_n21652_ | ~new_n21631_;
  assign new_n21673_ = ~new_n4225_ | ~new_n21628_;
  assign new_n21674_ = ~new_n3769_ | ~new_n21629_;
  assign new_n21675_ = ~pi0318;
  assign new_n21676_ = ~pi0319;
  assign new_n21677_ = ~pi0319 | ~pi0318;
  assign new_n21678_ = ~pi0320;
  assign new_n21679_ = ~pi0320 | ~new_n21765_;
  assign new_n21680_ = ~pi0321;
  assign new_n21681_ = ~pi0321 | ~new_n21766_;
  assign new_n21682_ = ~pi0322;
  assign new_n21683_ = ~pi0322 | ~new_n21767_;
  assign new_n21684_ = ~pi0323;
  assign new_n21685_ = ~pi0323 | ~new_n21768_;
  assign new_n21686_ = ~pi0324;
  assign new_n21687_ = ~pi0324 | ~new_n21769_;
  assign new_n21688_ = ~pi0325;
  assign new_n21689_ = ~pi0326;
  assign new_n21690_ = ~pi0325 | ~new_n21770_;
  assign new_n21691_ = ~new_n21771_ | ~pi0326;
  assign new_n21692_ = ~pi0327;
  assign new_n21693_ = ~pi0327 | ~new_n21772_;
  assign new_n21694_ = ~pi0328;
  assign new_n21695_ = ~pi0328 | ~new_n21773_;
  assign new_n21696_ = ~pi0329;
  assign new_n21697_ = ~pi0329 | ~new_n21774_;
  assign new_n21698_ = ~pi0330;
  assign new_n21699_ = ~pi0330 | ~new_n21775_;
  assign new_n21700_ = ~pi0331;
  assign new_n21701_ = ~pi0331 | ~new_n21776_;
  assign new_n21702_ = ~pi0332;
  assign new_n21703_ = ~pi0332 | ~new_n21777_;
  assign new_n21704_ = ~pi0333;
  assign new_n21705_ = ~pi0333 | ~new_n21778_;
  assign new_n21706_ = ~pi0334;
  assign new_n21707_ = ~pi0334 | ~new_n21779_;
  assign new_n21708_ = ~pi0335;
  assign new_n21709_ = ~pi0335 | ~new_n21780_;
  assign new_n21710_ = ~pi0336;
  assign new_n21711_ = ~pi0336 | ~new_n21781_;
  assign new_n21712_ = ~pi0337;
  assign new_n21713_ = ~pi0337 | ~new_n21782_;
  assign new_n21714_ = ~pi0338;
  assign new_n21715_ = ~pi0338 | ~new_n21783_;
  assign new_n21716_ = ~pi0339;
  assign new_n21717_ = ~pi0339 | ~new_n21784_;
  assign new_n21718_ = ~pi0340;
  assign new_n21719_ = ~pi0340 | ~new_n21785_;
  assign new_n21720_ = ~pi0341;
  assign new_n21721_ = ~pi0341 | ~new_n21786_;
  assign new_n21722_ = ~pi0342;
  assign new_n21723_ = ~pi0342 | ~new_n21787_;
  assign new_n21724_ = ~pi0343;
  assign new_n21725_ = ~pi0343 | ~new_n21788_;
  assign new_n21726_ = ~pi0344;
  assign new_n21727_ = ~pi0344 | ~new_n21789_;
  assign new_n21728_ = ~pi0345;
  assign new_n21729_ = ~pi0345 | ~new_n21790_;
  assign new_n21730_ = ~pi0346;
  assign new_n21731_ = ~pi0346 | ~new_n21791_;
  assign new_n21732_ = ~pi0347;
  assign new_n21733_ = ~new_n21795_ | ~new_n21794_;
  assign new_n21734_ = ~new_n21797_ | ~new_n21796_;
  assign new_n21735_ = ~new_n21799_ | ~new_n21798_;
  assign new_n21736_ = ~new_n21801_ | ~new_n21800_;
  assign new_n21737_ = ~new_n21803_ | ~new_n21802_;
  assign new_n21738_ = ~new_n21805_ | ~new_n21804_;
  assign new_n21739_ = ~new_n21807_ | ~new_n21806_;
  assign new_n21740_ = ~new_n21809_ | ~new_n21808_;
  assign new_n21741_ = ~new_n21811_ | ~new_n21810_;
  assign new_n21742_ = ~new_n21813_ | ~new_n21812_;
  assign new_n21743_ = ~new_n21815_ | ~new_n21814_;
  assign new_n21744_ = ~new_n21817_ | ~new_n21816_;
  assign new_n21745_ = ~new_n21819_ | ~new_n21818_;
  assign new_n21746_ = ~new_n21821_ | ~new_n21820_;
  assign new_n21747_ = ~new_n21823_ | ~new_n21822_;
  assign new_n21748_ = ~new_n21825_ | ~new_n21824_;
  assign new_n21749_ = ~new_n21827_ | ~new_n21826_;
  assign new_n21750_ = ~new_n21829_ | ~new_n21828_;
  assign new_n21751_ = ~new_n21831_ | ~new_n21830_;
  assign new_n21752_ = ~new_n21833_ | ~new_n21832_;
  assign new_n21753_ = ~new_n21835_ | ~new_n21834_;
  assign new_n21754_ = ~new_n21837_ | ~new_n21836_;
  assign new_n21755_ = ~new_n21839_ | ~new_n21838_;
  assign new_n21756_ = ~new_n21841_ | ~new_n21840_;
  assign new_n21757_ = ~new_n21843_ | ~new_n21842_;
  assign new_n21758_ = ~new_n21845_ | ~new_n21844_;
  assign new_n21759_ = ~new_n21847_ | ~new_n21846_;
  assign new_n21760_ = ~new_n21849_ | ~new_n21848_;
  assign new_n21761_ = ~new_n21851_ | ~new_n21850_;
  assign new_n21762_ = ~new_n21853_ | ~new_n21852_;
  assign new_n21763_ = ~pi0348;
  assign new_n21764_ = ~pi0347 | ~new_n21792_;
  assign new_n21765_ = ~new_n21677_;
  assign new_n21766_ = ~new_n21679_;
  assign new_n21767_ = ~new_n21681_;
  assign new_n21768_ = ~new_n21683_;
  assign new_n21769_ = ~new_n21685_;
  assign new_n21770_ = ~new_n21687_;
  assign new_n21771_ = ~new_n21690_;
  assign new_n21772_ = ~new_n21691_;
  assign new_n21773_ = ~new_n21693_;
  assign new_n21774_ = ~new_n21695_;
  assign new_n21775_ = ~new_n21697_;
  assign new_n21776_ = ~new_n21699_;
  assign new_n21777_ = ~new_n21701_;
  assign new_n21778_ = ~new_n21703_;
  assign new_n21779_ = ~new_n21705_;
  assign new_n21780_ = ~new_n21707_;
  assign new_n21781_ = ~new_n21709_;
  assign new_n21782_ = ~new_n21711_;
  assign new_n21783_ = ~new_n21713_;
  assign new_n21784_ = ~new_n21715_;
  assign new_n21785_ = ~new_n21717_;
  assign new_n21786_ = ~new_n21719_;
  assign new_n21787_ = ~new_n21721_;
  assign new_n21788_ = ~new_n21723_;
  assign new_n21789_ = ~new_n21725_;
  assign new_n21790_ = ~new_n21727_;
  assign new_n21791_ = ~new_n21729_;
  assign new_n21792_ = ~new_n21731_;
  assign new_n21793_ = ~new_n21764_;
  assign new_n21794_ = ~pi0326 | ~new_n21690_;
  assign new_n21795_ = ~new_n21771_ | ~new_n21689_;
  assign new_n21796_ = ~pi0325 | ~new_n21687_;
  assign new_n21797_ = ~new_n21770_ | ~new_n21688_;
  assign new_n21798_ = ~pi0324 | ~new_n21685_;
  assign new_n21799_ = ~new_n21769_ | ~new_n21686_;
  assign new_n21800_ = ~pi0323 | ~new_n21683_;
  assign new_n21801_ = ~new_n21768_ | ~new_n21684_;
  assign new_n21802_ = ~pi0322 | ~new_n21681_;
  assign new_n21803_ = ~new_n21767_ | ~new_n21682_;
  assign new_n21804_ = ~pi0321 | ~new_n21679_;
  assign new_n21805_ = ~new_n21766_ | ~new_n21680_;
  assign new_n21806_ = ~pi0320 | ~new_n21677_;
  assign new_n21807_ = ~new_n21765_ | ~new_n21678_;
  assign new_n21808_ = ~pi0348 | ~new_n21764_;
  assign new_n21809_ = ~new_n21793_ | ~new_n21763_;
  assign new_n21810_ = ~pi0347 | ~new_n21731_;
  assign new_n21811_ = ~new_n21792_ | ~new_n21732_;
  assign new_n21812_ = ~pi0319 | ~new_n21675_;
  assign new_n21813_ = ~pi0318 | ~new_n21676_;
  assign new_n21814_ = ~pi0346 | ~new_n21729_;
  assign new_n21815_ = ~new_n21791_ | ~new_n21730_;
  assign new_n21816_ = ~pi0345 | ~new_n21727_;
  assign new_n21817_ = ~new_n21790_ | ~new_n21728_;
  assign new_n21818_ = ~pi0344 | ~new_n21725_;
  assign new_n21819_ = ~new_n21789_ | ~new_n21726_;
  assign new_n21820_ = ~pi0343 | ~new_n21723_;
  assign new_n21821_ = ~new_n21788_ | ~new_n21724_;
  assign new_n21822_ = ~pi0342 | ~new_n21721_;
  assign new_n21823_ = ~new_n21787_ | ~new_n21722_;
  assign new_n21824_ = ~pi0341 | ~new_n21719_;
  assign new_n21825_ = ~new_n21786_ | ~new_n21720_;
  assign new_n21826_ = ~pi0340 | ~new_n21717_;
  assign new_n21827_ = ~new_n21785_ | ~new_n21718_;
  assign new_n21828_ = ~pi0339 | ~new_n21715_;
  assign new_n21829_ = ~new_n21784_ | ~new_n21716_;
  assign new_n21830_ = ~pi0338 | ~new_n21713_;
  assign new_n21831_ = ~new_n21783_ | ~new_n21714_;
  assign new_n21832_ = ~pi0337 | ~new_n21711_;
  assign new_n21833_ = ~new_n21782_ | ~new_n21712_;
  assign new_n21834_ = ~pi0336 | ~new_n21709_;
  assign new_n21835_ = ~new_n21781_ | ~new_n21710_;
  assign new_n21836_ = ~pi0335 | ~new_n21707_;
  assign new_n21837_ = ~new_n21780_ | ~new_n21708_;
  assign new_n21838_ = ~pi0334 | ~new_n21705_;
  assign new_n21839_ = ~new_n21779_ | ~new_n21706_;
  assign new_n21840_ = ~pi0333 | ~new_n21703_;
  assign new_n21841_ = ~new_n21778_ | ~new_n21704_;
  assign new_n21842_ = ~pi0332 | ~new_n21701_;
  assign new_n21843_ = ~new_n21777_ | ~new_n21702_;
  assign new_n21844_ = ~pi0331 | ~new_n21699_;
  assign new_n21845_ = ~new_n21776_ | ~new_n21700_;
  assign new_n21846_ = ~pi0330 | ~new_n21697_;
  assign new_n21847_ = ~new_n21775_ | ~new_n21698_;
  assign new_n21848_ = ~pi0329 | ~new_n21695_;
  assign new_n21849_ = ~new_n21774_ | ~new_n21696_;
  assign new_n21850_ = ~pi0328 | ~new_n21693_;
  assign new_n21851_ = ~new_n21773_ | ~new_n21694_;
  assign new_n21852_ = ~pi0327 | ~new_n21691_;
  assign new_n21853_ = ~new_n21772_ | ~new_n21692_;
  assign new_n21854_ = ~new_n27058_ & ~new_n21856_;
  assign new_n21855_ = new_n27073_ & new_n21857_;
  assign new_n21856_ = ~new_n27072_ & ~new_n21855_ & ~new_n27071_;
  assign new_n21857_ = new_n27059_ | new_n27074_;
  assign new_n21858_ = ~pi0317;
  assign new_n21859_ = ~pi0318;
  assign new_n21860_ = ~pi0318 | ~pi0317;
  assign new_n21861_ = ~pi0319;
  assign new_n21862_ = ~pi0319 | ~new_n21951_;
  assign new_n21863_ = ~pi0320;
  assign new_n21864_ = ~pi0320 | ~new_n21952_;
  assign new_n21865_ = ~pi0321;
  assign new_n21866_ = ~pi0321 | ~new_n21953_;
  assign new_n21867_ = ~pi0322;
  assign new_n21868_ = ~pi0322 | ~new_n21954_;
  assign new_n21869_ = ~pi0323;
  assign new_n21870_ = ~pi0323 | ~new_n21955_;
  assign new_n21871_ = ~pi0324;
  assign new_n21872_ = ~pi0324 | ~new_n21956_;
  assign new_n21873_ = ~pi0325;
  assign new_n21874_ = ~pi0326;
  assign new_n21875_ = ~pi0325 | ~new_n21957_;
  assign new_n21876_ = ~new_n21958_ | ~pi0326;
  assign new_n21877_ = ~pi0327;
  assign new_n21878_ = ~pi0327 | ~new_n21959_;
  assign new_n21879_ = ~pi0328;
  assign new_n21880_ = ~pi0328 | ~new_n21960_;
  assign new_n21881_ = ~pi0329;
  assign new_n21882_ = ~pi0329 | ~new_n21961_;
  assign new_n21883_ = ~pi0330;
  assign new_n21884_ = ~pi0330 | ~new_n21962_;
  assign new_n21885_ = ~pi0331;
  assign new_n21886_ = ~pi0331 | ~new_n21963_;
  assign new_n21887_ = ~pi0332;
  assign new_n21888_ = ~pi0332 | ~new_n21964_;
  assign new_n21889_ = ~pi0333;
  assign new_n21890_ = ~pi0333 | ~new_n21965_;
  assign new_n21891_ = ~pi0334;
  assign new_n21892_ = ~pi0334 | ~new_n21966_;
  assign new_n21893_ = ~pi0335;
  assign new_n21894_ = ~pi0335 | ~new_n21967_;
  assign new_n21895_ = ~pi0336;
  assign new_n21896_ = ~pi0336 | ~new_n21968_;
  assign new_n21897_ = ~pi0337;
  assign new_n21898_ = ~pi0337 | ~new_n21969_;
  assign new_n21899_ = ~pi0338;
  assign new_n21900_ = ~pi0338 | ~new_n21970_;
  assign new_n21901_ = ~pi0339;
  assign new_n21902_ = ~pi0339 | ~new_n21971_;
  assign new_n21903_ = ~pi0340;
  assign new_n21904_ = ~pi0340 | ~new_n21972_;
  assign new_n21905_ = ~pi0341;
  assign new_n21906_ = ~pi0341 | ~new_n21973_;
  assign new_n21907_ = ~pi0342;
  assign new_n21908_ = ~pi0342 | ~new_n21974_;
  assign new_n21909_ = ~pi0343;
  assign new_n21910_ = ~pi0343 | ~new_n21975_;
  assign new_n21911_ = ~pi0344;
  assign new_n21912_ = ~pi0344 | ~new_n21976_;
  assign new_n21913_ = ~pi0345;
  assign new_n21914_ = ~pi0345 | ~new_n21977_;
  assign new_n21915_ = ~pi0346;
  assign new_n21916_ = ~pi0346 | ~new_n21978_;
  assign new_n21917_ = ~pi0347;
  assign new_n21918_ = ~new_n21982_ | ~new_n21981_;
  assign new_n21919_ = ~new_n21984_ | ~new_n21983_;
  assign new_n21920_ = ~new_n21986_ | ~new_n21985_;
  assign new_n21921_ = ~new_n21988_ | ~new_n21987_;
  assign new_n21922_ = ~new_n21990_ | ~new_n21989_;
  assign new_n21923_ = ~new_n21992_ | ~new_n21991_;
  assign new_n21924_ = ~new_n21994_ | ~new_n21993_;
  assign new_n21925_ = ~new_n21996_ | ~new_n21995_;
  assign new_n21926_ = ~new_n21998_ | ~new_n21997_;
  assign new_n21927_ = ~new_n22000_ | ~new_n21999_;
  assign new_n21928_ = ~new_n22002_ | ~new_n22001_;
  assign new_n21929_ = ~new_n22004_ | ~new_n22003_;
  assign new_n21930_ = ~new_n22006_ | ~new_n22005_;
  assign new_n21931_ = ~new_n22008_ | ~new_n22007_;
  assign new_n21932_ = ~new_n22010_ | ~new_n22009_;
  assign new_n21933_ = ~new_n22012_ | ~new_n22011_;
  assign new_n21934_ = ~new_n22014_ | ~new_n22013_;
  assign new_n21935_ = ~new_n22016_ | ~new_n22015_;
  assign new_n21936_ = ~new_n22018_ | ~new_n22017_;
  assign new_n21937_ = ~new_n22020_ | ~new_n22019_;
  assign new_n21938_ = ~new_n22022_ | ~new_n22021_;
  assign new_n21939_ = ~new_n22024_ | ~new_n22023_;
  assign new_n21940_ = ~new_n22026_ | ~new_n22025_;
  assign new_n21941_ = ~new_n22028_ | ~new_n22027_;
  assign new_n21942_ = ~new_n22030_ | ~new_n22029_;
  assign new_n21943_ = ~new_n22032_ | ~new_n22031_;
  assign new_n21944_ = ~new_n22034_ | ~new_n22033_;
  assign new_n21945_ = ~new_n22036_ | ~new_n22035_;
  assign new_n21946_ = ~new_n22038_ | ~new_n22037_;
  assign new_n21947_ = ~new_n22040_ | ~new_n22039_;
  assign new_n21948_ = ~new_n22042_ | ~new_n22041_;
  assign new_n21949_ = ~pi0348;
  assign new_n21950_ = ~pi0347 | ~new_n21979_;
  assign new_n21951_ = ~new_n21860_;
  assign new_n21952_ = ~new_n21862_;
  assign new_n21953_ = ~new_n21864_;
  assign new_n21954_ = ~new_n21866_;
  assign new_n21955_ = ~new_n21868_;
  assign new_n21956_ = ~new_n21870_;
  assign new_n21957_ = ~new_n21872_;
  assign new_n21958_ = ~new_n21875_;
  assign new_n21959_ = ~new_n21876_;
  assign new_n21960_ = ~new_n21878_;
  assign new_n21961_ = ~new_n21880_;
  assign new_n21962_ = ~new_n21882_;
  assign new_n21963_ = ~new_n21884_;
  assign new_n21964_ = ~new_n21886_;
  assign new_n21965_ = ~new_n21888_;
  assign new_n21966_ = ~new_n21890_;
  assign new_n21967_ = ~new_n21892_;
  assign new_n21968_ = ~new_n21894_;
  assign new_n21969_ = ~new_n21896_;
  assign new_n21970_ = ~new_n21898_;
  assign new_n21971_ = ~new_n21900_;
  assign new_n21972_ = ~new_n21902_;
  assign new_n21973_ = ~new_n21904_;
  assign new_n21974_ = ~new_n21906_;
  assign new_n21975_ = ~new_n21908_;
  assign new_n21976_ = ~new_n21910_;
  assign new_n21977_ = ~new_n21912_;
  assign new_n21978_ = ~new_n21914_;
  assign new_n21979_ = ~new_n21916_;
  assign new_n21980_ = ~new_n21950_;
  assign new_n21981_ = ~pi0326 | ~new_n21875_;
  assign new_n21982_ = ~new_n21958_ | ~new_n21874_;
  assign new_n21983_ = ~pi0325 | ~new_n21872_;
  assign new_n21984_ = ~new_n21957_ | ~new_n21873_;
  assign new_n21985_ = ~pi0324 | ~new_n21870_;
  assign new_n21986_ = ~new_n21956_ | ~new_n21871_;
  assign new_n21987_ = ~pi0323 | ~new_n21868_;
  assign new_n21988_ = ~new_n21955_ | ~new_n21869_;
  assign new_n21989_ = ~pi0322 | ~new_n21866_;
  assign new_n21990_ = ~new_n21954_ | ~new_n21867_;
  assign new_n21991_ = ~pi0321 | ~new_n21864_;
  assign new_n21992_ = ~new_n21953_ | ~new_n21865_;
  assign new_n21993_ = ~pi0320 | ~new_n21862_;
  assign new_n21994_ = ~new_n21952_ | ~new_n21863_;
  assign new_n21995_ = ~pi0348 | ~new_n21950_;
  assign new_n21996_ = ~new_n21980_ | ~new_n21949_;
  assign new_n21997_ = ~pi0347 | ~new_n21916_;
  assign new_n21998_ = ~new_n21979_ | ~new_n21917_;
  assign new_n21999_ = ~pi0319 | ~new_n21860_;
  assign new_n22000_ = ~new_n21951_ | ~new_n21861_;
  assign new_n22001_ = ~pi0346 | ~new_n21914_;
  assign new_n22002_ = ~new_n21978_ | ~new_n21915_;
  assign new_n22003_ = ~pi0345 | ~new_n21912_;
  assign new_n22004_ = ~new_n21977_ | ~new_n21913_;
  assign new_n22005_ = ~pi0344 | ~new_n21910_;
  assign new_n22006_ = ~new_n21976_ | ~new_n21911_;
  assign new_n22007_ = ~pi0343 | ~new_n21908_;
  assign new_n22008_ = ~new_n21975_ | ~new_n21909_;
  assign new_n22009_ = ~pi0342 | ~new_n21906_;
  assign new_n22010_ = ~new_n21974_ | ~new_n21907_;
  assign new_n22011_ = ~pi0341 | ~new_n21904_;
  assign new_n22012_ = ~new_n21973_ | ~new_n21905_;
  assign new_n22013_ = ~pi0340 | ~new_n21902_;
  assign new_n22014_ = ~new_n21972_ | ~new_n21903_;
  assign new_n22015_ = ~pi0339 | ~new_n21900_;
  assign new_n22016_ = ~new_n21971_ | ~new_n21901_;
  assign new_n22017_ = ~pi0338 | ~new_n21898_;
  assign new_n22018_ = ~new_n21970_ | ~new_n21899_;
  assign new_n22019_ = ~pi0337 | ~new_n21896_;
  assign new_n22020_ = ~new_n21969_ | ~new_n21897_;
  assign new_n22021_ = ~pi0318 | ~new_n21858_;
  assign new_n22022_ = ~pi0317 | ~new_n21859_;
  assign new_n22023_ = ~pi0336 | ~new_n21894_;
  assign new_n22024_ = ~new_n21968_ | ~new_n21895_;
  assign new_n22025_ = ~pi0335 | ~new_n21892_;
  assign new_n22026_ = ~new_n21967_ | ~new_n21893_;
  assign new_n22027_ = ~pi0334 | ~new_n21890_;
  assign new_n22028_ = ~new_n21966_ | ~new_n21891_;
  assign new_n22029_ = ~pi0333 | ~new_n21888_;
  assign new_n22030_ = ~new_n21965_ | ~new_n21889_;
  assign new_n22031_ = ~pi0332 | ~new_n21886_;
  assign new_n22032_ = ~new_n21964_ | ~new_n21887_;
  assign new_n22033_ = ~pi0331 | ~new_n21884_;
  assign new_n22034_ = ~new_n21963_ | ~new_n21885_;
  assign new_n22035_ = ~pi0330 | ~new_n21882_;
  assign new_n22036_ = ~new_n21962_ | ~new_n21883_;
  assign new_n22037_ = ~pi0329 | ~new_n21880_;
  assign new_n22038_ = ~new_n21961_ | ~new_n21881_;
  assign new_n22039_ = ~pi0328 | ~new_n21878_;
  assign new_n22040_ = ~new_n21960_ | ~new_n21879_;
  assign new_n22041_ = ~pi0327 | ~new_n21876_;
  assign new_n22042_ = ~new_n21959_ | ~new_n21877_;
  assign new_n22043_ = new_n22163_ & new_n22065_;
  assign new_n22044_ = new_n22161_ & new_n22066_;
  assign new_n22045_ = new_n22159_ & new_n22067_;
  assign new_n22046_ = new_n22157_ & new_n22068_;
  assign new_n22047_ = new_n22155_ & new_n22069_;
  assign new_n22048_ = new_n22153_ & new_n22070_;
  assign new_n22049_ = new_n22151_ & new_n22071_;
  assign new_n22050_ = new_n22149_ & new_n22072_;
  assign new_n22051_ = new_n22147_ & new_n22073_;
  assign new_n22052_ = new_n22145_ & new_n22074_;
  assign new_n22053_ = new_n22143_ & new_n22075_;
  assign new_n22054_ = new_n22142_ & new_n22058_;
  assign new_n22055_ = new_n22129_ & new_n22059_;
  assign new_n22056_ = new_n22127_ & new_n22060_;
  assign new_n22057_ = new_n22125_ & new_n22061_;
  assign new_n22058_ = pi0349 | new_n22290_ | new_n22223_;
  assign new_n22059_ = ~new_n22120_ | ~new_n22064_ | ~new_n22095_;
  assign new_n22060_ = ~new_n22121_ | ~new_n22063_ | ~new_n22093_;
  assign new_n22061_ = ~new_n22122_ | ~new_n22062_ | ~new_n22091_;
  assign new_n22062_ = ~new_n22282_;
  assign new_n22063_ = ~new_n22284_;
  assign new_n22064_ = ~new_n22286_;
  assign new_n22065_ = ~new_n22123_ | ~new_n22089_ | ~new_n22086_;
  assign new_n22066_ = ~new_n22130_ | ~new_n22085_ | ~new_n22118_;
  assign new_n22067_ = ~new_n22131_ | ~new_n22084_ | ~new_n22116_;
  assign new_n22068_ = ~new_n22132_ | ~new_n22083_ | ~new_n22114_;
  assign new_n22069_ = ~new_n22133_ | ~new_n22082_ | ~new_n22112_;
  assign new_n22070_ = ~new_n22134_ | ~new_n22081_ | ~new_n22110_;
  assign new_n22071_ = ~new_n22135_ | ~new_n22080_ | ~new_n22106_;
  assign new_n22072_ = ~new_n22136_ | ~new_n22079_ | ~new_n22104_;
  assign new_n22073_ = ~new_n22137_ | ~new_n22078_ | ~new_n22102_;
  assign new_n22074_ = ~new_n22138_ | ~new_n22077_ | ~new_n22100_;
  assign new_n22075_ = ~new_n22139_ | ~new_n22076_;
  assign new_n22076_ = ~new_n22291_;
  assign new_n22077_ = ~new_n22292_;
  assign new_n22078_ = ~new_n22294_;
  assign new_n22079_ = ~new_n22296_;
  assign new_n22080_ = ~new_n22298_;
  assign new_n22081_ = ~new_n22300_;
  assign new_n22082_ = ~new_n22302_;
  assign new_n22083_ = ~new_n22304_;
  assign new_n22084_ = ~new_n22306_;
  assign new_n22085_ = ~new_n22308_;
  assign new_n22086_ = ~new_n22310_;
  assign new_n22087_ = ~new_n22186_ | ~new_n22185_;
  assign new_n22088_ = ~new_n22174_ | ~new_n22173_;
  assign new_n22089_ = ~new_n22281_;
  assign new_n22090_ = new_n22166_ & new_n22165_;
  assign new_n22091_ = ~new_n22283_;
  assign new_n22092_ = new_n22168_ & new_n22167_;
  assign new_n22093_ = ~new_n22285_;
  assign new_n22094_ = new_n22170_ & new_n22169_;
  assign new_n22095_ = ~new_n22287_;
  assign new_n22096_ = new_n22172_ & new_n22171_;
  assign new_n22097_ = ~new_n22288_;
  assign new_n22098_ = ~new_n22289_;
  assign new_n22099_ = new_n22176_ & new_n22175_;
  assign new_n22100_ = ~new_n22293_;
  assign new_n22101_ = new_n22178_ & new_n22177_;
  assign new_n22102_ = ~new_n22295_;
  assign new_n22103_ = new_n22180_ & new_n22179_;
  assign new_n22104_ = ~new_n22297_;
  assign new_n22105_ = new_n22182_ & new_n22181_;
  assign new_n22106_ = ~new_n22299_;
  assign new_n22107_ = new_n22184_ & new_n22183_;
  assign new_n22108_ = ~new_n22223_;
  assign new_n22109_ = ~pi0349;
  assign new_n22110_ = ~new_n22301_;
  assign new_n22111_ = new_n22188_ & new_n22187_;
  assign new_n22112_ = ~new_n22303_;
  assign new_n22113_ = new_n22190_ & new_n22189_;
  assign new_n22114_ = ~new_n22305_;
  assign new_n22115_ = new_n22192_ & new_n22191_;
  assign new_n22116_ = ~new_n22307_;
  assign new_n22117_ = new_n22194_ & new_n22193_;
  assign new_n22118_ = ~new_n22309_;
  assign new_n22119_ = new_n22196_ & new_n22195_;
  assign new_n22120_ = ~new_n22058_;
  assign new_n22121_ = ~new_n22059_;
  assign new_n22122_ = ~new_n22060_;
  assign new_n22123_ = ~new_n22061_;
  assign new_n22124_ = ~new_n22122_ | ~new_n22091_;
  assign new_n22125_ = ~new_n22282_ | ~new_n22124_;
  assign new_n22126_ = ~new_n22121_ | ~new_n22093_;
  assign new_n22127_ = ~new_n22284_ | ~new_n22126_;
  assign new_n22128_ = ~new_n22120_ | ~new_n22095_;
  assign new_n22129_ = ~new_n22286_ | ~new_n22128_;
  assign new_n22130_ = ~new_n22065_;
  assign new_n22131_ = ~new_n22066_;
  assign new_n22132_ = ~new_n22067_;
  assign new_n22133_ = ~new_n22068_;
  assign new_n22134_ = ~new_n22069_;
  assign new_n22135_ = ~new_n22070_;
  assign new_n22136_ = ~new_n22071_;
  assign new_n22137_ = ~new_n22072_;
  assign new_n22138_ = ~new_n22073_;
  assign new_n22139_ = ~new_n22074_;
  assign new_n22140_ = ~new_n22075_;
  assign new_n22141_ = new_n22223_ | pi0349;
  assign new_n22142_ = ~new_n22290_ | ~new_n22141_;
  assign new_n22143_ = ~new_n22291_ | ~new_n22074_;
  assign new_n22144_ = ~new_n22138_ | ~new_n22100_;
  assign new_n22145_ = ~new_n22292_ | ~new_n22144_;
  assign new_n22146_ = ~new_n22137_ | ~new_n22102_;
  assign new_n22147_ = ~new_n22294_ | ~new_n22146_;
  assign new_n22148_ = ~new_n22136_ | ~new_n22104_;
  assign new_n22149_ = ~new_n22296_ | ~new_n22148_;
  assign new_n22150_ = ~new_n22135_ | ~new_n22106_;
  assign new_n22151_ = ~new_n22298_ | ~new_n22150_;
  assign new_n22152_ = ~new_n22134_ | ~new_n22110_;
  assign new_n22153_ = ~new_n22300_ | ~new_n22152_;
  assign new_n22154_ = ~new_n22133_ | ~new_n22112_;
  assign new_n22155_ = ~new_n22302_ | ~new_n22154_;
  assign new_n22156_ = ~new_n22132_ | ~new_n22114_;
  assign new_n22157_ = ~new_n22304_ | ~new_n22156_;
  assign new_n22158_ = ~new_n22131_ | ~new_n22116_;
  assign new_n22159_ = ~new_n22306_ | ~new_n22158_;
  assign new_n22160_ = ~new_n22130_ | ~new_n22118_;
  assign new_n22161_ = ~new_n22308_ | ~new_n22160_;
  assign new_n22162_ = ~new_n22123_ | ~new_n22089_;
  assign new_n22163_ = ~new_n22310_ | ~new_n22162_;
  assign new_n22164_ = ~new_n22140_ | ~new_n22098_;
  assign new_n22165_ = ~new_n22281_ | ~new_n22061_;
  assign new_n22166_ = ~new_n22123_ | ~new_n22089_;
  assign new_n22167_ = ~new_n22283_ | ~new_n22060_;
  assign new_n22168_ = ~new_n22122_ | ~new_n22091_;
  assign new_n22169_ = ~new_n22285_ | ~new_n22059_;
  assign new_n22170_ = ~new_n22121_ | ~new_n22093_;
  assign new_n22171_ = ~new_n22287_ | ~new_n22058_;
  assign new_n22172_ = ~new_n22120_ | ~new_n22095_;
  assign new_n22173_ = ~new_n22164_ | ~new_n22097_;
  assign new_n22174_ = ~new_n22288_ | ~new_n22140_ | ~new_n22098_;
  assign new_n22175_ = ~new_n22289_ | ~new_n22075_;
  assign new_n22176_ = ~new_n22140_ | ~new_n22098_;
  assign new_n22177_ = ~new_n22293_ | ~new_n22073_;
  assign new_n22178_ = ~new_n22138_ | ~new_n22100_;
  assign new_n22179_ = ~new_n22295_ | ~new_n22072_;
  assign new_n22180_ = ~new_n22137_ | ~new_n22102_;
  assign new_n22181_ = ~new_n22297_ | ~new_n22071_;
  assign new_n22182_ = ~new_n22136_ | ~new_n22104_;
  assign new_n22183_ = ~new_n22299_ | ~new_n22070_;
  assign new_n22184_ = ~new_n22135_ | ~new_n22106_;
  assign new_n22185_ = ~new_n22223_ | ~new_n22109_;
  assign new_n22186_ = ~pi0349 | ~new_n22108_;
  assign new_n22187_ = ~new_n22301_ | ~new_n22069_;
  assign new_n22188_ = ~new_n22134_ | ~new_n22110_;
  assign new_n22189_ = ~new_n22303_ | ~new_n22068_;
  assign new_n22190_ = ~new_n22133_ | ~new_n22112_;
  assign new_n22191_ = ~new_n22305_ | ~new_n22067_;
  assign new_n22192_ = ~new_n22132_ | ~new_n22114_;
  assign new_n22193_ = ~new_n22307_ | ~new_n22066_;
  assign new_n22194_ = ~new_n22131_ | ~new_n22116_;
  assign new_n22195_ = ~new_n22309_ | ~new_n22065_;
  assign new_n22196_ = ~new_n22130_ | ~new_n22118_;
  assign new_n22197_ = ~pi0311;
  assign new_n22198_ = pi0307 & new_n22212_;
  assign new_n22199_ = ~pi0310;
  assign new_n22200_ = ~pi0310 | ~pi0311;
  assign new_n22201_ = ~pi0309;
  assign new_n22202_ = ~pi0309 | ~new_n22210_;
  assign new_n22203_ = ~pi0308;
  assign new_n22204_ = ~pi0308 | ~new_n22211_;
  assign new_n22205_ = ~pi0307;
  assign new_n22206_ = ~new_n22214_ | ~new_n22213_;
  assign new_n22207_ = ~new_n22216_ | ~new_n22215_;
  assign new_n22208_ = ~new_n22218_ | ~new_n22217_;
  assign new_n22209_ = ~new_n22220_ | ~new_n22219_;
  assign new_n22210_ = ~new_n22200_;
  assign new_n22211_ = ~new_n22202_;
  assign new_n22212_ = ~new_n22204_;
  assign new_n22213_ = ~pi0307 | ~new_n22204_;
  assign new_n22214_ = ~new_n22212_ | ~new_n22205_;
  assign new_n22215_ = ~pi0308 | ~new_n22202_;
  assign new_n22216_ = ~new_n22211_ | ~new_n22203_;
  assign new_n22217_ = ~pi0309 | ~new_n22200_;
  assign new_n22218_ = ~new_n22210_ | ~new_n22201_;
  assign new_n22219_ = ~pi0310 | ~new_n22197_;
  assign new_n22220_ = ~pi0311 | ~new_n22199_;
  assign new_n22221_ = ~new_n24683_ & ~new_n22222_;
  assign new_n22222_ = ~new_n24694_ & ~new_n24693_ & ~new_n24695_ & ~new_n24696_;
  assign new_n22223_ = ~pi0350;
  assign new_n22224_ = ~pi0351;
  assign new_n22225_ = ~pi0351 | ~pi0350;
  assign new_n22226_ = ~pi0352;
  assign new_n22227_ = ~pi0352 | ~new_n22313_;
  assign new_n22228_ = ~pi0353;
  assign new_n22229_ = ~pi0353 | ~new_n22314_;
  assign new_n22230_ = ~pi0354;
  assign new_n22231_ = ~pi0354 | ~new_n22315_;
  assign new_n22232_ = ~pi0355;
  assign new_n22233_ = ~pi0355 | ~new_n22316_;
  assign new_n22234_ = ~pi0356;
  assign new_n22235_ = ~pi0356 | ~new_n22317_;
  assign new_n22236_ = ~pi0357;
  assign new_n22237_ = ~pi0358;
  assign new_n22238_ = ~pi0357 | ~new_n22318_;
  assign new_n22239_ = ~new_n22319_ | ~pi0358;
  assign new_n22240_ = ~pi0359;
  assign new_n22241_ = ~pi0359 | ~new_n22320_;
  assign new_n22242_ = ~pi0360;
  assign new_n22243_ = ~pi0360 | ~new_n22321_;
  assign new_n22244_ = ~pi0361;
  assign new_n22245_ = ~pi0361 | ~new_n22322_;
  assign new_n22246_ = ~pi0362;
  assign new_n22247_ = ~pi0362 | ~new_n22323_;
  assign new_n22248_ = ~pi0363;
  assign new_n22249_ = ~pi0363 | ~new_n22324_;
  assign new_n22250_ = ~pi0364;
  assign new_n22251_ = ~pi0364 | ~new_n22325_;
  assign new_n22252_ = ~pi0365;
  assign new_n22253_ = ~pi0365 | ~new_n22326_;
  assign new_n22254_ = ~pi0366;
  assign new_n22255_ = ~pi0366 | ~new_n22327_;
  assign new_n22256_ = ~pi0367;
  assign new_n22257_ = ~pi0367 | ~new_n22328_;
  assign new_n22258_ = ~pi0368;
  assign new_n22259_ = ~pi0368 | ~new_n22329_;
  assign new_n22260_ = ~pi0369;
  assign new_n22261_ = ~pi0369 | ~new_n22330_;
  assign new_n22262_ = ~pi0370;
  assign new_n22263_ = ~pi0370 | ~new_n22331_;
  assign new_n22264_ = ~pi0371;
  assign new_n22265_ = ~pi0371 | ~new_n22332_;
  assign new_n22266_ = ~pi0372;
  assign new_n22267_ = ~pi0372 | ~new_n22333_;
  assign new_n22268_ = ~pi0373;
  assign new_n22269_ = ~pi0373 | ~new_n22334_;
  assign new_n22270_ = ~pi0374;
  assign new_n22271_ = ~pi0374 | ~new_n22335_;
  assign new_n22272_ = ~pi0375;
  assign new_n22273_ = ~pi0375 | ~new_n22336_;
  assign new_n22274_ = ~pi0376;
  assign new_n22275_ = ~pi0376 | ~new_n22337_;
  assign new_n22276_ = ~pi0377;
  assign new_n22277_ = ~pi0377 | ~new_n22338_;
  assign new_n22278_ = ~pi0378;
  assign new_n22279_ = ~pi0378 | ~new_n22339_;
  assign new_n22280_ = ~pi0379;
  assign new_n22281_ = ~new_n22343_ | ~new_n22342_;
  assign new_n22282_ = ~new_n22345_ | ~new_n22344_;
  assign new_n22283_ = ~new_n22347_ | ~new_n22346_;
  assign new_n22284_ = ~new_n22349_ | ~new_n22348_;
  assign new_n22285_ = ~new_n22351_ | ~new_n22350_;
  assign new_n22286_ = ~new_n22353_ | ~new_n22352_;
  assign new_n22287_ = ~new_n22355_ | ~new_n22354_;
  assign new_n22288_ = ~new_n22357_ | ~new_n22356_;
  assign new_n22289_ = ~new_n22359_ | ~new_n22358_;
  assign new_n22290_ = ~new_n22361_ | ~new_n22360_;
  assign new_n22291_ = ~new_n22363_ | ~new_n22362_;
  assign new_n22292_ = ~new_n22365_ | ~new_n22364_;
  assign new_n22293_ = ~new_n22367_ | ~new_n22366_;
  assign new_n22294_ = ~new_n22369_ | ~new_n22368_;
  assign new_n22295_ = ~new_n22371_ | ~new_n22370_;
  assign new_n22296_ = ~new_n22373_ | ~new_n22372_;
  assign new_n22297_ = ~new_n22375_ | ~new_n22374_;
  assign new_n22298_ = ~new_n22377_ | ~new_n22376_;
  assign new_n22299_ = ~new_n22379_ | ~new_n22378_;
  assign new_n22300_ = ~new_n22381_ | ~new_n22380_;
  assign new_n22301_ = ~new_n22383_ | ~new_n22382_;
  assign new_n22302_ = ~new_n22385_ | ~new_n22384_;
  assign new_n22303_ = ~new_n22387_ | ~new_n22386_;
  assign new_n22304_ = ~new_n22389_ | ~new_n22388_;
  assign new_n22305_ = ~new_n22391_ | ~new_n22390_;
  assign new_n22306_ = ~new_n22393_ | ~new_n22392_;
  assign new_n22307_ = ~new_n22395_ | ~new_n22394_;
  assign new_n22308_ = ~new_n22397_ | ~new_n22396_;
  assign new_n22309_ = ~new_n22399_ | ~new_n22398_;
  assign new_n22310_ = ~new_n22401_ | ~new_n22400_;
  assign new_n22311_ = ~pi0380;
  assign new_n22312_ = ~pi0379 | ~new_n22340_;
  assign new_n22313_ = ~new_n22225_;
  assign new_n22314_ = ~new_n22227_;
  assign new_n22315_ = ~new_n22229_;
  assign new_n22316_ = ~new_n22231_;
  assign new_n22317_ = ~new_n22233_;
  assign new_n22318_ = ~new_n22235_;
  assign new_n22319_ = ~new_n22238_;
  assign new_n22320_ = ~new_n22239_;
  assign new_n22321_ = ~new_n22241_;
  assign new_n22322_ = ~new_n22243_;
  assign new_n22323_ = ~new_n22245_;
  assign new_n22324_ = ~new_n22247_;
  assign new_n22325_ = ~new_n22249_;
  assign new_n22326_ = ~new_n22251_;
  assign new_n22327_ = ~new_n22253_;
  assign new_n22328_ = ~new_n22255_;
  assign new_n22329_ = ~new_n22257_;
  assign new_n22330_ = ~new_n22259_;
  assign new_n22331_ = ~new_n22261_;
  assign new_n22332_ = ~new_n22263_;
  assign new_n22333_ = ~new_n22265_;
  assign new_n22334_ = ~new_n22267_;
  assign new_n22335_ = ~new_n22269_;
  assign new_n22336_ = ~new_n22271_;
  assign new_n22337_ = ~new_n22273_;
  assign new_n22338_ = ~new_n22275_;
  assign new_n22339_ = ~new_n22277_;
  assign new_n22340_ = ~new_n22279_;
  assign new_n22341_ = ~new_n22312_;
  assign new_n22342_ = ~pi0358 | ~new_n22238_;
  assign new_n22343_ = ~new_n22319_ | ~new_n22237_;
  assign new_n22344_ = ~pi0357 | ~new_n22235_;
  assign new_n22345_ = ~new_n22318_ | ~new_n22236_;
  assign new_n22346_ = ~pi0356 | ~new_n22233_;
  assign new_n22347_ = ~new_n22317_ | ~new_n22234_;
  assign new_n22348_ = ~pi0355 | ~new_n22231_;
  assign new_n22349_ = ~new_n22316_ | ~new_n22232_;
  assign new_n22350_ = ~pi0354 | ~new_n22229_;
  assign new_n22351_ = ~new_n22315_ | ~new_n22230_;
  assign new_n22352_ = ~pi0353 | ~new_n22227_;
  assign new_n22353_ = ~new_n22314_ | ~new_n22228_;
  assign new_n22354_ = ~pi0352 | ~new_n22225_;
  assign new_n22355_ = ~new_n22313_ | ~new_n22226_;
  assign new_n22356_ = ~pi0380 | ~new_n22312_;
  assign new_n22357_ = ~new_n22341_ | ~new_n22311_;
  assign new_n22358_ = ~pi0379 | ~new_n22279_;
  assign new_n22359_ = ~new_n22340_ | ~new_n22280_;
  assign new_n22360_ = ~pi0351 | ~new_n22223_;
  assign new_n22361_ = ~pi0350 | ~new_n22224_;
  assign new_n22362_ = ~pi0378 | ~new_n22277_;
  assign new_n22363_ = ~new_n22339_ | ~new_n22278_;
  assign new_n22364_ = ~pi0377 | ~new_n22275_;
  assign new_n22365_ = ~new_n22338_ | ~new_n22276_;
  assign new_n22366_ = ~pi0376 | ~new_n22273_;
  assign new_n22367_ = ~new_n22337_ | ~new_n22274_;
  assign new_n22368_ = ~pi0375 | ~new_n22271_;
  assign new_n22369_ = ~new_n22336_ | ~new_n22272_;
  assign new_n22370_ = ~pi0374 | ~new_n22269_;
  assign new_n22371_ = ~new_n22335_ | ~new_n22270_;
  assign new_n22372_ = ~pi0373 | ~new_n22267_;
  assign new_n22373_ = ~new_n22334_ | ~new_n22268_;
  assign new_n22374_ = ~pi0372 | ~new_n22265_;
  assign new_n22375_ = ~new_n22333_ | ~new_n22266_;
  assign new_n22376_ = ~pi0371 | ~new_n22263_;
  assign new_n22377_ = ~new_n22332_ | ~new_n22264_;
  assign new_n22378_ = ~pi0370 | ~new_n22261_;
  assign new_n22379_ = ~new_n22331_ | ~new_n22262_;
  assign new_n22380_ = ~pi0369 | ~new_n22259_;
  assign new_n22381_ = ~new_n22330_ | ~new_n22260_;
  assign new_n22382_ = ~pi0368 | ~new_n22257_;
  assign new_n22383_ = ~new_n22329_ | ~new_n22258_;
  assign new_n22384_ = ~pi0367 | ~new_n22255_;
  assign new_n22385_ = ~new_n22328_ | ~new_n22256_;
  assign new_n22386_ = ~pi0366 | ~new_n22253_;
  assign new_n22387_ = ~new_n22327_ | ~new_n22254_;
  assign new_n22388_ = ~pi0365 | ~new_n22251_;
  assign new_n22389_ = ~new_n22326_ | ~new_n22252_;
  assign new_n22390_ = ~pi0364 | ~new_n22249_;
  assign new_n22391_ = ~new_n22325_ | ~new_n22250_;
  assign new_n22392_ = ~pi0363 | ~new_n22247_;
  assign new_n22393_ = ~new_n22324_ | ~new_n22248_;
  assign new_n22394_ = ~pi0362 | ~new_n22245_;
  assign new_n22395_ = ~new_n22323_ | ~new_n22246_;
  assign new_n22396_ = ~pi0361 | ~new_n22243_;
  assign new_n22397_ = ~new_n22322_ | ~new_n22244_;
  assign new_n22398_ = ~pi0360 | ~new_n22241_;
  assign new_n22399_ = ~new_n22321_ | ~new_n22242_;
  assign new_n22400_ = ~pi0359 | ~new_n22239_;
  assign new_n22401_ = ~new_n22320_ | ~new_n22240_;
  assign new_n22402_ = ~new_n22441_ | ~new_n22440_;
  assign new_n22403_ = ~new_n22405_ | ~new_n22442_;
  assign new_n22404_ = ~pi0311;
  assign new_n22405_ = ~pi0311 | ~new_n22414_;
  assign new_n22406_ = ~pi0315;
  assign new_n22407_ = ~pi0309;
  assign new_n22408_ = ~pi0314;
  assign new_n22409_ = ~pi0308;
  assign new_n22410_ = ~pi0313;
  assign new_n22411_ = ~pi0312;
  assign new_n22412_ = ~new_n22437_ | ~new_n22436_;
  assign new_n22413_ = ~pi0307;
  assign new_n22414_ = ~pi0316;
  assign new_n22415_ = ~new_n22447_ | ~new_n22446_;
  assign new_n22416_ = ~new_n22452_ | ~new_n22451_;
  assign new_n22417_ = ~new_n22457_ | ~new_n22456_;
  assign new_n22418_ = ~new_n22462_ | ~new_n22461_;
  assign new_n22419_ = ~new_n22444_ | ~new_n22443_;
  assign new_n22420_ = ~new_n22449_ | ~new_n22448_;
  assign new_n22421_ = ~new_n22454_ | ~new_n22453_;
  assign new_n22422_ = ~new_n22459_ | ~new_n22458_;
  assign new_n22423_ = ~new_n22433_ | ~new_n22432_;
  assign new_n22424_ = ~new_n22429_ | ~new_n22428_;
  assign new_n22425_ = ~pi0310;
  assign new_n22426_ = ~new_n22405_;
  assign new_n22427_ = ~new_n22426_ | ~new_n22406_;
  assign new_n22428_ = ~new_n22427_ | ~new_n22425_;
  assign new_n22429_ = ~pi0315 | ~new_n22405_;
  assign new_n22430_ = ~new_n22424_;
  assign new_n22431_ = ~pi0309 | ~new_n22408_;
  assign new_n22432_ = ~new_n22431_ | ~new_n22424_;
  assign new_n22433_ = ~pi0314 | ~new_n22407_;
  assign new_n22434_ = ~new_n22423_;
  assign new_n22435_ = ~pi0308 | ~new_n22410_;
  assign new_n22436_ = ~new_n22435_ | ~new_n22423_;
  assign new_n22437_ = ~pi0313 | ~new_n22409_;
  assign new_n22438_ = ~new_n22412_;
  assign new_n22439_ = ~pi0312 | ~new_n22413_;
  assign new_n22440_ = ~new_n22438_ | ~new_n22439_;
  assign new_n22441_ = ~pi0307 | ~new_n22411_;
  assign new_n22442_ = ~pi0316 | ~new_n22404_;
  assign new_n22443_ = ~pi0307 | ~new_n22411_;
  assign new_n22444_ = ~pi0312 | ~new_n22413_;
  assign new_n22445_ = ~new_n22419_;
  assign new_n22446_ = ~new_n22445_ | ~new_n22438_;
  assign new_n22447_ = ~new_n22419_ | ~new_n22412_;
  assign new_n22448_ = ~pi0308 | ~new_n22410_;
  assign new_n22449_ = ~pi0313 | ~new_n22409_;
  assign new_n22450_ = ~new_n22420_;
  assign new_n22451_ = ~new_n22434_ | ~new_n22450_;
  assign new_n22452_ = ~new_n22420_ | ~new_n22423_;
  assign new_n22453_ = ~pi0309 | ~new_n22408_;
  assign new_n22454_ = ~pi0314 | ~new_n22407_;
  assign new_n22455_ = ~new_n22421_;
  assign new_n22456_ = ~new_n22430_ | ~new_n22455_;
  assign new_n22457_ = ~new_n22421_ | ~new_n22424_;
  assign new_n22458_ = ~pi0310 | ~new_n22406_;
  assign new_n22459_ = ~pi0315 | ~new_n22425_;
  assign new_n22460_ = ~new_n22422_;
  assign new_n22461_ = ~new_n22460_ | ~new_n22426_;
  assign new_n22462_ = ~new_n22422_ | ~new_n22405_;
  assign new_n22463_ = ~pi0351;
  assign new_n22464_ = ~pi0352;
  assign new_n22465_ = ~pi0352 | ~pi0351;
  assign new_n22466_ = ~pi0353;
  assign new_n22467_ = ~pi0353 | ~new_n22550_;
  assign new_n22468_ = ~pi0354;
  assign new_n22469_ = ~pi0354 | ~new_n22551_;
  assign new_n22470_ = ~pi0355;
  assign new_n22471_ = ~pi0355 | ~new_n22552_;
  assign new_n22472_ = ~pi0356;
  assign new_n22473_ = ~pi0356 | ~new_n22553_;
  assign new_n22474_ = ~pi0357;
  assign new_n22475_ = ~pi0358;
  assign new_n22476_ = ~pi0357 | ~new_n22554_;
  assign new_n22477_ = ~new_n22555_ | ~pi0358;
  assign new_n22478_ = ~pi0359;
  assign new_n22479_ = ~pi0359 | ~new_n22556_;
  assign new_n22480_ = ~pi0360;
  assign new_n22481_ = ~pi0360 | ~new_n22557_;
  assign new_n22482_ = ~pi0361;
  assign new_n22483_ = ~pi0361 | ~new_n22558_;
  assign new_n22484_ = ~pi0362;
  assign new_n22485_ = ~pi0362 | ~new_n22559_;
  assign new_n22486_ = ~pi0363;
  assign new_n22487_ = ~pi0363 | ~new_n22560_;
  assign new_n22488_ = ~pi0364;
  assign new_n22489_ = ~pi0364 | ~new_n22561_;
  assign new_n22490_ = ~pi0365;
  assign new_n22491_ = ~pi0365 | ~new_n22562_;
  assign new_n22492_ = ~pi0366;
  assign new_n22493_ = ~pi0366 | ~new_n22563_;
  assign new_n22494_ = ~pi0367;
  assign new_n22495_ = ~pi0367 | ~new_n22564_;
  assign new_n22496_ = ~pi0368;
  assign new_n22497_ = ~pi0368 | ~new_n22565_;
  assign new_n22498_ = ~pi0369;
  assign new_n22499_ = ~pi0369 | ~new_n22566_;
  assign new_n22500_ = ~pi0370;
  assign new_n22501_ = ~pi0370 | ~new_n22567_;
  assign new_n22502_ = ~pi0371;
  assign new_n22503_ = ~pi0371 | ~new_n22568_;
  assign new_n22504_ = ~pi0372;
  assign new_n22505_ = ~pi0372 | ~new_n22569_;
  assign new_n22506_ = ~pi0373;
  assign new_n22507_ = ~pi0373 | ~new_n22570_;
  assign new_n22508_ = ~pi0374;
  assign new_n22509_ = ~pi0374 | ~new_n22571_;
  assign new_n22510_ = ~pi0375;
  assign new_n22511_ = ~pi0375 | ~new_n22572_;
  assign new_n22512_ = ~pi0376;
  assign new_n22513_ = ~pi0376 | ~new_n22573_;
  assign new_n22514_ = ~pi0377;
  assign new_n22515_ = ~pi0377 | ~new_n22574_;
  assign new_n22516_ = ~pi0378;
  assign new_n22517_ = ~pi0378 | ~new_n22575_;
  assign new_n22518_ = ~pi0379;
  assign new_n22519_ = ~new_n22579_ | ~new_n22578_;
  assign new_n22520_ = ~new_n22581_ | ~new_n22580_;
  assign new_n22521_ = ~new_n22583_ | ~new_n22582_;
  assign new_n22522_ = ~new_n22585_ | ~new_n22584_;
  assign new_n22523_ = ~new_n22587_ | ~new_n22586_;
  assign new_n22524_ = ~new_n22589_ | ~new_n22588_;
  assign new_n22525_ = ~new_n22591_ | ~new_n22590_;
  assign new_n22526_ = ~new_n22593_ | ~new_n22592_;
  assign new_n22527_ = ~new_n22595_ | ~new_n22594_;
  assign new_n22528_ = ~new_n22597_ | ~new_n22596_;
  assign new_n22529_ = ~new_n22599_ | ~new_n22598_;
  assign new_n22530_ = ~new_n22601_ | ~new_n22600_;
  assign new_n22531_ = ~new_n22603_ | ~new_n22602_;
  assign new_n22532_ = ~new_n22605_ | ~new_n22604_;
  assign new_n22533_ = ~new_n22607_ | ~new_n22606_;
  assign new_n22534_ = ~new_n22609_ | ~new_n22608_;
  assign new_n22535_ = ~new_n22611_ | ~new_n22610_;
  assign new_n22536_ = ~new_n22613_ | ~new_n22612_;
  assign new_n22537_ = ~new_n22615_ | ~new_n22614_;
  assign new_n22538_ = ~new_n22617_ | ~new_n22616_;
  assign new_n22539_ = ~new_n22619_ | ~new_n22618_;
  assign new_n22540_ = ~new_n22621_ | ~new_n22620_;
  assign new_n22541_ = ~new_n22623_ | ~new_n22622_;
  assign new_n22542_ = ~new_n22625_ | ~new_n22624_;
  assign new_n22543_ = ~new_n22627_ | ~new_n22626_;
  assign new_n22544_ = ~new_n22629_ | ~new_n22628_;
  assign new_n22545_ = ~new_n22631_ | ~new_n22630_;
  assign new_n22546_ = ~new_n22633_ | ~new_n22632_;
  assign new_n22547_ = ~new_n22635_ | ~new_n22634_;
  assign new_n22548_ = ~pi0380;
  assign new_n22549_ = ~pi0379 | ~new_n22576_;
  assign new_n22550_ = ~new_n22465_;
  assign new_n22551_ = ~new_n22467_;
  assign new_n22552_ = ~new_n22469_;
  assign new_n22553_ = ~new_n22471_;
  assign new_n22554_ = ~new_n22473_;
  assign new_n22555_ = ~new_n22476_;
  assign new_n22556_ = ~new_n22477_;
  assign new_n22557_ = ~new_n22479_;
  assign new_n22558_ = ~new_n22481_;
  assign new_n22559_ = ~new_n22483_;
  assign new_n22560_ = ~new_n22485_;
  assign new_n22561_ = ~new_n22487_;
  assign new_n22562_ = ~new_n22489_;
  assign new_n22563_ = ~new_n22491_;
  assign new_n22564_ = ~new_n22493_;
  assign new_n22565_ = ~new_n22495_;
  assign new_n22566_ = ~new_n22497_;
  assign new_n22567_ = ~new_n22499_;
  assign new_n22568_ = ~new_n22501_;
  assign new_n22569_ = ~new_n22503_;
  assign new_n22570_ = ~new_n22505_;
  assign new_n22571_ = ~new_n22507_;
  assign new_n22572_ = ~new_n22509_;
  assign new_n22573_ = ~new_n22511_;
  assign new_n22574_ = ~new_n22513_;
  assign new_n22575_ = ~new_n22515_;
  assign new_n22576_ = ~new_n22517_;
  assign new_n22577_ = ~new_n22549_;
  assign new_n22578_ = ~pi0358 | ~new_n22476_;
  assign new_n22579_ = ~new_n22555_ | ~new_n22475_;
  assign new_n22580_ = ~pi0357 | ~new_n22473_;
  assign new_n22581_ = ~new_n22554_ | ~new_n22474_;
  assign new_n22582_ = ~pi0356 | ~new_n22471_;
  assign new_n22583_ = ~new_n22553_ | ~new_n22472_;
  assign new_n22584_ = ~pi0355 | ~new_n22469_;
  assign new_n22585_ = ~new_n22552_ | ~new_n22470_;
  assign new_n22586_ = ~pi0354 | ~new_n22467_;
  assign new_n22587_ = ~new_n22551_ | ~new_n22468_;
  assign new_n22588_ = ~pi0353 | ~new_n22465_;
  assign new_n22589_ = ~new_n22550_ | ~new_n22466_;
  assign new_n22590_ = ~pi0352 | ~new_n22463_;
  assign new_n22591_ = ~pi0351 | ~new_n22464_;
  assign new_n22592_ = ~pi0380 | ~new_n22549_;
  assign new_n22593_ = ~new_n22577_ | ~new_n22548_;
  assign new_n22594_ = ~pi0379 | ~new_n22517_;
  assign new_n22595_ = ~new_n22576_ | ~new_n22518_;
  assign new_n22596_ = ~pi0378 | ~new_n22515_;
  assign new_n22597_ = ~new_n22575_ | ~new_n22516_;
  assign new_n22598_ = ~pi0377 | ~new_n22513_;
  assign new_n22599_ = ~new_n22574_ | ~new_n22514_;
  assign new_n22600_ = ~pi0376 | ~new_n22511_;
  assign new_n22601_ = ~new_n22573_ | ~new_n22512_;
  assign new_n22602_ = ~pi0375 | ~new_n22509_;
  assign new_n22603_ = ~new_n22572_ | ~new_n22510_;
  assign new_n22604_ = ~pi0374 | ~new_n22507_;
  assign new_n22605_ = ~new_n22571_ | ~new_n22508_;
  assign new_n22606_ = ~pi0373 | ~new_n22505_;
  assign new_n22607_ = ~new_n22570_ | ~new_n22506_;
  assign new_n22608_ = ~pi0372 | ~new_n22503_;
  assign new_n22609_ = ~new_n22569_ | ~new_n22504_;
  assign new_n22610_ = ~pi0371 | ~new_n22501_;
  assign new_n22611_ = ~new_n22568_ | ~new_n22502_;
  assign new_n22612_ = ~pi0370 | ~new_n22499_;
  assign new_n22613_ = ~new_n22567_ | ~new_n22500_;
  assign new_n22614_ = ~pi0369 | ~new_n22497_;
  assign new_n22615_ = ~new_n22566_ | ~new_n22498_;
  assign new_n22616_ = ~pi0368 | ~new_n22495_;
  assign new_n22617_ = ~new_n22565_ | ~new_n22496_;
  assign new_n22618_ = ~pi0367 | ~new_n22493_;
  assign new_n22619_ = ~new_n22564_ | ~new_n22494_;
  assign new_n22620_ = ~pi0366 | ~new_n22491_;
  assign new_n22621_ = ~new_n22563_ | ~new_n22492_;
  assign new_n22622_ = ~pi0365 | ~new_n22489_;
  assign new_n22623_ = ~new_n22562_ | ~new_n22490_;
  assign new_n22624_ = ~pi0364 | ~new_n22487_;
  assign new_n22625_ = ~new_n22561_ | ~new_n22488_;
  assign new_n22626_ = ~pi0363 | ~new_n22485_;
  assign new_n22627_ = ~new_n22560_ | ~new_n22486_;
  assign new_n22628_ = ~pi0362 | ~new_n22483_;
  assign new_n22629_ = ~new_n22559_ | ~new_n22484_;
  assign new_n22630_ = ~pi0361 | ~new_n22481_;
  assign new_n22631_ = ~new_n22558_ | ~new_n22482_;
  assign new_n22632_ = ~pi0360 | ~new_n22479_;
  assign new_n22633_ = ~new_n22557_ | ~new_n22480_;
  assign new_n22634_ = ~pi0359 | ~new_n22477_;
  assign new_n22635_ = ~new_n22556_ | ~new_n22478_;
  assign new_n22636_ = ~new_n24059_ & ~new_n22638_;
  assign new_n22637_ = new_n24060_ & new_n24075_;
  assign new_n22638_ = ~new_n24073_ & ~new_n24072_ & ~new_n24074_ & ~new_n22637_;
  assign new_n22639_ = new_n22821_ & new_n22680_;
  assign new_n22640_ = new_n22819_ & new_n22681_;
  assign new_n22641_ = new_n22817_ & new_n22711_;
  assign new_n22642_ = new_n22816_ & new_n22685_;
  assign new_n22643_ = new_n22814_ & new_n22688_;
  assign new_n22644_ = new_n22812_ & new_n22691_;
  assign new_n22645_ = new_n22810_ & new_n22693_;
  assign new_n22646_ = new_n22809_ & new_n22695_;
  assign new_n22647_ = new_n22808_ & new_n22698_;
  assign new_n22648_ = new_n22806_ & new_n22701_;
  assign new_n22649_ = new_n22804_ & new_n22703_;
  assign new_n22650_ = new_n22803_ & new_n22706_;
  assign new_n22651_ = new_n22801_ & new_n22708_;
  assign new_n22652_ = new_n22788_ & new_n22787_;
  assign new_n22653_ = new_n22786_ & new_n22784_;
  assign new_n22654_ = ~new_n22827_ | ~new_n22883_ | ~new_n22882_;
  assign new_n22655_ = ~new_n23849_;
  assign new_n22656_ = ~pi0321;
  assign new_n22657_ = ~new_n23850_;
  assign new_n22658_ = ~pi0320;
  assign new_n22659_ = ~new_n3777_;
  assign new_n22660_ = ~pi0317;
  assign new_n22661_ = ~pi0318;
  assign new_n22662_ = ~pi0317 | ~new_n3777_;
  assign new_n22663_ = ~new_n23834_;
  assign new_n22664_ = ~new_n23851_;
  assign new_n22665_ = ~pi0319;
  assign new_n22666_ = ~pi0322;
  assign new_n22667_ = ~new_n23848_;
  assign new_n22668_ = ~new_n23847_;
  assign new_n22669_ = ~pi0323;
  assign new_n22670_ = ~pi0324;
  assign new_n22671_ = ~new_n23846_;
  assign new_n22672_ = ~new_n23835_;
  assign new_n22673_ = ~pi0325;
  assign new_n22674_ = ~pi0326;
  assign new_n22675_ = ~new_n22766_ | ~new_n22765_;
  assign new_n22676_ = ~new_n22675_ | ~new_n22768_;
  assign new_n22677_ = ~pi0327;
  assign new_n22678_ = ~pi0328;
  assign new_n22679_ = ~pi0329;
  assign new_n22680_ = ~new_n22732_ | ~new_n22740_;
  assign new_n22681_ = ~new_n22733_ | ~new_n22754_;
  assign new_n22682_ = ~pi0330;
  assign new_n22683_ = ~pi0332;
  assign new_n22684_ = ~pi0331;
  assign new_n22685_ = ~new_n22789_ | ~new_n22734_;
  assign new_n22686_ = ~pi0334;
  assign new_n22687_ = ~pi0333;
  assign new_n22688_ = ~new_n22735_ | ~new_n22791_;
  assign new_n22689_ = ~pi0335;
  assign new_n22690_ = ~pi0336;
  assign new_n22691_ = ~new_n22736_ | ~new_n22792_;
  assign new_n22692_ = ~pi0337;
  assign new_n22693_ = ~pi0337 | ~new_n22793_;
  assign new_n22694_ = ~pi0338;
  assign new_n22695_ = ~pi0338 | ~new_n22794_;
  assign new_n22696_ = ~pi0340;
  assign new_n22697_ = ~pi0339;
  assign new_n22698_ = ~new_n22737_ | ~new_n22795_;
  assign new_n22699_ = ~pi0342;
  assign new_n22700_ = ~pi0341;
  assign new_n22701_ = ~new_n22738_ | ~new_n22796_;
  assign new_n22702_ = ~pi0343;
  assign new_n22703_ = ~pi0343 | ~new_n22797_;
  assign new_n22704_ = ~pi0345;
  assign new_n22705_ = ~pi0344;
  assign new_n22706_ = ~new_n22739_ | ~new_n22798_;
  assign new_n22707_ = ~pi0346;
  assign new_n22708_ = ~pi0346 | ~new_n22799_;
  assign new_n22709_ = ~pi0347;
  assign new_n22710_ = ~new_n23834_ | ~new_n22759_;
  assign new_n22711_ = ~pi0330 | ~new_n22789_;
  assign new_n22712_ = ~new_n22865_ | ~new_n22864_;
  assign new_n22713_ = ~new_n22874_ | ~new_n22873_;
  assign new_n22714_ = ~new_n22876_ | ~new_n22875_;
  assign new_n22715_ = ~new_n22878_ | ~new_n22877_;
  assign new_n22716_ = ~new_n22885_ | ~new_n22884_;
  assign new_n22717_ = ~new_n22887_ | ~new_n22886_;
  assign new_n22718_ = ~new_n22889_ | ~new_n22888_;
  assign new_n22719_ = ~new_n22891_ | ~new_n22890_;
  assign new_n22720_ = ~new_n22893_ | ~new_n22892_;
  assign new_n22721_ = ~new_n22836_ | ~new_n22835_;
  assign new_n22722_ = ~new_n22843_ | ~new_n22842_;
  assign new_n22723_ = ~new_n22850_ | ~new_n22849_;
  assign new_n22724_ = ~new_n22857_ | ~new_n22856_;
  assign new_n22725_ = ~new_n22863_ | ~new_n22862_;
  assign new_n22726_ = ~new_n22872_ | ~new_n22871_;
  assign new_n22727_ = new_n23850_ & pi0320;
  assign new_n22728_ = new_n22768_ & new_n22758_;
  assign new_n22729_ = new_n22825_ & new_n22760_;
  assign new_n22730_ = new_n22770_ & new_n22859_ & new_n22858_;
  assign new_n22731_ = new_n22760_ & new_n22758_;
  assign new_n22732_ = pi0326 & pi0327;
  assign new_n22733_ = pi0329 & pi0328;
  assign new_n22734_ = pi0330 & pi0331 & pi0332;
  assign new_n22735_ = pi0334 & pi0333;
  assign new_n22736_ = pi0335 & pi0336;
  assign new_n22737_ = pi0340 & pi0339;
  assign new_n22738_ = pi0342 & pi0341;
  assign new_n22739_ = pi0345 & pi0344;
  assign new_n22740_ = ~new_n22782_ | ~new_n22781_;
  assign new_n22741_ = new_n22829_ & new_n22828_;
  assign new_n22742_ = new_n22831_ & new_n22830_;
  assign new_n22743_ = ~new_n22824_ | ~new_n22778_ | ~new_n22755_;
  assign new_n22744_ = new_n22838_ & new_n22837_;
  assign new_n22745_ = ~new_n22776_ | ~new_n22775_;
  assign new_n22746_ = new_n22845_ & new_n22844_;
  assign new_n22747_ = ~new_n22823_ | ~new_n22772_ | ~new_n22756_;
  assign new_n22748_ = new_n22852_ & new_n22851_;
  assign new_n22749_ = ~new_n22729_ | ~new_n22826_;
  assign new_n22750_ = new_n22861_ & new_n22860_;
  assign new_n22751_ = ~pi0348;
  assign new_n22752_ = new_n22867_ & new_n22866_;
  assign new_n22753_ = ~new_n22710_ | ~new_n22762_;
  assign new_n22754_ = ~new_n22680_;
  assign new_n22755_ = ~pi0324 | ~new_n22745_;
  assign new_n22756_ = ~pi0322 | ~new_n22749_;
  assign new_n22757_ = ~new_n22710_;
  assign new_n22758_ = pi0321 | new_n23849_;
  assign new_n22759_ = ~new_n22662_;
  assign new_n22760_ = ~pi0321 | ~new_n23849_;
  assign new_n22761_ = ~new_n22663_ | ~new_n22662_;
  assign new_n22762_ = ~pi0318 | ~new_n22761_;
  assign new_n22763_ = ~new_n22753_;
  assign new_n22764_ = new_n23851_ | pi0319;
  assign new_n22765_ = ~new_n22764_ | ~new_n22753_;
  assign new_n22766_ = ~pi0319 | ~new_n23851_;
  assign new_n22767_ = ~new_n22675_;
  assign new_n22768_ = pi0320 | new_n23850_;
  assign new_n22769_ = ~new_n22676_;
  assign new_n22770_ = ~pi0320 | ~new_n23850_;
  assign new_n22771_ = ~new_n22749_;
  assign new_n22772_ = ~new_n23848_ | ~new_n22749_;
  assign new_n22773_ = ~new_n22747_;
  assign new_n22774_ = new_n23847_ | pi0323;
  assign new_n22775_ = ~new_n22774_ | ~new_n22747_;
  assign new_n22776_ = ~pi0323 | ~new_n23847_;
  assign new_n22777_ = ~new_n22745_;
  assign new_n22778_ = ~new_n23846_ | ~new_n22745_;
  assign new_n22779_ = ~new_n22743_;
  assign new_n22780_ = new_n23835_ | pi0325;
  assign new_n22781_ = ~new_n22780_ | ~new_n22743_;
  assign new_n22782_ = ~pi0325 | ~new_n23835_;
  assign new_n22783_ = ~new_n22740_;
  assign new_n22784_ = ~new_n22730_ | ~new_n22676_;
  assign new_n22785_ = ~new_n22770_ | ~new_n22676_;
  assign new_n22786_ = ~new_n22731_ | ~new_n22785_;
  assign new_n22787_ = ~new_n22750_ | ~new_n22767_;
  assign new_n22788_ = ~new_n22769_ | ~new_n22770_;
  assign new_n22789_ = ~new_n22681_;
  assign new_n22790_ = ~new_n22711_;
  assign new_n22791_ = ~new_n22685_;
  assign new_n22792_ = ~new_n22688_;
  assign new_n22793_ = ~new_n22691_;
  assign new_n22794_ = ~new_n22693_;
  assign new_n22795_ = ~new_n22695_;
  assign new_n22796_ = ~new_n22698_;
  assign new_n22797_ = ~new_n22701_;
  assign new_n22798_ = ~new_n22703_;
  assign new_n22799_ = ~new_n22706_;
  assign new_n22800_ = ~new_n22708_;
  assign new_n22801_ = ~new_n22707_ | ~new_n22706_;
  assign new_n22802_ = ~pi0344 | ~new_n22798_;
  assign new_n22803_ = ~new_n22704_ | ~new_n22802_;
  assign new_n22804_ = ~new_n22702_ | ~new_n22701_;
  assign new_n22805_ = ~pi0341 | ~new_n22796_;
  assign new_n22806_ = ~new_n22699_ | ~new_n22805_;
  assign new_n22807_ = ~pi0339 | ~new_n22795_;
  assign new_n22808_ = ~new_n22696_ | ~new_n22807_;
  assign new_n22809_ = ~new_n22694_ | ~new_n22693_;
  assign new_n22810_ = ~new_n22692_ | ~new_n22691_;
  assign new_n22811_ = ~pi0335 | ~new_n22792_;
  assign new_n22812_ = ~new_n22690_ | ~new_n22811_;
  assign new_n22813_ = ~pi0333 | ~new_n22791_;
  assign new_n22814_ = ~new_n22686_ | ~new_n22813_;
  assign new_n22815_ = ~new_n22790_ | ~pi0331;
  assign new_n22816_ = ~new_n22683_ | ~new_n22815_;
  assign new_n22817_ = ~new_n22682_ | ~new_n22681_;
  assign new_n22818_ = ~new_n22754_ | ~pi0328;
  assign new_n22819_ = ~new_n22679_ | ~new_n22818_;
  assign new_n22820_ = ~pi0326 | ~new_n22740_;
  assign new_n22821_ = ~new_n22677_ | ~new_n22820_;
  assign new_n22822_ = ~pi0347 | ~new_n22800_;
  assign new_n22823_ = ~new_n23848_ | ~pi0322;
  assign new_n22824_ = ~new_n23846_ | ~pi0324;
  assign new_n22825_ = ~new_n22727_ | ~new_n22758_;
  assign new_n22826_ = ~new_n22728_ | ~new_n22675_;
  assign new_n22827_ = ~new_n22757_ | ~pi0318;
  assign new_n22828_ = ~pi0326 | ~new_n22740_;
  assign new_n22829_ = ~new_n22783_ | ~new_n22674_;
  assign new_n22830_ = ~pi0325 | ~new_n22672_;
  assign new_n22831_ = ~new_n23835_ | ~new_n22673_;
  assign new_n22832_ = ~pi0325 | ~new_n22672_;
  assign new_n22833_ = ~new_n23835_ | ~new_n22673_;
  assign new_n22834_ = ~new_n22833_ | ~new_n22832_;
  assign new_n22835_ = ~new_n22742_ | ~new_n22743_;
  assign new_n22836_ = ~new_n22779_ | ~new_n22834_;
  assign new_n22837_ = ~pi0324 | ~new_n22671_;
  assign new_n22838_ = ~new_n23846_ | ~new_n22670_;
  assign new_n22839_ = ~pi0324 | ~new_n22671_;
  assign new_n22840_ = ~new_n23846_ | ~new_n22670_;
  assign new_n22841_ = ~new_n22840_ | ~new_n22839_;
  assign new_n22842_ = ~new_n22744_ | ~new_n22745_;
  assign new_n22843_ = ~new_n22777_ | ~new_n22841_;
  assign new_n22844_ = ~pi0323 | ~new_n22668_;
  assign new_n22845_ = ~new_n23847_ | ~new_n22669_;
  assign new_n22846_ = ~pi0323 | ~new_n22668_;
  assign new_n22847_ = ~new_n23847_ | ~new_n22669_;
  assign new_n22848_ = ~new_n22847_ | ~new_n22846_;
  assign new_n22849_ = ~new_n22746_ | ~new_n22747_;
  assign new_n22850_ = ~new_n22773_ | ~new_n22848_;
  assign new_n22851_ = ~pi0322 | ~new_n22667_;
  assign new_n22852_ = ~new_n23848_ | ~new_n22666_;
  assign new_n22853_ = ~pi0322 | ~new_n22667_;
  assign new_n22854_ = ~new_n23848_ | ~new_n22666_;
  assign new_n22855_ = ~new_n22854_ | ~new_n22853_;
  assign new_n22856_ = ~new_n22748_ | ~new_n22749_;
  assign new_n22857_ = ~new_n22771_ | ~new_n22855_;
  assign new_n22858_ = ~pi0321 | ~new_n22655_;
  assign new_n22859_ = ~new_n23849_ | ~new_n22656_;
  assign new_n22860_ = ~pi0320 | ~new_n22657_;
  assign new_n22861_ = ~new_n23850_ | ~new_n22658_;
  assign new_n22862_ = ~pi0348 | ~new_n22822_;
  assign new_n22863_ = ~new_n22751_ | ~pi0347 | ~new_n22800_;
  assign new_n22864_ = ~pi0347 | ~new_n22708_;
  assign new_n22865_ = ~new_n22800_ | ~new_n22709_;
  assign new_n22866_ = ~pi0319 | ~new_n22664_;
  assign new_n22867_ = ~new_n23851_ | ~new_n22665_;
  assign new_n22868_ = ~pi0319 | ~new_n22664_;
  assign new_n22869_ = ~new_n23851_ | ~new_n22665_;
  assign new_n22870_ = ~new_n22869_ | ~new_n22868_;
  assign new_n22871_ = ~new_n22752_ | ~new_n22753_;
  assign new_n22872_ = ~new_n22763_ | ~new_n22870_;
  assign new_n22873_ = ~pi0344 | ~new_n22703_;
  assign new_n22874_ = ~new_n22798_ | ~new_n22705_;
  assign new_n22875_ = ~pi0341 | ~new_n22698_;
  assign new_n22876_ = ~new_n22796_ | ~new_n22700_;
  assign new_n22877_ = ~pi0339 | ~new_n22695_;
  assign new_n22878_ = ~new_n22795_ | ~new_n22697_;
  assign new_n22879_ = ~pi0318 | ~new_n22662_;
  assign new_n22880_ = ~new_n22759_ | ~new_n22661_;
  assign new_n22881_ = ~new_n22880_ | ~new_n22879_;
  assign new_n22882_ = ~new_n23834_ | ~new_n22662_ | ~new_n22661_;
  assign new_n22883_ = ~new_n22881_ | ~new_n22663_;
  assign new_n22884_ = ~pi0335 | ~new_n22688_;
  assign new_n22885_ = ~new_n22792_ | ~new_n22689_;
  assign new_n22886_ = ~pi0333 | ~new_n22685_;
  assign new_n22887_ = ~new_n22791_ | ~new_n22687_;
  assign new_n22888_ = ~pi0331 | ~new_n22711_;
  assign new_n22889_ = ~new_n22790_ | ~new_n22684_;
  assign new_n22890_ = ~new_n22754_ | ~new_n22678_;
  assign new_n22891_ = ~pi0328 | ~new_n22680_;
  assign new_n22892_ = ~pi0317 | ~new_n22659_;
  assign new_n22893_ = ~new_n3777_ | ~new_n22660_;
  assign new_n22894_ = new_n22895_ | new_n4460_;
  assign new_n22895_ = ~new_n24742_ & ~new_n24741_;
  assign new_n22896_ = ~new_n4457_;
  assign new_n22897_ = ~new_n4458_;
  assign new_n22898_ = ~new_n3788_;
  assign new_n22899_ = ~new_n4456_;
  assign new_n22900_ = ~pi0509;
  assign new_n22901_ = ~pi0510;
  assign new_n22902_ = ~pi0510 | ~pi0509;
  assign new_n22903_ = ~pi0511;
  assign new_n22904_ = ~pi0511 | ~new_n22990_;
  assign new_n22905_ = ~pi0512;
  assign new_n22906_ = ~pi0512 | ~new_n22991_;
  assign new_n22907_ = ~pi0513;
  assign new_n22908_ = ~pi0513 | ~new_n22992_;
  assign new_n22909_ = ~pi0514;
  assign new_n22910_ = ~pi0514 | ~new_n22993_;
  assign new_n22911_ = ~pi0515;
  assign new_n22912_ = ~pi0515 | ~new_n22994_;
  assign new_n22913_ = ~pi0516;
  assign new_n22914_ = ~pi0517;
  assign new_n22915_ = ~pi0516 | ~new_n22995_;
  assign new_n22916_ = ~new_n22996_ | ~pi0517;
  assign new_n22917_ = ~pi0518;
  assign new_n22918_ = ~pi0518 | ~new_n22997_;
  assign new_n22919_ = ~pi0519;
  assign new_n22920_ = ~pi0519 | ~new_n22998_;
  assign new_n22921_ = ~pi0520;
  assign new_n22922_ = ~pi0520 | ~new_n22999_;
  assign new_n22923_ = ~pi0521;
  assign new_n22924_ = ~pi0521 | ~new_n23000_;
  assign new_n22925_ = ~pi0522;
  assign new_n22926_ = ~pi0522 | ~new_n23001_;
  assign new_n22927_ = ~pi0523;
  assign new_n22928_ = ~pi0523 | ~new_n23002_;
  assign new_n22929_ = ~pi0524;
  assign new_n22930_ = ~pi0524 | ~new_n23003_;
  assign new_n22931_ = ~pi0525;
  assign new_n22932_ = ~pi0525 | ~new_n23004_;
  assign new_n22933_ = ~pi0526;
  assign new_n22934_ = ~pi0526 | ~new_n23005_;
  assign new_n22935_ = ~pi0527;
  assign new_n22936_ = ~pi0527 | ~new_n23006_;
  assign new_n22937_ = ~pi0528;
  assign new_n22938_ = ~pi0528 | ~new_n23007_;
  assign new_n22939_ = ~pi0529;
  assign new_n22940_ = ~pi0529 | ~new_n23008_;
  assign new_n22941_ = ~pi0530;
  assign new_n22942_ = ~pi0530 | ~new_n23009_;
  assign new_n22943_ = ~pi0531;
  assign new_n22944_ = ~pi0531 | ~new_n23010_;
  assign new_n22945_ = ~pi0532;
  assign new_n22946_ = ~pi0532 | ~new_n23011_;
  assign new_n22947_ = ~pi0533;
  assign new_n22948_ = ~pi0533 | ~new_n23012_;
  assign new_n22949_ = ~pi0534;
  assign new_n22950_ = ~pi0534 | ~new_n23013_;
  assign new_n22951_ = ~pi0535;
  assign new_n22952_ = ~pi0535 | ~new_n23014_;
  assign new_n22953_ = ~pi0536;
  assign new_n22954_ = ~pi0536 | ~new_n23015_;
  assign new_n22955_ = ~pi0537;
  assign new_n22956_ = ~pi0537 | ~new_n23016_;
  assign new_n22957_ = ~pi0538;
  assign new_n22958_ = ~new_n23020_ | ~new_n23019_;
  assign new_n22959_ = ~new_n23022_ | ~new_n23021_;
  assign new_n22960_ = ~new_n23024_ | ~new_n23023_;
  assign new_n22961_ = ~new_n23026_ | ~new_n23025_;
  assign new_n22962_ = ~new_n23028_ | ~new_n23027_;
  assign new_n22963_ = ~new_n23030_ | ~new_n23029_;
  assign new_n22964_ = ~new_n23032_ | ~new_n23031_;
  assign new_n22965_ = ~new_n23034_ | ~new_n23033_;
  assign new_n22966_ = ~new_n23036_ | ~new_n23035_;
  assign new_n22967_ = ~new_n23038_ | ~new_n23037_;
  assign new_n22968_ = ~new_n23040_ | ~new_n23039_;
  assign new_n22969_ = ~new_n23042_ | ~new_n23041_;
  assign new_n22970_ = ~new_n23044_ | ~new_n23043_;
  assign new_n22971_ = ~new_n23046_ | ~new_n23045_;
  assign new_n22972_ = ~new_n23048_ | ~new_n23047_;
  assign new_n22973_ = ~new_n23050_ | ~new_n23049_;
  assign new_n22974_ = ~new_n23052_ | ~new_n23051_;
  assign new_n22975_ = ~new_n23054_ | ~new_n23053_;
  assign new_n22976_ = ~new_n23056_ | ~new_n23055_;
  assign new_n22977_ = ~new_n23058_ | ~new_n23057_;
  assign new_n22978_ = ~new_n23060_ | ~new_n23059_;
  assign new_n22979_ = ~new_n23062_ | ~new_n23061_;
  assign new_n22980_ = ~new_n23064_ | ~new_n23063_;
  assign new_n22981_ = ~new_n23066_ | ~new_n23065_;
  assign new_n22982_ = ~new_n23068_ | ~new_n23067_;
  assign new_n22983_ = ~new_n23070_ | ~new_n23069_;
  assign new_n22984_ = ~new_n23072_ | ~new_n23071_;
  assign new_n22985_ = ~new_n23074_ | ~new_n23073_;
  assign new_n22986_ = ~new_n23076_ | ~new_n23075_;
  assign new_n22987_ = ~new_n23078_ | ~new_n23077_;
  assign new_n22988_ = ~pi0539;
  assign new_n22989_ = ~pi0538 | ~new_n23017_;
  assign new_n22990_ = ~new_n22902_;
  assign new_n22991_ = ~new_n22904_;
  assign new_n22992_ = ~new_n22906_;
  assign new_n22993_ = ~new_n22908_;
  assign new_n22994_ = ~new_n22910_;
  assign new_n22995_ = ~new_n22912_;
  assign new_n22996_ = ~new_n22915_;
  assign new_n22997_ = ~new_n22916_;
  assign new_n22998_ = ~new_n22918_;
  assign new_n22999_ = ~new_n22920_;
  assign new_n23000_ = ~new_n22922_;
  assign new_n23001_ = ~new_n22924_;
  assign new_n23002_ = ~new_n22926_;
  assign new_n23003_ = ~new_n22928_;
  assign new_n23004_ = ~new_n22930_;
  assign new_n23005_ = ~new_n22932_;
  assign new_n23006_ = ~new_n22934_;
  assign new_n23007_ = ~new_n22936_;
  assign new_n23008_ = ~new_n22938_;
  assign new_n23009_ = ~new_n22940_;
  assign new_n23010_ = ~new_n22942_;
  assign new_n23011_ = ~new_n22944_;
  assign new_n23012_ = ~new_n22946_;
  assign new_n23013_ = ~new_n22948_;
  assign new_n23014_ = ~new_n22950_;
  assign new_n23015_ = ~new_n22952_;
  assign new_n23016_ = ~new_n22954_;
  assign new_n23017_ = ~new_n22956_;
  assign new_n23018_ = ~new_n22989_;
  assign new_n23019_ = ~pi0517 | ~new_n22915_;
  assign new_n23020_ = ~new_n22996_ | ~new_n22914_;
  assign new_n23021_ = ~pi0516 | ~new_n22912_;
  assign new_n23022_ = ~new_n22995_ | ~new_n22913_;
  assign new_n23023_ = ~pi0515 | ~new_n22910_;
  assign new_n23024_ = ~new_n22994_ | ~new_n22911_;
  assign new_n23025_ = ~pi0514 | ~new_n22908_;
  assign new_n23026_ = ~new_n22993_ | ~new_n22909_;
  assign new_n23027_ = ~pi0513 | ~new_n22906_;
  assign new_n23028_ = ~new_n22992_ | ~new_n22907_;
  assign new_n23029_ = ~pi0512 | ~new_n22904_;
  assign new_n23030_ = ~new_n22991_ | ~new_n22905_;
  assign new_n23031_ = ~pi0511 | ~new_n22902_;
  assign new_n23032_ = ~new_n22990_ | ~new_n22903_;
  assign new_n23033_ = ~pi0539 | ~new_n22989_;
  assign new_n23034_ = ~new_n23018_ | ~new_n22988_;
  assign new_n23035_ = ~pi0538 | ~new_n22956_;
  assign new_n23036_ = ~new_n23017_ | ~new_n22957_;
  assign new_n23037_ = ~pi0510 | ~new_n22900_;
  assign new_n23038_ = ~pi0509 | ~new_n22901_;
  assign new_n23039_ = ~pi0537 | ~new_n22954_;
  assign new_n23040_ = ~new_n23016_ | ~new_n22955_;
  assign new_n23041_ = ~pi0536 | ~new_n22952_;
  assign new_n23042_ = ~new_n23015_ | ~new_n22953_;
  assign new_n23043_ = ~pi0535 | ~new_n22950_;
  assign new_n23044_ = ~new_n23014_ | ~new_n22951_;
  assign new_n23045_ = ~pi0534 | ~new_n22948_;
  assign new_n23046_ = ~new_n23013_ | ~new_n22949_;
  assign new_n23047_ = ~pi0533 | ~new_n22946_;
  assign new_n23048_ = ~new_n23012_ | ~new_n22947_;
  assign new_n23049_ = ~pi0532 | ~new_n22944_;
  assign new_n23050_ = ~new_n23011_ | ~new_n22945_;
  assign new_n23051_ = ~pi0531 | ~new_n22942_;
  assign new_n23052_ = ~new_n23010_ | ~new_n22943_;
  assign new_n23053_ = ~pi0530 | ~new_n22940_;
  assign new_n23054_ = ~new_n23009_ | ~new_n22941_;
  assign new_n23055_ = ~pi0529 | ~new_n22938_;
  assign new_n23056_ = ~new_n23008_ | ~new_n22939_;
  assign new_n23057_ = ~pi0528 | ~new_n22936_;
  assign new_n23058_ = ~new_n23007_ | ~new_n22937_;
  assign new_n23059_ = ~pi0527 | ~new_n22934_;
  assign new_n23060_ = ~new_n23006_ | ~new_n22935_;
  assign new_n23061_ = ~pi0526 | ~new_n22932_;
  assign new_n23062_ = ~new_n23005_ | ~new_n22933_;
  assign new_n23063_ = ~pi0525 | ~new_n22930_;
  assign new_n23064_ = ~new_n23004_ | ~new_n22931_;
  assign new_n23065_ = ~pi0524 | ~new_n22928_;
  assign new_n23066_ = ~new_n23003_ | ~new_n22929_;
  assign new_n23067_ = ~pi0523 | ~new_n22926_;
  assign new_n23068_ = ~new_n23002_ | ~new_n22927_;
  assign new_n23069_ = ~pi0522 | ~new_n22924_;
  assign new_n23070_ = ~new_n23001_ | ~new_n22925_;
  assign new_n23071_ = ~pi0521 | ~new_n22922_;
  assign new_n23072_ = ~new_n23000_ | ~new_n22923_;
  assign new_n23073_ = ~pi0520 | ~new_n22920_;
  assign new_n23074_ = ~new_n22999_ | ~new_n22921_;
  assign new_n23075_ = ~pi0519 | ~new_n22918_;
  assign new_n23076_ = ~new_n22998_ | ~new_n22919_;
  assign new_n23077_ = ~pi0518 | ~new_n22916_;
  assign new_n23078_ = ~new_n22997_ | ~new_n22917_;
  assign new_n23079_ = ~pi0509;
  assign new_n23080_ = ~pi0510;
  assign new_n23081_ = ~pi0510 | ~pi0509;
  assign new_n23082_ = ~pi0511;
  assign new_n23083_ = ~pi0511 | ~new_n23169_;
  assign new_n23084_ = ~pi0512;
  assign new_n23085_ = ~pi0512 | ~new_n23170_;
  assign new_n23086_ = ~pi0513;
  assign new_n23087_ = ~pi0513 | ~new_n23171_;
  assign new_n23088_ = ~pi0514;
  assign new_n23089_ = ~pi0514 | ~new_n23172_;
  assign new_n23090_ = ~pi0515;
  assign new_n23091_ = ~pi0515 | ~new_n23173_;
  assign new_n23092_ = ~pi0516;
  assign new_n23093_ = ~pi0517;
  assign new_n23094_ = ~pi0516 | ~new_n23174_;
  assign new_n23095_ = ~new_n23175_ | ~pi0517;
  assign new_n23096_ = ~pi0518;
  assign new_n23097_ = ~pi0518 | ~new_n23176_;
  assign new_n23098_ = ~pi0519;
  assign new_n23099_ = ~pi0519 | ~new_n23177_;
  assign new_n23100_ = ~pi0520;
  assign new_n23101_ = ~pi0520 | ~new_n23178_;
  assign new_n23102_ = ~pi0521;
  assign new_n23103_ = ~pi0521 | ~new_n23179_;
  assign new_n23104_ = ~pi0522;
  assign new_n23105_ = ~pi0522 | ~new_n23180_;
  assign new_n23106_ = ~pi0523;
  assign new_n23107_ = ~pi0523 | ~new_n23181_;
  assign new_n23108_ = ~pi0524;
  assign new_n23109_ = ~pi0524 | ~new_n23182_;
  assign new_n23110_ = ~pi0525;
  assign new_n23111_ = ~pi0525 | ~new_n23183_;
  assign new_n23112_ = ~pi0526;
  assign new_n23113_ = ~pi0526 | ~new_n23184_;
  assign new_n23114_ = ~pi0527;
  assign new_n23115_ = ~pi0527 | ~new_n23185_;
  assign new_n23116_ = ~pi0528;
  assign new_n23117_ = ~pi0528 | ~new_n23186_;
  assign new_n23118_ = ~pi0529;
  assign new_n23119_ = ~pi0529 | ~new_n23187_;
  assign new_n23120_ = ~pi0530;
  assign new_n23121_ = ~pi0530 | ~new_n23188_;
  assign new_n23122_ = ~pi0531;
  assign new_n23123_ = ~pi0531 | ~new_n23189_;
  assign new_n23124_ = ~pi0532;
  assign new_n23125_ = ~pi0532 | ~new_n23190_;
  assign new_n23126_ = ~pi0533;
  assign new_n23127_ = ~pi0533 | ~new_n23191_;
  assign new_n23128_ = ~pi0534;
  assign new_n23129_ = ~pi0534 | ~new_n23192_;
  assign new_n23130_ = ~pi0535;
  assign new_n23131_ = ~pi0535 | ~new_n23193_;
  assign new_n23132_ = ~pi0536;
  assign new_n23133_ = ~pi0536 | ~new_n23194_;
  assign new_n23134_ = ~pi0537;
  assign new_n23135_ = ~pi0537 | ~new_n23195_;
  assign new_n23136_ = ~pi0538;
  assign new_n23137_ = ~new_n23199_ | ~new_n23198_;
  assign new_n23138_ = ~new_n23201_ | ~new_n23200_;
  assign new_n23139_ = ~new_n23203_ | ~new_n23202_;
  assign new_n23140_ = ~new_n23205_ | ~new_n23204_;
  assign new_n23141_ = ~new_n23207_ | ~new_n23206_;
  assign new_n23142_ = ~new_n23209_ | ~new_n23208_;
  assign new_n23143_ = ~new_n23211_ | ~new_n23210_;
  assign new_n23144_ = ~new_n23213_ | ~new_n23212_;
  assign new_n23145_ = ~new_n23215_ | ~new_n23214_;
  assign new_n23146_ = ~new_n23217_ | ~new_n23216_;
  assign new_n23147_ = ~new_n23219_ | ~new_n23218_;
  assign new_n23148_ = ~new_n23221_ | ~new_n23220_;
  assign new_n23149_ = ~new_n23223_ | ~new_n23222_;
  assign new_n23150_ = ~new_n23225_ | ~new_n23224_;
  assign new_n23151_ = ~new_n23227_ | ~new_n23226_;
  assign new_n23152_ = ~new_n23229_ | ~new_n23228_;
  assign new_n23153_ = ~new_n23231_ | ~new_n23230_;
  assign new_n23154_ = ~new_n23233_ | ~new_n23232_;
  assign new_n23155_ = ~new_n23235_ | ~new_n23234_;
  assign new_n23156_ = ~new_n23237_ | ~new_n23236_;
  assign new_n23157_ = ~new_n23239_ | ~new_n23238_;
  assign new_n23158_ = ~new_n23241_ | ~new_n23240_;
  assign new_n23159_ = ~new_n23243_ | ~new_n23242_;
  assign new_n23160_ = ~new_n23245_ | ~new_n23244_;
  assign new_n23161_ = ~new_n23247_ | ~new_n23246_;
  assign new_n23162_ = ~new_n23249_ | ~new_n23248_;
  assign new_n23163_ = ~new_n23251_ | ~new_n23250_;
  assign new_n23164_ = ~new_n23253_ | ~new_n23252_;
  assign new_n23165_ = ~new_n23255_ | ~new_n23254_;
  assign new_n23166_ = ~new_n23257_ | ~new_n23256_;
  assign new_n23167_ = ~pi0539;
  assign new_n23168_ = ~pi0538 | ~new_n23196_;
  assign new_n23169_ = ~new_n23081_;
  assign new_n23170_ = ~new_n23083_;
  assign new_n23171_ = ~new_n23085_;
  assign new_n23172_ = ~new_n23087_;
  assign new_n23173_ = ~new_n23089_;
  assign new_n23174_ = ~new_n23091_;
  assign new_n23175_ = ~new_n23094_;
  assign new_n23176_ = ~new_n23095_;
  assign new_n23177_ = ~new_n23097_;
  assign new_n23178_ = ~new_n23099_;
  assign new_n23179_ = ~new_n23101_;
  assign new_n23180_ = ~new_n23103_;
  assign new_n23181_ = ~new_n23105_;
  assign new_n23182_ = ~new_n23107_;
  assign new_n23183_ = ~new_n23109_;
  assign new_n23184_ = ~new_n23111_;
  assign new_n23185_ = ~new_n23113_;
  assign new_n23186_ = ~new_n23115_;
  assign new_n23187_ = ~new_n23117_;
  assign new_n23188_ = ~new_n23119_;
  assign new_n23189_ = ~new_n23121_;
  assign new_n23190_ = ~new_n23123_;
  assign new_n23191_ = ~new_n23125_;
  assign new_n23192_ = ~new_n23127_;
  assign new_n23193_ = ~new_n23129_;
  assign new_n23194_ = ~new_n23131_;
  assign new_n23195_ = ~new_n23133_;
  assign new_n23196_ = ~new_n23135_;
  assign new_n23197_ = ~new_n23168_;
  assign new_n23198_ = ~pi0517 | ~new_n23094_;
  assign new_n23199_ = ~new_n23175_ | ~new_n23093_;
  assign new_n23200_ = ~pi0516 | ~new_n23091_;
  assign new_n23201_ = ~new_n23174_ | ~new_n23092_;
  assign new_n23202_ = ~pi0515 | ~new_n23089_;
  assign new_n23203_ = ~new_n23173_ | ~new_n23090_;
  assign new_n23204_ = ~pi0514 | ~new_n23087_;
  assign new_n23205_ = ~new_n23172_ | ~new_n23088_;
  assign new_n23206_ = ~pi0513 | ~new_n23085_;
  assign new_n23207_ = ~new_n23171_ | ~new_n23086_;
  assign new_n23208_ = ~pi0512 | ~new_n23083_;
  assign new_n23209_ = ~new_n23170_ | ~new_n23084_;
  assign new_n23210_ = ~pi0511 | ~new_n23081_;
  assign new_n23211_ = ~new_n23169_ | ~new_n23082_;
  assign new_n23212_ = ~pi0539 | ~new_n23168_;
  assign new_n23213_ = ~new_n23197_ | ~new_n23167_;
  assign new_n23214_ = ~pi0538 | ~new_n23135_;
  assign new_n23215_ = ~new_n23196_ | ~new_n23136_;
  assign new_n23216_ = ~pi0510 | ~new_n23079_;
  assign new_n23217_ = ~pi0509 | ~new_n23080_;
  assign new_n23218_ = ~pi0537 | ~new_n23133_;
  assign new_n23219_ = ~new_n23195_ | ~new_n23134_;
  assign new_n23220_ = ~pi0536 | ~new_n23131_;
  assign new_n23221_ = ~new_n23194_ | ~new_n23132_;
  assign new_n23222_ = ~pi0535 | ~new_n23129_;
  assign new_n23223_ = ~new_n23193_ | ~new_n23130_;
  assign new_n23224_ = ~pi0534 | ~new_n23127_;
  assign new_n23225_ = ~new_n23192_ | ~new_n23128_;
  assign new_n23226_ = ~pi0533 | ~new_n23125_;
  assign new_n23227_ = ~new_n23191_ | ~new_n23126_;
  assign new_n23228_ = ~pi0532 | ~new_n23123_;
  assign new_n23229_ = ~new_n23190_ | ~new_n23124_;
  assign new_n23230_ = ~pi0531 | ~new_n23121_;
  assign new_n23231_ = ~new_n23189_ | ~new_n23122_;
  assign new_n23232_ = ~pi0530 | ~new_n23119_;
  assign new_n23233_ = ~new_n23188_ | ~new_n23120_;
  assign new_n23234_ = ~pi0529 | ~new_n23117_;
  assign new_n23235_ = ~new_n23187_ | ~new_n23118_;
  assign new_n23236_ = ~pi0528 | ~new_n23115_;
  assign new_n23237_ = ~new_n23186_ | ~new_n23116_;
  assign new_n23238_ = ~pi0527 | ~new_n23113_;
  assign new_n23239_ = ~new_n23185_ | ~new_n23114_;
  assign new_n23240_ = ~pi0526 | ~new_n23111_;
  assign new_n23241_ = ~new_n23184_ | ~new_n23112_;
  assign new_n23242_ = ~pi0525 | ~new_n23109_;
  assign new_n23243_ = ~new_n23183_ | ~new_n23110_;
  assign new_n23244_ = ~pi0524 | ~new_n23107_;
  assign new_n23245_ = ~new_n23182_ | ~new_n23108_;
  assign new_n23246_ = ~pi0523 | ~new_n23105_;
  assign new_n23247_ = ~new_n23181_ | ~new_n23106_;
  assign new_n23248_ = ~pi0522 | ~new_n23103_;
  assign new_n23249_ = ~new_n23180_ | ~new_n23104_;
  assign new_n23250_ = ~pi0521 | ~new_n23101_;
  assign new_n23251_ = ~new_n23179_ | ~new_n23102_;
  assign new_n23252_ = ~pi0520 | ~new_n23099_;
  assign new_n23253_ = ~new_n23178_ | ~new_n23100_;
  assign new_n23254_ = ~pi0519 | ~new_n23097_;
  assign new_n23255_ = ~new_n23177_ | ~new_n23098_;
  assign new_n23256_ = ~pi0518 | ~new_n23095_;
  assign new_n23257_ = ~new_n23176_ | ~new_n23096_;
  assign new_n23258_ = ~pi0317;
  assign new_n23259_ = ~pi0318;
  assign new_n23260_ = ~pi0318 | ~pi0317;
  assign new_n23261_ = ~pi0319;
  assign new_n23262_ = ~pi0319 | ~new_n23351_;
  assign new_n23263_ = ~pi0320;
  assign new_n23264_ = ~pi0320 | ~new_n23352_;
  assign new_n23265_ = ~pi0321;
  assign new_n23266_ = ~pi0321 | ~new_n23353_;
  assign new_n23267_ = ~pi0322;
  assign new_n23268_ = ~pi0322 | ~new_n23354_;
  assign new_n23269_ = ~pi0323;
  assign new_n23270_ = ~pi0323 | ~new_n23355_;
  assign new_n23271_ = ~pi0324;
  assign new_n23272_ = ~pi0324 | ~new_n23356_;
  assign new_n23273_ = ~pi0325;
  assign new_n23274_ = ~pi0326;
  assign new_n23275_ = ~pi0325 | ~new_n23357_;
  assign new_n23276_ = ~new_n23358_ | ~pi0326;
  assign new_n23277_ = ~pi0327;
  assign new_n23278_ = ~pi0327 | ~new_n23359_;
  assign new_n23279_ = ~pi0328;
  assign new_n23280_ = ~pi0328 | ~new_n23360_;
  assign new_n23281_ = ~pi0329;
  assign new_n23282_ = ~pi0329 | ~new_n23361_;
  assign new_n23283_ = ~pi0330;
  assign new_n23284_ = ~pi0330 | ~new_n23362_;
  assign new_n23285_ = ~pi0331;
  assign new_n23286_ = ~pi0331 | ~new_n23363_;
  assign new_n23287_ = ~pi0332;
  assign new_n23288_ = ~pi0332 | ~new_n23364_;
  assign new_n23289_ = ~pi0333;
  assign new_n23290_ = ~pi0333 | ~new_n23365_;
  assign new_n23291_ = ~pi0334;
  assign new_n23292_ = ~pi0334 | ~new_n23366_;
  assign new_n23293_ = ~pi0335;
  assign new_n23294_ = ~pi0335 | ~new_n23367_;
  assign new_n23295_ = ~pi0336;
  assign new_n23296_ = ~pi0336 | ~new_n23368_;
  assign new_n23297_ = ~pi0337;
  assign new_n23298_ = ~pi0337 | ~new_n23369_;
  assign new_n23299_ = ~pi0338;
  assign new_n23300_ = ~pi0338 | ~new_n23370_;
  assign new_n23301_ = ~pi0339;
  assign new_n23302_ = ~pi0339 | ~new_n23371_;
  assign new_n23303_ = ~pi0340;
  assign new_n23304_ = ~pi0340 | ~new_n23372_;
  assign new_n23305_ = ~pi0341;
  assign new_n23306_ = ~pi0341 | ~new_n23373_;
  assign new_n23307_ = ~pi0342;
  assign new_n23308_ = ~pi0342 | ~new_n23374_;
  assign new_n23309_ = ~pi0343;
  assign new_n23310_ = ~pi0343 | ~new_n23375_;
  assign new_n23311_ = ~pi0344;
  assign new_n23312_ = ~pi0344 | ~new_n23376_;
  assign new_n23313_ = ~pi0345;
  assign new_n23314_ = ~pi0345 | ~new_n23377_;
  assign new_n23315_ = ~pi0346;
  assign new_n23316_ = ~pi0346 | ~new_n23378_;
  assign new_n23317_ = ~pi0347;
  assign new_n23318_ = ~new_n23382_ | ~new_n23381_;
  assign new_n23319_ = ~new_n23384_ | ~new_n23383_;
  assign new_n23320_ = ~new_n23386_ | ~new_n23385_;
  assign new_n23321_ = ~new_n23388_ | ~new_n23387_;
  assign new_n23322_ = ~new_n23390_ | ~new_n23389_;
  assign new_n23323_ = ~new_n23392_ | ~new_n23391_;
  assign new_n23324_ = ~new_n23394_ | ~new_n23393_;
  assign new_n23325_ = ~new_n23396_ | ~new_n23395_;
  assign new_n23326_ = ~new_n23398_ | ~new_n23397_;
  assign new_n23327_ = ~new_n23400_ | ~new_n23399_;
  assign new_n23328_ = ~new_n23402_ | ~new_n23401_;
  assign new_n23329_ = ~new_n23404_ | ~new_n23403_;
  assign new_n23330_ = ~new_n23406_ | ~new_n23405_;
  assign new_n23331_ = ~new_n23408_ | ~new_n23407_;
  assign new_n23332_ = ~new_n23410_ | ~new_n23409_;
  assign new_n23333_ = ~new_n23412_ | ~new_n23411_;
  assign new_n23334_ = ~new_n23414_ | ~new_n23413_;
  assign new_n23335_ = ~new_n23416_ | ~new_n23415_;
  assign new_n23336_ = ~new_n23418_ | ~new_n23417_;
  assign new_n23337_ = ~new_n23420_ | ~new_n23419_;
  assign new_n23338_ = ~new_n23422_ | ~new_n23421_;
  assign new_n23339_ = ~new_n23424_ | ~new_n23423_;
  assign new_n23340_ = ~new_n23426_ | ~new_n23425_;
  assign new_n23341_ = ~new_n23428_ | ~new_n23427_;
  assign new_n23342_ = ~new_n23430_ | ~new_n23429_;
  assign new_n23343_ = ~new_n23432_ | ~new_n23431_;
  assign new_n23344_ = ~new_n23434_ | ~new_n23433_;
  assign new_n23345_ = ~new_n23436_ | ~new_n23435_;
  assign new_n23346_ = ~new_n23438_ | ~new_n23437_;
  assign new_n23347_ = ~new_n23440_ | ~new_n23439_;
  assign new_n23348_ = ~new_n23442_ | ~new_n23441_;
  assign new_n23349_ = ~pi0348;
  assign new_n23350_ = ~pi0347 | ~new_n23379_;
  assign new_n23351_ = ~new_n23260_;
  assign new_n23352_ = ~new_n23262_;
  assign new_n23353_ = ~new_n23264_;
  assign new_n23354_ = ~new_n23266_;
  assign new_n23355_ = ~new_n23268_;
  assign new_n23356_ = ~new_n23270_;
  assign new_n23357_ = ~new_n23272_;
  assign new_n23358_ = ~new_n23275_;
  assign new_n23359_ = ~new_n23276_;
  assign new_n23360_ = ~new_n23278_;
  assign new_n23361_ = ~new_n23280_;
  assign new_n23362_ = ~new_n23282_;
  assign new_n23363_ = ~new_n23284_;
  assign new_n23364_ = ~new_n23286_;
  assign new_n23365_ = ~new_n23288_;
  assign new_n23366_ = ~new_n23290_;
  assign new_n23367_ = ~new_n23292_;
  assign new_n23368_ = ~new_n23294_;
  assign new_n23369_ = ~new_n23296_;
  assign new_n23370_ = ~new_n23298_;
  assign new_n23371_ = ~new_n23300_;
  assign new_n23372_ = ~new_n23302_;
  assign new_n23373_ = ~new_n23304_;
  assign new_n23374_ = ~new_n23306_;
  assign new_n23375_ = ~new_n23308_;
  assign new_n23376_ = ~new_n23310_;
  assign new_n23377_ = ~new_n23312_;
  assign new_n23378_ = ~new_n23314_;
  assign new_n23379_ = ~new_n23316_;
  assign new_n23380_ = ~new_n23350_;
  assign new_n23381_ = ~pi0326 | ~new_n23275_;
  assign new_n23382_ = ~new_n23358_ | ~new_n23274_;
  assign new_n23383_ = ~pi0325 | ~new_n23272_;
  assign new_n23384_ = ~new_n23357_ | ~new_n23273_;
  assign new_n23385_ = ~pi0324 | ~new_n23270_;
  assign new_n23386_ = ~new_n23356_ | ~new_n23271_;
  assign new_n23387_ = ~pi0323 | ~new_n23268_;
  assign new_n23388_ = ~new_n23355_ | ~new_n23269_;
  assign new_n23389_ = ~pi0322 | ~new_n23266_;
  assign new_n23390_ = ~new_n23354_ | ~new_n23267_;
  assign new_n23391_ = ~pi0321 | ~new_n23264_;
  assign new_n23392_ = ~new_n23353_ | ~new_n23265_;
  assign new_n23393_ = ~pi0320 | ~new_n23262_;
  assign new_n23394_ = ~new_n23352_ | ~new_n23263_;
  assign new_n23395_ = ~pi0348 | ~new_n23350_;
  assign new_n23396_ = ~new_n23380_ | ~new_n23349_;
  assign new_n23397_ = ~pi0347 | ~new_n23316_;
  assign new_n23398_ = ~new_n23379_ | ~new_n23317_;
  assign new_n23399_ = ~pi0319 | ~new_n23260_;
  assign new_n23400_ = ~new_n23351_ | ~new_n23261_;
  assign new_n23401_ = ~pi0346 | ~new_n23314_;
  assign new_n23402_ = ~new_n23378_ | ~new_n23315_;
  assign new_n23403_ = ~pi0345 | ~new_n23312_;
  assign new_n23404_ = ~new_n23377_ | ~new_n23313_;
  assign new_n23405_ = ~pi0344 | ~new_n23310_;
  assign new_n23406_ = ~new_n23376_ | ~new_n23311_;
  assign new_n23407_ = ~pi0343 | ~new_n23308_;
  assign new_n23408_ = ~new_n23375_ | ~new_n23309_;
  assign new_n23409_ = ~pi0342 | ~new_n23306_;
  assign new_n23410_ = ~new_n23374_ | ~new_n23307_;
  assign new_n23411_ = ~pi0341 | ~new_n23304_;
  assign new_n23412_ = ~new_n23373_ | ~new_n23305_;
  assign new_n23413_ = ~pi0340 | ~new_n23302_;
  assign new_n23414_ = ~new_n23372_ | ~new_n23303_;
  assign new_n23415_ = ~pi0339 | ~new_n23300_;
  assign new_n23416_ = ~new_n23371_ | ~new_n23301_;
  assign new_n23417_ = ~pi0338 | ~new_n23298_;
  assign new_n23418_ = ~new_n23370_ | ~new_n23299_;
  assign new_n23419_ = ~pi0337 | ~new_n23296_;
  assign new_n23420_ = ~new_n23369_ | ~new_n23297_;
  assign new_n23421_ = ~pi0318 | ~new_n23258_;
  assign new_n23422_ = ~pi0317 | ~new_n23259_;
  assign new_n23423_ = ~pi0336 | ~new_n23294_;
  assign new_n23424_ = ~new_n23368_ | ~new_n23295_;
  assign new_n23425_ = ~pi0335 | ~new_n23292_;
  assign new_n23426_ = ~new_n23367_ | ~new_n23293_;
  assign new_n23427_ = ~pi0334 | ~new_n23290_;
  assign new_n23428_ = ~new_n23366_ | ~new_n23291_;
  assign new_n23429_ = ~pi0333 | ~new_n23288_;
  assign new_n23430_ = ~new_n23365_ | ~new_n23289_;
  assign new_n23431_ = ~pi0332 | ~new_n23286_;
  assign new_n23432_ = ~new_n23364_ | ~new_n23287_;
  assign new_n23433_ = ~pi0331 | ~new_n23284_;
  assign new_n23434_ = ~new_n23363_ | ~new_n23285_;
  assign new_n23435_ = ~pi0330 | ~new_n23282_;
  assign new_n23436_ = ~new_n23362_ | ~new_n23283_;
  assign new_n23437_ = ~pi0329 | ~new_n23280_;
  assign new_n23438_ = ~new_n23361_ | ~new_n23281_;
  assign new_n23439_ = ~pi0328 | ~new_n23278_;
  assign new_n23440_ = ~new_n23360_ | ~new_n23279_;
  assign new_n23441_ = ~pi0327 | ~new_n23276_;
  assign new_n23442_ = ~new_n23359_ | ~new_n23277_;
  assign new_n23443_ = ~new_n22402_ & ~new_n23445_;
  assign new_n23444_ = new_n22417_ & new_n23446_;
  assign new_n23445_ = ~new_n23444_ & ~new_n22416_ & ~new_n22415_;
  assign new_n23446_ = new_n22403_ | new_n22418_;
  assign new_n23447_ = ~pi0317;
  assign new_n23448_ = ~pi0318;
  assign new_n23449_ = ~pi0318 | ~pi0317;
  assign new_n23450_ = ~pi0319;
  assign new_n23451_ = ~pi0319 | ~new_n23540_;
  assign new_n23452_ = ~pi0320;
  assign new_n23453_ = ~pi0320 | ~new_n23541_;
  assign new_n23454_ = ~pi0321;
  assign new_n23455_ = ~pi0321 | ~new_n23542_;
  assign new_n23456_ = ~pi0322;
  assign new_n23457_ = ~pi0322 | ~new_n23543_;
  assign new_n23458_ = ~pi0323;
  assign new_n23459_ = ~pi0323 | ~new_n23544_;
  assign new_n23460_ = ~pi0324;
  assign new_n23461_ = ~pi0324 | ~new_n23545_;
  assign new_n23462_ = ~pi0325;
  assign new_n23463_ = ~pi0326;
  assign new_n23464_ = ~pi0325 | ~new_n23546_;
  assign new_n23465_ = ~new_n23547_ | ~pi0326;
  assign new_n23466_ = ~pi0327;
  assign new_n23467_ = ~pi0327 | ~new_n23548_;
  assign new_n23468_ = ~pi0328;
  assign new_n23469_ = ~pi0328 | ~new_n23549_;
  assign new_n23470_ = ~pi0329;
  assign new_n23471_ = ~pi0329 | ~new_n23550_;
  assign new_n23472_ = ~pi0330;
  assign new_n23473_ = ~pi0330 | ~new_n23551_;
  assign new_n23474_ = ~pi0331;
  assign new_n23475_ = ~pi0331 | ~new_n23552_;
  assign new_n23476_ = ~pi0332;
  assign new_n23477_ = ~pi0332 | ~new_n23553_;
  assign new_n23478_ = ~pi0333;
  assign new_n23479_ = ~pi0333 | ~new_n23554_;
  assign new_n23480_ = ~pi0334;
  assign new_n23481_ = ~pi0334 | ~new_n23555_;
  assign new_n23482_ = ~pi0335;
  assign new_n23483_ = ~pi0335 | ~new_n23556_;
  assign new_n23484_ = ~pi0336;
  assign new_n23485_ = ~pi0336 | ~new_n23557_;
  assign new_n23486_ = ~pi0337;
  assign new_n23487_ = ~pi0337 | ~new_n23558_;
  assign new_n23488_ = ~pi0338;
  assign new_n23489_ = ~pi0338 | ~new_n23559_;
  assign new_n23490_ = ~pi0339;
  assign new_n23491_ = ~pi0339 | ~new_n23560_;
  assign new_n23492_ = ~pi0340;
  assign new_n23493_ = ~pi0340 | ~new_n23561_;
  assign new_n23494_ = ~pi0341;
  assign new_n23495_ = ~pi0341 | ~new_n23562_;
  assign new_n23496_ = ~pi0342;
  assign new_n23497_ = ~pi0342 | ~new_n23563_;
  assign new_n23498_ = ~pi0343;
  assign new_n23499_ = ~pi0343 | ~new_n23564_;
  assign new_n23500_ = ~pi0344;
  assign new_n23501_ = ~pi0344 | ~new_n23565_;
  assign new_n23502_ = ~pi0345;
  assign new_n23503_ = ~pi0345 | ~new_n23566_;
  assign new_n23504_ = ~pi0346;
  assign new_n23505_ = ~pi0346 | ~new_n23567_;
  assign new_n23506_ = ~pi0347;
  assign new_n23507_ = ~new_n23571_ | ~new_n23570_;
  assign new_n23508_ = ~new_n23573_ | ~new_n23572_;
  assign new_n23509_ = ~new_n23575_ | ~new_n23574_;
  assign new_n23510_ = ~new_n23577_ | ~new_n23576_;
  assign new_n23511_ = ~new_n23579_ | ~new_n23578_;
  assign new_n23512_ = ~new_n23581_ | ~new_n23580_;
  assign new_n23513_ = ~new_n23583_ | ~new_n23582_;
  assign new_n23514_ = ~new_n23585_ | ~new_n23584_;
  assign new_n23515_ = ~new_n23587_ | ~new_n23586_;
  assign new_n23516_ = ~new_n23589_ | ~new_n23588_;
  assign new_n23517_ = ~new_n23591_ | ~new_n23590_;
  assign new_n23518_ = ~new_n23593_ | ~new_n23592_;
  assign new_n23519_ = ~new_n23595_ | ~new_n23594_;
  assign new_n23520_ = ~new_n23597_ | ~new_n23596_;
  assign new_n23521_ = ~new_n23599_ | ~new_n23598_;
  assign new_n23522_ = ~new_n23601_ | ~new_n23600_;
  assign new_n23523_ = ~new_n23603_ | ~new_n23602_;
  assign new_n23524_ = ~new_n23605_ | ~new_n23604_;
  assign new_n23525_ = ~new_n23607_ | ~new_n23606_;
  assign new_n23526_ = ~new_n23609_ | ~new_n23608_;
  assign new_n23527_ = ~new_n23611_ | ~new_n23610_;
  assign new_n23528_ = ~new_n23613_ | ~new_n23612_;
  assign new_n23529_ = ~new_n23615_ | ~new_n23614_;
  assign new_n23530_ = ~new_n23617_ | ~new_n23616_;
  assign new_n23531_ = ~new_n23619_ | ~new_n23618_;
  assign new_n23532_ = ~new_n23621_ | ~new_n23620_;
  assign new_n23533_ = ~new_n23623_ | ~new_n23622_;
  assign new_n23534_ = ~new_n23625_ | ~new_n23624_;
  assign new_n23535_ = ~new_n23627_ | ~new_n23626_;
  assign new_n23536_ = ~new_n23629_ | ~new_n23628_;
  assign new_n23537_ = ~new_n23631_ | ~new_n23630_;
  assign new_n23538_ = ~pi0348;
  assign new_n23539_ = ~pi0347 | ~new_n23568_;
  assign new_n23540_ = ~new_n23449_;
  assign new_n23541_ = ~new_n23451_;
  assign new_n23542_ = ~new_n23453_;
  assign new_n23543_ = ~new_n23455_;
  assign new_n23544_ = ~new_n23457_;
  assign new_n23545_ = ~new_n23459_;
  assign new_n23546_ = ~new_n23461_;
  assign new_n23547_ = ~new_n23464_;
  assign new_n23548_ = ~new_n23465_;
  assign new_n23549_ = ~new_n23467_;
  assign new_n23550_ = ~new_n23469_;
  assign new_n23551_ = ~new_n23471_;
  assign new_n23552_ = ~new_n23473_;
  assign new_n23553_ = ~new_n23475_;
  assign new_n23554_ = ~new_n23477_;
  assign new_n23555_ = ~new_n23479_;
  assign new_n23556_ = ~new_n23481_;
  assign new_n23557_ = ~new_n23483_;
  assign new_n23558_ = ~new_n23485_;
  assign new_n23559_ = ~new_n23487_;
  assign new_n23560_ = ~new_n23489_;
  assign new_n23561_ = ~new_n23491_;
  assign new_n23562_ = ~new_n23493_;
  assign new_n23563_ = ~new_n23495_;
  assign new_n23564_ = ~new_n23497_;
  assign new_n23565_ = ~new_n23499_;
  assign new_n23566_ = ~new_n23501_;
  assign new_n23567_ = ~new_n23503_;
  assign new_n23568_ = ~new_n23505_;
  assign new_n23569_ = ~new_n23539_;
  assign new_n23570_ = ~pi0326 | ~new_n23464_;
  assign new_n23571_ = ~new_n23547_ | ~new_n23463_;
  assign new_n23572_ = ~pi0325 | ~new_n23461_;
  assign new_n23573_ = ~new_n23546_ | ~new_n23462_;
  assign new_n23574_ = ~pi0324 | ~new_n23459_;
  assign new_n23575_ = ~new_n23545_ | ~new_n23460_;
  assign new_n23576_ = ~pi0323 | ~new_n23457_;
  assign new_n23577_ = ~new_n23544_ | ~new_n23458_;
  assign new_n23578_ = ~pi0322 | ~new_n23455_;
  assign new_n23579_ = ~new_n23543_ | ~new_n23456_;
  assign new_n23580_ = ~pi0321 | ~new_n23453_;
  assign new_n23581_ = ~new_n23542_ | ~new_n23454_;
  assign new_n23582_ = ~pi0320 | ~new_n23451_;
  assign new_n23583_ = ~new_n23541_ | ~new_n23452_;
  assign new_n23584_ = ~pi0348 | ~new_n23539_;
  assign new_n23585_ = ~new_n23569_ | ~new_n23538_;
  assign new_n23586_ = ~pi0347 | ~new_n23505_;
  assign new_n23587_ = ~new_n23568_ | ~new_n23506_;
  assign new_n23588_ = ~pi0319 | ~new_n23449_;
  assign new_n23589_ = ~new_n23540_ | ~new_n23450_;
  assign new_n23590_ = ~pi0346 | ~new_n23503_;
  assign new_n23591_ = ~new_n23567_ | ~new_n23504_;
  assign new_n23592_ = ~pi0345 | ~new_n23501_;
  assign new_n23593_ = ~new_n23566_ | ~new_n23502_;
  assign new_n23594_ = ~pi0344 | ~new_n23499_;
  assign new_n23595_ = ~new_n23565_ | ~new_n23500_;
  assign new_n23596_ = ~pi0343 | ~new_n23497_;
  assign new_n23597_ = ~new_n23564_ | ~new_n23498_;
  assign new_n23598_ = ~pi0342 | ~new_n23495_;
  assign new_n23599_ = ~new_n23563_ | ~new_n23496_;
  assign new_n23600_ = ~pi0341 | ~new_n23493_;
  assign new_n23601_ = ~new_n23562_ | ~new_n23494_;
  assign new_n23602_ = ~pi0340 | ~new_n23491_;
  assign new_n23603_ = ~new_n23561_ | ~new_n23492_;
  assign new_n23604_ = ~pi0339 | ~new_n23489_;
  assign new_n23605_ = ~new_n23560_ | ~new_n23490_;
  assign new_n23606_ = ~pi0338 | ~new_n23487_;
  assign new_n23607_ = ~new_n23559_ | ~new_n23488_;
  assign new_n23608_ = ~pi0337 | ~new_n23485_;
  assign new_n23609_ = ~new_n23558_ | ~new_n23486_;
  assign new_n23610_ = ~pi0318 | ~new_n23447_;
  assign new_n23611_ = ~pi0317 | ~new_n23448_;
  assign new_n23612_ = ~pi0336 | ~new_n23483_;
  assign new_n23613_ = ~new_n23557_ | ~new_n23484_;
  assign new_n23614_ = ~pi0335 | ~new_n23481_;
  assign new_n23615_ = ~new_n23556_ | ~new_n23482_;
  assign new_n23616_ = ~pi0334 | ~new_n23479_;
  assign new_n23617_ = ~new_n23555_ | ~new_n23480_;
  assign new_n23618_ = ~pi0333 | ~new_n23477_;
  assign new_n23619_ = ~new_n23554_ | ~new_n23478_;
  assign new_n23620_ = ~pi0332 | ~new_n23475_;
  assign new_n23621_ = ~new_n23553_ | ~new_n23476_;
  assign new_n23622_ = ~pi0331 | ~new_n23473_;
  assign new_n23623_ = ~new_n23552_ | ~new_n23474_;
  assign new_n23624_ = ~pi0330 | ~new_n23471_;
  assign new_n23625_ = ~new_n23551_ | ~new_n23472_;
  assign new_n23626_ = ~pi0329 | ~new_n23469_;
  assign new_n23627_ = ~new_n23550_ | ~new_n23470_;
  assign new_n23628_ = ~pi0328 | ~new_n23467_;
  assign new_n23629_ = ~new_n23549_ | ~new_n23468_;
  assign new_n23630_ = ~pi0327 | ~new_n23465_;
  assign new_n23631_ = ~new_n23548_ | ~new_n23466_;
  assign new_n23632_ = ~new_n23653_ | ~new_n23654_;
  assign new_n23633_ = ~pi0312;
  assign new_n23634_ = ~pi0316 | ~new_n23641_;
  assign new_n23635_ = ~pi0315;
  assign new_n23636_ = ~new_n4462_;
  assign new_n23637_ = ~pi0314;
  assign new_n23638_ = ~pi0313;
  assign new_n23639_ = ~new_n4461_;
  assign new_n23640_ = ~new_n4460_;
  assign new_n23641_ = ~new_n4464_;
  assign new_n23642_ = ~new_n23634_;
  assign new_n23643_ = ~pi0315 | ~new_n23642_;
  assign new_n23644_ = ~new_n4463_ | ~new_n23643_;
  assign new_n23645_ = ~new_n23634_ | ~new_n23635_;
  assign new_n23646_ = ~new_n4462_ | ~new_n23637_;
  assign new_n23647_ = ~new_n23644_ | ~new_n23645_ | ~new_n23646_;
  assign new_n23648_ = ~pi0314 | ~new_n23636_;
  assign new_n23649_ = ~pi0313 | ~new_n23639_;
  assign new_n23650_ = ~new_n23647_ | ~new_n23648_ | ~new_n23649_;
  assign new_n23651_ = ~new_n4461_ | ~new_n23638_;
  assign new_n23652_ = ~new_n4460_ | ~new_n23633_;
  assign new_n23653_ = ~new_n23650_ | ~new_n23651_ | ~new_n23652_;
  assign new_n23654_ = ~pi0312 | ~new_n23640_;
  assign new_n23655_ = ~pi0350;
  assign new_n23656_ = ~pi0351;
  assign new_n23657_ = ~pi0351 | ~pi0350;
  assign new_n23658_ = ~pi0352;
  assign new_n23659_ = ~pi0352 | ~new_n23745_;
  assign new_n23660_ = ~pi0353;
  assign new_n23661_ = ~pi0353 | ~new_n23746_;
  assign new_n23662_ = ~pi0354;
  assign new_n23663_ = ~pi0354 | ~new_n23747_;
  assign new_n23664_ = ~pi0355;
  assign new_n23665_ = ~pi0355 | ~new_n23748_;
  assign new_n23666_ = ~pi0356;
  assign new_n23667_ = ~pi0356 | ~new_n23749_;
  assign new_n23668_ = ~pi0357;
  assign new_n23669_ = ~pi0358;
  assign new_n23670_ = ~pi0357 | ~new_n23750_;
  assign new_n23671_ = ~new_n23751_ | ~pi0358;
  assign new_n23672_ = ~pi0359;
  assign new_n23673_ = ~pi0359 | ~new_n23752_;
  assign new_n23674_ = ~pi0360;
  assign new_n23675_ = ~pi0360 | ~new_n23753_;
  assign new_n23676_ = ~pi0361;
  assign new_n23677_ = ~pi0361 | ~new_n23754_;
  assign new_n23678_ = ~pi0362;
  assign new_n23679_ = ~pi0362 | ~new_n23755_;
  assign new_n23680_ = ~pi0363;
  assign new_n23681_ = ~pi0363 | ~new_n23756_;
  assign new_n23682_ = ~pi0364;
  assign new_n23683_ = ~pi0364 | ~new_n23757_;
  assign new_n23684_ = ~pi0365;
  assign new_n23685_ = ~pi0365 | ~new_n23758_;
  assign new_n23686_ = ~pi0366;
  assign new_n23687_ = ~pi0366 | ~new_n23759_;
  assign new_n23688_ = ~pi0367;
  assign new_n23689_ = ~pi0367 | ~new_n23760_;
  assign new_n23690_ = ~pi0368;
  assign new_n23691_ = ~pi0368 | ~new_n23761_;
  assign new_n23692_ = ~pi0369;
  assign new_n23693_ = ~pi0369 | ~new_n23762_;
  assign new_n23694_ = ~pi0370;
  assign new_n23695_ = ~pi0370 | ~new_n23763_;
  assign new_n23696_ = ~pi0371;
  assign new_n23697_ = ~pi0371 | ~new_n23764_;
  assign new_n23698_ = ~pi0372;
  assign new_n23699_ = ~pi0372 | ~new_n23765_;
  assign new_n23700_ = ~pi0373;
  assign new_n23701_ = ~pi0373 | ~new_n23766_;
  assign new_n23702_ = ~pi0374;
  assign new_n23703_ = ~pi0374 | ~new_n23767_;
  assign new_n23704_ = ~pi0375;
  assign new_n23705_ = ~pi0375 | ~new_n23768_;
  assign new_n23706_ = ~pi0376;
  assign new_n23707_ = ~pi0376 | ~new_n23769_;
  assign new_n23708_ = ~pi0377;
  assign new_n23709_ = ~pi0377 | ~new_n23770_;
  assign new_n23710_ = ~pi0378;
  assign new_n23711_ = ~pi0378 | ~new_n23771_;
  assign new_n23712_ = ~pi0379;
  assign new_n23713_ = ~new_n23775_ | ~new_n23774_;
  assign new_n23714_ = ~new_n23777_ | ~new_n23776_;
  assign new_n23715_ = ~new_n23779_ | ~new_n23778_;
  assign new_n23716_ = ~new_n23781_ | ~new_n23780_;
  assign new_n23717_ = ~new_n23783_ | ~new_n23782_;
  assign new_n23718_ = ~new_n23785_ | ~new_n23784_;
  assign new_n23719_ = ~new_n23787_ | ~new_n23786_;
  assign new_n23720_ = ~new_n23789_ | ~new_n23788_;
  assign new_n23721_ = ~new_n23791_ | ~new_n23790_;
  assign new_n23722_ = ~new_n23793_ | ~new_n23792_;
  assign new_n23723_ = ~new_n23795_ | ~new_n23794_;
  assign new_n23724_ = ~new_n23797_ | ~new_n23796_;
  assign new_n23725_ = ~new_n23799_ | ~new_n23798_;
  assign new_n23726_ = ~new_n23801_ | ~new_n23800_;
  assign new_n23727_ = ~new_n23803_ | ~new_n23802_;
  assign new_n23728_ = ~new_n23805_ | ~new_n23804_;
  assign new_n23729_ = ~new_n23807_ | ~new_n23806_;
  assign new_n23730_ = ~new_n23809_ | ~new_n23808_;
  assign new_n23731_ = ~new_n23811_ | ~new_n23810_;
  assign new_n23732_ = ~new_n23813_ | ~new_n23812_;
  assign new_n23733_ = ~new_n23815_ | ~new_n23814_;
  assign new_n23734_ = ~new_n23817_ | ~new_n23816_;
  assign new_n23735_ = ~new_n23819_ | ~new_n23818_;
  assign new_n23736_ = ~new_n23821_ | ~new_n23820_;
  assign new_n23737_ = ~new_n23823_ | ~new_n23822_;
  assign new_n23738_ = ~new_n23825_ | ~new_n23824_;
  assign new_n23739_ = ~new_n23827_ | ~new_n23826_;
  assign new_n23740_ = ~new_n23829_ | ~new_n23828_;
  assign new_n23741_ = ~new_n23831_ | ~new_n23830_;
  assign new_n23742_ = ~new_n23833_ | ~new_n23832_;
  assign new_n23743_ = ~pi0380;
  assign new_n23744_ = ~pi0379 | ~new_n23772_;
  assign new_n23745_ = ~new_n23657_;
  assign new_n23746_ = ~new_n23659_;
  assign new_n23747_ = ~new_n23661_;
  assign new_n23748_ = ~new_n23663_;
  assign new_n23749_ = ~new_n23665_;
  assign new_n23750_ = ~new_n23667_;
  assign new_n23751_ = ~new_n23670_;
  assign new_n23752_ = ~new_n23671_;
  assign new_n23753_ = ~new_n23673_;
  assign new_n23754_ = ~new_n23675_;
  assign new_n23755_ = ~new_n23677_;
  assign new_n23756_ = ~new_n23679_;
  assign new_n23757_ = ~new_n23681_;
  assign new_n23758_ = ~new_n23683_;
  assign new_n23759_ = ~new_n23685_;
  assign new_n23760_ = ~new_n23687_;
  assign new_n23761_ = ~new_n23689_;
  assign new_n23762_ = ~new_n23691_;
  assign new_n23763_ = ~new_n23693_;
  assign new_n23764_ = ~new_n23695_;
  assign new_n23765_ = ~new_n23697_;
  assign new_n23766_ = ~new_n23699_;
  assign new_n23767_ = ~new_n23701_;
  assign new_n23768_ = ~new_n23703_;
  assign new_n23769_ = ~new_n23705_;
  assign new_n23770_ = ~new_n23707_;
  assign new_n23771_ = ~new_n23709_;
  assign new_n23772_ = ~new_n23711_;
  assign new_n23773_ = ~new_n23744_;
  assign new_n23774_ = ~pi0358 | ~new_n23670_;
  assign new_n23775_ = ~new_n23751_ | ~new_n23669_;
  assign new_n23776_ = ~pi0357 | ~new_n23667_;
  assign new_n23777_ = ~new_n23750_ | ~new_n23668_;
  assign new_n23778_ = ~pi0356 | ~new_n23665_;
  assign new_n23779_ = ~new_n23749_ | ~new_n23666_;
  assign new_n23780_ = ~pi0355 | ~new_n23663_;
  assign new_n23781_ = ~new_n23748_ | ~new_n23664_;
  assign new_n23782_ = ~pi0354 | ~new_n23661_;
  assign new_n23783_ = ~new_n23747_ | ~new_n23662_;
  assign new_n23784_ = ~pi0353 | ~new_n23659_;
  assign new_n23785_ = ~new_n23746_ | ~new_n23660_;
  assign new_n23786_ = ~pi0352 | ~new_n23657_;
  assign new_n23787_ = ~new_n23745_ | ~new_n23658_;
  assign new_n23788_ = ~pi0380 | ~new_n23744_;
  assign new_n23789_ = ~new_n23773_ | ~new_n23743_;
  assign new_n23790_ = ~pi0379 | ~new_n23711_;
  assign new_n23791_ = ~new_n23772_ | ~new_n23712_;
  assign new_n23792_ = ~pi0351 | ~new_n23655_;
  assign new_n23793_ = ~pi0350 | ~new_n23656_;
  assign new_n23794_ = ~pi0378 | ~new_n23709_;
  assign new_n23795_ = ~new_n23771_ | ~new_n23710_;
  assign new_n23796_ = ~pi0377 | ~new_n23707_;
  assign new_n23797_ = ~new_n23770_ | ~new_n23708_;
  assign new_n23798_ = ~pi0376 | ~new_n23705_;
  assign new_n23799_ = ~new_n23769_ | ~new_n23706_;
  assign new_n23800_ = ~pi0375 | ~new_n23703_;
  assign new_n23801_ = ~new_n23768_ | ~new_n23704_;
  assign new_n23802_ = ~pi0374 | ~new_n23701_;
  assign new_n23803_ = ~new_n23767_ | ~new_n23702_;
  assign new_n23804_ = ~pi0373 | ~new_n23699_;
  assign new_n23805_ = ~new_n23766_ | ~new_n23700_;
  assign new_n23806_ = ~pi0372 | ~new_n23697_;
  assign new_n23807_ = ~new_n23765_ | ~new_n23698_;
  assign new_n23808_ = ~pi0371 | ~new_n23695_;
  assign new_n23809_ = ~new_n23764_ | ~new_n23696_;
  assign new_n23810_ = ~pi0370 | ~new_n23693_;
  assign new_n23811_ = ~new_n23763_ | ~new_n23694_;
  assign new_n23812_ = ~pi0369 | ~new_n23691_;
  assign new_n23813_ = ~new_n23762_ | ~new_n23692_;
  assign new_n23814_ = ~pi0368 | ~new_n23689_;
  assign new_n23815_ = ~new_n23761_ | ~new_n23690_;
  assign new_n23816_ = ~pi0367 | ~new_n23687_;
  assign new_n23817_ = ~new_n23760_ | ~new_n23688_;
  assign new_n23818_ = ~pi0366 | ~new_n23685_;
  assign new_n23819_ = ~new_n23759_ | ~new_n23686_;
  assign new_n23820_ = ~pi0365 | ~new_n23683_;
  assign new_n23821_ = ~new_n23758_ | ~new_n23684_;
  assign new_n23822_ = ~pi0364 | ~new_n23681_;
  assign new_n23823_ = ~new_n23757_ | ~new_n23682_;
  assign new_n23824_ = ~pi0363 | ~new_n23679_;
  assign new_n23825_ = ~new_n23756_ | ~new_n23680_;
  assign new_n23826_ = ~pi0362 | ~new_n23677_;
  assign new_n23827_ = ~new_n23755_ | ~new_n23678_;
  assign new_n23828_ = ~pi0361 | ~new_n23675_;
  assign new_n23829_ = ~new_n23754_ | ~new_n23676_;
  assign new_n23830_ = ~pi0360 | ~new_n23673_;
  assign new_n23831_ = ~new_n23753_ | ~new_n23674_;
  assign new_n23832_ = ~pi0359 | ~new_n23671_;
  assign new_n23833_ = ~new_n23752_ | ~new_n23672_;
  assign new_n23834_ = ~new_n3778_;
  assign new_n23835_ = new_n23852_ & new_n23857_;
  assign new_n23836_ = ~new_n3779_;
  assign new_n23837_ = ~new_n3779_ | ~new_n3778_;
  assign new_n23838_ = ~new_n3780_;
  assign new_n23839_ = ~new_n3780_ | ~new_n23854_;
  assign new_n23840_ = ~new_n3781_;
  assign new_n23841_ = ~new_n3781_ | ~new_n23855_;
  assign new_n23842_ = ~new_n3782_;
  assign new_n23843_ = ~new_n3782_ | ~new_n23856_;
  assign new_n23844_ = ~new_n3784_;
  assign new_n23845_ = ~new_n3783_;
  assign new_n23846_ = ~new_n23860_ | ~new_n23859_;
  assign new_n23847_ = ~new_n23862_ | ~new_n23861_;
  assign new_n23848_ = ~new_n23864_ | ~new_n23863_;
  assign new_n23849_ = ~new_n23866_ | ~new_n23865_;
  assign new_n23850_ = ~new_n23868_ | ~new_n23867_;
  assign new_n23851_ = ~new_n23870_ | ~new_n23869_;
  assign new_n23852_ = new_n3784_ & new_n3783_;
  assign new_n23853_ = ~new_n3783_ | ~new_n23857_;
  assign new_n23854_ = ~new_n23837_;
  assign new_n23855_ = ~new_n23839_;
  assign new_n23856_ = ~new_n23841_;
  assign new_n23857_ = ~new_n23843_;
  assign new_n23858_ = ~new_n23853_;
  assign new_n23859_ = ~new_n3784_ | ~new_n23853_;
  assign new_n23860_ = ~new_n23858_ | ~new_n23844_;
  assign new_n23861_ = ~new_n3783_ | ~new_n23843_;
  assign new_n23862_ = ~new_n23857_ | ~new_n23845_;
  assign new_n23863_ = ~new_n3782_ | ~new_n23841_;
  assign new_n23864_ = ~new_n23856_ | ~new_n23842_;
  assign new_n23865_ = ~new_n3781_ | ~new_n23839_;
  assign new_n23866_ = ~new_n23855_ | ~new_n23840_;
  assign new_n23867_ = ~new_n3780_ | ~new_n23837_;
  assign new_n23868_ = ~new_n23854_ | ~new_n23838_;
  assign new_n23869_ = ~new_n3779_ | ~new_n23834_;
  assign new_n23870_ = ~new_n3778_ | ~new_n23836_;
  assign new_n23871_ = ~pi0307;
  assign new_n23872_ = ~new_n23876_ | ~new_n23875_;
  assign new_n23873_ = ~pi0318;
  assign new_n23874_ = ~pi0317;
  assign new_n23875_ = ~pi0318 | ~new_n23874_;
  assign new_n23876_ = ~pi0317 | ~new_n23873_;
  assign new_n23877_ = new_n23879_ | new_n3785_;
  assign new_n23878_ = new_n22897_ & new_n22896_;
  assign new_n23879_ = ~new_n22898_ & ~new_n22899_ & ~new_n23878_;
  assign new_n23880_ = ~pi0318;
  assign new_n23881_ = ~pi0319;
  assign new_n23882_ = ~pi0319 | ~pi0318;
  assign new_n23883_ = ~pi0320;
  assign new_n23884_ = ~pi0320 | ~new_n23970_;
  assign new_n23885_ = ~pi0321;
  assign new_n23886_ = ~pi0321 | ~new_n23971_;
  assign new_n23887_ = ~pi0322;
  assign new_n23888_ = ~pi0322 | ~new_n23972_;
  assign new_n23889_ = ~pi0323;
  assign new_n23890_ = ~pi0323 | ~new_n23973_;
  assign new_n23891_ = ~pi0324;
  assign new_n23892_ = ~pi0324 | ~new_n23974_;
  assign new_n23893_ = ~pi0325;
  assign new_n23894_ = ~pi0326;
  assign new_n23895_ = ~pi0325 | ~new_n23975_;
  assign new_n23896_ = ~new_n23976_ | ~pi0326;
  assign new_n23897_ = ~pi0327;
  assign new_n23898_ = ~pi0327 | ~new_n23977_;
  assign new_n23899_ = ~pi0328;
  assign new_n23900_ = ~pi0328 | ~new_n23978_;
  assign new_n23901_ = ~pi0329;
  assign new_n23902_ = ~pi0329 | ~new_n23979_;
  assign new_n23903_ = ~pi0330;
  assign new_n23904_ = ~pi0330 | ~new_n23980_;
  assign new_n23905_ = ~pi0331;
  assign new_n23906_ = ~pi0331 | ~new_n23981_;
  assign new_n23907_ = ~pi0332;
  assign new_n23908_ = ~pi0332 | ~new_n23982_;
  assign new_n23909_ = ~pi0333;
  assign new_n23910_ = ~pi0333 | ~new_n23983_;
  assign new_n23911_ = ~pi0334;
  assign new_n23912_ = ~pi0334 | ~new_n23984_;
  assign new_n23913_ = ~pi0335;
  assign new_n23914_ = ~pi0335 | ~new_n23985_;
  assign new_n23915_ = ~pi0336;
  assign new_n23916_ = ~pi0336 | ~new_n23986_;
  assign new_n23917_ = ~pi0337;
  assign new_n23918_ = ~pi0337 | ~new_n23987_;
  assign new_n23919_ = ~pi0338;
  assign new_n23920_ = ~pi0338 | ~new_n23988_;
  assign new_n23921_ = ~pi0339;
  assign new_n23922_ = ~pi0339 | ~new_n23989_;
  assign new_n23923_ = ~pi0340;
  assign new_n23924_ = ~pi0340 | ~new_n23990_;
  assign new_n23925_ = ~pi0341;
  assign new_n23926_ = ~pi0341 | ~new_n23991_;
  assign new_n23927_ = ~pi0342;
  assign new_n23928_ = ~pi0342 | ~new_n23992_;
  assign new_n23929_ = ~pi0343;
  assign new_n23930_ = ~pi0343 | ~new_n23993_;
  assign new_n23931_ = ~pi0344;
  assign new_n23932_ = ~pi0344 | ~new_n23994_;
  assign new_n23933_ = ~pi0345;
  assign new_n23934_ = ~pi0345 | ~new_n23995_;
  assign new_n23935_ = ~pi0346;
  assign new_n23936_ = ~pi0346 | ~new_n23996_;
  assign new_n23937_ = ~pi0347;
  assign new_n23938_ = ~new_n24000_ | ~new_n23999_;
  assign new_n23939_ = ~new_n24002_ | ~new_n24001_;
  assign new_n23940_ = ~new_n24004_ | ~new_n24003_;
  assign new_n23941_ = ~new_n24006_ | ~new_n24005_;
  assign new_n23942_ = ~new_n24008_ | ~new_n24007_;
  assign new_n23943_ = ~new_n24010_ | ~new_n24009_;
  assign new_n23944_ = ~new_n24012_ | ~new_n24011_;
  assign new_n23945_ = ~new_n24014_ | ~new_n24013_;
  assign new_n23946_ = ~new_n24016_ | ~new_n24015_;
  assign new_n23947_ = ~new_n24018_ | ~new_n24017_;
  assign new_n23948_ = ~new_n24020_ | ~new_n24019_;
  assign new_n23949_ = ~new_n24022_ | ~new_n24021_;
  assign new_n23950_ = ~new_n24024_ | ~new_n24023_;
  assign new_n23951_ = ~new_n24026_ | ~new_n24025_;
  assign new_n23952_ = ~new_n24028_ | ~new_n24027_;
  assign new_n23953_ = ~new_n24030_ | ~new_n24029_;
  assign new_n23954_ = ~new_n24032_ | ~new_n24031_;
  assign new_n23955_ = ~new_n24034_ | ~new_n24033_;
  assign new_n23956_ = ~new_n24036_ | ~new_n24035_;
  assign new_n23957_ = ~new_n24038_ | ~new_n24037_;
  assign new_n23958_ = ~new_n24040_ | ~new_n24039_;
  assign new_n23959_ = ~new_n24042_ | ~new_n24041_;
  assign new_n23960_ = ~new_n24044_ | ~new_n24043_;
  assign new_n23961_ = ~new_n24046_ | ~new_n24045_;
  assign new_n23962_ = ~new_n24048_ | ~new_n24047_;
  assign new_n23963_ = ~new_n24050_ | ~new_n24049_;
  assign new_n23964_ = ~new_n24052_ | ~new_n24051_;
  assign new_n23965_ = ~new_n24054_ | ~new_n24053_;
  assign new_n23966_ = ~new_n24056_ | ~new_n24055_;
  assign new_n23967_ = ~new_n24058_ | ~new_n24057_;
  assign new_n23968_ = ~pi0348;
  assign new_n23969_ = ~pi0347 | ~new_n23997_;
  assign new_n23970_ = ~new_n23882_;
  assign new_n23971_ = ~new_n23884_;
  assign new_n23972_ = ~new_n23886_;
  assign new_n23973_ = ~new_n23888_;
  assign new_n23974_ = ~new_n23890_;
  assign new_n23975_ = ~new_n23892_;
  assign new_n23976_ = ~new_n23895_;
  assign new_n23977_ = ~new_n23896_;
  assign new_n23978_ = ~new_n23898_;
  assign new_n23979_ = ~new_n23900_;
  assign new_n23980_ = ~new_n23902_;
  assign new_n23981_ = ~new_n23904_;
  assign new_n23982_ = ~new_n23906_;
  assign new_n23983_ = ~new_n23908_;
  assign new_n23984_ = ~new_n23910_;
  assign new_n23985_ = ~new_n23912_;
  assign new_n23986_ = ~new_n23914_;
  assign new_n23987_ = ~new_n23916_;
  assign new_n23988_ = ~new_n23918_;
  assign new_n23989_ = ~new_n23920_;
  assign new_n23990_ = ~new_n23922_;
  assign new_n23991_ = ~new_n23924_;
  assign new_n23992_ = ~new_n23926_;
  assign new_n23993_ = ~new_n23928_;
  assign new_n23994_ = ~new_n23930_;
  assign new_n23995_ = ~new_n23932_;
  assign new_n23996_ = ~new_n23934_;
  assign new_n23997_ = ~new_n23936_;
  assign new_n23998_ = ~new_n23969_;
  assign new_n23999_ = ~pi0326 | ~new_n23895_;
  assign new_n24000_ = ~new_n23976_ | ~new_n23894_;
  assign new_n24001_ = ~pi0325 | ~new_n23892_;
  assign new_n24002_ = ~new_n23975_ | ~new_n23893_;
  assign new_n24003_ = ~pi0324 | ~new_n23890_;
  assign new_n24004_ = ~new_n23974_ | ~new_n23891_;
  assign new_n24005_ = ~pi0323 | ~new_n23888_;
  assign new_n24006_ = ~new_n23973_ | ~new_n23889_;
  assign new_n24007_ = ~pi0322 | ~new_n23886_;
  assign new_n24008_ = ~new_n23972_ | ~new_n23887_;
  assign new_n24009_ = ~pi0321 | ~new_n23884_;
  assign new_n24010_ = ~new_n23971_ | ~new_n23885_;
  assign new_n24011_ = ~pi0320 | ~new_n23882_;
  assign new_n24012_ = ~new_n23970_ | ~new_n23883_;
  assign new_n24013_ = ~pi0348 | ~new_n23969_;
  assign new_n24014_ = ~new_n23998_ | ~new_n23968_;
  assign new_n24015_ = ~pi0347 | ~new_n23936_;
  assign new_n24016_ = ~new_n23997_ | ~new_n23937_;
  assign new_n24017_ = ~pi0319 | ~new_n23880_;
  assign new_n24018_ = ~pi0318 | ~new_n23881_;
  assign new_n24019_ = ~pi0346 | ~new_n23934_;
  assign new_n24020_ = ~new_n23996_ | ~new_n23935_;
  assign new_n24021_ = ~pi0345 | ~new_n23932_;
  assign new_n24022_ = ~new_n23995_ | ~new_n23933_;
  assign new_n24023_ = ~pi0344 | ~new_n23930_;
  assign new_n24024_ = ~new_n23994_ | ~new_n23931_;
  assign new_n24025_ = ~pi0343 | ~new_n23928_;
  assign new_n24026_ = ~new_n23993_ | ~new_n23929_;
  assign new_n24027_ = ~pi0342 | ~new_n23926_;
  assign new_n24028_ = ~new_n23992_ | ~new_n23927_;
  assign new_n24029_ = ~pi0341 | ~new_n23924_;
  assign new_n24030_ = ~new_n23991_ | ~new_n23925_;
  assign new_n24031_ = ~pi0340 | ~new_n23922_;
  assign new_n24032_ = ~new_n23990_ | ~new_n23923_;
  assign new_n24033_ = ~pi0339 | ~new_n23920_;
  assign new_n24034_ = ~new_n23989_ | ~new_n23921_;
  assign new_n24035_ = ~pi0338 | ~new_n23918_;
  assign new_n24036_ = ~new_n23988_ | ~new_n23919_;
  assign new_n24037_ = ~pi0337 | ~new_n23916_;
  assign new_n24038_ = ~new_n23987_ | ~new_n23917_;
  assign new_n24039_ = ~pi0336 | ~new_n23914_;
  assign new_n24040_ = ~new_n23986_ | ~new_n23915_;
  assign new_n24041_ = ~pi0335 | ~new_n23912_;
  assign new_n24042_ = ~new_n23985_ | ~new_n23913_;
  assign new_n24043_ = ~pi0334 | ~new_n23910_;
  assign new_n24044_ = ~new_n23984_ | ~new_n23911_;
  assign new_n24045_ = ~pi0333 | ~new_n23908_;
  assign new_n24046_ = ~new_n23983_ | ~new_n23909_;
  assign new_n24047_ = ~pi0332 | ~new_n23906_;
  assign new_n24048_ = ~new_n23982_ | ~new_n23907_;
  assign new_n24049_ = ~pi0331 | ~new_n23904_;
  assign new_n24050_ = ~new_n23981_ | ~new_n23905_;
  assign new_n24051_ = ~pi0330 | ~new_n23902_;
  assign new_n24052_ = ~new_n23980_ | ~new_n23903_;
  assign new_n24053_ = ~pi0329 | ~new_n23900_;
  assign new_n24054_ = ~new_n23979_ | ~new_n23901_;
  assign new_n24055_ = ~pi0328 | ~new_n23898_;
  assign new_n24056_ = ~new_n23978_ | ~new_n23899_;
  assign new_n24057_ = ~pi0327 | ~new_n23896_;
  assign new_n24058_ = ~new_n23977_ | ~new_n23897_;
  assign new_n24059_ = ~new_n24098_ | ~new_n24097_;
  assign new_n24060_ = ~new_n24062_ | ~new_n24099_;
  assign new_n24061_ = ~pi0311;
  assign new_n24062_ = ~pi0311 | ~new_n24071_;
  assign new_n24063_ = ~pi0315;
  assign new_n24064_ = ~pi0309;
  assign new_n24065_ = ~pi0314;
  assign new_n24066_ = ~pi0308;
  assign new_n24067_ = ~pi0313;
  assign new_n24068_ = ~pi0312;
  assign new_n24069_ = ~new_n24094_ | ~new_n24093_;
  assign new_n24070_ = ~pi0307;
  assign new_n24071_ = ~pi0316;
  assign new_n24072_ = ~new_n24104_ | ~new_n24103_;
  assign new_n24073_ = ~new_n24109_ | ~new_n24108_;
  assign new_n24074_ = ~new_n24114_ | ~new_n24113_;
  assign new_n24075_ = ~new_n24119_ | ~new_n24118_;
  assign new_n24076_ = ~new_n24101_ | ~new_n24100_;
  assign new_n24077_ = ~new_n24106_ | ~new_n24105_;
  assign new_n24078_ = ~new_n24111_ | ~new_n24110_;
  assign new_n24079_ = ~new_n24116_ | ~new_n24115_;
  assign new_n24080_ = ~new_n24090_ | ~new_n24089_;
  assign new_n24081_ = ~new_n24086_ | ~new_n24085_;
  assign new_n24082_ = ~pi0310;
  assign new_n24083_ = ~new_n24062_;
  assign new_n24084_ = ~new_n24083_ | ~new_n24063_;
  assign new_n24085_ = ~new_n24084_ | ~new_n24082_;
  assign new_n24086_ = ~pi0315 | ~new_n24062_;
  assign new_n24087_ = ~new_n24081_;
  assign new_n24088_ = ~pi0309 | ~new_n24065_;
  assign new_n24089_ = ~new_n24088_ | ~new_n24081_;
  assign new_n24090_ = ~pi0314 | ~new_n24064_;
  assign new_n24091_ = ~new_n24080_;
  assign new_n24092_ = ~pi0308 | ~new_n24067_;
  assign new_n24093_ = ~new_n24092_ | ~new_n24080_;
  assign new_n24094_ = ~pi0313 | ~new_n24066_;
  assign new_n24095_ = ~new_n24069_;
  assign new_n24096_ = ~pi0312 | ~new_n24070_;
  assign new_n24097_ = ~new_n24095_ | ~new_n24096_;
  assign new_n24098_ = ~pi0307 | ~new_n24068_;
  assign new_n24099_ = ~pi0316 | ~new_n24061_;
  assign new_n24100_ = ~pi0307 | ~new_n24068_;
  assign new_n24101_ = ~pi0312 | ~new_n24070_;
  assign new_n24102_ = ~new_n24076_;
  assign new_n24103_ = ~new_n24102_ | ~new_n24095_;
  assign new_n24104_ = ~new_n24076_ | ~new_n24069_;
  assign new_n24105_ = ~pi0308 | ~new_n24067_;
  assign new_n24106_ = ~pi0313 | ~new_n24066_;
  assign new_n24107_ = ~new_n24077_;
  assign new_n24108_ = ~new_n24091_ | ~new_n24107_;
  assign new_n24109_ = ~new_n24077_ | ~new_n24080_;
  assign new_n24110_ = ~pi0309 | ~new_n24065_;
  assign new_n24111_ = ~pi0314 | ~new_n24064_;
  assign new_n24112_ = ~new_n24078_;
  assign new_n24113_ = ~new_n24087_ | ~new_n24112_;
  assign new_n24114_ = ~new_n24078_ | ~new_n24081_;
  assign new_n24115_ = ~pi0310 | ~new_n24063_;
  assign new_n24116_ = ~pi0315 | ~new_n24082_;
  assign new_n24117_ = ~new_n24079_;
  assign new_n24118_ = ~new_n24117_ | ~new_n24083_;
  assign new_n24119_ = ~new_n24079_ | ~new_n24062_;
  assign new_n24120_ = ~new_n24157_ | ~new_n24156_;
  assign new_n24121_ = ~pi0311 | ~new_n24141_;
  assign new_n24122_ = ~pi0315;
  assign new_n24123_ = ~pi0309;
  assign new_n24124_ = ~pi0314;
  assign new_n24125_ = ~pi0308;
  assign new_n24126_ = ~pi0313;
  assign new_n24127_ = ~pi0312;
  assign new_n24128_ = ~new_n24153_ | ~new_n24152_;
  assign new_n24129_ = ~pi0307;
  assign new_n24130_ = ~new_n24162_ | ~new_n24161_;
  assign new_n24131_ = ~new_n24167_ | ~new_n24166_;
  assign new_n24132_ = ~new_n24172_ | ~new_n24171_;
  assign new_n24133_ = ~new_n24177_ | ~new_n24176_;
  assign new_n24134_ = ~new_n24159_ | ~new_n24158_;
  assign new_n24135_ = ~new_n24164_ | ~new_n24163_;
  assign new_n24136_ = ~new_n24169_ | ~new_n24168_;
  assign new_n24137_ = ~new_n24174_ | ~new_n24173_;
  assign new_n24138_ = ~new_n24149_ | ~new_n24148_;
  assign new_n24139_ = ~new_n24145_ | ~new_n24144_;
  assign new_n24140_ = ~pi0310;
  assign new_n24141_ = ~pi0316;
  assign new_n24142_ = ~new_n24121_;
  assign new_n24143_ = ~new_n24142_ | ~new_n24122_;
  assign new_n24144_ = ~new_n24143_ | ~new_n24140_;
  assign new_n24145_ = ~pi0315 | ~new_n24121_;
  assign new_n24146_ = ~new_n24139_;
  assign new_n24147_ = ~pi0309 | ~new_n24124_;
  assign new_n24148_ = ~new_n24147_ | ~new_n24139_;
  assign new_n24149_ = ~pi0314 | ~new_n24123_;
  assign new_n24150_ = ~new_n24138_;
  assign new_n24151_ = ~pi0308 | ~new_n24126_;
  assign new_n24152_ = ~new_n24151_ | ~new_n24138_;
  assign new_n24153_ = ~pi0313 | ~new_n24125_;
  assign new_n24154_ = ~new_n24128_;
  assign new_n24155_ = ~pi0312 | ~new_n24129_;
  assign new_n24156_ = ~new_n24154_ | ~new_n24155_;
  assign new_n24157_ = ~pi0307 | ~new_n24127_;
  assign new_n24158_ = ~pi0307 | ~new_n24127_;
  assign new_n24159_ = ~pi0312 | ~new_n24129_;
  assign new_n24160_ = ~new_n24134_;
  assign new_n24161_ = ~new_n24160_ | ~new_n24154_;
  assign new_n24162_ = ~new_n24134_ | ~new_n24128_;
  assign new_n24163_ = ~pi0308 | ~new_n24126_;
  assign new_n24164_ = ~pi0313 | ~new_n24125_;
  assign new_n24165_ = ~new_n24135_;
  assign new_n24166_ = ~new_n24150_ | ~new_n24165_;
  assign new_n24167_ = ~new_n24135_ | ~new_n24138_;
  assign new_n24168_ = ~pi0309 | ~new_n24124_;
  assign new_n24169_ = ~pi0314 | ~new_n24123_;
  assign new_n24170_ = ~new_n24136_;
  assign new_n24171_ = ~new_n24146_ | ~new_n24170_;
  assign new_n24172_ = ~new_n24136_ | ~new_n24139_;
  assign new_n24173_ = ~pi0310 | ~new_n24122_;
  assign new_n24174_ = ~pi0315 | ~new_n24140_;
  assign new_n24175_ = ~new_n24137_;
  assign new_n24176_ = ~new_n24175_ | ~new_n24142_;
  assign new_n24177_ = ~new_n24137_ | ~new_n24121_;
  assign new_n24178_ = pi0344 & pi0345;
  assign new_n24179_ = new_n24362_ & new_n24360_;
  assign new_n24180_ = new_n24361_ & new_n24352_;
  assign new_n24181_ = new_n24180_ & new_n24363_;
  assign new_n24182_ = new_n24179_ & new_n24364_;
  assign new_n24183_ = new_n24383_ & new_n24378_;
  assign new_n24184_ = new_n24379_ & new_n24330_ & new_n24380_ & new_n24384_;
  assign new_n24185_ = new_n24183_ & new_n24385_;
  assign new_n24186_ = new_n24184_ & new_n24386_;
  assign new_n24187_ = new_n24185_ & new_n24387_;
  assign new_n24188_ = new_n24186_ & new_n24388_;
  assign new_n24189_ = new_n24429_ & new_n24426_;
  assign new_n24190_ = new_n24423_ & new_n24422_;
  assign new_n24191_ = new_n24418_ & new_n24415_;
  assign new_n24192_ = new_n24407_ & new_n24404_;
  assign new_n24193_ = new_n24401_ & new_n24477_;
  assign new_n24194_ = new_n24399_ & new_n24470_;
  assign new_n24195_ = ~new_n24481_ | ~new_n24600_ | ~new_n24599_;
  assign new_n24196_ = ~new_n26366_;
  assign new_n24197_ = ~pi0324;
  assign new_n24198_ = ~new_n26365_;
  assign new_n24199_ = ~pi0322;
  assign new_n24200_ = ~new_n26376_;
  assign new_n24201_ = ~pi0321;
  assign new_n24202_ = ~new_n26367_;
  assign new_n24203_ = ~pi0317;
  assign new_n24204_ = ~pi0317 | ~new_n26367_;
  assign new_n24205_ = ~new_n27120_;
  assign new_n24206_ = ~new_n26370_;
  assign new_n24207_ = ~pi0319;
  assign new_n24208_ = ~pi0318;
  assign new_n24209_ = ~new_n26364_;
  assign new_n24210_ = ~pi0320;
  assign new_n24211_ = ~new_n26374_;
  assign new_n24212_ = ~pi0323;
  assign new_n24213_ = ~new_n26363_;
  assign new_n24214_ = ~pi0325;
  assign new_n24215_ = ~pi0326;
  assign new_n24216_ = ~pi0342;
  assign new_n24217_ = ~pi0343;
  assign new_n24218_ = ~pi0341;
  assign new_n24219_ = ~pi0340;
  assign new_n24220_ = ~pi0339;
  assign new_n24221_ = ~pi0336;
  assign new_n24222_ = ~pi0338;
  assign new_n24223_ = ~pi0335;
  assign new_n24224_ = ~pi0329;
  assign new_n24225_ = ~pi0330;
  assign new_n24226_ = ~pi0328;
  assign new_n24227_ = ~pi0327;
  assign new_n24228_ = ~pi0331;
  assign new_n24229_ = ~pi0332;
  assign new_n24230_ = ~pi0333;
  assign new_n24231_ = ~pi0336 | ~pi0337;
  assign new_n24232_ = ~pi0344;
  assign new_n24233_ = ~pi0346;
  assign new_n24234_ = ~pi0347;
  assign new_n24235_ = ~new_n24443_ | ~new_n24396_ | ~new_n24325_;
  assign new_n24236_ = ~new_n24279_ | ~new_n24392_;
  assign new_n24237_ = ~new_n24278_ | ~new_n24458_;
  assign new_n24238_ = ~new_n24450_ | ~new_n24379_;
  assign new_n24239_ = ~new_n24451_ | ~new_n24221_;
  assign new_n24240_ = ~new_n27120_ | ~new_n24335_;
  assign new_n24241_ = ~new_n24276_ | ~new_n24372_;
  assign new_n24242_ = ~new_n24464_ | ~new_n24182_;
  assign new_n24243_ = ~new_n24658_ | ~new_n24657_;
  assign new_n24244_ = ~new_n24486_ | ~new_n24485_;
  assign new_n24245_ = ~new_n24493_ | ~new_n24492_;
  assign new_n24246_ = ~new_n24500_ | ~new_n24499_;
  assign new_n24247_ = ~new_n24507_ | ~new_n24506_;
  assign new_n24248_ = ~new_n24514_ | ~new_n24513_;
  assign new_n24249_ = ~new_n24519_ | ~new_n24518_;
  assign new_n24250_ = ~new_n24524_ | ~new_n24523_;
  assign new_n24251_ = ~new_n24535_ | ~new_n24534_;
  assign new_n24252_ = ~new_n24540_ | ~new_n24539_;
  assign new_n24253_ = ~new_n24547_ | ~new_n24546_;
  assign new_n24254_ = ~new_n24558_ | ~new_n24557_;
  assign new_n24255_ = ~new_n24565_ | ~new_n24564_;
  assign new_n24256_ = ~new_n24572_ | ~new_n24571_;
  assign new_n24257_ = ~new_n24579_ | ~new_n24578_;
  assign new_n24258_ = ~new_n24586_ | ~new_n24585_;
  assign new_n24259_ = ~new_n24593_ | ~new_n24592_;
  assign new_n24260_ = ~new_n24605_ | ~new_n24604_;
  assign new_n24261_ = ~new_n24612_ | ~new_n24611_;
  assign new_n24262_ = ~new_n24623_ | ~new_n24622_;
  assign new_n24263_ = ~new_n24630_ | ~new_n24629_;
  assign new_n24264_ = ~new_n24637_ | ~new_n24636_;
  assign new_n24265_ = ~new_n24644_ | ~new_n24643_;
  assign new_n24266_ = ~new_n24651_ | ~new_n24650_;
  assign new_n24267_ = ~new_n24656_ | ~new_n24655_;
  assign new_n24268_ = new_n24334_ & new_n24337_ & new_n24338_;
  assign new_n24269_ = new_n26364_ & pi0320;
  assign new_n24270_ = new_n24342_ & new_n24336_;
  assign new_n24271_ = new_n24338_ & new_n24337_;
  assign new_n24272_ = new_n24181_ & new_n24328_;
  assign new_n24273_ = new_n24366_ & new_n24329_;
  assign new_n24274_ = new_n24273_ & new_n24182_;
  assign new_n24275_ = pi0334 & pi0333;
  assign new_n24276_ = new_n24373_ & new_n24230_;
  assign new_n24277_ = new_n24389_ & new_n24187_;
  assign new_n24278_ = new_n24188_ & new_n24390_;
  assign new_n24279_ = new_n24393_ & new_n24331_ & new_n24232_;
  assign new_n24280_ = new_n24393_ & new_n24331_;
  assign new_n24281_ = new_n24443_ & pi0348 & new_n24234_;
  assign new_n24282_ = pi0347 & pi0348;
  assign new_n24283_ = new_n24331_ & new_n24560_ & new_n24559_;
  assign new_n24284_ = new_n24406_ & new_n24327_;
  assign new_n24285_ = new_n24411_ & new_n24330_;
  assign new_n24286_ = new_n24417_ & new_n24330_;
  assign new_n24287_ = new_n24329_ & new_n24639_ & new_n24638_;
  assign new_n24288_ = new_n24428_ & new_n24328_;
  assign new_n24289_ = ~new_n24442_ | ~new_n24350_ | ~new_n24326_;
  assign new_n24290_ = new_n24488_ & new_n24487_;
  assign new_n24291_ = ~new_n24474_ | ~new_n24441_;
  assign new_n24292_ = new_n24495_ & new_n24494_;
  assign new_n24293_ = ~new_n24347_ | ~new_n24346_;
  assign new_n24294_ = new_n24502_ & new_n24501_;
  assign new_n24295_ = ~new_n24472_ | ~new_n24440_;
  assign new_n24296_ = new_n24509_ & new_n24508_;
  assign new_n24297_ = ~new_n24270_ | ~new_n24341_;
  assign new_n24298_ = ~new_n24355_ | ~new_n24354_;
  assign new_n24299_ = ~new_n24333_ | ~new_n24357_;
  assign new_n24300_ = new_n24530_ & new_n24529_;
  assign new_n24301_ = ~new_n24445_ | ~new_n24444_ | ~new_n24240_;
  assign new_n24302_ = new_n24542_ & new_n24541_;
  assign new_n24303_ = ~new_n24478_ | ~new_n24449_ | ~new_n24448_;
  assign new_n24304_ = new_n24553_ & new_n24552_;
  assign new_n24305_ = ~new_n24280_ | ~new_n24392_;
  assign new_n24306_ = new_n24567_ & new_n24566_;
  assign new_n24307_ = ~new_n24456_ | ~new_n24188_;
  assign new_n24308_ = new_n24574_ & new_n24573_;
  assign new_n24309_ = ~new_n24454_ | ~new_n24186_;
  assign new_n24310_ = new_n24581_ & new_n24580_;
  assign new_n24311_ = ~new_n24452_ | ~new_n24184_;
  assign new_n24312_ = new_n24588_ & new_n24587_;
  assign new_n24313_ = ~new_n24285_ | ~new_n24410_;
  assign new_n24314_ = new_n24607_ & new_n24606_;
  assign new_n24315_ = ~new_n24447_ | ~new_n24446_ | ~new_n24375_;
  assign new_n24316_ = new_n24618_ & new_n24617_;
  assign new_n24317_ = ~new_n24373_ | ~new_n24372_;
  assign new_n24318_ = new_n24625_ & new_n24624_;
  assign new_n24319_ = ~new_n24369_ | ~new_n24368_;
  assign new_n24320_ = new_n24632_ & new_n24631_;
  assign new_n24321_ = ~new_n24274_ | ~new_n24466_;
  assign new_n24322_ = new_n24646_ & new_n24645_;
  assign new_n24323_ = ~new_n24462_ | ~new_n24179_;
  assign new_n24324_ = ~new_n24460_ | ~new_n24360_;
  assign new_n24325_ = ~new_n26363_ | ~new_n24303_;
  assign new_n24326_ = ~new_n26363_ | ~new_n24291_;
  assign new_n24327_ = ~new_n24391_ | ~new_n24213_;
  assign new_n24328_ = ~new_n24365_ | ~new_n24213_;
  assign new_n24329_ = ~pi0329 | ~new_n26363_;
  assign new_n24330_ = ~pi0337 | ~new_n26363_;
  assign new_n24331_ = ~pi0342 | ~new_n26363_;
  assign new_n24332_ = ~new_n24240_;
  assign new_n24333_ = ~pi0319 | ~new_n26370_;
  assign new_n24334_ = pi0321 | new_n26376_;
  assign new_n24335_ = ~new_n24204_;
  assign new_n24336_ = ~pi0321 | ~new_n26376_;
  assign new_n24337_ = new_n26364_ | pi0320;
  assign new_n24338_ = new_n26370_ | pi0319;
  assign new_n24339_ = ~new_n24301_;
  assign new_n24340_ = ~new_n24444_ | ~new_n24240_ | ~new_n24333_ | ~new_n24445_;
  assign new_n24341_ = ~new_n24268_ | ~new_n24340_;
  assign new_n24342_ = ~new_n24269_ | ~new_n24334_;
  assign new_n24343_ = ~new_n24297_;
  assign new_n24344_ = pi0322 | new_n26365_;
  assign new_n24345_ = new_n26374_ | pi0323;
  assign new_n24346_ = ~new_n24345_ | ~new_n24295_;
  assign new_n24347_ = ~pi0323 | ~new_n26374_;
  assign new_n24348_ = ~new_n24293_;
  assign new_n24349_ = pi0324 | new_n26366_;
  assign new_n24350_ = ~pi0325 | ~new_n24291_;
  assign new_n24351_ = ~new_n24289_;
  assign new_n24352_ = pi0326 | new_n26363_;
  assign new_n24353_ = ~pi0326 | ~new_n26363_;
  assign new_n24354_ = ~new_n24271_ | ~new_n24340_;
  assign new_n24355_ = ~pi0320 | ~new_n26364_;
  assign new_n24356_ = ~new_n24298_;
  assign new_n24357_ = ~new_n24301_ | ~new_n24338_;
  assign new_n24358_ = ~new_n24299_;
  assign new_n24359_ = ~pi0320 | ~new_n26364_;
  assign new_n24360_ = ~pi0326 | ~new_n26363_;
  assign new_n24361_ = new_n26363_ | pi0327;
  assign new_n24362_ = ~pi0327 | ~new_n26363_;
  assign new_n24363_ = new_n26363_ | pi0328;
  assign new_n24364_ = ~pi0328 | ~new_n26363_;
  assign new_n24365_ = ~pi0330 | ~pi0329;
  assign new_n24366_ = ~pi0330 | ~new_n26363_;
  assign new_n24367_ = new_n26363_ | pi0331;
  assign new_n24368_ = ~new_n24367_ | ~new_n24321_;
  assign new_n24369_ = ~pi0331 | ~new_n26363_;
  assign new_n24370_ = ~new_n24319_;
  assign new_n24371_ = new_n26363_ | pi0332;
  assign new_n24372_ = ~new_n24371_ | ~new_n24319_;
  assign new_n24373_ = ~pi0332 | ~new_n26363_;
  assign new_n24374_ = ~new_n24317_;
  assign new_n24375_ = ~new_n24275_ | ~new_n24317_;
  assign new_n24376_ = ~new_n24241_;
  assign new_n24377_ = ~new_n24315_;
  assign new_n24378_ = new_n26363_ | pi0335;
  assign new_n24379_ = ~pi0335 | ~new_n26363_;
  assign new_n24380_ = ~pi0336 | ~new_n26363_;
  assign new_n24381_ = ~new_n24231_;
  assign new_n24382_ = ~new_n24381_ | ~pi0338;
  assign new_n24383_ = ~new_n24213_ | ~new_n24382_;
  assign new_n24384_ = ~pi0338 | ~new_n26363_;
  assign new_n24385_ = new_n26363_ | pi0339;
  assign new_n24386_ = ~pi0339 | ~new_n26363_;
  assign new_n24387_ = new_n26363_ | pi0340;
  assign new_n24388_ = ~pi0340 | ~new_n26363_;
  assign new_n24389_ = new_n26363_ | pi0341;
  assign new_n24390_ = ~pi0341 | ~new_n26363_;
  assign new_n24391_ = ~pi0343 | ~pi0342;
  assign new_n24392_ = ~new_n24237_ | ~new_n24327_;
  assign new_n24393_ = ~pi0343 | ~new_n26363_;
  assign new_n24394_ = ~new_n24305_;
  assign new_n24395_ = ~new_n24236_;
  assign new_n24396_ = ~pi0346 | ~new_n24303_;
  assign new_n24397_ = ~new_n24235_;
  assign new_n24398_ = ~new_n24325_ | ~new_n24281_;
  assign new_n24399_ = ~new_n24468_ | ~new_n24528_ | ~new_n24527_;
  assign new_n24400_ = ~new_n24395_ | ~pi0345;
  assign new_n24401_ = ~new_n24236_ | ~new_n24551_ | ~new_n24550_;
  assign new_n24402_ = new_n26363_ | pi0342;
  assign new_n24403_ = ~new_n24402_ | ~new_n24237_;
  assign new_n24404_ = ~new_n24283_ | ~new_n24403_;
  assign new_n24405_ = ~new_n24459_ | ~new_n24331_;
  assign new_n24406_ = ~pi0343 | ~new_n26363_;
  assign new_n24407_ = ~new_n24284_ | ~new_n24405_;
  assign new_n24408_ = pi0342 | new_n26363_;
  assign new_n24409_ = ~new_n24239_;
  assign new_n24410_ = ~new_n26363_ | ~new_n24239_;
  assign new_n24411_ = ~new_n24381_ | ~new_n24238_;
  assign new_n24412_ = ~new_n24313_;
  assign new_n24413_ = ~new_n24409_ | ~pi0337;
  assign new_n24414_ = ~pi0336 | ~new_n24238_;
  assign new_n24415_ = ~new_n24414_ | ~new_n24595_ | ~new_n24594_;
  assign new_n24416_ = ~new_n24451_ | ~new_n24380_;
  assign new_n24417_ = ~new_n24231_ | ~new_n24213_;
  assign new_n24418_ = ~new_n24286_ | ~new_n24416_;
  assign new_n24419_ = pi0336 | new_n26363_;
  assign new_n24420_ = ~new_n24376_ | ~pi0334;
  assign new_n24421_ = ~pi0333 | ~new_n24317_;
  assign new_n24422_ = ~new_n24421_ | ~new_n24614_ | ~new_n24613_;
  assign new_n24423_ = ~new_n24241_ | ~new_n24616_ | ~new_n24615_;
  assign new_n24424_ = new_n26363_ | pi0329;
  assign new_n24425_ = ~new_n24424_ | ~new_n24242_;
  assign new_n24426_ = ~new_n24287_ | ~new_n24425_;
  assign new_n24427_ = ~new_n24465_ | ~new_n24329_;
  assign new_n24428_ = ~pi0330 | ~new_n26363_;
  assign new_n24429_ = ~new_n24288_ | ~new_n24427_;
  assign new_n24430_ = pi0329 | new_n26363_;
  assign new_n24431_ = ~pi0327 | ~new_n26363_;
  assign new_n24432_ = ~new_n24353_ | ~new_n24352_;
  assign new_n24433_ = ~new_n24336_ | ~new_n24334_;
  assign new_n24434_ = ~new_n24359_ | ~new_n24337_;
  assign new_n24435_ = ~new_n24338_ | ~new_n24333_;
  assign new_n24436_ = ~new_n24408_ | ~new_n24331_;
  assign new_n24437_ = ~new_n24419_ | ~new_n24380_;
  assign new_n24438_ = ~new_n24430_ | ~new_n24329_;
  assign new_n24439_ = ~new_n24431_ | ~new_n24361_;
  assign new_n24440_ = ~pi0322 | ~new_n26365_;
  assign new_n24441_ = ~pi0324 | ~new_n26366_;
  assign new_n24442_ = ~pi0325 | ~new_n26363_;
  assign new_n24443_ = ~pi0346 | ~new_n26363_;
  assign new_n24444_ = ~pi0318 | ~new_n24335_;
  assign new_n24445_ = ~pi0318 | ~new_n27120_;
  assign new_n24446_ = ~new_n26363_ | ~new_n24241_;
  assign new_n24447_ = ~pi0334 | ~new_n26363_;
  assign new_n24448_ = ~new_n26363_ | ~new_n24236_;
  assign new_n24449_ = ~pi0345 | ~new_n26363_;
  assign new_n24450_ = ~new_n24378_ | ~new_n24315_;
  assign new_n24451_ = ~new_n24238_;
  assign new_n24452_ = ~new_n24183_ | ~new_n24315_;
  assign new_n24453_ = ~new_n24311_;
  assign new_n24454_ = ~new_n24185_ | ~new_n24315_;
  assign new_n24455_ = ~new_n24309_;
  assign new_n24456_ = ~new_n24187_ | ~new_n24315_;
  assign new_n24457_ = ~new_n24307_;
  assign new_n24458_ = ~new_n24277_ | ~new_n24315_;
  assign new_n24459_ = ~new_n24237_;
  assign new_n24460_ = ~new_n24352_ | ~new_n24289_;
  assign new_n24461_ = ~new_n24324_;
  assign new_n24462_ = ~new_n24180_ | ~new_n24289_;
  assign new_n24463_ = ~new_n24323_;
  assign new_n24464_ = ~new_n24181_ | ~new_n24289_;
  assign new_n24465_ = ~new_n24242_;
  assign new_n24466_ = ~new_n24272_ | ~new_n24289_;
  assign new_n24467_ = ~new_n24321_;
  assign new_n24468_ = ~new_n24397_ | ~new_n24234_;
  assign new_n24469_ = ~pi0347 | ~new_n24235_;
  assign new_n24470_ = ~new_n24469_ | ~new_n24526_ | ~new_n24525_;
  assign new_n24471_ = ~new_n24282_ | ~new_n24235_;
  assign new_n24472_ = ~new_n24344_ | ~new_n24297_;
  assign new_n24473_ = ~new_n24295_;
  assign new_n24474_ = ~new_n24349_ | ~new_n24293_;
  assign new_n24475_ = ~new_n24291_;
  assign new_n24476_ = ~pi0344 | ~new_n24305_;
  assign new_n24477_ = ~new_n24476_ | ~new_n24549_ | ~new_n24548_;
  assign new_n24478_ = ~new_n24178_ | ~new_n24305_;
  assign new_n24479_ = ~new_n24303_;
  assign new_n24480_ = ~new_n24178_ | ~new_n24305_;
  assign new_n24481_ = ~new_n24332_ | ~pi0318;
  assign new_n24482_ = ~new_n26363_ | ~new_n24215_;
  assign new_n24483_ = ~pi0326 | ~new_n24213_;
  assign new_n24484_ = ~new_n24483_ | ~new_n24482_;
  assign new_n24485_ = ~new_n24432_ | ~new_n24289_;
  assign new_n24486_ = ~new_n24351_ | ~new_n24484_;
  assign new_n24487_ = ~new_n26363_ | ~new_n24214_;
  assign new_n24488_ = ~pi0325 | ~new_n24213_;
  assign new_n24489_ = ~new_n26363_ | ~new_n24214_;
  assign new_n24490_ = ~pi0325 | ~new_n24213_;
  assign new_n24491_ = ~new_n24490_ | ~new_n24489_;
  assign new_n24492_ = ~new_n24290_ | ~new_n24291_;
  assign new_n24493_ = ~new_n24475_ | ~new_n24491_;
  assign new_n24494_ = ~pi0324 | ~new_n24196_;
  assign new_n24495_ = ~new_n26366_ | ~new_n24197_;
  assign new_n24496_ = ~pi0324 | ~new_n24196_;
  assign new_n24497_ = ~new_n26366_ | ~new_n24197_;
  assign new_n24498_ = ~new_n24497_ | ~new_n24496_;
  assign new_n24499_ = ~new_n24292_ | ~new_n24293_;
  assign new_n24500_ = ~new_n24348_ | ~new_n24498_;
  assign new_n24501_ = ~pi0323 | ~new_n24211_;
  assign new_n24502_ = ~new_n26374_ | ~new_n24212_;
  assign new_n24503_ = ~pi0323 | ~new_n24211_;
  assign new_n24504_ = ~new_n26374_ | ~new_n24212_;
  assign new_n24505_ = ~new_n24504_ | ~new_n24503_;
  assign new_n24506_ = ~new_n24294_ | ~new_n24295_;
  assign new_n24507_ = ~new_n24473_ | ~new_n24505_;
  assign new_n24508_ = ~pi0322 | ~new_n24198_;
  assign new_n24509_ = ~new_n26365_ | ~new_n24199_;
  assign new_n24510_ = ~pi0322 | ~new_n24198_;
  assign new_n24511_ = ~new_n26365_ | ~new_n24199_;
  assign new_n24512_ = ~new_n24511_ | ~new_n24510_;
  assign new_n24513_ = ~new_n24296_ | ~new_n24297_;
  assign new_n24514_ = ~new_n24343_ | ~new_n24512_;
  assign new_n24515_ = ~pi0321 | ~new_n24200_;
  assign new_n24516_ = ~new_n26376_ | ~new_n24201_;
  assign new_n24517_ = ~new_n24516_ | ~new_n24515_;
  assign new_n24518_ = ~new_n24433_ | ~new_n24298_;
  assign new_n24519_ = ~new_n24356_ | ~new_n24517_;
  assign new_n24520_ = ~pi0320 | ~new_n24209_;
  assign new_n24521_ = ~new_n26364_ | ~new_n24210_;
  assign new_n24522_ = ~new_n24521_ | ~new_n24520_;
  assign new_n24523_ = ~new_n24434_ | ~new_n24299_;
  assign new_n24524_ = ~new_n24358_ | ~new_n24522_;
  assign new_n24525_ = ~pi0348 | ~new_n24213_;
  assign new_n24526_ = ~new_n26363_ | ~new_n24398_;
  assign new_n24527_ = ~pi0348 | ~new_n26363_;
  assign new_n24528_ = ~new_n24471_ | ~new_n24213_;
  assign new_n24529_ = ~new_n26363_ | ~new_n24234_;
  assign new_n24530_ = ~pi0347 | ~new_n24213_;
  assign new_n24531_ = ~new_n26363_ | ~new_n24234_;
  assign new_n24532_ = ~pi0347 | ~new_n24213_;
  assign new_n24533_ = ~new_n24532_ | ~new_n24531_;
  assign new_n24534_ = ~new_n24300_ | ~new_n24235_;
  assign new_n24535_ = ~new_n24533_ | ~new_n24397_;
  assign new_n24536_ = ~pi0319 | ~new_n24206_;
  assign new_n24537_ = ~new_n26370_ | ~new_n24207_;
  assign new_n24538_ = ~new_n24537_ | ~new_n24536_;
  assign new_n24539_ = ~new_n24435_ | ~new_n24301_;
  assign new_n24540_ = ~new_n24339_ | ~new_n24538_;
  assign new_n24541_ = ~new_n26363_ | ~new_n24233_;
  assign new_n24542_ = ~pi0346 | ~new_n24213_;
  assign new_n24543_ = ~new_n26363_ | ~new_n24233_;
  assign new_n24544_ = ~pi0346 | ~new_n24213_;
  assign new_n24545_ = ~new_n24544_ | ~new_n24543_;
  assign new_n24546_ = ~new_n24302_ | ~new_n24303_;
  assign new_n24547_ = ~new_n24479_ | ~new_n24545_;
  assign new_n24548_ = ~pi0345 | ~new_n24213_;
  assign new_n24549_ = ~new_n26363_ | ~new_n24400_;
  assign new_n24550_ = ~pi0345 | ~new_n26363_;
  assign new_n24551_ = ~new_n24480_ | ~new_n24213_;
  assign new_n24552_ = ~pi0344 | ~new_n24213_;
  assign new_n24553_ = ~new_n26363_ | ~new_n24232_;
  assign new_n24554_ = ~pi0344 | ~new_n24213_;
  assign new_n24555_ = ~new_n26363_ | ~new_n24232_;
  assign new_n24556_ = ~new_n24555_ | ~new_n24554_;
  assign new_n24557_ = ~new_n24304_ | ~new_n24305_;
  assign new_n24558_ = ~new_n24394_ | ~new_n24556_;
  assign new_n24559_ = ~pi0343 | ~new_n24213_;
  assign new_n24560_ = ~new_n26363_ | ~new_n24217_;
  assign new_n24561_ = ~pi0342 | ~new_n24213_;
  assign new_n24562_ = ~new_n26363_ | ~new_n24216_;
  assign new_n24563_ = ~new_n24562_ | ~new_n24561_;
  assign new_n24564_ = ~new_n24237_ | ~new_n24436_;
  assign new_n24565_ = ~new_n24563_ | ~new_n24459_;
  assign new_n24566_ = ~pi0341 | ~new_n24213_;
  assign new_n24567_ = ~new_n26363_ | ~new_n24218_;
  assign new_n24568_ = ~pi0341 | ~new_n24213_;
  assign new_n24569_ = ~new_n26363_ | ~new_n24218_;
  assign new_n24570_ = ~new_n24569_ | ~new_n24568_;
  assign new_n24571_ = ~new_n24306_ | ~new_n24307_;
  assign new_n24572_ = ~new_n24457_ | ~new_n24570_;
  assign new_n24573_ = ~pi0340 | ~new_n24213_;
  assign new_n24574_ = ~new_n26363_ | ~new_n24219_;
  assign new_n24575_ = ~pi0340 | ~new_n24213_;
  assign new_n24576_ = ~new_n26363_ | ~new_n24219_;
  assign new_n24577_ = ~new_n24576_ | ~new_n24575_;
  assign new_n24578_ = ~new_n24308_ | ~new_n24309_;
  assign new_n24579_ = ~new_n24455_ | ~new_n24577_;
  assign new_n24580_ = ~pi0339 | ~new_n24213_;
  assign new_n24581_ = ~new_n26363_ | ~new_n24220_;
  assign new_n24582_ = ~pi0339 | ~new_n24213_;
  assign new_n24583_ = ~new_n26363_ | ~new_n24220_;
  assign new_n24584_ = ~new_n24583_ | ~new_n24582_;
  assign new_n24585_ = ~new_n24310_ | ~new_n24311_;
  assign new_n24586_ = ~new_n24453_ | ~new_n24584_;
  assign new_n24587_ = ~pi0338 | ~new_n24213_;
  assign new_n24588_ = ~new_n26363_ | ~new_n24222_;
  assign new_n24589_ = ~pi0338 | ~new_n24213_;
  assign new_n24590_ = ~new_n26363_ | ~new_n24222_;
  assign new_n24591_ = ~new_n24590_ | ~new_n24589_;
  assign new_n24592_ = ~new_n24312_ | ~new_n24313_;
  assign new_n24593_ = ~new_n24412_ | ~new_n24591_;
  assign new_n24594_ = ~pi0337 | ~new_n24213_;
  assign new_n24595_ = ~new_n26363_ | ~new_n24413_;
  assign new_n24596_ = ~pi0318 | ~new_n24204_;
  assign new_n24597_ = ~new_n24335_ | ~new_n24208_;
  assign new_n24598_ = ~new_n24597_ | ~new_n24596_;
  assign new_n24599_ = ~new_n27120_ | ~new_n24204_ | ~new_n24208_;
  assign new_n24600_ = ~new_n24598_ | ~new_n24205_;
  assign new_n24601_ = ~pi0336 | ~new_n24213_;
  assign new_n24602_ = ~new_n26363_ | ~new_n24221_;
  assign new_n24603_ = ~new_n24602_ | ~new_n24601_;
  assign new_n24604_ = ~new_n24238_ | ~new_n24437_;
  assign new_n24605_ = ~new_n24603_ | ~new_n24451_;
  assign new_n24606_ = ~pi0335 | ~new_n24213_;
  assign new_n24607_ = ~new_n26363_ | ~new_n24223_;
  assign new_n24608_ = ~pi0335 | ~new_n24213_;
  assign new_n24609_ = ~new_n26363_ | ~new_n24223_;
  assign new_n24610_ = ~new_n24609_ | ~new_n24608_;
  assign new_n24611_ = ~new_n24314_ | ~new_n24315_;
  assign new_n24612_ = ~new_n24377_ | ~new_n24610_;
  assign new_n24613_ = ~pi0334 | ~new_n24213_;
  assign new_n24614_ = ~new_n26363_ | ~new_n24420_;
  assign new_n24615_ = ~pi0334 | ~new_n26363_;
  assign new_n24616_ = ~new_n24375_ | ~new_n24213_;
  assign new_n24617_ = ~pi0333 | ~new_n24213_;
  assign new_n24618_ = ~new_n26363_ | ~new_n24230_;
  assign new_n24619_ = ~pi0333 | ~new_n24213_;
  assign new_n24620_ = ~new_n26363_ | ~new_n24230_;
  assign new_n24621_ = ~new_n24620_ | ~new_n24619_;
  assign new_n24622_ = ~new_n24316_ | ~new_n24317_;
  assign new_n24623_ = ~new_n24374_ | ~new_n24621_;
  assign new_n24624_ = ~pi0332 | ~new_n24213_;
  assign new_n24625_ = ~new_n26363_ | ~new_n24229_;
  assign new_n24626_ = ~pi0332 | ~new_n24213_;
  assign new_n24627_ = ~new_n26363_ | ~new_n24229_;
  assign new_n24628_ = ~new_n24627_ | ~new_n24626_;
  assign new_n24629_ = ~new_n24318_ | ~new_n24319_;
  assign new_n24630_ = ~new_n24370_ | ~new_n24628_;
  assign new_n24631_ = ~pi0331 | ~new_n24213_;
  assign new_n24632_ = ~new_n26363_ | ~new_n24228_;
  assign new_n24633_ = ~pi0331 | ~new_n24213_;
  assign new_n24634_ = ~new_n26363_ | ~new_n24228_;
  assign new_n24635_ = ~new_n24634_ | ~new_n24633_;
  assign new_n24636_ = ~new_n24320_ | ~new_n24321_;
  assign new_n24637_ = ~new_n24467_ | ~new_n24635_;
  assign new_n24638_ = ~pi0330 | ~new_n24213_;
  assign new_n24639_ = ~new_n26363_ | ~new_n24225_;
  assign new_n24640_ = ~pi0329 | ~new_n24213_;
  assign new_n24641_ = ~new_n26363_ | ~new_n24224_;
  assign new_n24642_ = ~new_n24641_ | ~new_n24640_;
  assign new_n24643_ = ~new_n24242_ | ~new_n24438_;
  assign new_n24644_ = ~new_n24642_ | ~new_n24465_;
  assign new_n24645_ = ~pi0328 | ~new_n24213_;
  assign new_n24646_ = ~new_n26363_ | ~new_n24226_;
  assign new_n24647_ = ~pi0328 | ~new_n24213_;
  assign new_n24648_ = ~new_n26363_ | ~new_n24226_;
  assign new_n24649_ = ~new_n24648_ | ~new_n24647_;
  assign new_n24650_ = ~new_n24322_ | ~new_n24323_;
  assign new_n24651_ = ~new_n24463_ | ~new_n24649_;
  assign new_n24652_ = ~pi0327 | ~new_n24213_;
  assign new_n24653_ = ~new_n26363_ | ~new_n24227_;
  assign new_n24654_ = ~new_n24653_ | ~new_n24652_;
  assign new_n24655_ = ~new_n24324_ | ~new_n24439_;
  assign new_n24656_ = ~new_n24461_ | ~new_n24654_;
  assign new_n24657_ = ~pi0317 | ~new_n24202_;
  assign new_n24658_ = ~new_n26367_ | ~new_n24203_;
  assign new_n24659_ = ~pi0311;
  assign new_n24660_ = pi0307 & new_n24674_;
  assign new_n24661_ = ~pi0310;
  assign new_n24662_ = ~pi0310 | ~pi0311;
  assign new_n24663_ = ~pi0309;
  assign new_n24664_ = ~pi0309 | ~new_n24672_;
  assign new_n24665_ = ~pi0308;
  assign new_n24666_ = ~pi0308 | ~new_n24673_;
  assign new_n24667_ = ~pi0307;
  assign new_n24668_ = ~new_n24676_ | ~new_n24675_;
  assign new_n24669_ = ~new_n24678_ | ~new_n24677_;
  assign new_n24670_ = ~new_n24680_ | ~new_n24679_;
  assign new_n24671_ = ~new_n24682_ | ~new_n24681_;
  assign new_n24672_ = ~new_n24662_;
  assign new_n24673_ = ~new_n24664_;
  assign new_n24674_ = ~new_n24666_;
  assign new_n24675_ = ~pi0307 | ~new_n24666_;
  assign new_n24676_ = ~new_n24674_ | ~new_n24667_;
  assign new_n24677_ = ~pi0308 | ~new_n24664_;
  assign new_n24678_ = ~new_n24673_ | ~new_n24665_;
  assign new_n24679_ = ~pi0309 | ~new_n24662_;
  assign new_n24680_ = ~new_n24672_ | ~new_n24663_;
  assign new_n24681_ = ~pi0310 | ~new_n24659_;
  assign new_n24682_ = ~pi0311 | ~new_n24661_;
  assign new_n24683_ = ~new_n24720_ | ~new_n24719_;
  assign new_n24684_ = ~pi0311 | ~new_n24704_;
  assign new_n24685_ = ~pi0315;
  assign new_n24686_ = ~pi0309;
  assign new_n24687_ = ~pi0314;
  assign new_n24688_ = ~pi0308;
  assign new_n24689_ = ~pi0313;
  assign new_n24690_ = ~pi0312;
  assign new_n24691_ = ~new_n24716_ | ~new_n24715_;
  assign new_n24692_ = ~pi0307;
  assign new_n24693_ = ~new_n24725_ | ~new_n24724_;
  assign new_n24694_ = ~new_n24730_ | ~new_n24729_;
  assign new_n24695_ = ~new_n24735_ | ~new_n24734_;
  assign new_n24696_ = ~new_n24740_ | ~new_n24739_;
  assign new_n24697_ = ~new_n24722_ | ~new_n24721_;
  assign new_n24698_ = ~new_n24727_ | ~new_n24726_;
  assign new_n24699_ = ~new_n24732_ | ~new_n24731_;
  assign new_n24700_ = ~new_n24737_ | ~new_n24736_;
  assign new_n24701_ = ~new_n24712_ | ~new_n24711_;
  assign new_n24702_ = ~new_n24708_ | ~new_n24707_;
  assign new_n24703_ = ~pi0310;
  assign new_n24704_ = ~pi0316;
  assign new_n24705_ = ~new_n24684_;
  assign new_n24706_ = ~new_n24705_ | ~new_n24685_;
  assign new_n24707_ = ~new_n24706_ | ~new_n24703_;
  assign new_n24708_ = ~pi0315 | ~new_n24684_;
  assign new_n24709_ = ~new_n24702_;
  assign new_n24710_ = ~pi0309 | ~new_n24687_;
  assign new_n24711_ = ~new_n24710_ | ~new_n24702_;
  assign new_n24712_ = ~pi0314 | ~new_n24686_;
  assign new_n24713_ = ~new_n24701_;
  assign new_n24714_ = ~pi0308 | ~new_n24689_;
  assign new_n24715_ = ~new_n24714_ | ~new_n24701_;
  assign new_n24716_ = ~pi0313 | ~new_n24688_;
  assign new_n24717_ = ~new_n24691_;
  assign new_n24718_ = ~pi0312 | ~new_n24692_;
  assign new_n24719_ = ~new_n24717_ | ~new_n24718_;
  assign new_n24720_ = ~pi0307 | ~new_n24690_;
  assign new_n24721_ = ~pi0307 | ~new_n24690_;
  assign new_n24722_ = ~pi0312 | ~new_n24692_;
  assign new_n24723_ = ~new_n24697_;
  assign new_n24724_ = ~new_n24723_ | ~new_n24717_;
  assign new_n24725_ = ~new_n24697_ | ~new_n24691_;
  assign new_n24726_ = ~pi0308 | ~new_n24689_;
  assign new_n24727_ = ~pi0313 | ~new_n24688_;
  assign new_n24728_ = ~new_n24698_;
  assign new_n24729_ = ~new_n24713_ | ~new_n24728_;
  assign new_n24730_ = ~new_n24698_ | ~new_n24701_;
  assign new_n24731_ = ~pi0309 | ~new_n24687_;
  assign new_n24732_ = ~pi0314 | ~new_n24686_;
  assign new_n24733_ = ~new_n24699_;
  assign new_n24734_ = ~new_n24709_ | ~new_n24733_;
  assign new_n24735_ = ~new_n24699_ | ~new_n24702_;
  assign new_n24736_ = ~pi0310 | ~new_n24685_;
  assign new_n24737_ = ~pi0315 | ~new_n24703_;
  assign new_n24738_ = ~new_n24700_;
  assign new_n24739_ = ~new_n24738_ | ~new_n24705_;
  assign new_n24740_ = ~new_n24700_ | ~new_n24684_;
  assign new_n24741_ = ~new_n4461_;
  assign new_n24742_ = ~new_n4462_;
  assign new_n24743_ = ~pi0318;
  assign new_n24744_ = ~pi0319;
  assign new_n24745_ = ~pi0319 | ~pi0318;
  assign new_n24746_ = ~pi0320;
  assign new_n24747_ = ~pi0320 | ~new_n24833_;
  assign new_n24748_ = ~pi0321;
  assign new_n24749_ = ~pi0321 | ~new_n24834_;
  assign new_n24750_ = ~pi0322;
  assign new_n24751_ = ~pi0322 | ~new_n24835_;
  assign new_n24752_ = ~pi0323;
  assign new_n24753_ = ~pi0323 | ~new_n24836_;
  assign new_n24754_ = ~pi0324;
  assign new_n24755_ = ~pi0324 | ~new_n24837_;
  assign new_n24756_ = ~pi0325;
  assign new_n24757_ = ~pi0326;
  assign new_n24758_ = ~pi0325 | ~new_n24838_;
  assign new_n24759_ = ~new_n24839_ | ~pi0326;
  assign new_n24760_ = ~pi0327;
  assign new_n24761_ = ~pi0327 | ~new_n24840_;
  assign new_n24762_ = ~pi0328;
  assign new_n24763_ = ~pi0328 | ~new_n24841_;
  assign new_n24764_ = ~pi0329;
  assign new_n24765_ = ~pi0329 | ~new_n24842_;
  assign new_n24766_ = ~pi0330;
  assign new_n24767_ = ~pi0330 | ~new_n24843_;
  assign new_n24768_ = ~pi0331;
  assign new_n24769_ = ~pi0331 | ~new_n24844_;
  assign new_n24770_ = ~pi0332;
  assign new_n24771_ = ~pi0332 | ~new_n24845_;
  assign new_n24772_ = ~pi0333;
  assign new_n24773_ = ~pi0333 | ~new_n24846_;
  assign new_n24774_ = ~pi0334;
  assign new_n24775_ = ~pi0334 | ~new_n24847_;
  assign new_n24776_ = ~pi0335;
  assign new_n24777_ = ~pi0335 | ~new_n24848_;
  assign new_n24778_ = ~pi0336;
  assign new_n24779_ = ~pi0336 | ~new_n24849_;
  assign new_n24780_ = ~pi0337;
  assign new_n24781_ = ~pi0337 | ~new_n24850_;
  assign new_n24782_ = ~pi0338;
  assign new_n24783_ = ~pi0338 | ~new_n24851_;
  assign new_n24784_ = ~pi0339;
  assign new_n24785_ = ~pi0339 | ~new_n24852_;
  assign new_n24786_ = ~pi0340;
  assign new_n24787_ = ~pi0340 | ~new_n24853_;
  assign new_n24788_ = ~pi0341;
  assign new_n24789_ = ~pi0341 | ~new_n24854_;
  assign new_n24790_ = ~pi0342;
  assign new_n24791_ = ~pi0342 | ~new_n24855_;
  assign new_n24792_ = ~pi0343;
  assign new_n24793_ = ~pi0343 | ~new_n24856_;
  assign new_n24794_ = ~pi0344;
  assign new_n24795_ = ~pi0344 | ~new_n24857_;
  assign new_n24796_ = ~pi0345;
  assign new_n24797_ = ~pi0345 | ~new_n24858_;
  assign new_n24798_ = ~pi0346;
  assign new_n24799_ = ~pi0346 | ~new_n24859_;
  assign new_n24800_ = ~pi0347;
  assign new_n24801_ = ~new_n24863_ | ~new_n24862_;
  assign new_n24802_ = ~new_n24865_ | ~new_n24864_;
  assign new_n24803_ = ~new_n24867_ | ~new_n24866_;
  assign new_n24804_ = ~new_n24869_ | ~new_n24868_;
  assign new_n24805_ = ~new_n24871_ | ~new_n24870_;
  assign new_n24806_ = ~new_n24873_ | ~new_n24872_;
  assign new_n24807_ = ~new_n24875_ | ~new_n24874_;
  assign new_n24808_ = ~new_n24877_ | ~new_n24876_;
  assign new_n24809_ = ~new_n24879_ | ~new_n24878_;
  assign new_n24810_ = ~new_n24881_ | ~new_n24880_;
  assign new_n24811_ = ~new_n24883_ | ~new_n24882_;
  assign new_n24812_ = ~new_n24885_ | ~new_n24884_;
  assign new_n24813_ = ~new_n24887_ | ~new_n24886_;
  assign new_n24814_ = ~new_n24889_ | ~new_n24888_;
  assign new_n24815_ = ~new_n24891_ | ~new_n24890_;
  assign new_n24816_ = ~new_n24893_ | ~new_n24892_;
  assign new_n24817_ = ~new_n24895_ | ~new_n24894_;
  assign new_n24818_ = ~new_n24897_ | ~new_n24896_;
  assign new_n24819_ = ~new_n24899_ | ~new_n24898_;
  assign new_n24820_ = ~new_n24901_ | ~new_n24900_;
  assign new_n24821_ = ~new_n24903_ | ~new_n24902_;
  assign new_n24822_ = ~new_n24905_ | ~new_n24904_;
  assign new_n24823_ = ~new_n24907_ | ~new_n24906_;
  assign new_n24824_ = ~new_n24909_ | ~new_n24908_;
  assign new_n24825_ = ~new_n24911_ | ~new_n24910_;
  assign new_n24826_ = ~new_n24913_ | ~new_n24912_;
  assign new_n24827_ = ~new_n24915_ | ~new_n24914_;
  assign new_n24828_ = ~new_n24917_ | ~new_n24916_;
  assign new_n24829_ = ~new_n24919_ | ~new_n24918_;
  assign new_n24830_ = ~new_n24921_ | ~new_n24920_;
  assign new_n24831_ = ~pi0348;
  assign new_n24832_ = ~pi0347 | ~new_n24860_;
  assign new_n24833_ = ~new_n24745_;
  assign new_n24834_ = ~new_n24747_;
  assign new_n24835_ = ~new_n24749_;
  assign new_n24836_ = ~new_n24751_;
  assign new_n24837_ = ~new_n24753_;
  assign new_n24838_ = ~new_n24755_;
  assign new_n24839_ = ~new_n24758_;
  assign new_n24840_ = ~new_n24759_;
  assign new_n24841_ = ~new_n24761_;
  assign new_n24842_ = ~new_n24763_;
  assign new_n24843_ = ~new_n24765_;
  assign new_n24844_ = ~new_n24767_;
  assign new_n24845_ = ~new_n24769_;
  assign new_n24846_ = ~new_n24771_;
  assign new_n24847_ = ~new_n24773_;
  assign new_n24848_ = ~new_n24775_;
  assign new_n24849_ = ~new_n24777_;
  assign new_n24850_ = ~new_n24779_;
  assign new_n24851_ = ~new_n24781_;
  assign new_n24852_ = ~new_n24783_;
  assign new_n24853_ = ~new_n24785_;
  assign new_n24854_ = ~new_n24787_;
  assign new_n24855_ = ~new_n24789_;
  assign new_n24856_ = ~new_n24791_;
  assign new_n24857_ = ~new_n24793_;
  assign new_n24858_ = ~new_n24795_;
  assign new_n24859_ = ~new_n24797_;
  assign new_n24860_ = ~new_n24799_;
  assign new_n24861_ = ~new_n24832_;
  assign new_n24862_ = ~pi0326 | ~new_n24758_;
  assign new_n24863_ = ~new_n24839_ | ~new_n24757_;
  assign new_n24864_ = ~pi0325 | ~new_n24755_;
  assign new_n24865_ = ~new_n24838_ | ~new_n24756_;
  assign new_n24866_ = ~pi0324 | ~new_n24753_;
  assign new_n24867_ = ~new_n24837_ | ~new_n24754_;
  assign new_n24868_ = ~pi0323 | ~new_n24751_;
  assign new_n24869_ = ~new_n24836_ | ~new_n24752_;
  assign new_n24870_ = ~pi0322 | ~new_n24749_;
  assign new_n24871_ = ~new_n24835_ | ~new_n24750_;
  assign new_n24872_ = ~pi0321 | ~new_n24747_;
  assign new_n24873_ = ~new_n24834_ | ~new_n24748_;
  assign new_n24874_ = ~pi0320 | ~new_n24745_;
  assign new_n24875_ = ~new_n24833_ | ~new_n24746_;
  assign new_n24876_ = ~pi0348 | ~new_n24832_;
  assign new_n24877_ = ~new_n24861_ | ~new_n24831_;
  assign new_n24878_ = ~pi0347 | ~new_n24799_;
  assign new_n24879_ = ~new_n24860_ | ~new_n24800_;
  assign new_n24880_ = ~pi0319 | ~new_n24743_;
  assign new_n24881_ = ~pi0318 | ~new_n24744_;
  assign new_n24882_ = ~pi0346 | ~new_n24797_;
  assign new_n24883_ = ~new_n24859_ | ~new_n24798_;
  assign new_n24884_ = ~pi0345 | ~new_n24795_;
  assign new_n24885_ = ~new_n24858_ | ~new_n24796_;
  assign new_n24886_ = ~pi0344 | ~new_n24793_;
  assign new_n24887_ = ~new_n24857_ | ~new_n24794_;
  assign new_n24888_ = ~pi0343 | ~new_n24791_;
  assign new_n24889_ = ~new_n24856_ | ~new_n24792_;
  assign new_n24890_ = ~pi0342 | ~new_n24789_;
  assign new_n24891_ = ~new_n24855_ | ~new_n24790_;
  assign new_n24892_ = ~pi0341 | ~new_n24787_;
  assign new_n24893_ = ~new_n24854_ | ~new_n24788_;
  assign new_n24894_ = ~pi0340 | ~new_n24785_;
  assign new_n24895_ = ~new_n24853_ | ~new_n24786_;
  assign new_n24896_ = ~pi0339 | ~new_n24783_;
  assign new_n24897_ = ~new_n24852_ | ~new_n24784_;
  assign new_n24898_ = ~pi0338 | ~new_n24781_;
  assign new_n24899_ = ~new_n24851_ | ~new_n24782_;
  assign new_n24900_ = ~pi0337 | ~new_n24779_;
  assign new_n24901_ = ~new_n24850_ | ~new_n24780_;
  assign new_n24902_ = ~pi0336 | ~new_n24777_;
  assign new_n24903_ = ~new_n24849_ | ~new_n24778_;
  assign new_n24904_ = ~pi0335 | ~new_n24775_;
  assign new_n24905_ = ~new_n24848_ | ~new_n24776_;
  assign new_n24906_ = ~pi0334 | ~new_n24773_;
  assign new_n24907_ = ~new_n24847_ | ~new_n24774_;
  assign new_n24908_ = ~pi0333 | ~new_n24771_;
  assign new_n24909_ = ~new_n24846_ | ~new_n24772_;
  assign new_n24910_ = ~pi0332 | ~new_n24769_;
  assign new_n24911_ = ~new_n24845_ | ~new_n24770_;
  assign new_n24912_ = ~pi0331 | ~new_n24767_;
  assign new_n24913_ = ~new_n24844_ | ~new_n24768_;
  assign new_n24914_ = ~pi0330 | ~new_n24765_;
  assign new_n24915_ = ~new_n24843_ | ~new_n24766_;
  assign new_n24916_ = ~pi0329 | ~new_n24763_;
  assign new_n24917_ = ~new_n24842_ | ~new_n24764_;
  assign new_n24918_ = ~pi0328 | ~new_n24761_;
  assign new_n24919_ = ~new_n24841_ | ~new_n24762_;
  assign new_n24920_ = ~pi0327 | ~new_n24759_;
  assign new_n24921_ = ~new_n24840_ | ~new_n24760_;
  assign new_n24922_ = ~pi0317;
  assign new_n24923_ = ~new_n25010_ | ~new_n25044_;
  assign new_n24924_ = ~pi0318;
  assign new_n24925_ = ~pi0320;
  assign new_n24926_ = ~pi0320 | ~new_n25010_;
  assign new_n24927_ = ~pi0321;
  assign new_n24928_ = ~pi0321 | ~new_n25016_;
  assign new_n24929_ = ~pi0322;
  assign new_n24930_ = ~pi0322 | ~new_n25017_;
  assign new_n24931_ = ~pi0323;
  assign new_n24932_ = ~pi0323 | ~new_n25018_;
  assign new_n24933_ = ~pi0324;
  assign new_n24934_ = ~pi0324 | ~new_n25019_;
  assign new_n24935_ = ~pi0325;
  assign new_n24936_ = ~pi0326;
  assign new_n24937_ = ~pi0325 | ~new_n25020_;
  assign new_n24938_ = ~new_n25021_ | ~pi0326;
  assign new_n24939_ = ~pi0327;
  assign new_n24940_ = ~pi0327 | ~new_n25022_;
  assign new_n24941_ = ~pi0328;
  assign new_n24942_ = ~pi0328 | ~new_n25023_;
  assign new_n24943_ = ~pi0329;
  assign new_n24944_ = ~pi0329 | ~new_n25024_;
  assign new_n24945_ = ~pi0330;
  assign new_n24946_ = ~pi0330 | ~new_n25025_;
  assign new_n24947_ = ~pi0331;
  assign new_n24948_ = ~pi0331 | ~new_n25026_;
  assign new_n24949_ = ~pi0332;
  assign new_n24950_ = ~pi0332 | ~new_n25027_;
  assign new_n24951_ = ~pi0333;
  assign new_n24952_ = ~pi0333 | ~new_n25028_;
  assign new_n24953_ = ~pi0334;
  assign new_n24954_ = ~pi0334 | ~new_n25029_;
  assign new_n24955_ = ~pi0335;
  assign new_n24956_ = ~pi0335 | ~new_n25030_;
  assign new_n24957_ = ~pi0336;
  assign new_n24958_ = ~pi0336 | ~new_n25031_;
  assign new_n24959_ = ~pi0337;
  assign new_n24960_ = ~pi0337 | ~new_n25032_;
  assign new_n24961_ = ~pi0338;
  assign new_n24962_ = ~pi0338 | ~new_n25033_;
  assign new_n24963_ = ~pi0339;
  assign new_n24964_ = ~pi0339 | ~new_n25034_;
  assign new_n24965_ = ~pi0340;
  assign new_n24966_ = ~pi0340 | ~new_n25035_;
  assign new_n24967_ = ~pi0341;
  assign new_n24968_ = ~pi0341 | ~new_n25036_;
  assign new_n24969_ = ~pi0342;
  assign new_n24970_ = ~pi0342 | ~new_n25037_;
  assign new_n24971_ = ~pi0343;
  assign new_n24972_ = ~pi0343 | ~new_n25038_;
  assign new_n24973_ = ~pi0344;
  assign new_n24974_ = ~pi0344 | ~new_n25039_;
  assign new_n24975_ = ~pi0345;
  assign new_n24976_ = ~pi0345 | ~new_n25040_;
  assign new_n24977_ = ~pi0346;
  assign new_n24978_ = ~pi0346 | ~new_n25041_;
  assign new_n24979_ = ~pi0347;
  assign new_n24980_ = ~pi0319;
  assign new_n24981_ = ~new_n25046_ | ~new_n25045_;
  assign new_n24982_ = ~new_n25048_ | ~new_n25047_;
  assign new_n24983_ = ~new_n25050_ | ~new_n25049_;
  assign new_n24984_ = ~new_n25052_ | ~new_n25051_;
  assign new_n24985_ = ~new_n25054_ | ~new_n25053_;
  assign new_n24986_ = ~new_n25056_ | ~new_n25055_;
  assign new_n24987_ = ~new_n25060_ | ~new_n25059_;
  assign new_n24988_ = ~new_n25062_ | ~new_n25061_;
  assign new_n24989_ = ~new_n25064_ | ~new_n25063_;
  assign new_n24990_ = ~new_n25066_ | ~new_n25065_;
  assign new_n24991_ = ~new_n25068_ | ~new_n25067_;
  assign new_n24992_ = ~new_n25070_ | ~new_n25069_;
  assign new_n24993_ = ~new_n25072_ | ~new_n25071_;
  assign new_n24994_ = ~new_n25074_ | ~new_n25073_;
  assign new_n24995_ = ~new_n25076_ | ~new_n25075_;
  assign new_n24996_ = ~new_n25078_ | ~new_n25077_;
  assign new_n24997_ = ~new_n25080_ | ~new_n25079_;
  assign new_n24998_ = ~new_n25082_ | ~new_n25081_;
  assign new_n24999_ = ~new_n25084_ | ~new_n25083_;
  assign new_n25000_ = ~new_n25086_ | ~new_n25085_;
  assign new_n25001_ = ~new_n25088_ | ~new_n25087_;
  assign new_n25002_ = ~new_n25090_ | ~new_n25089_;
  assign new_n25003_ = ~new_n25092_ | ~new_n25091_;
  assign new_n25004_ = ~new_n25094_ | ~new_n25093_;
  assign new_n25005_ = ~new_n25096_ | ~new_n25095_;
  assign new_n25006_ = ~new_n25098_ | ~new_n25097_;
  assign new_n25007_ = ~new_n25100_ | ~new_n25099_;
  assign new_n25008_ = ~new_n25102_ | ~new_n25101_;
  assign new_n25009_ = ~new_n25104_ | ~new_n25103_;
  assign new_n25010_ = ~new_n24980_ | ~new_n25014_;
  assign new_n25011_ = new_n25058_ & new_n25057_;
  assign new_n25012_ = ~pi0348;
  assign new_n25013_ = ~pi0347 | ~new_n25042_;
  assign new_n25014_ = ~pi0318 | ~pi0317;
  assign new_n25015_ = ~new_n25010_;
  assign new_n25016_ = ~new_n24926_;
  assign new_n25017_ = ~new_n24928_;
  assign new_n25018_ = ~new_n24930_;
  assign new_n25019_ = ~new_n24932_;
  assign new_n25020_ = ~new_n24934_;
  assign new_n25021_ = ~new_n24937_;
  assign new_n25022_ = ~new_n24938_;
  assign new_n25023_ = ~new_n24940_;
  assign new_n25024_ = ~new_n24942_;
  assign new_n25025_ = ~new_n24944_;
  assign new_n25026_ = ~new_n24946_;
  assign new_n25027_ = ~new_n24948_;
  assign new_n25028_ = ~new_n24950_;
  assign new_n25029_ = ~new_n24952_;
  assign new_n25030_ = ~new_n24954_;
  assign new_n25031_ = ~new_n24956_;
  assign new_n25032_ = ~new_n24958_;
  assign new_n25033_ = ~new_n24960_;
  assign new_n25034_ = ~new_n24962_;
  assign new_n25035_ = ~new_n24964_;
  assign new_n25036_ = ~new_n24966_;
  assign new_n25037_ = ~new_n24968_;
  assign new_n25038_ = ~new_n24970_;
  assign new_n25039_ = ~new_n24972_;
  assign new_n25040_ = ~new_n24974_;
  assign new_n25041_ = ~new_n24976_;
  assign new_n25042_ = ~new_n24978_;
  assign new_n25043_ = ~new_n25013_;
  assign new_n25044_ = ~pi0319 | ~pi0318 | ~pi0317;
  assign new_n25045_ = ~pi0326 | ~new_n24937_;
  assign new_n25046_ = ~new_n25021_ | ~new_n24936_;
  assign new_n25047_ = ~pi0325 | ~new_n24934_;
  assign new_n25048_ = ~new_n25020_ | ~new_n24935_;
  assign new_n25049_ = ~pi0324 | ~new_n24932_;
  assign new_n25050_ = ~new_n25019_ | ~new_n24933_;
  assign new_n25051_ = ~pi0323 | ~new_n24930_;
  assign new_n25052_ = ~new_n25018_ | ~new_n24931_;
  assign new_n25053_ = ~pi0322 | ~new_n24928_;
  assign new_n25054_ = ~new_n25017_ | ~new_n24929_;
  assign new_n25055_ = ~pi0321 | ~new_n24926_;
  assign new_n25056_ = ~new_n25016_ | ~new_n24927_;
  assign new_n25057_ = ~pi0320 | ~new_n25010_;
  assign new_n25058_ = ~new_n25015_ | ~new_n24925_;
  assign new_n25059_ = ~pi0348 | ~new_n25013_;
  assign new_n25060_ = ~new_n25043_ | ~new_n25012_;
  assign new_n25061_ = ~pi0347 | ~new_n24978_;
  assign new_n25062_ = ~new_n25042_ | ~new_n24979_;
  assign new_n25063_ = ~pi0346 | ~new_n24976_;
  assign new_n25064_ = ~new_n25041_ | ~new_n24977_;
  assign new_n25065_ = ~pi0345 | ~new_n24974_;
  assign new_n25066_ = ~new_n25040_ | ~new_n24975_;
  assign new_n25067_ = ~pi0344 | ~new_n24972_;
  assign new_n25068_ = ~new_n25039_ | ~new_n24973_;
  assign new_n25069_ = ~pi0343 | ~new_n24970_;
  assign new_n25070_ = ~new_n25038_ | ~new_n24971_;
  assign new_n25071_ = ~pi0342 | ~new_n24968_;
  assign new_n25072_ = ~new_n25037_ | ~new_n24969_;
  assign new_n25073_ = ~pi0341 | ~new_n24966_;
  assign new_n25074_ = ~new_n25036_ | ~new_n24967_;
  assign new_n25075_ = ~pi0340 | ~new_n24964_;
  assign new_n25076_ = ~new_n25035_ | ~new_n24965_;
  assign new_n25077_ = ~pi0339 | ~new_n24962_;
  assign new_n25078_ = ~new_n25034_ | ~new_n24963_;
  assign new_n25079_ = ~pi0338 | ~new_n24960_;
  assign new_n25080_ = ~new_n25033_ | ~new_n24961_;
  assign new_n25081_ = ~pi0337 | ~new_n24958_;
  assign new_n25082_ = ~new_n25032_ | ~new_n24959_;
  assign new_n25083_ = ~pi0318 | ~new_n24922_;
  assign new_n25084_ = ~pi0317 | ~new_n24924_;
  assign new_n25085_ = ~pi0336 | ~new_n24956_;
  assign new_n25086_ = ~new_n25031_ | ~new_n24957_;
  assign new_n25087_ = ~pi0335 | ~new_n24954_;
  assign new_n25088_ = ~new_n25030_ | ~new_n24955_;
  assign new_n25089_ = ~pi0334 | ~new_n24952_;
  assign new_n25090_ = ~new_n25029_ | ~new_n24953_;
  assign new_n25091_ = ~pi0333 | ~new_n24950_;
  assign new_n25092_ = ~new_n25028_ | ~new_n24951_;
  assign new_n25093_ = ~pi0332 | ~new_n24948_;
  assign new_n25094_ = ~new_n25027_ | ~new_n24949_;
  assign new_n25095_ = ~pi0331 | ~new_n24946_;
  assign new_n25096_ = ~new_n25026_ | ~new_n24947_;
  assign new_n25097_ = ~pi0330 | ~new_n24944_;
  assign new_n25098_ = ~new_n25025_ | ~new_n24945_;
  assign new_n25099_ = ~pi0329 | ~new_n24942_;
  assign new_n25100_ = ~new_n25024_ | ~new_n24943_;
  assign new_n25101_ = ~pi0328 | ~new_n24940_;
  assign new_n25102_ = ~new_n25023_ | ~new_n24941_;
  assign new_n25103_ = ~pi0327 | ~new_n24938_;
  assign new_n25104_ = ~new_n25022_ | ~new_n24939_;
  assign new_n25105_ = ~new_n24120_ & ~new_n25106_;
  assign new_n25106_ = ~new_n24131_ & ~new_n24130_ & ~new_n24132_ & ~new_n24133_;
  assign new_n25107_ = new_n25227_ & new_n25129_;
  assign new_n25108_ = new_n25225_ & new_n25130_;
  assign new_n25109_ = new_n25223_ & new_n25131_;
  assign new_n25110_ = new_n25221_ & new_n25132_;
  assign new_n25111_ = new_n25219_ & new_n25133_;
  assign new_n25112_ = new_n25217_ & new_n25134_;
  assign new_n25113_ = new_n25215_ & new_n25135_;
  assign new_n25114_ = new_n25213_ & new_n25136_;
  assign new_n25115_ = new_n25211_ & new_n25137_;
  assign new_n25116_ = new_n25209_ & new_n25138_;
  assign new_n25117_ = new_n25207_ & new_n25139_;
  assign new_n25118_ = new_n25206_ & new_n25122_;
  assign new_n25119_ = new_n25193_ & new_n25123_;
  assign new_n25120_ = new_n25191_ & new_n25124_;
  assign new_n25121_ = new_n25189_ & new_n25125_;
  assign new_n25122_ = pi0476 | pi0478 | pi0477;
  assign new_n25123_ = ~new_n25184_ | ~new_n25128_ | ~new_n25159_;
  assign new_n25124_ = ~new_n25185_ | ~new_n25127_ | ~new_n25157_;
  assign new_n25125_ = ~new_n25186_ | ~new_n25126_ | ~new_n25155_;
  assign new_n25126_ = ~pi0484;
  assign new_n25127_ = ~pi0482;
  assign new_n25128_ = ~pi0480;
  assign new_n25129_ = ~new_n25187_ | ~new_n25153_ | ~new_n25150_;
  assign new_n25130_ = ~new_n25194_ | ~new_n25149_ | ~new_n25182_;
  assign new_n25131_ = ~new_n25195_ | ~new_n25148_ | ~new_n25180_;
  assign new_n25132_ = ~new_n25196_ | ~new_n25147_ | ~new_n25178_;
  assign new_n25133_ = ~new_n25197_ | ~new_n25146_ | ~new_n25176_;
  assign new_n25134_ = ~new_n25198_ | ~new_n25145_ | ~new_n25174_;
  assign new_n25135_ = ~new_n25199_ | ~new_n25144_ | ~new_n25170_;
  assign new_n25136_ = ~new_n25200_ | ~new_n25143_ | ~new_n25168_;
  assign new_n25137_ = ~new_n25201_ | ~new_n25142_ | ~new_n25166_;
  assign new_n25138_ = ~new_n25202_ | ~new_n25141_ | ~new_n25164_;
  assign new_n25139_ = ~new_n25203_ | ~new_n25140_;
  assign new_n25140_ = ~pi0505;
  assign new_n25141_ = ~pi0504;
  assign new_n25142_ = ~pi0502;
  assign new_n25143_ = ~pi0500;
  assign new_n25144_ = ~pi0498;
  assign new_n25145_ = ~pi0496;
  assign new_n25146_ = ~pi0494;
  assign new_n25147_ = ~pi0492;
  assign new_n25148_ = ~pi0490;
  assign new_n25149_ = ~pi0488;
  assign new_n25150_ = ~pi0486;
  assign new_n25151_ = ~new_n25250_ | ~new_n25249_;
  assign new_n25152_ = ~new_n25238_ | ~new_n25237_;
  assign new_n25153_ = ~pi0485;
  assign new_n25154_ = new_n25230_ & new_n25229_;
  assign new_n25155_ = ~pi0483;
  assign new_n25156_ = new_n25232_ & new_n25231_;
  assign new_n25157_ = ~pi0481;
  assign new_n25158_ = new_n25234_ & new_n25233_;
  assign new_n25159_ = ~pi0479;
  assign new_n25160_ = new_n25236_ & new_n25235_;
  assign new_n25161_ = ~pi0507;
  assign new_n25162_ = ~pi0506;
  assign new_n25163_ = new_n25240_ & new_n25239_;
  assign new_n25164_ = ~pi0503;
  assign new_n25165_ = new_n25242_ & new_n25241_;
  assign new_n25166_ = ~pi0501;
  assign new_n25167_ = new_n25244_ & new_n25243_;
  assign new_n25168_ = ~pi0499;
  assign new_n25169_ = new_n25246_ & new_n25245_;
  assign new_n25170_ = ~pi0497;
  assign new_n25171_ = new_n25248_ & new_n25247_;
  assign new_n25172_ = ~pi0477;
  assign new_n25173_ = ~pi0476;
  assign new_n25174_ = ~pi0495;
  assign new_n25175_ = new_n25252_ & new_n25251_;
  assign new_n25176_ = ~pi0493;
  assign new_n25177_ = new_n25254_ & new_n25253_;
  assign new_n25178_ = ~pi0491;
  assign new_n25179_ = new_n25256_ & new_n25255_;
  assign new_n25180_ = ~pi0489;
  assign new_n25181_ = new_n25258_ & new_n25257_;
  assign new_n25182_ = ~pi0487;
  assign new_n25183_ = new_n25260_ & new_n25259_;
  assign new_n25184_ = ~new_n25122_;
  assign new_n25185_ = ~new_n25123_;
  assign new_n25186_ = ~new_n25124_;
  assign new_n25187_ = ~new_n25125_;
  assign new_n25188_ = ~new_n25186_ | ~new_n25155_;
  assign new_n25189_ = ~pi0484 | ~new_n25188_;
  assign new_n25190_ = ~new_n25185_ | ~new_n25157_;
  assign new_n25191_ = ~pi0482 | ~new_n25190_;
  assign new_n25192_ = ~new_n25184_ | ~new_n25159_;
  assign new_n25193_ = ~pi0480 | ~new_n25192_;
  assign new_n25194_ = ~new_n25129_;
  assign new_n25195_ = ~new_n25130_;
  assign new_n25196_ = ~new_n25131_;
  assign new_n25197_ = ~new_n25132_;
  assign new_n25198_ = ~new_n25133_;
  assign new_n25199_ = ~new_n25134_;
  assign new_n25200_ = ~new_n25135_;
  assign new_n25201_ = ~new_n25136_;
  assign new_n25202_ = ~new_n25137_;
  assign new_n25203_ = ~new_n25138_;
  assign new_n25204_ = ~new_n25139_;
  assign new_n25205_ = pi0477 | pi0476;
  assign new_n25206_ = ~pi0478 | ~new_n25205_;
  assign new_n25207_ = ~pi0505 | ~new_n25138_;
  assign new_n25208_ = ~new_n25202_ | ~new_n25164_;
  assign new_n25209_ = ~pi0504 | ~new_n25208_;
  assign new_n25210_ = ~new_n25201_ | ~new_n25166_;
  assign new_n25211_ = ~pi0502 | ~new_n25210_;
  assign new_n25212_ = ~new_n25200_ | ~new_n25168_;
  assign new_n25213_ = ~pi0500 | ~new_n25212_;
  assign new_n25214_ = ~new_n25199_ | ~new_n25170_;
  assign new_n25215_ = ~pi0498 | ~new_n25214_;
  assign new_n25216_ = ~new_n25198_ | ~new_n25174_;
  assign new_n25217_ = ~pi0496 | ~new_n25216_;
  assign new_n25218_ = ~new_n25197_ | ~new_n25176_;
  assign new_n25219_ = ~pi0494 | ~new_n25218_;
  assign new_n25220_ = ~new_n25196_ | ~new_n25178_;
  assign new_n25221_ = ~pi0492 | ~new_n25220_;
  assign new_n25222_ = ~new_n25195_ | ~new_n25180_;
  assign new_n25223_ = ~pi0490 | ~new_n25222_;
  assign new_n25224_ = ~new_n25194_ | ~new_n25182_;
  assign new_n25225_ = ~pi0488 | ~new_n25224_;
  assign new_n25226_ = ~new_n25187_ | ~new_n25153_;
  assign new_n25227_ = ~pi0486 | ~new_n25226_;
  assign new_n25228_ = ~new_n25204_ | ~new_n25162_;
  assign new_n25229_ = ~pi0485 | ~new_n25125_;
  assign new_n25230_ = ~new_n25187_ | ~new_n25153_;
  assign new_n25231_ = ~pi0483 | ~new_n25124_;
  assign new_n25232_ = ~new_n25186_ | ~new_n25155_;
  assign new_n25233_ = ~pi0481 | ~new_n25123_;
  assign new_n25234_ = ~new_n25185_ | ~new_n25157_;
  assign new_n25235_ = ~pi0479 | ~new_n25122_;
  assign new_n25236_ = ~new_n25184_ | ~new_n25159_;
  assign new_n25237_ = ~new_n25228_ | ~new_n25161_;
  assign new_n25238_ = ~pi0507 | ~new_n25204_ | ~new_n25162_;
  assign new_n25239_ = ~pi0506 | ~new_n25139_;
  assign new_n25240_ = ~new_n25204_ | ~new_n25162_;
  assign new_n25241_ = ~pi0503 | ~new_n25137_;
  assign new_n25242_ = ~new_n25202_ | ~new_n25164_;
  assign new_n25243_ = ~pi0501 | ~new_n25136_;
  assign new_n25244_ = ~new_n25201_ | ~new_n25166_;
  assign new_n25245_ = ~pi0499 | ~new_n25135_;
  assign new_n25246_ = ~new_n25200_ | ~new_n25168_;
  assign new_n25247_ = ~pi0497 | ~new_n25134_;
  assign new_n25248_ = ~new_n25199_ | ~new_n25170_;
  assign new_n25249_ = ~pi0477 | ~new_n25173_;
  assign new_n25250_ = ~pi0476 | ~new_n25172_;
  assign new_n25251_ = ~pi0495 | ~new_n25133_;
  assign new_n25252_ = ~new_n25198_ | ~new_n25174_;
  assign new_n25253_ = ~pi0493 | ~new_n25132_;
  assign new_n25254_ = ~new_n25197_ | ~new_n25176_;
  assign new_n25255_ = ~pi0491 | ~new_n25131_;
  assign new_n25256_ = ~new_n25196_ | ~new_n25178_;
  assign new_n25257_ = ~pi0489 | ~new_n25130_;
  assign new_n25258_ = ~new_n25195_ | ~new_n25180_;
  assign new_n25259_ = ~pi0487 | ~new_n25129_;
  assign new_n25260_ = ~new_n25194_ | ~new_n25182_;
  assign new_n25261_ = ~pi0318;
  assign new_n25262_ = ~pi0319;
  assign new_n25263_ = ~pi0319 | ~pi0318;
  assign new_n25264_ = ~pi0320;
  assign new_n25265_ = ~pi0320 | ~new_n25351_;
  assign new_n25266_ = ~pi0321;
  assign new_n25267_ = ~pi0321 | ~new_n25352_;
  assign new_n25268_ = ~pi0322;
  assign new_n25269_ = ~pi0322 | ~new_n25353_;
  assign new_n25270_ = ~pi0323;
  assign new_n25271_ = ~pi0323 | ~new_n25354_;
  assign new_n25272_ = ~pi0324;
  assign new_n25273_ = ~pi0324 | ~new_n25355_;
  assign new_n25274_ = ~pi0325;
  assign new_n25275_ = ~pi0326;
  assign new_n25276_ = ~pi0325 | ~new_n25356_;
  assign new_n25277_ = ~new_n25357_ | ~pi0326;
  assign new_n25278_ = ~pi0327;
  assign new_n25279_ = ~pi0327 | ~new_n25358_;
  assign new_n25280_ = ~pi0328;
  assign new_n25281_ = ~pi0328 | ~new_n25359_;
  assign new_n25282_ = ~pi0329;
  assign new_n25283_ = ~pi0329 | ~new_n25360_;
  assign new_n25284_ = ~pi0330;
  assign new_n25285_ = ~pi0330 | ~new_n25361_;
  assign new_n25286_ = ~pi0331;
  assign new_n25287_ = ~pi0331 | ~new_n25362_;
  assign new_n25288_ = ~pi0332;
  assign new_n25289_ = ~pi0332 | ~new_n25363_;
  assign new_n25290_ = ~pi0333;
  assign new_n25291_ = ~pi0333 | ~new_n25364_;
  assign new_n25292_ = ~pi0334;
  assign new_n25293_ = ~pi0334 | ~new_n25365_;
  assign new_n25294_ = ~pi0335;
  assign new_n25295_ = ~pi0335 | ~new_n25366_;
  assign new_n25296_ = ~pi0336;
  assign new_n25297_ = ~pi0336 | ~new_n25367_;
  assign new_n25298_ = ~pi0337;
  assign new_n25299_ = ~pi0337 | ~new_n25368_;
  assign new_n25300_ = ~pi0338;
  assign new_n25301_ = ~pi0338 | ~new_n25369_;
  assign new_n25302_ = ~pi0339;
  assign new_n25303_ = ~pi0339 | ~new_n25370_;
  assign new_n25304_ = ~pi0340;
  assign new_n25305_ = ~pi0340 | ~new_n25371_;
  assign new_n25306_ = ~pi0341;
  assign new_n25307_ = ~pi0341 | ~new_n25372_;
  assign new_n25308_ = ~pi0342;
  assign new_n25309_ = ~pi0342 | ~new_n25373_;
  assign new_n25310_ = ~pi0343;
  assign new_n25311_ = ~pi0343 | ~new_n25374_;
  assign new_n25312_ = ~pi0344;
  assign new_n25313_ = ~pi0344 | ~new_n25375_;
  assign new_n25314_ = ~pi0345;
  assign new_n25315_ = ~pi0345 | ~new_n25376_;
  assign new_n25316_ = ~pi0346;
  assign new_n25317_ = ~pi0346 | ~new_n25377_;
  assign new_n25318_ = ~pi0347;
  assign new_n25319_ = ~new_n25381_ | ~new_n25380_;
  assign new_n25320_ = ~new_n25383_ | ~new_n25382_;
  assign new_n25321_ = ~new_n25385_ | ~new_n25384_;
  assign new_n25322_ = ~new_n25387_ | ~new_n25386_;
  assign new_n25323_ = ~new_n25389_ | ~new_n25388_;
  assign new_n25324_ = ~new_n25391_ | ~new_n25390_;
  assign new_n25325_ = ~new_n25393_ | ~new_n25392_;
  assign new_n25326_ = ~new_n25395_ | ~new_n25394_;
  assign new_n25327_ = ~new_n25397_ | ~new_n25396_;
  assign new_n25328_ = ~new_n25399_ | ~new_n25398_;
  assign new_n25329_ = ~new_n25401_ | ~new_n25400_;
  assign new_n25330_ = ~new_n25403_ | ~new_n25402_;
  assign new_n25331_ = ~new_n25405_ | ~new_n25404_;
  assign new_n25332_ = ~new_n25407_ | ~new_n25406_;
  assign new_n25333_ = ~new_n25409_ | ~new_n25408_;
  assign new_n25334_ = ~new_n25411_ | ~new_n25410_;
  assign new_n25335_ = ~new_n25413_ | ~new_n25412_;
  assign new_n25336_ = ~new_n25415_ | ~new_n25414_;
  assign new_n25337_ = ~new_n25417_ | ~new_n25416_;
  assign new_n25338_ = ~new_n25419_ | ~new_n25418_;
  assign new_n25339_ = ~new_n25421_ | ~new_n25420_;
  assign new_n25340_ = ~new_n25423_ | ~new_n25422_;
  assign new_n25341_ = ~new_n25425_ | ~new_n25424_;
  assign new_n25342_ = ~new_n25427_ | ~new_n25426_;
  assign new_n25343_ = ~new_n25429_ | ~new_n25428_;
  assign new_n25344_ = ~new_n25431_ | ~new_n25430_;
  assign new_n25345_ = ~new_n25433_ | ~new_n25432_;
  assign new_n25346_ = ~new_n25435_ | ~new_n25434_;
  assign new_n25347_ = ~new_n25437_ | ~new_n25436_;
  assign new_n25348_ = ~new_n25439_ | ~new_n25438_;
  assign new_n25349_ = ~pi0348;
  assign new_n25350_ = ~pi0347 | ~new_n25378_;
  assign new_n25351_ = ~new_n25263_;
  assign new_n25352_ = ~new_n25265_;
  assign new_n25353_ = ~new_n25267_;
  assign new_n25354_ = ~new_n25269_;
  assign new_n25355_ = ~new_n25271_;
  assign new_n25356_ = ~new_n25273_;
  assign new_n25357_ = ~new_n25276_;
  assign new_n25358_ = ~new_n25277_;
  assign new_n25359_ = ~new_n25279_;
  assign new_n25360_ = ~new_n25281_;
  assign new_n25361_ = ~new_n25283_;
  assign new_n25362_ = ~new_n25285_;
  assign new_n25363_ = ~new_n25287_;
  assign new_n25364_ = ~new_n25289_;
  assign new_n25365_ = ~new_n25291_;
  assign new_n25366_ = ~new_n25293_;
  assign new_n25367_ = ~new_n25295_;
  assign new_n25368_ = ~new_n25297_;
  assign new_n25369_ = ~new_n25299_;
  assign new_n25370_ = ~new_n25301_;
  assign new_n25371_ = ~new_n25303_;
  assign new_n25372_ = ~new_n25305_;
  assign new_n25373_ = ~new_n25307_;
  assign new_n25374_ = ~new_n25309_;
  assign new_n25375_ = ~new_n25311_;
  assign new_n25376_ = ~new_n25313_;
  assign new_n25377_ = ~new_n25315_;
  assign new_n25378_ = ~new_n25317_;
  assign new_n25379_ = ~new_n25350_;
  assign new_n25380_ = ~pi0326 | ~new_n25276_;
  assign new_n25381_ = ~new_n25357_ | ~new_n25275_;
  assign new_n25382_ = ~pi0325 | ~new_n25273_;
  assign new_n25383_ = ~new_n25356_ | ~new_n25274_;
  assign new_n25384_ = ~pi0324 | ~new_n25271_;
  assign new_n25385_ = ~new_n25355_ | ~new_n25272_;
  assign new_n25386_ = ~pi0323 | ~new_n25269_;
  assign new_n25387_ = ~new_n25354_ | ~new_n25270_;
  assign new_n25388_ = ~pi0322 | ~new_n25267_;
  assign new_n25389_ = ~new_n25353_ | ~new_n25268_;
  assign new_n25390_ = ~pi0321 | ~new_n25265_;
  assign new_n25391_ = ~new_n25352_ | ~new_n25266_;
  assign new_n25392_ = ~pi0320 | ~new_n25263_;
  assign new_n25393_ = ~new_n25351_ | ~new_n25264_;
  assign new_n25394_ = ~pi0348 | ~new_n25350_;
  assign new_n25395_ = ~new_n25379_ | ~new_n25349_;
  assign new_n25396_ = ~pi0347 | ~new_n25317_;
  assign new_n25397_ = ~new_n25378_ | ~new_n25318_;
  assign new_n25398_ = ~pi0319 | ~new_n25261_;
  assign new_n25399_ = ~pi0318 | ~new_n25262_;
  assign new_n25400_ = ~pi0346 | ~new_n25315_;
  assign new_n25401_ = ~new_n25377_ | ~new_n25316_;
  assign new_n25402_ = ~pi0345 | ~new_n25313_;
  assign new_n25403_ = ~new_n25376_ | ~new_n25314_;
  assign new_n25404_ = ~pi0344 | ~new_n25311_;
  assign new_n25405_ = ~new_n25375_ | ~new_n25312_;
  assign new_n25406_ = ~pi0343 | ~new_n25309_;
  assign new_n25407_ = ~new_n25374_ | ~new_n25310_;
  assign new_n25408_ = ~pi0342 | ~new_n25307_;
  assign new_n25409_ = ~new_n25373_ | ~new_n25308_;
  assign new_n25410_ = ~pi0341 | ~new_n25305_;
  assign new_n25411_ = ~new_n25372_ | ~new_n25306_;
  assign new_n25412_ = ~pi0340 | ~new_n25303_;
  assign new_n25413_ = ~new_n25371_ | ~new_n25304_;
  assign new_n25414_ = ~pi0339 | ~new_n25301_;
  assign new_n25415_ = ~new_n25370_ | ~new_n25302_;
  assign new_n25416_ = ~pi0338 | ~new_n25299_;
  assign new_n25417_ = ~new_n25369_ | ~new_n25300_;
  assign new_n25418_ = ~pi0337 | ~new_n25297_;
  assign new_n25419_ = ~new_n25368_ | ~new_n25298_;
  assign new_n25420_ = ~pi0336 | ~new_n25295_;
  assign new_n25421_ = ~new_n25367_ | ~new_n25296_;
  assign new_n25422_ = ~pi0335 | ~new_n25293_;
  assign new_n25423_ = ~new_n25366_ | ~new_n25294_;
  assign new_n25424_ = ~pi0334 | ~new_n25291_;
  assign new_n25425_ = ~new_n25365_ | ~new_n25292_;
  assign new_n25426_ = ~pi0333 | ~new_n25289_;
  assign new_n25427_ = ~new_n25364_ | ~new_n25290_;
  assign new_n25428_ = ~pi0332 | ~new_n25287_;
  assign new_n25429_ = ~new_n25363_ | ~new_n25288_;
  assign new_n25430_ = ~pi0331 | ~new_n25285_;
  assign new_n25431_ = ~new_n25362_ | ~new_n25286_;
  assign new_n25432_ = ~pi0330 | ~new_n25283_;
  assign new_n25433_ = ~new_n25361_ | ~new_n25284_;
  assign new_n25434_ = ~pi0329 | ~new_n25281_;
  assign new_n25435_ = ~new_n25360_ | ~new_n25282_;
  assign new_n25436_ = ~pi0328 | ~new_n25279_;
  assign new_n25437_ = ~new_n25359_ | ~new_n25280_;
  assign new_n25438_ = ~pi0327 | ~new_n25277_;
  assign new_n25439_ = ~new_n25358_ | ~new_n25278_;
  assign new_n25440_ = ~pi0317;
  assign new_n25441_ = ~pi0318;
  assign new_n25442_ = ~pi0318 | ~pi0317;
  assign new_n25443_ = ~pi0319;
  assign new_n25444_ = ~pi0319 | ~new_n25533_;
  assign new_n25445_ = ~pi0320;
  assign new_n25446_ = ~pi0320 | ~new_n25534_;
  assign new_n25447_ = ~pi0321;
  assign new_n25448_ = ~pi0321 | ~new_n25535_;
  assign new_n25449_ = ~pi0322;
  assign new_n25450_ = ~pi0322 | ~new_n25536_;
  assign new_n25451_ = ~pi0323;
  assign new_n25452_ = ~pi0323 | ~new_n25537_;
  assign new_n25453_ = ~pi0324;
  assign new_n25454_ = ~pi0324 | ~new_n25538_;
  assign new_n25455_ = ~pi0325;
  assign new_n25456_ = ~pi0326;
  assign new_n25457_ = ~pi0325 | ~new_n25539_;
  assign new_n25458_ = ~new_n25540_ | ~pi0326;
  assign new_n25459_ = ~pi0327;
  assign new_n25460_ = ~pi0327 | ~new_n25541_;
  assign new_n25461_ = ~pi0328;
  assign new_n25462_ = ~pi0328 | ~new_n25542_;
  assign new_n25463_ = ~pi0329;
  assign new_n25464_ = ~pi0329 | ~new_n25543_;
  assign new_n25465_ = ~pi0330;
  assign new_n25466_ = ~pi0330 | ~new_n25544_;
  assign new_n25467_ = ~pi0331;
  assign new_n25468_ = ~pi0331 | ~new_n25545_;
  assign new_n25469_ = ~pi0332;
  assign new_n25470_ = ~pi0332 | ~new_n25546_;
  assign new_n25471_ = ~pi0333;
  assign new_n25472_ = ~pi0333 | ~new_n25547_;
  assign new_n25473_ = ~pi0334;
  assign new_n25474_ = ~pi0334 | ~new_n25548_;
  assign new_n25475_ = ~pi0335;
  assign new_n25476_ = ~pi0335 | ~new_n25549_;
  assign new_n25477_ = ~pi0336;
  assign new_n25478_ = ~pi0336 | ~new_n25550_;
  assign new_n25479_ = ~pi0337;
  assign new_n25480_ = ~pi0337 | ~new_n25551_;
  assign new_n25481_ = ~pi0338;
  assign new_n25482_ = ~pi0338 | ~new_n25552_;
  assign new_n25483_ = ~pi0339;
  assign new_n25484_ = ~pi0339 | ~new_n25553_;
  assign new_n25485_ = ~pi0340;
  assign new_n25486_ = ~pi0340 | ~new_n25554_;
  assign new_n25487_ = ~pi0341;
  assign new_n25488_ = ~pi0341 | ~new_n25555_;
  assign new_n25489_ = ~pi0342;
  assign new_n25490_ = ~pi0342 | ~new_n25556_;
  assign new_n25491_ = ~pi0343;
  assign new_n25492_ = ~pi0343 | ~new_n25557_;
  assign new_n25493_ = ~pi0344;
  assign new_n25494_ = ~pi0344 | ~new_n25558_;
  assign new_n25495_ = ~pi0345;
  assign new_n25496_ = ~pi0345 | ~new_n25559_;
  assign new_n25497_ = ~pi0346;
  assign new_n25498_ = ~pi0346 | ~new_n25560_;
  assign new_n25499_ = ~pi0347;
  assign new_n25500_ = ~new_n25564_ | ~new_n25563_;
  assign new_n25501_ = ~new_n25566_ | ~new_n25565_;
  assign new_n25502_ = ~new_n25568_ | ~new_n25567_;
  assign new_n25503_ = ~new_n25570_ | ~new_n25569_;
  assign new_n25504_ = ~new_n25572_ | ~new_n25571_;
  assign new_n25505_ = ~new_n25574_ | ~new_n25573_;
  assign new_n25506_ = ~new_n25576_ | ~new_n25575_;
  assign new_n25507_ = ~new_n25578_ | ~new_n25577_;
  assign new_n25508_ = ~new_n25580_ | ~new_n25579_;
  assign new_n25509_ = ~new_n25582_ | ~new_n25581_;
  assign new_n25510_ = ~new_n25584_ | ~new_n25583_;
  assign new_n25511_ = ~new_n25586_ | ~new_n25585_;
  assign new_n25512_ = ~new_n25588_ | ~new_n25587_;
  assign new_n25513_ = ~new_n25590_ | ~new_n25589_;
  assign new_n25514_ = ~new_n25592_ | ~new_n25591_;
  assign new_n25515_ = ~new_n25594_ | ~new_n25593_;
  assign new_n25516_ = ~new_n25596_ | ~new_n25595_;
  assign new_n25517_ = ~new_n25598_ | ~new_n25597_;
  assign new_n25518_ = ~new_n25600_ | ~new_n25599_;
  assign new_n25519_ = ~new_n25602_ | ~new_n25601_;
  assign new_n25520_ = ~new_n25604_ | ~new_n25603_;
  assign new_n25521_ = ~new_n25606_ | ~new_n25605_;
  assign new_n25522_ = ~new_n25608_ | ~new_n25607_;
  assign new_n25523_ = ~new_n25610_ | ~new_n25609_;
  assign new_n25524_ = ~new_n25612_ | ~new_n25611_;
  assign new_n25525_ = ~new_n25614_ | ~new_n25613_;
  assign new_n25526_ = ~new_n25616_ | ~new_n25615_;
  assign new_n25527_ = ~new_n25618_ | ~new_n25617_;
  assign new_n25528_ = ~new_n25620_ | ~new_n25619_;
  assign new_n25529_ = ~new_n25622_ | ~new_n25621_;
  assign new_n25530_ = ~new_n25624_ | ~new_n25623_;
  assign new_n25531_ = ~pi0348;
  assign new_n25532_ = ~pi0347 | ~new_n25561_;
  assign new_n25533_ = ~new_n25442_;
  assign new_n25534_ = ~new_n25444_;
  assign new_n25535_ = ~new_n25446_;
  assign new_n25536_ = ~new_n25448_;
  assign new_n25537_ = ~new_n25450_;
  assign new_n25538_ = ~new_n25452_;
  assign new_n25539_ = ~new_n25454_;
  assign new_n25540_ = ~new_n25457_;
  assign new_n25541_ = ~new_n25458_;
  assign new_n25542_ = ~new_n25460_;
  assign new_n25543_ = ~new_n25462_;
  assign new_n25544_ = ~new_n25464_;
  assign new_n25545_ = ~new_n25466_;
  assign new_n25546_ = ~new_n25468_;
  assign new_n25547_ = ~new_n25470_;
  assign new_n25548_ = ~new_n25472_;
  assign new_n25549_ = ~new_n25474_;
  assign new_n25550_ = ~new_n25476_;
  assign new_n25551_ = ~new_n25478_;
  assign new_n25552_ = ~new_n25480_;
  assign new_n25553_ = ~new_n25482_;
  assign new_n25554_ = ~new_n25484_;
  assign new_n25555_ = ~new_n25486_;
  assign new_n25556_ = ~new_n25488_;
  assign new_n25557_ = ~new_n25490_;
  assign new_n25558_ = ~new_n25492_;
  assign new_n25559_ = ~new_n25494_;
  assign new_n25560_ = ~new_n25496_;
  assign new_n25561_ = ~new_n25498_;
  assign new_n25562_ = ~new_n25532_;
  assign new_n25563_ = ~pi0326 | ~new_n25457_;
  assign new_n25564_ = ~new_n25540_ | ~new_n25456_;
  assign new_n25565_ = ~pi0325 | ~new_n25454_;
  assign new_n25566_ = ~new_n25539_ | ~new_n25455_;
  assign new_n25567_ = ~pi0324 | ~new_n25452_;
  assign new_n25568_ = ~new_n25538_ | ~new_n25453_;
  assign new_n25569_ = ~pi0323 | ~new_n25450_;
  assign new_n25570_ = ~new_n25537_ | ~new_n25451_;
  assign new_n25571_ = ~pi0322 | ~new_n25448_;
  assign new_n25572_ = ~new_n25536_ | ~new_n25449_;
  assign new_n25573_ = ~pi0321 | ~new_n25446_;
  assign new_n25574_ = ~new_n25535_ | ~new_n25447_;
  assign new_n25575_ = ~pi0320 | ~new_n25444_;
  assign new_n25576_ = ~new_n25534_ | ~new_n25445_;
  assign new_n25577_ = ~pi0348 | ~new_n25532_;
  assign new_n25578_ = ~new_n25562_ | ~new_n25531_;
  assign new_n25579_ = ~pi0347 | ~new_n25498_;
  assign new_n25580_ = ~new_n25561_ | ~new_n25499_;
  assign new_n25581_ = ~pi0319 | ~new_n25442_;
  assign new_n25582_ = ~new_n25533_ | ~new_n25443_;
  assign new_n25583_ = ~pi0346 | ~new_n25496_;
  assign new_n25584_ = ~new_n25560_ | ~new_n25497_;
  assign new_n25585_ = ~pi0345 | ~new_n25494_;
  assign new_n25586_ = ~new_n25559_ | ~new_n25495_;
  assign new_n25587_ = ~pi0344 | ~new_n25492_;
  assign new_n25588_ = ~new_n25558_ | ~new_n25493_;
  assign new_n25589_ = ~pi0343 | ~new_n25490_;
  assign new_n25590_ = ~new_n25557_ | ~new_n25491_;
  assign new_n25591_ = ~pi0342 | ~new_n25488_;
  assign new_n25592_ = ~new_n25556_ | ~new_n25489_;
  assign new_n25593_ = ~pi0341 | ~new_n25486_;
  assign new_n25594_ = ~new_n25555_ | ~new_n25487_;
  assign new_n25595_ = ~pi0340 | ~new_n25484_;
  assign new_n25596_ = ~new_n25554_ | ~new_n25485_;
  assign new_n25597_ = ~pi0339 | ~new_n25482_;
  assign new_n25598_ = ~new_n25553_ | ~new_n25483_;
  assign new_n25599_ = ~pi0338 | ~new_n25480_;
  assign new_n25600_ = ~new_n25552_ | ~new_n25481_;
  assign new_n25601_ = ~pi0337 | ~new_n25478_;
  assign new_n25602_ = ~new_n25551_ | ~new_n25479_;
  assign new_n25603_ = ~pi0318 | ~new_n25440_;
  assign new_n25604_ = ~pi0317 | ~new_n25441_;
  assign new_n25605_ = ~pi0336 | ~new_n25476_;
  assign new_n25606_ = ~new_n25550_ | ~new_n25477_;
  assign new_n25607_ = ~pi0335 | ~new_n25474_;
  assign new_n25608_ = ~new_n25549_ | ~new_n25475_;
  assign new_n25609_ = ~pi0334 | ~new_n25472_;
  assign new_n25610_ = ~new_n25548_ | ~new_n25473_;
  assign new_n25611_ = ~pi0333 | ~new_n25470_;
  assign new_n25612_ = ~new_n25547_ | ~new_n25471_;
  assign new_n25613_ = ~pi0332 | ~new_n25468_;
  assign new_n25614_ = ~new_n25546_ | ~new_n25469_;
  assign new_n25615_ = ~pi0331 | ~new_n25466_;
  assign new_n25616_ = ~new_n25545_ | ~new_n25467_;
  assign new_n25617_ = ~pi0330 | ~new_n25464_;
  assign new_n25618_ = ~new_n25544_ | ~new_n25465_;
  assign new_n25619_ = ~pi0329 | ~new_n25462_;
  assign new_n25620_ = ~new_n25543_ | ~new_n25463_;
  assign new_n25621_ = ~pi0328 | ~new_n25460_;
  assign new_n25622_ = ~new_n25542_ | ~new_n25461_;
  assign new_n25623_ = ~pi0327 | ~new_n25458_;
  assign new_n25624_ = ~new_n25541_ | ~new_n25459_;
  assign new_n25625_ = ~pi0317;
  assign new_n25626_ = ~new_n25713_ | ~new_n25747_;
  assign new_n25627_ = ~pi0318;
  assign new_n25628_ = ~pi0320;
  assign new_n25629_ = ~pi0320 | ~new_n25713_;
  assign new_n25630_ = ~pi0321;
  assign new_n25631_ = ~pi0321 | ~new_n25719_;
  assign new_n25632_ = ~pi0322;
  assign new_n25633_ = ~pi0322 | ~new_n25720_;
  assign new_n25634_ = ~pi0323;
  assign new_n25635_ = ~pi0323 | ~new_n25721_;
  assign new_n25636_ = ~pi0324;
  assign new_n25637_ = ~pi0324 | ~new_n25722_;
  assign new_n25638_ = ~pi0325;
  assign new_n25639_ = ~pi0326;
  assign new_n25640_ = ~pi0325 | ~new_n25723_;
  assign new_n25641_ = ~new_n25724_ | ~pi0326;
  assign new_n25642_ = ~pi0327;
  assign new_n25643_ = ~pi0327 | ~new_n25725_;
  assign new_n25644_ = ~pi0328;
  assign new_n25645_ = ~pi0328 | ~new_n25726_;
  assign new_n25646_ = ~pi0329;
  assign new_n25647_ = ~pi0329 | ~new_n25727_;
  assign new_n25648_ = ~pi0330;
  assign new_n25649_ = ~pi0330 | ~new_n25728_;
  assign new_n25650_ = ~pi0331;
  assign new_n25651_ = ~pi0331 | ~new_n25729_;
  assign new_n25652_ = ~pi0332;
  assign new_n25653_ = ~pi0332 | ~new_n25730_;
  assign new_n25654_ = ~pi0333;
  assign new_n25655_ = ~pi0333 | ~new_n25731_;
  assign new_n25656_ = ~pi0334;
  assign new_n25657_ = ~pi0334 | ~new_n25732_;
  assign new_n25658_ = ~pi0335;
  assign new_n25659_ = ~pi0335 | ~new_n25733_;
  assign new_n25660_ = ~pi0336;
  assign new_n25661_ = ~pi0336 | ~new_n25734_;
  assign new_n25662_ = ~pi0337;
  assign new_n25663_ = ~pi0337 | ~new_n25735_;
  assign new_n25664_ = ~pi0338;
  assign new_n25665_ = ~pi0338 | ~new_n25736_;
  assign new_n25666_ = ~pi0339;
  assign new_n25667_ = ~pi0339 | ~new_n25737_;
  assign new_n25668_ = ~pi0340;
  assign new_n25669_ = ~pi0340 | ~new_n25738_;
  assign new_n25670_ = ~pi0341;
  assign new_n25671_ = ~pi0341 | ~new_n25739_;
  assign new_n25672_ = ~pi0342;
  assign new_n25673_ = ~pi0342 | ~new_n25740_;
  assign new_n25674_ = ~pi0343;
  assign new_n25675_ = ~pi0343 | ~new_n25741_;
  assign new_n25676_ = ~pi0344;
  assign new_n25677_ = ~pi0344 | ~new_n25742_;
  assign new_n25678_ = ~pi0345;
  assign new_n25679_ = ~pi0345 | ~new_n25743_;
  assign new_n25680_ = ~pi0346;
  assign new_n25681_ = ~pi0346 | ~new_n25744_;
  assign new_n25682_ = ~pi0347;
  assign new_n25683_ = ~pi0319;
  assign new_n25684_ = ~new_n25749_ | ~new_n25748_;
  assign new_n25685_ = ~new_n25751_ | ~new_n25750_;
  assign new_n25686_ = ~new_n25753_ | ~new_n25752_;
  assign new_n25687_ = ~new_n25755_ | ~new_n25754_;
  assign new_n25688_ = ~new_n25757_ | ~new_n25756_;
  assign new_n25689_ = ~new_n25759_ | ~new_n25758_;
  assign new_n25690_ = ~new_n25763_ | ~new_n25762_;
  assign new_n25691_ = ~new_n25765_ | ~new_n25764_;
  assign new_n25692_ = ~new_n25767_ | ~new_n25766_;
  assign new_n25693_ = ~new_n25769_ | ~new_n25768_;
  assign new_n25694_ = ~new_n25771_ | ~new_n25770_;
  assign new_n25695_ = ~new_n25773_ | ~new_n25772_;
  assign new_n25696_ = ~new_n25775_ | ~new_n25774_;
  assign new_n25697_ = ~new_n25777_ | ~new_n25776_;
  assign new_n25698_ = ~new_n25779_ | ~new_n25778_;
  assign new_n25699_ = ~new_n25781_ | ~new_n25780_;
  assign new_n25700_ = ~new_n25783_ | ~new_n25782_;
  assign new_n25701_ = ~new_n25785_ | ~new_n25784_;
  assign new_n25702_ = ~new_n25787_ | ~new_n25786_;
  assign new_n25703_ = ~new_n25789_ | ~new_n25788_;
  assign new_n25704_ = ~new_n25791_ | ~new_n25790_;
  assign new_n25705_ = ~new_n25793_ | ~new_n25792_;
  assign new_n25706_ = ~new_n25795_ | ~new_n25794_;
  assign new_n25707_ = ~new_n25797_ | ~new_n25796_;
  assign new_n25708_ = ~new_n25799_ | ~new_n25798_;
  assign new_n25709_ = ~new_n25801_ | ~new_n25800_;
  assign new_n25710_ = ~new_n25803_ | ~new_n25802_;
  assign new_n25711_ = ~new_n25805_ | ~new_n25804_;
  assign new_n25712_ = ~new_n25807_ | ~new_n25806_;
  assign new_n25713_ = ~new_n25683_ | ~new_n25717_;
  assign new_n25714_ = new_n25761_ & new_n25760_;
  assign new_n25715_ = ~pi0348;
  assign new_n25716_ = ~pi0347 | ~new_n25745_;
  assign new_n25717_ = ~pi0318 | ~pi0317;
  assign new_n25718_ = ~new_n25713_;
  assign new_n25719_ = ~new_n25629_;
  assign new_n25720_ = ~new_n25631_;
  assign new_n25721_ = ~new_n25633_;
  assign new_n25722_ = ~new_n25635_;
  assign new_n25723_ = ~new_n25637_;
  assign new_n25724_ = ~new_n25640_;
  assign new_n25725_ = ~new_n25641_;
  assign new_n25726_ = ~new_n25643_;
  assign new_n25727_ = ~new_n25645_;
  assign new_n25728_ = ~new_n25647_;
  assign new_n25729_ = ~new_n25649_;
  assign new_n25730_ = ~new_n25651_;
  assign new_n25731_ = ~new_n25653_;
  assign new_n25732_ = ~new_n25655_;
  assign new_n25733_ = ~new_n25657_;
  assign new_n25734_ = ~new_n25659_;
  assign new_n25735_ = ~new_n25661_;
  assign new_n25736_ = ~new_n25663_;
  assign new_n25737_ = ~new_n25665_;
  assign new_n25738_ = ~new_n25667_;
  assign new_n25739_ = ~new_n25669_;
  assign new_n25740_ = ~new_n25671_;
  assign new_n25741_ = ~new_n25673_;
  assign new_n25742_ = ~new_n25675_;
  assign new_n25743_ = ~new_n25677_;
  assign new_n25744_ = ~new_n25679_;
  assign new_n25745_ = ~new_n25681_;
  assign new_n25746_ = ~new_n25716_;
  assign new_n25747_ = ~pi0319 | ~pi0318 | ~pi0317;
  assign new_n25748_ = ~pi0326 | ~new_n25640_;
  assign new_n25749_ = ~new_n25724_ | ~new_n25639_;
  assign new_n25750_ = ~pi0325 | ~new_n25637_;
  assign new_n25751_ = ~new_n25723_ | ~new_n25638_;
  assign new_n25752_ = ~pi0324 | ~new_n25635_;
  assign new_n25753_ = ~new_n25722_ | ~new_n25636_;
  assign new_n25754_ = ~pi0323 | ~new_n25633_;
  assign new_n25755_ = ~new_n25721_ | ~new_n25634_;
  assign new_n25756_ = ~pi0322 | ~new_n25631_;
  assign new_n25757_ = ~new_n25720_ | ~new_n25632_;
  assign new_n25758_ = ~pi0321 | ~new_n25629_;
  assign new_n25759_ = ~new_n25719_ | ~new_n25630_;
  assign new_n25760_ = ~pi0320 | ~new_n25713_;
  assign new_n25761_ = ~new_n25718_ | ~new_n25628_;
  assign new_n25762_ = ~pi0348 | ~new_n25716_;
  assign new_n25763_ = ~new_n25746_ | ~new_n25715_;
  assign new_n25764_ = ~pi0347 | ~new_n25681_;
  assign new_n25765_ = ~new_n25745_ | ~new_n25682_;
  assign new_n25766_ = ~pi0346 | ~new_n25679_;
  assign new_n25767_ = ~new_n25744_ | ~new_n25680_;
  assign new_n25768_ = ~pi0345 | ~new_n25677_;
  assign new_n25769_ = ~new_n25743_ | ~new_n25678_;
  assign new_n25770_ = ~pi0344 | ~new_n25675_;
  assign new_n25771_ = ~new_n25742_ | ~new_n25676_;
  assign new_n25772_ = ~pi0343 | ~new_n25673_;
  assign new_n25773_ = ~new_n25741_ | ~new_n25674_;
  assign new_n25774_ = ~pi0342 | ~new_n25671_;
  assign new_n25775_ = ~new_n25740_ | ~new_n25672_;
  assign new_n25776_ = ~pi0341 | ~new_n25669_;
  assign new_n25777_ = ~new_n25739_ | ~new_n25670_;
  assign new_n25778_ = ~pi0340 | ~new_n25667_;
  assign new_n25779_ = ~new_n25738_ | ~new_n25668_;
  assign new_n25780_ = ~pi0339 | ~new_n25665_;
  assign new_n25781_ = ~new_n25737_ | ~new_n25666_;
  assign new_n25782_ = ~pi0338 | ~new_n25663_;
  assign new_n25783_ = ~new_n25736_ | ~new_n25664_;
  assign new_n25784_ = ~pi0337 | ~new_n25661_;
  assign new_n25785_ = ~new_n25735_ | ~new_n25662_;
  assign new_n25786_ = ~pi0318 | ~new_n25625_;
  assign new_n25787_ = ~pi0317 | ~new_n25627_;
  assign new_n25788_ = ~pi0336 | ~new_n25659_;
  assign new_n25789_ = ~new_n25734_ | ~new_n25660_;
  assign new_n25790_ = ~pi0335 | ~new_n25657_;
  assign new_n25791_ = ~new_n25733_ | ~new_n25658_;
  assign new_n25792_ = ~pi0334 | ~new_n25655_;
  assign new_n25793_ = ~new_n25732_ | ~new_n25656_;
  assign new_n25794_ = ~pi0333 | ~new_n25653_;
  assign new_n25795_ = ~new_n25731_ | ~new_n25654_;
  assign new_n25796_ = ~pi0332 | ~new_n25651_;
  assign new_n25797_ = ~new_n25730_ | ~new_n25652_;
  assign new_n25798_ = ~pi0331 | ~new_n25649_;
  assign new_n25799_ = ~new_n25729_ | ~new_n25650_;
  assign new_n25800_ = ~pi0330 | ~new_n25647_;
  assign new_n25801_ = ~new_n25728_ | ~new_n25648_;
  assign new_n25802_ = ~pi0329 | ~new_n25645_;
  assign new_n25803_ = ~new_n25727_ | ~new_n25646_;
  assign new_n25804_ = ~pi0328 | ~new_n25643_;
  assign new_n25805_ = ~new_n25726_ | ~new_n25644_;
  assign new_n25806_ = ~pi0327 | ~new_n25641_;
  assign new_n25807_ = ~new_n25725_ | ~new_n25642_;
  assign new_n25808_ = ~pi0317;
  assign new_n25809_ = ~pi0318;
  assign new_n25810_ = ~pi0318 | ~pi0317;
  assign new_n25811_ = ~pi0319;
  assign new_n25812_ = ~pi0319 | ~new_n25901_;
  assign new_n25813_ = ~pi0320;
  assign new_n25814_ = ~pi0320 | ~new_n25902_;
  assign new_n25815_ = ~pi0321;
  assign new_n25816_ = ~pi0321 | ~new_n25903_;
  assign new_n25817_ = ~pi0322;
  assign new_n25818_ = ~pi0322 | ~new_n25904_;
  assign new_n25819_ = ~pi0323;
  assign new_n25820_ = ~pi0323 | ~new_n25905_;
  assign new_n25821_ = ~pi0324;
  assign new_n25822_ = ~pi0324 | ~new_n25906_;
  assign new_n25823_ = ~pi0325;
  assign new_n25824_ = ~pi0326;
  assign new_n25825_ = ~pi0325 | ~new_n25907_;
  assign new_n25826_ = ~new_n25908_ | ~pi0326;
  assign new_n25827_ = ~pi0327;
  assign new_n25828_ = ~pi0327 | ~new_n25909_;
  assign new_n25829_ = ~pi0328;
  assign new_n25830_ = ~pi0328 | ~new_n25910_;
  assign new_n25831_ = ~pi0329;
  assign new_n25832_ = ~pi0329 | ~new_n25911_;
  assign new_n25833_ = ~pi0330;
  assign new_n25834_ = ~pi0330 | ~new_n25912_;
  assign new_n25835_ = ~pi0331;
  assign new_n25836_ = ~pi0331 | ~new_n25913_;
  assign new_n25837_ = ~pi0332;
  assign new_n25838_ = ~pi0332 | ~new_n25914_;
  assign new_n25839_ = ~pi0333;
  assign new_n25840_ = ~pi0333 | ~new_n25915_;
  assign new_n25841_ = ~pi0334;
  assign new_n25842_ = ~pi0334 | ~new_n25916_;
  assign new_n25843_ = ~pi0335;
  assign new_n25844_ = ~pi0335 | ~new_n25917_;
  assign new_n25845_ = ~pi0336;
  assign new_n25846_ = ~pi0336 | ~new_n25918_;
  assign new_n25847_ = ~pi0337;
  assign new_n25848_ = ~pi0337 | ~new_n25919_;
  assign new_n25849_ = ~pi0338;
  assign new_n25850_ = ~pi0338 | ~new_n25920_;
  assign new_n25851_ = ~pi0339;
  assign new_n25852_ = ~pi0339 | ~new_n25921_;
  assign new_n25853_ = ~pi0340;
  assign new_n25854_ = ~pi0340 | ~new_n25922_;
  assign new_n25855_ = ~pi0341;
  assign new_n25856_ = ~pi0341 | ~new_n25923_;
  assign new_n25857_ = ~pi0342;
  assign new_n25858_ = ~pi0342 | ~new_n25924_;
  assign new_n25859_ = ~pi0343;
  assign new_n25860_ = ~pi0343 | ~new_n25925_;
  assign new_n25861_ = ~pi0344;
  assign new_n25862_ = ~pi0344 | ~new_n25926_;
  assign new_n25863_ = ~pi0345;
  assign new_n25864_ = ~pi0345 | ~new_n25927_;
  assign new_n25865_ = ~pi0346;
  assign new_n25866_ = ~pi0346 | ~new_n25928_;
  assign new_n25867_ = ~pi0347;
  assign new_n25868_ = ~new_n25932_ | ~new_n25931_;
  assign new_n25869_ = ~new_n25934_ | ~new_n25933_;
  assign new_n25870_ = ~new_n25936_ | ~new_n25935_;
  assign new_n25871_ = ~new_n25938_ | ~new_n25937_;
  assign new_n25872_ = ~new_n25940_ | ~new_n25939_;
  assign new_n25873_ = ~new_n25942_ | ~new_n25941_;
  assign new_n25874_ = ~new_n25944_ | ~new_n25943_;
  assign new_n25875_ = ~new_n25946_ | ~new_n25945_;
  assign new_n25876_ = ~new_n25948_ | ~new_n25947_;
  assign new_n25877_ = ~new_n25950_ | ~new_n25949_;
  assign new_n25878_ = ~new_n25952_ | ~new_n25951_;
  assign new_n25879_ = ~new_n25954_ | ~new_n25953_;
  assign new_n25880_ = ~new_n25956_ | ~new_n25955_;
  assign new_n25881_ = ~new_n25958_ | ~new_n25957_;
  assign new_n25882_ = ~new_n25960_ | ~new_n25959_;
  assign new_n25883_ = ~new_n25962_ | ~new_n25961_;
  assign new_n25884_ = ~new_n25964_ | ~new_n25963_;
  assign new_n25885_ = ~new_n25966_ | ~new_n25965_;
  assign new_n25886_ = ~new_n25968_ | ~new_n25967_;
  assign new_n25887_ = ~new_n25970_ | ~new_n25969_;
  assign new_n25888_ = ~new_n25972_ | ~new_n25971_;
  assign new_n25889_ = ~new_n25974_ | ~new_n25973_;
  assign new_n25890_ = ~new_n25976_ | ~new_n25975_;
  assign new_n25891_ = ~new_n25978_ | ~new_n25977_;
  assign new_n25892_ = ~new_n25980_ | ~new_n25979_;
  assign new_n25893_ = ~new_n25982_ | ~new_n25981_;
  assign new_n25894_ = ~new_n25984_ | ~new_n25983_;
  assign new_n25895_ = ~new_n25986_ | ~new_n25985_;
  assign new_n25896_ = ~new_n25988_ | ~new_n25987_;
  assign new_n25897_ = ~new_n25990_ | ~new_n25989_;
  assign new_n25898_ = ~new_n25992_ | ~new_n25991_;
  assign new_n25899_ = ~pi0348;
  assign new_n25900_ = ~pi0347 | ~new_n25929_;
  assign new_n25901_ = ~new_n25810_;
  assign new_n25902_ = ~new_n25812_;
  assign new_n25903_ = ~new_n25814_;
  assign new_n25904_ = ~new_n25816_;
  assign new_n25905_ = ~new_n25818_;
  assign new_n25906_ = ~new_n25820_;
  assign new_n25907_ = ~new_n25822_;
  assign new_n25908_ = ~new_n25825_;
  assign new_n25909_ = ~new_n25826_;
  assign new_n25910_ = ~new_n25828_;
  assign new_n25911_ = ~new_n25830_;
  assign new_n25912_ = ~new_n25832_;
  assign new_n25913_ = ~new_n25834_;
  assign new_n25914_ = ~new_n25836_;
  assign new_n25915_ = ~new_n25838_;
  assign new_n25916_ = ~new_n25840_;
  assign new_n25917_ = ~new_n25842_;
  assign new_n25918_ = ~new_n25844_;
  assign new_n25919_ = ~new_n25846_;
  assign new_n25920_ = ~new_n25848_;
  assign new_n25921_ = ~new_n25850_;
  assign new_n25922_ = ~new_n25852_;
  assign new_n25923_ = ~new_n25854_;
  assign new_n25924_ = ~new_n25856_;
  assign new_n25925_ = ~new_n25858_;
  assign new_n25926_ = ~new_n25860_;
  assign new_n25927_ = ~new_n25862_;
  assign new_n25928_ = ~new_n25864_;
  assign new_n25929_ = ~new_n25866_;
  assign new_n25930_ = ~new_n25900_;
  assign new_n25931_ = ~pi0326 | ~new_n25825_;
  assign new_n25932_ = ~new_n25908_ | ~new_n25824_;
  assign new_n25933_ = ~pi0325 | ~new_n25822_;
  assign new_n25934_ = ~new_n25907_ | ~new_n25823_;
  assign new_n25935_ = ~pi0324 | ~new_n25820_;
  assign new_n25936_ = ~new_n25906_ | ~new_n25821_;
  assign new_n25937_ = ~pi0323 | ~new_n25818_;
  assign new_n25938_ = ~new_n25905_ | ~new_n25819_;
  assign new_n25939_ = ~pi0322 | ~new_n25816_;
  assign new_n25940_ = ~new_n25904_ | ~new_n25817_;
  assign new_n25941_ = ~pi0321 | ~new_n25814_;
  assign new_n25942_ = ~new_n25903_ | ~new_n25815_;
  assign new_n25943_ = ~pi0320 | ~new_n25812_;
  assign new_n25944_ = ~new_n25902_ | ~new_n25813_;
  assign new_n25945_ = ~pi0348 | ~new_n25900_;
  assign new_n25946_ = ~new_n25930_ | ~new_n25899_;
  assign new_n25947_ = ~pi0347 | ~new_n25866_;
  assign new_n25948_ = ~new_n25929_ | ~new_n25867_;
  assign new_n25949_ = ~pi0319 | ~new_n25810_;
  assign new_n25950_ = ~new_n25901_ | ~new_n25811_;
  assign new_n25951_ = ~pi0346 | ~new_n25864_;
  assign new_n25952_ = ~new_n25928_ | ~new_n25865_;
  assign new_n25953_ = ~pi0345 | ~new_n25862_;
  assign new_n25954_ = ~new_n25927_ | ~new_n25863_;
  assign new_n25955_ = ~pi0344 | ~new_n25860_;
  assign new_n25956_ = ~new_n25926_ | ~new_n25861_;
  assign new_n25957_ = ~pi0343 | ~new_n25858_;
  assign new_n25958_ = ~new_n25925_ | ~new_n25859_;
  assign new_n25959_ = ~pi0342 | ~new_n25856_;
  assign new_n25960_ = ~new_n25924_ | ~new_n25857_;
  assign new_n25961_ = ~pi0341 | ~new_n25854_;
  assign new_n25962_ = ~new_n25923_ | ~new_n25855_;
  assign new_n25963_ = ~pi0340 | ~new_n25852_;
  assign new_n25964_ = ~new_n25922_ | ~new_n25853_;
  assign new_n25965_ = ~pi0339 | ~new_n25850_;
  assign new_n25966_ = ~new_n25921_ | ~new_n25851_;
  assign new_n25967_ = ~pi0338 | ~new_n25848_;
  assign new_n25968_ = ~new_n25920_ | ~new_n25849_;
  assign new_n25969_ = ~pi0337 | ~new_n25846_;
  assign new_n25970_ = ~new_n25919_ | ~new_n25847_;
  assign new_n25971_ = ~pi0318 | ~new_n25808_;
  assign new_n25972_ = ~pi0317 | ~new_n25809_;
  assign new_n25973_ = ~pi0336 | ~new_n25844_;
  assign new_n25974_ = ~new_n25918_ | ~new_n25845_;
  assign new_n25975_ = ~pi0335 | ~new_n25842_;
  assign new_n25976_ = ~new_n25917_ | ~new_n25843_;
  assign new_n25977_ = ~pi0334 | ~new_n25840_;
  assign new_n25978_ = ~new_n25916_ | ~new_n25841_;
  assign new_n25979_ = ~pi0333 | ~new_n25838_;
  assign new_n25980_ = ~new_n25915_ | ~new_n25839_;
  assign new_n25981_ = ~pi0332 | ~new_n25836_;
  assign new_n25982_ = ~new_n25914_ | ~new_n25837_;
  assign new_n25983_ = ~pi0331 | ~new_n25834_;
  assign new_n25984_ = ~new_n25913_ | ~new_n25835_;
  assign new_n25985_ = ~pi0330 | ~new_n25832_;
  assign new_n25986_ = ~new_n25912_ | ~new_n25833_;
  assign new_n25987_ = ~pi0329 | ~new_n25830_;
  assign new_n25988_ = ~new_n25911_ | ~new_n25831_;
  assign new_n25989_ = ~pi0328 | ~new_n25828_;
  assign new_n25990_ = ~new_n25910_ | ~new_n25829_;
  assign new_n25991_ = ~pi0327 | ~new_n25826_;
  assign new_n25992_ = ~new_n25909_ | ~new_n25827_;
  assign new_n25993_ = ~pi0317;
  assign new_n25994_ = ~pi0318;
  assign new_n25995_ = ~pi0318 | ~pi0317;
  assign new_n25996_ = ~pi0319;
  assign new_n25997_ = ~pi0319 | ~new_n26086_;
  assign new_n25998_ = ~pi0320;
  assign new_n25999_ = ~pi0320 | ~new_n26087_;
  assign new_n26000_ = ~pi0321;
  assign new_n26001_ = ~pi0321 | ~new_n26088_;
  assign new_n26002_ = ~pi0322;
  assign new_n26003_ = ~pi0322 | ~new_n26089_;
  assign new_n26004_ = ~pi0323;
  assign new_n26005_ = ~pi0323 | ~new_n26090_;
  assign new_n26006_ = ~pi0324;
  assign new_n26007_ = ~pi0324 | ~new_n26091_;
  assign new_n26008_ = ~pi0325;
  assign new_n26009_ = ~pi0326;
  assign new_n26010_ = ~pi0325 | ~new_n26092_;
  assign new_n26011_ = ~new_n26093_ | ~pi0326;
  assign new_n26012_ = ~pi0327;
  assign new_n26013_ = ~pi0327 | ~new_n26094_;
  assign new_n26014_ = ~pi0328;
  assign new_n26015_ = ~pi0328 | ~new_n26095_;
  assign new_n26016_ = ~pi0329;
  assign new_n26017_ = ~pi0329 | ~new_n26096_;
  assign new_n26018_ = ~pi0330;
  assign new_n26019_ = ~pi0330 | ~new_n26097_;
  assign new_n26020_ = ~pi0331;
  assign new_n26021_ = ~pi0331 | ~new_n26098_;
  assign new_n26022_ = ~pi0332;
  assign new_n26023_ = ~pi0332 | ~new_n26099_;
  assign new_n26024_ = ~pi0333;
  assign new_n26025_ = ~pi0333 | ~new_n26100_;
  assign new_n26026_ = ~pi0334;
  assign new_n26027_ = ~pi0334 | ~new_n26101_;
  assign new_n26028_ = ~pi0335;
  assign new_n26029_ = ~pi0335 | ~new_n26102_;
  assign new_n26030_ = ~pi0336;
  assign new_n26031_ = ~pi0336 | ~new_n26103_;
  assign new_n26032_ = ~pi0337;
  assign new_n26033_ = ~pi0337 | ~new_n26104_;
  assign new_n26034_ = ~pi0338;
  assign new_n26035_ = ~pi0338 | ~new_n26105_;
  assign new_n26036_ = ~pi0339;
  assign new_n26037_ = ~pi0339 | ~new_n26106_;
  assign new_n26038_ = ~pi0340;
  assign new_n26039_ = ~pi0340 | ~new_n26107_;
  assign new_n26040_ = ~pi0341;
  assign new_n26041_ = ~pi0341 | ~new_n26108_;
  assign new_n26042_ = ~pi0342;
  assign new_n26043_ = ~pi0342 | ~new_n26109_;
  assign new_n26044_ = ~pi0343;
  assign new_n26045_ = ~pi0343 | ~new_n26110_;
  assign new_n26046_ = ~pi0344;
  assign new_n26047_ = ~pi0344 | ~new_n26111_;
  assign new_n26048_ = ~pi0345;
  assign new_n26049_ = ~pi0345 | ~new_n26112_;
  assign new_n26050_ = ~pi0346;
  assign new_n26051_ = ~pi0346 | ~new_n26113_;
  assign new_n26052_ = ~pi0347;
  assign new_n26053_ = ~new_n26117_ | ~new_n26116_;
  assign new_n26054_ = ~new_n26119_ | ~new_n26118_;
  assign new_n26055_ = ~new_n26121_ | ~new_n26120_;
  assign new_n26056_ = ~new_n26123_ | ~new_n26122_;
  assign new_n26057_ = ~new_n26125_ | ~new_n26124_;
  assign new_n26058_ = ~new_n26127_ | ~new_n26126_;
  assign new_n26059_ = ~new_n26129_ | ~new_n26128_;
  assign new_n26060_ = ~new_n26131_ | ~new_n26130_;
  assign new_n26061_ = ~new_n26133_ | ~new_n26132_;
  assign new_n26062_ = ~new_n26135_ | ~new_n26134_;
  assign new_n26063_ = ~new_n26137_ | ~new_n26136_;
  assign new_n26064_ = ~new_n26139_ | ~new_n26138_;
  assign new_n26065_ = ~new_n26141_ | ~new_n26140_;
  assign new_n26066_ = ~new_n26143_ | ~new_n26142_;
  assign new_n26067_ = ~new_n26145_ | ~new_n26144_;
  assign new_n26068_ = ~new_n26147_ | ~new_n26146_;
  assign new_n26069_ = ~new_n26149_ | ~new_n26148_;
  assign new_n26070_ = ~new_n26151_ | ~new_n26150_;
  assign new_n26071_ = ~new_n26153_ | ~new_n26152_;
  assign new_n26072_ = ~new_n26155_ | ~new_n26154_;
  assign new_n26073_ = ~new_n26157_ | ~new_n26156_;
  assign new_n26074_ = ~new_n26159_ | ~new_n26158_;
  assign new_n26075_ = ~new_n26161_ | ~new_n26160_;
  assign new_n26076_ = ~new_n26163_ | ~new_n26162_;
  assign new_n26077_ = ~new_n26165_ | ~new_n26164_;
  assign new_n26078_ = ~new_n26167_ | ~new_n26166_;
  assign new_n26079_ = ~new_n26169_ | ~new_n26168_;
  assign new_n26080_ = ~new_n26171_ | ~new_n26170_;
  assign new_n26081_ = ~new_n26173_ | ~new_n26172_;
  assign new_n26082_ = ~new_n26175_ | ~new_n26174_;
  assign new_n26083_ = ~new_n26177_ | ~new_n26176_;
  assign new_n26084_ = ~pi0348;
  assign new_n26085_ = ~pi0347 | ~new_n26114_;
  assign new_n26086_ = ~new_n25995_;
  assign new_n26087_ = ~new_n25997_;
  assign new_n26088_ = ~new_n25999_;
  assign new_n26089_ = ~new_n26001_;
  assign new_n26090_ = ~new_n26003_;
  assign new_n26091_ = ~new_n26005_;
  assign new_n26092_ = ~new_n26007_;
  assign new_n26093_ = ~new_n26010_;
  assign new_n26094_ = ~new_n26011_;
  assign new_n26095_ = ~new_n26013_;
  assign new_n26096_ = ~new_n26015_;
  assign new_n26097_ = ~new_n26017_;
  assign new_n26098_ = ~new_n26019_;
  assign new_n26099_ = ~new_n26021_;
  assign new_n26100_ = ~new_n26023_;
  assign new_n26101_ = ~new_n26025_;
  assign new_n26102_ = ~new_n26027_;
  assign new_n26103_ = ~new_n26029_;
  assign new_n26104_ = ~new_n26031_;
  assign new_n26105_ = ~new_n26033_;
  assign new_n26106_ = ~new_n26035_;
  assign new_n26107_ = ~new_n26037_;
  assign new_n26108_ = ~new_n26039_;
  assign new_n26109_ = ~new_n26041_;
  assign new_n26110_ = ~new_n26043_;
  assign new_n26111_ = ~new_n26045_;
  assign new_n26112_ = ~new_n26047_;
  assign new_n26113_ = ~new_n26049_;
  assign new_n26114_ = ~new_n26051_;
  assign new_n26115_ = ~new_n26085_;
  assign new_n26116_ = ~pi0326 | ~new_n26010_;
  assign new_n26117_ = ~new_n26093_ | ~new_n26009_;
  assign new_n26118_ = ~pi0325 | ~new_n26007_;
  assign new_n26119_ = ~new_n26092_ | ~new_n26008_;
  assign new_n26120_ = ~pi0324 | ~new_n26005_;
  assign new_n26121_ = ~new_n26091_ | ~new_n26006_;
  assign new_n26122_ = ~pi0323 | ~new_n26003_;
  assign new_n26123_ = ~new_n26090_ | ~new_n26004_;
  assign new_n26124_ = ~pi0322 | ~new_n26001_;
  assign new_n26125_ = ~new_n26089_ | ~new_n26002_;
  assign new_n26126_ = ~pi0321 | ~new_n25999_;
  assign new_n26127_ = ~new_n26088_ | ~new_n26000_;
  assign new_n26128_ = ~pi0320 | ~new_n25997_;
  assign new_n26129_ = ~new_n26087_ | ~new_n25998_;
  assign new_n26130_ = ~pi0348 | ~new_n26085_;
  assign new_n26131_ = ~new_n26115_ | ~new_n26084_;
  assign new_n26132_ = ~pi0347 | ~new_n26051_;
  assign new_n26133_ = ~new_n26114_ | ~new_n26052_;
  assign new_n26134_ = ~pi0319 | ~new_n25995_;
  assign new_n26135_ = ~new_n26086_ | ~new_n25996_;
  assign new_n26136_ = ~pi0346 | ~new_n26049_;
  assign new_n26137_ = ~new_n26113_ | ~new_n26050_;
  assign new_n26138_ = ~pi0345 | ~new_n26047_;
  assign new_n26139_ = ~new_n26112_ | ~new_n26048_;
  assign new_n26140_ = ~pi0344 | ~new_n26045_;
  assign new_n26141_ = ~new_n26111_ | ~new_n26046_;
  assign new_n26142_ = ~pi0343 | ~new_n26043_;
  assign new_n26143_ = ~new_n26110_ | ~new_n26044_;
  assign new_n26144_ = ~pi0342 | ~new_n26041_;
  assign new_n26145_ = ~new_n26109_ | ~new_n26042_;
  assign new_n26146_ = ~pi0341 | ~new_n26039_;
  assign new_n26147_ = ~new_n26108_ | ~new_n26040_;
  assign new_n26148_ = ~pi0340 | ~new_n26037_;
  assign new_n26149_ = ~new_n26107_ | ~new_n26038_;
  assign new_n26150_ = ~pi0339 | ~new_n26035_;
  assign new_n26151_ = ~new_n26106_ | ~new_n26036_;
  assign new_n26152_ = ~pi0338 | ~new_n26033_;
  assign new_n26153_ = ~new_n26105_ | ~new_n26034_;
  assign new_n26154_ = ~pi0337 | ~new_n26031_;
  assign new_n26155_ = ~new_n26104_ | ~new_n26032_;
  assign new_n26156_ = ~pi0318 | ~new_n25993_;
  assign new_n26157_ = ~pi0317 | ~new_n25994_;
  assign new_n26158_ = ~pi0336 | ~new_n26029_;
  assign new_n26159_ = ~new_n26103_ | ~new_n26030_;
  assign new_n26160_ = ~pi0335 | ~new_n26027_;
  assign new_n26161_ = ~new_n26102_ | ~new_n26028_;
  assign new_n26162_ = ~pi0334 | ~new_n26025_;
  assign new_n26163_ = ~new_n26101_ | ~new_n26026_;
  assign new_n26164_ = ~pi0333 | ~new_n26023_;
  assign new_n26165_ = ~new_n26100_ | ~new_n26024_;
  assign new_n26166_ = ~pi0332 | ~new_n26021_;
  assign new_n26167_ = ~new_n26099_ | ~new_n26022_;
  assign new_n26168_ = ~pi0331 | ~new_n26019_;
  assign new_n26169_ = ~new_n26098_ | ~new_n26020_;
  assign new_n26170_ = ~pi0330 | ~new_n26017_;
  assign new_n26171_ = ~new_n26097_ | ~new_n26018_;
  assign new_n26172_ = ~pi0329 | ~new_n26015_;
  assign new_n26173_ = ~new_n26096_ | ~new_n26016_;
  assign new_n26174_ = ~pi0328 | ~new_n26013_;
  assign new_n26175_ = ~new_n26095_ | ~new_n26014_;
  assign new_n26176_ = ~pi0327 | ~new_n26011_;
  assign new_n26177_ = ~new_n26094_ | ~new_n26012_;
  assign new_n26178_ = ~pi0317;
  assign new_n26179_ = ~pi0318;
  assign new_n26180_ = ~pi0318 | ~pi0317;
  assign new_n26181_ = ~pi0319;
  assign new_n26182_ = ~pi0319 | ~new_n26271_;
  assign new_n26183_ = ~pi0320;
  assign new_n26184_ = ~pi0320 | ~new_n26272_;
  assign new_n26185_ = ~pi0321;
  assign new_n26186_ = ~pi0321 | ~new_n26273_;
  assign new_n26187_ = ~pi0322;
  assign new_n26188_ = ~pi0322 | ~new_n26274_;
  assign new_n26189_ = ~pi0323;
  assign new_n26190_ = ~pi0323 | ~new_n26275_;
  assign new_n26191_ = ~pi0324;
  assign new_n26192_ = ~pi0324 | ~new_n26276_;
  assign new_n26193_ = ~pi0325;
  assign new_n26194_ = ~pi0326;
  assign new_n26195_ = ~pi0325 | ~new_n26277_;
  assign new_n26196_ = ~new_n26278_ | ~pi0326;
  assign new_n26197_ = ~pi0327;
  assign new_n26198_ = ~pi0327 | ~new_n26279_;
  assign new_n26199_ = ~pi0328;
  assign new_n26200_ = ~pi0328 | ~new_n26280_;
  assign new_n26201_ = ~pi0329;
  assign new_n26202_ = ~pi0329 | ~new_n26281_;
  assign new_n26203_ = ~pi0330;
  assign new_n26204_ = ~pi0330 | ~new_n26282_;
  assign new_n26205_ = ~pi0331;
  assign new_n26206_ = ~pi0331 | ~new_n26283_;
  assign new_n26207_ = ~pi0332;
  assign new_n26208_ = ~pi0332 | ~new_n26284_;
  assign new_n26209_ = ~pi0333;
  assign new_n26210_ = ~pi0333 | ~new_n26285_;
  assign new_n26211_ = ~pi0334;
  assign new_n26212_ = ~pi0334 | ~new_n26286_;
  assign new_n26213_ = ~pi0335;
  assign new_n26214_ = ~pi0335 | ~new_n26287_;
  assign new_n26215_ = ~pi0336;
  assign new_n26216_ = ~pi0336 | ~new_n26288_;
  assign new_n26217_ = ~pi0337;
  assign new_n26218_ = ~pi0337 | ~new_n26289_;
  assign new_n26219_ = ~pi0338;
  assign new_n26220_ = ~pi0338 | ~new_n26290_;
  assign new_n26221_ = ~pi0339;
  assign new_n26222_ = ~pi0339 | ~new_n26291_;
  assign new_n26223_ = ~pi0340;
  assign new_n26224_ = ~pi0340 | ~new_n26292_;
  assign new_n26225_ = ~pi0341;
  assign new_n26226_ = ~pi0341 | ~new_n26293_;
  assign new_n26227_ = ~pi0342;
  assign new_n26228_ = ~pi0342 | ~new_n26294_;
  assign new_n26229_ = ~pi0343;
  assign new_n26230_ = ~pi0343 | ~new_n26295_;
  assign new_n26231_ = ~pi0344;
  assign new_n26232_ = ~pi0344 | ~new_n26296_;
  assign new_n26233_ = ~pi0345;
  assign new_n26234_ = ~pi0345 | ~new_n26297_;
  assign new_n26235_ = ~pi0346;
  assign new_n26236_ = ~pi0346 | ~new_n26298_;
  assign new_n26237_ = ~pi0347;
  assign new_n26238_ = ~new_n26302_ | ~new_n26301_;
  assign new_n26239_ = ~new_n26304_ | ~new_n26303_;
  assign new_n26240_ = ~new_n26306_ | ~new_n26305_;
  assign new_n26241_ = ~new_n26308_ | ~new_n26307_;
  assign new_n26242_ = ~new_n26310_ | ~new_n26309_;
  assign new_n26243_ = ~new_n26312_ | ~new_n26311_;
  assign new_n26244_ = ~new_n26314_ | ~new_n26313_;
  assign new_n26245_ = ~new_n26316_ | ~new_n26315_;
  assign new_n26246_ = ~new_n26318_ | ~new_n26317_;
  assign new_n26247_ = ~new_n26320_ | ~new_n26319_;
  assign new_n26248_ = ~new_n26322_ | ~new_n26321_;
  assign new_n26249_ = ~new_n26324_ | ~new_n26323_;
  assign new_n26250_ = ~new_n26326_ | ~new_n26325_;
  assign new_n26251_ = ~new_n26328_ | ~new_n26327_;
  assign new_n26252_ = ~new_n26330_ | ~new_n26329_;
  assign new_n26253_ = ~new_n26332_ | ~new_n26331_;
  assign new_n26254_ = ~new_n26334_ | ~new_n26333_;
  assign new_n26255_ = ~new_n26336_ | ~new_n26335_;
  assign new_n26256_ = ~new_n26338_ | ~new_n26337_;
  assign new_n26257_ = ~new_n26340_ | ~new_n26339_;
  assign new_n26258_ = ~new_n26342_ | ~new_n26341_;
  assign new_n26259_ = ~new_n26344_ | ~new_n26343_;
  assign new_n26260_ = ~new_n26346_ | ~new_n26345_;
  assign new_n26261_ = ~new_n26348_ | ~new_n26347_;
  assign new_n26262_ = ~new_n26350_ | ~new_n26349_;
  assign new_n26263_ = ~new_n26352_ | ~new_n26351_;
  assign new_n26264_ = ~new_n26354_ | ~new_n26353_;
  assign new_n26265_ = ~new_n26356_ | ~new_n26355_;
  assign new_n26266_ = ~new_n26358_ | ~new_n26357_;
  assign new_n26267_ = ~new_n26360_ | ~new_n26359_;
  assign new_n26268_ = ~new_n26362_ | ~new_n26361_;
  assign new_n26269_ = ~pi0348;
  assign new_n26270_ = ~pi0347 | ~new_n26299_;
  assign new_n26271_ = ~new_n26180_;
  assign new_n26272_ = ~new_n26182_;
  assign new_n26273_ = ~new_n26184_;
  assign new_n26274_ = ~new_n26186_;
  assign new_n26275_ = ~new_n26188_;
  assign new_n26276_ = ~new_n26190_;
  assign new_n26277_ = ~new_n26192_;
  assign new_n26278_ = ~new_n26195_;
  assign new_n26279_ = ~new_n26196_;
  assign new_n26280_ = ~new_n26198_;
  assign new_n26281_ = ~new_n26200_;
  assign new_n26282_ = ~new_n26202_;
  assign new_n26283_ = ~new_n26204_;
  assign new_n26284_ = ~new_n26206_;
  assign new_n26285_ = ~new_n26208_;
  assign new_n26286_ = ~new_n26210_;
  assign new_n26287_ = ~new_n26212_;
  assign new_n26288_ = ~new_n26214_;
  assign new_n26289_ = ~new_n26216_;
  assign new_n26290_ = ~new_n26218_;
  assign new_n26291_ = ~new_n26220_;
  assign new_n26292_ = ~new_n26222_;
  assign new_n26293_ = ~new_n26224_;
  assign new_n26294_ = ~new_n26226_;
  assign new_n26295_ = ~new_n26228_;
  assign new_n26296_ = ~new_n26230_;
  assign new_n26297_ = ~new_n26232_;
  assign new_n26298_ = ~new_n26234_;
  assign new_n26299_ = ~new_n26236_;
  assign new_n26300_ = ~new_n26270_;
  assign new_n26301_ = ~pi0326 | ~new_n26195_;
  assign new_n26302_ = ~new_n26278_ | ~new_n26194_;
  assign new_n26303_ = ~pi0325 | ~new_n26192_;
  assign new_n26304_ = ~new_n26277_ | ~new_n26193_;
  assign new_n26305_ = ~pi0324 | ~new_n26190_;
  assign new_n26306_ = ~new_n26276_ | ~new_n26191_;
  assign new_n26307_ = ~pi0323 | ~new_n26188_;
  assign new_n26308_ = ~new_n26275_ | ~new_n26189_;
  assign new_n26309_ = ~pi0322 | ~new_n26186_;
  assign new_n26310_ = ~new_n26274_ | ~new_n26187_;
  assign new_n26311_ = ~pi0321 | ~new_n26184_;
  assign new_n26312_ = ~new_n26273_ | ~new_n26185_;
  assign new_n26313_ = ~pi0320 | ~new_n26182_;
  assign new_n26314_ = ~new_n26272_ | ~new_n26183_;
  assign new_n26315_ = ~pi0348 | ~new_n26270_;
  assign new_n26316_ = ~new_n26300_ | ~new_n26269_;
  assign new_n26317_ = ~pi0347 | ~new_n26236_;
  assign new_n26318_ = ~new_n26299_ | ~new_n26237_;
  assign new_n26319_ = ~pi0319 | ~new_n26180_;
  assign new_n26320_ = ~new_n26271_ | ~new_n26181_;
  assign new_n26321_ = ~pi0346 | ~new_n26234_;
  assign new_n26322_ = ~new_n26298_ | ~new_n26235_;
  assign new_n26323_ = ~pi0345 | ~new_n26232_;
  assign new_n26324_ = ~new_n26297_ | ~new_n26233_;
  assign new_n26325_ = ~pi0344 | ~new_n26230_;
  assign new_n26326_ = ~new_n26296_ | ~new_n26231_;
  assign new_n26327_ = ~pi0343 | ~new_n26228_;
  assign new_n26328_ = ~new_n26295_ | ~new_n26229_;
  assign new_n26329_ = ~pi0342 | ~new_n26226_;
  assign new_n26330_ = ~new_n26294_ | ~new_n26227_;
  assign new_n26331_ = ~pi0341 | ~new_n26224_;
  assign new_n26332_ = ~new_n26293_ | ~new_n26225_;
  assign new_n26333_ = ~pi0340 | ~new_n26222_;
  assign new_n26334_ = ~new_n26292_ | ~new_n26223_;
  assign new_n26335_ = ~pi0339 | ~new_n26220_;
  assign new_n26336_ = ~new_n26291_ | ~new_n26221_;
  assign new_n26337_ = ~pi0338 | ~new_n26218_;
  assign new_n26338_ = ~new_n26290_ | ~new_n26219_;
  assign new_n26339_ = ~pi0337 | ~new_n26216_;
  assign new_n26340_ = ~new_n26289_ | ~new_n26217_;
  assign new_n26341_ = ~pi0318 | ~new_n26178_;
  assign new_n26342_ = ~pi0317 | ~new_n26179_;
  assign new_n26343_ = ~pi0336 | ~new_n26214_;
  assign new_n26344_ = ~new_n26288_ | ~new_n26215_;
  assign new_n26345_ = ~pi0335 | ~new_n26212_;
  assign new_n26346_ = ~new_n26287_ | ~new_n26213_;
  assign new_n26347_ = ~pi0334 | ~new_n26210_;
  assign new_n26348_ = ~new_n26286_ | ~new_n26211_;
  assign new_n26349_ = ~pi0333 | ~new_n26208_;
  assign new_n26350_ = ~new_n26285_ | ~new_n26209_;
  assign new_n26351_ = ~pi0332 | ~new_n26206_;
  assign new_n26352_ = ~new_n26284_ | ~new_n26207_;
  assign new_n26353_ = ~pi0331 | ~new_n26204_;
  assign new_n26354_ = ~new_n26283_ | ~new_n26205_;
  assign new_n26355_ = ~pi0330 | ~new_n26202_;
  assign new_n26356_ = ~new_n26282_ | ~new_n26203_;
  assign new_n26357_ = ~pi0329 | ~new_n26200_;
  assign new_n26358_ = ~new_n26281_ | ~new_n26201_;
  assign new_n26359_ = ~pi0328 | ~new_n26198_;
  assign new_n26360_ = ~new_n26280_ | ~new_n26199_;
  assign new_n26361_ = ~pi0327 | ~new_n26196_;
  assign new_n26362_ = ~new_n26279_ | ~new_n26197_;
  assign new_n26363_ = ~new_n26372_ | ~new_n26380_;
  assign new_n26364_ = new_n26386_ & new_n26368_;
  assign new_n26365_ = new_n26384_ & new_n26369_;
  assign new_n26366_ = new_n26382_ & new_n26363_;
  assign new_n26367_ = ~new_n27123_;
  assign new_n26368_ = new_n27125_ | new_n27124_ | new_n27120_;
  assign new_n26369_ = ~new_n26371_ | ~new_n26379_;
  assign new_n26370_ = ~new_n26392_ | ~new_n26391_;
  assign new_n26371_ = ~new_n27126_ & ~new_n27122_;
  assign new_n26372_ = ~new_n27119_ & ~new_n27121_;
  assign new_n26373_ = ~new_n27119_;
  assign new_n26374_ = new_n26388_ & new_n26387_;
  assign new_n26375_ = ~new_n27126_;
  assign new_n26376_ = new_n26390_ & new_n26389_;
  assign new_n26377_ = ~new_n27120_;
  assign new_n26378_ = ~new_n27125_;
  assign new_n26379_ = ~new_n26368_;
  assign new_n26380_ = ~new_n26369_;
  assign new_n26381_ = ~new_n26380_ | ~new_n26373_;
  assign new_n26382_ = ~new_n27121_ | ~new_n26381_;
  assign new_n26383_ = ~new_n26379_ | ~new_n26375_;
  assign new_n26384_ = ~new_n27122_ | ~new_n26383_;
  assign new_n26385_ = new_n27120_ | new_n27125_;
  assign new_n26386_ = ~new_n27124_ | ~new_n26385_;
  assign new_n26387_ = ~new_n27119_ | ~new_n26369_;
  assign new_n26388_ = ~new_n26380_ | ~new_n26373_;
  assign new_n26389_ = ~new_n27126_ | ~new_n26368_;
  assign new_n26390_ = ~new_n26379_ | ~new_n26375_;
  assign new_n26391_ = ~new_n27120_ | ~new_n26378_;
  assign new_n26392_ = ~new_n27125_ | ~new_n26377_;
  assign new_n26393_ = ~pi0317;
  assign new_n26394_ = ~pi0318;
  assign new_n26395_ = ~pi0318 | ~pi0317;
  assign new_n26396_ = ~pi0319;
  assign new_n26397_ = ~pi0319 | ~new_n26486_;
  assign new_n26398_ = ~pi0320;
  assign new_n26399_ = ~pi0320 | ~new_n26487_;
  assign new_n26400_ = ~pi0321;
  assign new_n26401_ = ~pi0321 | ~new_n26488_;
  assign new_n26402_ = ~pi0322;
  assign new_n26403_ = ~pi0322 | ~new_n26489_;
  assign new_n26404_ = ~pi0323;
  assign new_n26405_ = ~pi0323 | ~new_n26490_;
  assign new_n26406_ = ~pi0324;
  assign new_n26407_ = ~pi0324 | ~new_n26491_;
  assign new_n26408_ = ~pi0325;
  assign new_n26409_ = ~pi0326;
  assign new_n26410_ = ~pi0325 | ~new_n26492_;
  assign new_n26411_ = ~new_n26493_ | ~pi0326;
  assign new_n26412_ = ~pi0327;
  assign new_n26413_ = ~pi0327 | ~new_n26494_;
  assign new_n26414_ = ~pi0328;
  assign new_n26415_ = ~pi0328 | ~new_n26495_;
  assign new_n26416_ = ~pi0329;
  assign new_n26417_ = ~pi0329 | ~new_n26496_;
  assign new_n26418_ = ~pi0330;
  assign new_n26419_ = ~pi0330 | ~new_n26497_;
  assign new_n26420_ = ~pi0331;
  assign new_n26421_ = ~pi0331 | ~new_n26498_;
  assign new_n26422_ = ~pi0332;
  assign new_n26423_ = ~pi0332 | ~new_n26499_;
  assign new_n26424_ = ~pi0333;
  assign new_n26425_ = ~pi0333 | ~new_n26500_;
  assign new_n26426_ = ~pi0334;
  assign new_n26427_ = ~pi0334 | ~new_n26501_;
  assign new_n26428_ = ~pi0335;
  assign new_n26429_ = ~pi0335 | ~new_n26502_;
  assign new_n26430_ = ~pi0336;
  assign new_n26431_ = ~pi0336 | ~new_n26503_;
  assign new_n26432_ = ~pi0337;
  assign new_n26433_ = ~pi0337 | ~new_n26504_;
  assign new_n26434_ = ~pi0338;
  assign new_n26435_ = ~pi0338 | ~new_n26505_;
  assign new_n26436_ = ~pi0339;
  assign new_n26437_ = ~pi0339 | ~new_n26506_;
  assign new_n26438_ = ~pi0340;
  assign new_n26439_ = ~pi0340 | ~new_n26507_;
  assign new_n26440_ = ~pi0341;
  assign new_n26441_ = ~pi0341 | ~new_n26508_;
  assign new_n26442_ = ~pi0342;
  assign new_n26443_ = ~pi0342 | ~new_n26509_;
  assign new_n26444_ = ~pi0343;
  assign new_n26445_ = ~pi0343 | ~new_n26510_;
  assign new_n26446_ = ~pi0344;
  assign new_n26447_ = ~pi0344 | ~new_n26511_;
  assign new_n26448_ = ~pi0345;
  assign new_n26449_ = ~pi0345 | ~new_n26512_;
  assign new_n26450_ = ~pi0346;
  assign new_n26451_ = ~pi0346 | ~new_n26513_;
  assign new_n26452_ = ~pi0347;
  assign new_n26453_ = ~new_n26517_ | ~new_n26516_;
  assign new_n26454_ = ~new_n26519_ | ~new_n26518_;
  assign new_n26455_ = ~new_n26521_ | ~new_n26520_;
  assign new_n26456_ = ~new_n26523_ | ~new_n26522_;
  assign new_n26457_ = ~new_n26525_ | ~new_n26524_;
  assign new_n26458_ = ~new_n26527_ | ~new_n26526_;
  assign new_n26459_ = ~new_n26529_ | ~new_n26528_;
  assign new_n26460_ = ~new_n26531_ | ~new_n26530_;
  assign new_n26461_ = ~new_n26533_ | ~new_n26532_;
  assign new_n26462_ = ~new_n26535_ | ~new_n26534_;
  assign new_n26463_ = ~new_n26537_ | ~new_n26536_;
  assign new_n26464_ = ~new_n26539_ | ~new_n26538_;
  assign new_n26465_ = ~new_n26541_ | ~new_n26540_;
  assign new_n26466_ = ~new_n26543_ | ~new_n26542_;
  assign new_n26467_ = ~new_n26545_ | ~new_n26544_;
  assign new_n26468_ = ~new_n26547_ | ~new_n26546_;
  assign new_n26469_ = ~new_n26549_ | ~new_n26548_;
  assign new_n26470_ = ~new_n26551_ | ~new_n26550_;
  assign new_n26471_ = ~new_n26553_ | ~new_n26552_;
  assign new_n26472_ = ~new_n26555_ | ~new_n26554_;
  assign new_n26473_ = ~new_n26557_ | ~new_n26556_;
  assign new_n26474_ = ~new_n26559_ | ~new_n26558_;
  assign new_n26475_ = ~new_n26561_ | ~new_n26560_;
  assign new_n26476_ = ~new_n26563_ | ~new_n26562_;
  assign new_n26477_ = ~new_n26565_ | ~new_n26564_;
  assign new_n26478_ = ~new_n26567_ | ~new_n26566_;
  assign new_n26479_ = ~new_n26569_ | ~new_n26568_;
  assign new_n26480_ = ~new_n26571_ | ~new_n26570_;
  assign new_n26481_ = ~new_n26573_ | ~new_n26572_;
  assign new_n26482_ = ~new_n26575_ | ~new_n26574_;
  assign new_n26483_ = ~new_n26577_ | ~new_n26576_;
  assign new_n26484_ = ~pi0348;
  assign new_n26485_ = ~pi0347 | ~new_n26514_;
  assign new_n26486_ = ~new_n26395_;
  assign new_n26487_ = ~new_n26397_;
  assign new_n26488_ = ~new_n26399_;
  assign new_n26489_ = ~new_n26401_;
  assign new_n26490_ = ~new_n26403_;
  assign new_n26491_ = ~new_n26405_;
  assign new_n26492_ = ~new_n26407_;
  assign new_n26493_ = ~new_n26410_;
  assign new_n26494_ = ~new_n26411_;
  assign new_n26495_ = ~new_n26413_;
  assign new_n26496_ = ~new_n26415_;
  assign new_n26497_ = ~new_n26417_;
  assign new_n26498_ = ~new_n26419_;
  assign new_n26499_ = ~new_n26421_;
  assign new_n26500_ = ~new_n26423_;
  assign new_n26501_ = ~new_n26425_;
  assign new_n26502_ = ~new_n26427_;
  assign new_n26503_ = ~new_n26429_;
  assign new_n26504_ = ~new_n26431_;
  assign new_n26505_ = ~new_n26433_;
  assign new_n26506_ = ~new_n26435_;
  assign new_n26507_ = ~new_n26437_;
  assign new_n26508_ = ~new_n26439_;
  assign new_n26509_ = ~new_n26441_;
  assign new_n26510_ = ~new_n26443_;
  assign new_n26511_ = ~new_n26445_;
  assign new_n26512_ = ~new_n26447_;
  assign new_n26513_ = ~new_n26449_;
  assign new_n26514_ = ~new_n26451_;
  assign new_n26515_ = ~new_n26485_;
  assign new_n26516_ = ~pi0326 | ~new_n26410_;
  assign new_n26517_ = ~new_n26493_ | ~new_n26409_;
  assign new_n26518_ = ~pi0325 | ~new_n26407_;
  assign new_n26519_ = ~new_n26492_ | ~new_n26408_;
  assign new_n26520_ = ~pi0324 | ~new_n26405_;
  assign new_n26521_ = ~new_n26491_ | ~new_n26406_;
  assign new_n26522_ = ~pi0323 | ~new_n26403_;
  assign new_n26523_ = ~new_n26490_ | ~new_n26404_;
  assign new_n26524_ = ~pi0322 | ~new_n26401_;
  assign new_n26525_ = ~new_n26489_ | ~new_n26402_;
  assign new_n26526_ = ~pi0321 | ~new_n26399_;
  assign new_n26527_ = ~new_n26488_ | ~new_n26400_;
  assign new_n26528_ = ~pi0320 | ~new_n26397_;
  assign new_n26529_ = ~new_n26487_ | ~new_n26398_;
  assign new_n26530_ = ~pi0348 | ~new_n26485_;
  assign new_n26531_ = ~new_n26515_ | ~new_n26484_;
  assign new_n26532_ = ~pi0347 | ~new_n26451_;
  assign new_n26533_ = ~new_n26514_ | ~new_n26452_;
  assign new_n26534_ = ~pi0319 | ~new_n26395_;
  assign new_n26535_ = ~new_n26486_ | ~new_n26396_;
  assign new_n26536_ = ~pi0346 | ~new_n26449_;
  assign new_n26537_ = ~new_n26513_ | ~new_n26450_;
  assign new_n26538_ = ~pi0345 | ~new_n26447_;
  assign new_n26539_ = ~new_n26512_ | ~new_n26448_;
  assign new_n26540_ = ~pi0344 | ~new_n26445_;
  assign new_n26541_ = ~new_n26511_ | ~new_n26446_;
  assign new_n26542_ = ~pi0343 | ~new_n26443_;
  assign new_n26543_ = ~new_n26510_ | ~new_n26444_;
  assign new_n26544_ = ~pi0342 | ~new_n26441_;
  assign new_n26545_ = ~new_n26509_ | ~new_n26442_;
  assign new_n26546_ = ~pi0341 | ~new_n26439_;
  assign new_n26547_ = ~new_n26508_ | ~new_n26440_;
  assign new_n26548_ = ~pi0340 | ~new_n26437_;
  assign new_n26549_ = ~new_n26507_ | ~new_n26438_;
  assign new_n26550_ = ~pi0339 | ~new_n26435_;
  assign new_n26551_ = ~new_n26506_ | ~new_n26436_;
  assign new_n26552_ = ~pi0338 | ~new_n26433_;
  assign new_n26553_ = ~new_n26505_ | ~new_n26434_;
  assign new_n26554_ = ~pi0337 | ~new_n26431_;
  assign new_n26555_ = ~new_n26504_ | ~new_n26432_;
  assign new_n26556_ = ~pi0318 | ~new_n26393_;
  assign new_n26557_ = ~pi0317 | ~new_n26394_;
  assign new_n26558_ = ~pi0336 | ~new_n26429_;
  assign new_n26559_ = ~new_n26503_ | ~new_n26430_;
  assign new_n26560_ = ~pi0335 | ~new_n26427_;
  assign new_n26561_ = ~new_n26502_ | ~new_n26428_;
  assign new_n26562_ = ~pi0334 | ~new_n26425_;
  assign new_n26563_ = ~new_n26501_ | ~new_n26426_;
  assign new_n26564_ = ~pi0333 | ~new_n26423_;
  assign new_n26565_ = ~new_n26500_ | ~new_n26424_;
  assign new_n26566_ = ~pi0332 | ~new_n26421_;
  assign new_n26567_ = ~new_n26499_ | ~new_n26422_;
  assign new_n26568_ = ~pi0331 | ~new_n26419_;
  assign new_n26569_ = ~new_n26498_ | ~new_n26420_;
  assign new_n26570_ = ~pi0330 | ~new_n26417_;
  assign new_n26571_ = ~new_n26497_ | ~new_n26418_;
  assign new_n26572_ = ~pi0329 | ~new_n26415_;
  assign new_n26573_ = ~new_n26496_ | ~new_n26416_;
  assign new_n26574_ = ~pi0328 | ~new_n26413_;
  assign new_n26575_ = ~new_n26495_ | ~new_n26414_;
  assign new_n26576_ = ~pi0327 | ~new_n26411_;
  assign new_n26577_ = ~new_n26494_ | ~new_n26412_;
  assign new_n26578_ = ~new_n26615_ | ~new_n26614_;
  assign new_n26579_ = ~pi0311 | ~new_n26599_;
  assign new_n26580_ = ~pi0315;
  assign new_n26581_ = ~pi0309;
  assign new_n26582_ = ~pi0314;
  assign new_n26583_ = ~pi0308;
  assign new_n26584_ = ~pi0313;
  assign new_n26585_ = ~pi0312;
  assign new_n26586_ = ~new_n26611_ | ~new_n26610_;
  assign new_n26587_ = ~pi0307;
  assign new_n26588_ = ~new_n26620_ | ~new_n26619_;
  assign new_n26589_ = ~new_n26625_ | ~new_n26624_;
  assign new_n26590_ = ~new_n26630_ | ~new_n26629_;
  assign new_n26591_ = ~new_n26635_ | ~new_n26634_;
  assign new_n26592_ = ~new_n26617_ | ~new_n26616_;
  assign new_n26593_ = ~new_n26622_ | ~new_n26621_;
  assign new_n26594_ = ~new_n26627_ | ~new_n26626_;
  assign new_n26595_ = ~new_n26632_ | ~new_n26631_;
  assign new_n26596_ = ~new_n26607_ | ~new_n26606_;
  assign new_n26597_ = ~new_n26603_ | ~new_n26602_;
  assign new_n26598_ = ~pi0310;
  assign new_n26599_ = ~pi0316;
  assign new_n26600_ = ~new_n26579_;
  assign new_n26601_ = ~new_n26600_ | ~new_n26580_;
  assign new_n26602_ = ~new_n26601_ | ~new_n26598_;
  assign new_n26603_ = ~pi0315 | ~new_n26579_;
  assign new_n26604_ = ~new_n26597_;
  assign new_n26605_ = ~pi0309 | ~new_n26582_;
  assign new_n26606_ = ~new_n26605_ | ~new_n26597_;
  assign new_n26607_ = ~pi0314 | ~new_n26581_;
  assign new_n26608_ = ~new_n26596_;
  assign new_n26609_ = ~pi0308 | ~new_n26584_;
  assign new_n26610_ = ~new_n26609_ | ~new_n26596_;
  assign new_n26611_ = ~pi0313 | ~new_n26583_;
  assign new_n26612_ = ~new_n26586_;
  assign new_n26613_ = ~pi0312 | ~new_n26587_;
  assign new_n26614_ = ~new_n26612_ | ~new_n26613_;
  assign new_n26615_ = ~pi0307 | ~new_n26585_;
  assign new_n26616_ = ~pi0307 | ~new_n26585_;
  assign new_n26617_ = ~pi0312 | ~new_n26587_;
  assign new_n26618_ = ~new_n26592_;
  assign new_n26619_ = ~new_n26618_ | ~new_n26612_;
  assign new_n26620_ = ~new_n26592_ | ~new_n26586_;
  assign new_n26621_ = ~pi0308 | ~new_n26584_;
  assign new_n26622_ = ~pi0313 | ~new_n26583_;
  assign new_n26623_ = ~new_n26593_;
  assign new_n26624_ = ~new_n26608_ | ~new_n26623_;
  assign new_n26625_ = ~new_n26593_ | ~new_n26596_;
  assign new_n26626_ = ~pi0309 | ~new_n26582_;
  assign new_n26627_ = ~pi0314 | ~new_n26581_;
  assign new_n26628_ = ~new_n26594_;
  assign new_n26629_ = ~new_n26604_ | ~new_n26628_;
  assign new_n26630_ = ~new_n26594_ | ~new_n26597_;
  assign new_n26631_ = ~pi0310 | ~new_n26580_;
  assign new_n26632_ = ~pi0315 | ~new_n26598_;
  assign new_n26633_ = ~new_n26595_;
  assign new_n26634_ = ~new_n26633_ | ~new_n26600_;
  assign new_n26635_ = ~new_n26595_ | ~new_n26579_;
  assign new_n26636_ = new_n26765_ & new_n26764_;
  assign new_n26637_ = new_n26828_ & new_n26680_;
  assign new_n26638_ = new_n26826_ & new_n26681_;
  assign new_n26639_ = new_n26824_ & new_n26710_;
  assign new_n26640_ = new_n26823_ & new_n26685_;
  assign new_n26641_ = new_n26821_ & new_n26688_;
  assign new_n26642_ = new_n26819_ & new_n26691_;
  assign new_n26643_ = new_n26817_ & new_n26800_;
  assign new_n26644_ = new_n26816_ & new_n26694_;
  assign new_n26645_ = new_n26815_ & new_n26697_;
  assign new_n26646_ = new_n26813_ & new_n26700_;
  assign new_n26647_ = new_n26811_ & new_n26702_;
  assign new_n26648_ = new_n26810_ & new_n26705_;
  assign new_n26649_ = new_n26808_ & new_n26707_;
  assign new_n26650_ = new_n26794_ & new_n26791_;
  assign new_n26651_ = new_n26787_ & new_n26784_;
  assign new_n26652_ = ~new_n26835_ | ~new_n26887_ | ~new_n26886_;
  assign new_n26653_ = ~new_n27033_;
  assign new_n26654_ = ~pi0321;
  assign new_n26655_ = ~pi0322;
  assign new_n26656_ = ~pi0321 | ~new_n27033_;
  assign new_n26657_ = ~new_n27032_;
  assign new_n26658_ = ~new_n27018_;
  assign new_n26659_ = ~pi0319;
  assign new_n26660_ = ~pi0320;
  assign new_n26661_ = ~pi0319 | ~new_n27018_;
  assign new_n26662_ = ~new_n27038_;
  assign new_n26663_ = ~new_n27017_;
  assign new_n26664_ = ~pi0317;
  assign new_n26665_ = ~pi0318;
  assign new_n26666_ = ~pi0317 | ~new_n27017_;
  assign new_n26667_ = ~new_n27034_;
  assign new_n26668_ = ~new_n27031_;
  assign new_n26669_ = ~pi0323;
  assign new_n26670_ = ~pi0324;
  assign new_n26671_ = ~new_n27030_;
  assign new_n26672_ = ~new_n27019_;
  assign new_n26673_ = ~pi0325;
  assign new_n26674_ = ~pi0326;
  assign new_n26675_ = ~new_n26726_ | ~new_n26762_;
  assign new_n26676_ = ~new_n26709_ | ~new_n26755_;
  assign new_n26677_ = ~pi0327;
  assign new_n26678_ = ~pi0328;
  assign new_n26679_ = ~pi0329;
  assign new_n26680_ = ~new_n26731_ | ~new_n26740_;
  assign new_n26681_ = ~new_n26732_ | ~new_n26749_;
  assign new_n26682_ = ~pi0330;
  assign new_n26683_ = ~pi0332;
  assign new_n26684_ = ~pi0331;
  assign new_n26685_ = ~new_n26795_ | ~new_n26733_;
  assign new_n26686_ = ~pi0334;
  assign new_n26687_ = ~pi0333;
  assign new_n26688_ = ~new_n26734_ | ~new_n26797_;
  assign new_n26689_ = ~pi0335;
  assign new_n26690_ = ~pi0336;
  assign new_n26691_ = ~new_n26735_ | ~new_n26798_;
  assign new_n26692_ = ~pi0337;
  assign new_n26693_ = ~pi0338;
  assign new_n26694_ = ~new_n26736_ | ~new_n26799_;
  assign new_n26695_ = ~pi0340;
  assign new_n26696_ = ~pi0339;
  assign new_n26697_ = ~new_n26737_ | ~new_n26801_;
  assign new_n26698_ = ~pi0342;
  assign new_n26699_ = ~pi0341;
  assign new_n26700_ = ~new_n26738_ | ~new_n26802_;
  assign new_n26701_ = ~pi0343;
  assign new_n26702_ = ~pi0343 | ~new_n26803_;
  assign new_n26703_ = ~pi0345;
  assign new_n26704_ = ~pi0344;
  assign new_n26705_ = ~new_n26739_ | ~new_n26804_;
  assign new_n26706_ = ~pi0346;
  assign new_n26707_ = ~pi0346 | ~new_n26805_;
  assign new_n26708_ = ~pi0347;
  assign new_n26709_ = ~new_n27034_ | ~new_n26753_;
  assign new_n26710_ = ~pi0330 | ~new_n26795_;
  assign new_n26711_ = ~new_n26871_ | ~new_n26870_;
  assign new_n26712_ = ~new_n26878_ | ~new_n26877_;
  assign new_n26713_ = ~new_n26880_ | ~new_n26879_;
  assign new_n26714_ = ~new_n26882_ | ~new_n26881_;
  assign new_n26715_ = ~new_n26889_ | ~new_n26888_;
  assign new_n26716_ = ~new_n26891_ | ~new_n26890_;
  assign new_n26717_ = ~new_n26893_ | ~new_n26892_;
  assign new_n26718_ = ~new_n26895_ | ~new_n26894_;
  assign new_n26719_ = ~new_n26897_ | ~new_n26896_;
  assign new_n26720_ = ~new_n26844_ | ~new_n26843_;
  assign new_n26721_ = ~new_n26851_ | ~new_n26850_;
  assign new_n26722_ = ~new_n26858_ | ~new_n26857_;
  assign new_n26723_ = ~new_n26865_ | ~new_n26864_;
  assign new_n26724_ = ~new_n26869_ | ~new_n26868_;
  assign new_n26725_ = ~new_n26876_ | ~new_n26875_;
  assign new_n26726_ = new_n26761_ & new_n26760_;
  assign new_n26727_ = new_n26769_ & new_n26768_;
  assign new_n26728_ = new_n26656_ & new_n26860_ & new_n26859_;
  assign new_n26729_ = new_n26786_ & new_n26636_;
  assign new_n26730_ = new_n26661_ & new_n26867_ & new_n26866_;
  assign new_n26731_ = pi0326 & pi0327;
  assign new_n26732_ = pi0329 & pi0328;
  assign new_n26733_ = pi0330 & pi0331 & pi0332;
  assign new_n26734_ = pi0334 & pi0333;
  assign new_n26735_ = pi0335 & pi0336;
  assign new_n26736_ = pi0337 & pi0338;
  assign new_n26737_ = pi0340 & pi0339;
  assign new_n26738_ = pi0342 & pi0341;
  assign new_n26739_ = pi0345 & pi0344;
  assign new_n26740_ = ~new_n26780_ | ~new_n26779_;
  assign new_n26741_ = new_n26837_ & new_n26836_;
  assign new_n26742_ = new_n26839_ & new_n26838_;
  assign new_n26743_ = ~new_n26832_ | ~new_n26776_ | ~new_n26750_;
  assign new_n26744_ = new_n26846_ & new_n26845_;
  assign new_n26745_ = ~new_n26774_ | ~new_n26773_;
  assign new_n26746_ = new_n26853_ & new_n26852_;
  assign new_n26747_ = ~new_n26727_ | ~new_n26770_;
  assign new_n26748_ = ~pi0348;
  assign new_n26749_ = ~new_n26680_;
  assign new_n26750_ = ~pi0324 | ~new_n26745_;
  assign new_n26751_ = ~new_n26834_ | ~new_n26833_;
  assign new_n26752_ = ~new_n26709_;
  assign new_n26753_ = ~new_n26666_;
  assign new_n26754_ = ~new_n26667_ | ~new_n26666_;
  assign new_n26755_ = ~pi0318 | ~new_n26754_;
  assign new_n26756_ = ~new_n26676_;
  assign new_n26757_ = pi0319 | new_n27018_;
  assign new_n26758_ = ~new_n26661_;
  assign new_n26759_ = ~new_n26662_ | ~new_n26661_;
  assign new_n26760_ = ~pi0320 | ~new_n26759_;
  assign new_n26761_ = ~new_n27038_ | ~new_n26758_;
  assign new_n26762_ = ~new_n26676_ | ~new_n26751_;
  assign new_n26763_ = ~new_n26675_;
  assign new_n26764_ = pi0322 | new_n27032_;
  assign new_n26765_ = pi0321 | new_n27033_;
  assign new_n26766_ = ~new_n26656_;
  assign new_n26767_ = ~new_n26657_ | ~new_n26656_;
  assign new_n26768_ = ~pi0322 | ~new_n26767_;
  assign new_n26769_ = ~new_n27032_ | ~new_n26766_;
  assign new_n26770_ = ~new_n26636_ | ~new_n26675_;
  assign new_n26771_ = ~new_n26747_;
  assign new_n26772_ = new_n27031_ | pi0323;
  assign new_n26773_ = ~new_n26772_ | ~new_n26747_;
  assign new_n26774_ = ~pi0323 | ~new_n27031_;
  assign new_n26775_ = ~new_n26745_;
  assign new_n26776_ = ~new_n27030_ | ~new_n26745_;
  assign new_n26777_ = ~new_n26743_;
  assign new_n26778_ = new_n27019_ | pi0325;
  assign new_n26779_ = ~new_n26778_ | ~new_n26743_;
  assign new_n26780_ = ~pi0325 | ~new_n27019_;
  assign new_n26781_ = ~new_n26740_;
  assign new_n26782_ = new_n27033_ | pi0321;
  assign new_n26783_ = ~new_n26782_ | ~new_n26675_;
  assign new_n26784_ = ~new_n26728_ | ~new_n26783_;
  assign new_n26785_ = ~new_n26763_ | ~new_n26656_;
  assign new_n26786_ = ~new_n27032_ | ~pi0322;
  assign new_n26787_ = ~new_n26729_ | ~new_n26785_;
  assign new_n26788_ = pi0321 | new_n27033_;
  assign new_n26789_ = new_n27018_ | pi0319;
  assign new_n26790_ = ~new_n26789_ | ~new_n26676_;
  assign new_n26791_ = ~new_n26730_ | ~new_n26790_;
  assign new_n26792_ = ~new_n26756_ | ~new_n26661_;
  assign new_n26793_ = ~new_n27038_ | ~pi0320;
  assign new_n26794_ = ~new_n26751_ | ~new_n26792_ | ~new_n26793_;
  assign new_n26795_ = ~new_n26681_;
  assign new_n26796_ = ~new_n26710_;
  assign new_n26797_ = ~new_n26685_;
  assign new_n26798_ = ~new_n26688_;
  assign new_n26799_ = ~new_n26691_;
  assign new_n26800_ = ~pi0337 | ~new_n26799_;
  assign new_n26801_ = ~new_n26694_;
  assign new_n26802_ = ~new_n26697_;
  assign new_n26803_ = ~new_n26700_;
  assign new_n26804_ = ~new_n26702_;
  assign new_n26805_ = ~new_n26705_;
  assign new_n26806_ = ~new_n26707_;
  assign new_n26807_ = pi0319 | new_n27018_;
  assign new_n26808_ = ~new_n26706_ | ~new_n26705_;
  assign new_n26809_ = ~pi0344 | ~new_n26804_;
  assign new_n26810_ = ~new_n26703_ | ~new_n26809_;
  assign new_n26811_ = ~new_n26701_ | ~new_n26700_;
  assign new_n26812_ = ~pi0341 | ~new_n26802_;
  assign new_n26813_ = ~new_n26698_ | ~new_n26812_;
  assign new_n26814_ = ~pi0339 | ~new_n26801_;
  assign new_n26815_ = ~new_n26695_ | ~new_n26814_;
  assign new_n26816_ = ~new_n26693_ | ~new_n26800_;
  assign new_n26817_ = ~new_n26692_ | ~new_n26691_;
  assign new_n26818_ = ~pi0335 | ~new_n26798_;
  assign new_n26819_ = ~new_n26690_ | ~new_n26818_;
  assign new_n26820_ = ~pi0333 | ~new_n26797_;
  assign new_n26821_ = ~new_n26686_ | ~new_n26820_;
  assign new_n26822_ = ~new_n26796_ | ~pi0331;
  assign new_n26823_ = ~new_n26683_ | ~new_n26822_;
  assign new_n26824_ = ~new_n26682_ | ~new_n26681_;
  assign new_n26825_ = ~new_n26749_ | ~pi0328;
  assign new_n26826_ = ~new_n26679_ | ~new_n26825_;
  assign new_n26827_ = ~pi0326 | ~new_n26740_;
  assign new_n26828_ = ~new_n26677_ | ~new_n26827_;
  assign new_n26829_ = ~new_n26788_ | ~new_n26656_;
  assign new_n26830_ = ~pi0347 | ~new_n26806_;
  assign new_n26831_ = ~new_n26807_ | ~new_n26661_;
  assign new_n26832_ = ~new_n27030_ | ~pi0324;
  assign new_n26833_ = ~pi0320 | ~new_n26757_;
  assign new_n26834_ = ~new_n27038_ | ~new_n26757_;
  assign new_n26835_ = ~new_n26752_ | ~pi0318;
  assign new_n26836_ = ~pi0326 | ~new_n26740_;
  assign new_n26837_ = ~new_n26781_ | ~new_n26674_;
  assign new_n26838_ = ~pi0325 | ~new_n26672_;
  assign new_n26839_ = ~new_n27019_ | ~new_n26673_;
  assign new_n26840_ = ~pi0325 | ~new_n26672_;
  assign new_n26841_ = ~new_n27019_ | ~new_n26673_;
  assign new_n26842_ = ~new_n26841_ | ~new_n26840_;
  assign new_n26843_ = ~new_n26742_ | ~new_n26743_;
  assign new_n26844_ = ~new_n26777_ | ~new_n26842_;
  assign new_n26845_ = ~pi0324 | ~new_n26671_;
  assign new_n26846_ = ~new_n27030_ | ~new_n26670_;
  assign new_n26847_ = ~pi0324 | ~new_n26671_;
  assign new_n26848_ = ~new_n27030_ | ~new_n26670_;
  assign new_n26849_ = ~new_n26848_ | ~new_n26847_;
  assign new_n26850_ = ~new_n26744_ | ~new_n26745_;
  assign new_n26851_ = ~new_n26775_ | ~new_n26849_;
  assign new_n26852_ = ~pi0323 | ~new_n26668_;
  assign new_n26853_ = ~new_n27031_ | ~new_n26669_;
  assign new_n26854_ = ~pi0323 | ~new_n26668_;
  assign new_n26855_ = ~new_n27031_ | ~new_n26669_;
  assign new_n26856_ = ~new_n26855_ | ~new_n26854_;
  assign new_n26857_ = ~new_n26746_ | ~new_n26747_;
  assign new_n26858_ = ~new_n26771_ | ~new_n26856_;
  assign new_n26859_ = ~pi0322 | ~new_n26657_;
  assign new_n26860_ = ~new_n27032_ | ~new_n26655_;
  assign new_n26861_ = ~pi0321 | ~new_n26653_;
  assign new_n26862_ = ~new_n27033_ | ~new_n26654_;
  assign new_n26863_ = ~new_n26862_ | ~new_n26861_;
  assign new_n26864_ = ~new_n26829_ | ~new_n26675_;
  assign new_n26865_ = ~new_n26863_ | ~new_n26763_;
  assign new_n26866_ = ~pi0320 | ~new_n26662_;
  assign new_n26867_ = ~new_n27038_ | ~new_n26660_;
  assign new_n26868_ = ~pi0348 | ~new_n26830_;
  assign new_n26869_ = ~new_n26748_ | ~pi0347 | ~new_n26806_;
  assign new_n26870_ = ~pi0347 | ~new_n26707_;
  assign new_n26871_ = ~new_n26806_ | ~new_n26708_;
  assign new_n26872_ = ~pi0319 | ~new_n26658_;
  assign new_n26873_ = ~new_n27018_ | ~new_n26659_;
  assign new_n26874_ = ~new_n26873_ | ~new_n26872_;
  assign new_n26875_ = ~new_n26831_ | ~new_n26676_;
  assign new_n26876_ = ~new_n26874_ | ~new_n26756_;
  assign new_n26877_ = ~pi0344 | ~new_n26702_;
  assign new_n26878_ = ~new_n26804_ | ~new_n26704_;
  assign new_n26879_ = ~pi0341 | ~new_n26697_;
  assign new_n26880_ = ~new_n26802_ | ~new_n26699_;
  assign new_n26881_ = ~pi0339 | ~new_n26694_;
  assign new_n26882_ = ~new_n26801_ | ~new_n26696_;
  assign new_n26883_ = ~pi0318 | ~new_n26666_;
  assign new_n26884_ = ~new_n26753_ | ~new_n26665_;
  assign new_n26885_ = ~new_n26884_ | ~new_n26883_;
  assign new_n26886_ = ~new_n27034_ | ~new_n26666_ | ~new_n26665_;
  assign new_n26887_ = ~new_n26885_ | ~new_n26667_;
  assign new_n26888_ = ~pi0335 | ~new_n26688_;
  assign new_n26889_ = ~new_n26798_ | ~new_n26689_;
  assign new_n26890_ = ~pi0333 | ~new_n26685_;
  assign new_n26891_ = ~new_n26797_ | ~new_n26687_;
  assign new_n26892_ = ~pi0331 | ~new_n26710_;
  assign new_n26893_ = ~new_n26796_ | ~new_n26684_;
  assign new_n26894_ = ~new_n26749_ | ~new_n26678_;
  assign new_n26895_ = ~pi0328 | ~new_n26680_;
  assign new_n26896_ = ~pi0317 | ~new_n26663_;
  assign new_n26897_ = ~new_n27017_ | ~new_n26664_;
  assign new_n26898_ = ~new_n26935_ | ~new_n26934_;
  assign new_n26899_ = ~pi0311 | ~new_n26919_;
  assign new_n26900_ = ~pi0315;
  assign new_n26901_ = ~pi0309;
  assign new_n26902_ = ~pi0314;
  assign new_n26903_ = ~pi0308;
  assign new_n26904_ = ~pi0313;
  assign new_n26905_ = ~pi0312;
  assign new_n26906_ = ~new_n26931_ | ~new_n26930_;
  assign new_n26907_ = ~pi0307;
  assign new_n26908_ = ~new_n26940_ | ~new_n26939_;
  assign new_n26909_ = ~new_n26945_ | ~new_n26944_;
  assign new_n26910_ = ~new_n26950_ | ~new_n26949_;
  assign new_n26911_ = ~new_n26955_ | ~new_n26954_;
  assign new_n26912_ = ~new_n26937_ | ~new_n26936_;
  assign new_n26913_ = ~new_n26942_ | ~new_n26941_;
  assign new_n26914_ = ~new_n26947_ | ~new_n26946_;
  assign new_n26915_ = ~new_n26952_ | ~new_n26951_;
  assign new_n26916_ = ~new_n26927_ | ~new_n26926_;
  assign new_n26917_ = ~new_n26923_ | ~new_n26922_;
  assign new_n26918_ = ~pi0310;
  assign new_n26919_ = ~pi0316;
  assign new_n26920_ = ~new_n26899_;
  assign new_n26921_ = ~new_n26920_ | ~new_n26900_;
  assign new_n26922_ = ~new_n26921_ | ~new_n26918_;
  assign new_n26923_ = ~pi0315 | ~new_n26899_;
  assign new_n26924_ = ~new_n26917_;
  assign new_n26925_ = ~pi0309 | ~new_n26902_;
  assign new_n26926_ = ~new_n26925_ | ~new_n26917_;
  assign new_n26927_ = ~pi0314 | ~new_n26901_;
  assign new_n26928_ = ~new_n26916_;
  assign new_n26929_ = ~pi0308 | ~new_n26904_;
  assign new_n26930_ = ~new_n26929_ | ~new_n26916_;
  assign new_n26931_ = ~pi0313 | ~new_n26903_;
  assign new_n26932_ = ~new_n26906_;
  assign new_n26933_ = ~pi0312 | ~new_n26907_;
  assign new_n26934_ = ~new_n26932_ | ~new_n26933_;
  assign new_n26935_ = ~pi0307 | ~new_n26905_;
  assign new_n26936_ = ~pi0307 | ~new_n26905_;
  assign new_n26937_ = ~pi0312 | ~new_n26907_;
  assign new_n26938_ = ~new_n26912_;
  assign new_n26939_ = ~new_n26938_ | ~new_n26932_;
  assign new_n26940_ = ~new_n26912_ | ~new_n26906_;
  assign new_n26941_ = ~pi0308 | ~new_n26904_;
  assign new_n26942_ = ~pi0313 | ~new_n26903_;
  assign new_n26943_ = ~new_n26913_;
  assign new_n26944_ = ~new_n26928_ | ~new_n26943_;
  assign new_n26945_ = ~new_n26913_ | ~new_n26916_;
  assign new_n26946_ = ~pi0309 | ~new_n26902_;
  assign new_n26947_ = ~pi0314 | ~new_n26901_;
  assign new_n26948_ = ~new_n26914_;
  assign new_n26949_ = ~new_n26924_ | ~new_n26948_;
  assign new_n26950_ = ~new_n26914_ | ~new_n26917_;
  assign new_n26951_ = ~pi0310 | ~new_n26900_;
  assign new_n26952_ = ~pi0315 | ~new_n26918_;
  assign new_n26953_ = ~new_n26915_;
  assign new_n26954_ = ~new_n26953_ | ~new_n26920_;
  assign new_n26955_ = ~new_n26915_ | ~new_n26899_;
  assign new_n26956_ = ~new_n26995_ | ~new_n26994_;
  assign new_n26957_ = ~new_n26959_ | ~new_n26996_;
  assign new_n26958_ = ~pi0311;
  assign new_n26959_ = ~pi0311 | ~new_n26968_;
  assign new_n26960_ = ~pi0315;
  assign new_n26961_ = ~pi0309;
  assign new_n26962_ = ~pi0314;
  assign new_n26963_ = ~pi0308;
  assign new_n26964_ = ~pi0313;
  assign new_n26965_ = ~pi0312;
  assign new_n26966_ = ~new_n26991_ | ~new_n26990_;
  assign new_n26967_ = ~pi0307;
  assign new_n26968_ = ~pi0316;
  assign new_n26969_ = ~new_n27001_ | ~new_n27000_;
  assign new_n26970_ = ~new_n27006_ | ~new_n27005_;
  assign new_n26971_ = ~new_n27011_ | ~new_n27010_;
  assign new_n26972_ = ~new_n27016_ | ~new_n27015_;
  assign new_n26973_ = ~new_n26998_ | ~new_n26997_;
  assign new_n26974_ = ~new_n27003_ | ~new_n27002_;
  assign new_n26975_ = ~new_n27008_ | ~new_n27007_;
  assign new_n26976_ = ~new_n27013_ | ~new_n27012_;
  assign new_n26977_ = ~new_n26987_ | ~new_n26986_;
  assign new_n26978_ = ~new_n26983_ | ~new_n26982_;
  assign new_n26979_ = ~pi0310;
  assign new_n26980_ = ~new_n26959_;
  assign new_n26981_ = ~new_n26980_ | ~new_n26960_;
  assign new_n26982_ = ~new_n26981_ | ~new_n26979_;
  assign new_n26983_ = ~pi0315 | ~new_n26959_;
  assign new_n26984_ = ~new_n26978_;
  assign new_n26985_ = ~pi0309 | ~new_n26962_;
  assign new_n26986_ = ~new_n26985_ | ~new_n26978_;
  assign new_n26987_ = ~pi0314 | ~new_n26961_;
  assign new_n26988_ = ~new_n26977_;
  assign new_n26989_ = ~pi0308 | ~new_n26964_;
  assign new_n26990_ = ~new_n26989_ | ~new_n26977_;
  assign new_n26991_ = ~pi0313 | ~new_n26963_;
  assign new_n26992_ = ~new_n26966_;
  assign new_n26993_ = ~pi0312 | ~new_n26967_;
  assign new_n26994_ = ~new_n26992_ | ~new_n26993_;
  assign new_n26995_ = ~pi0307 | ~new_n26965_;
  assign new_n26996_ = ~pi0316 | ~new_n26958_;
  assign new_n26997_ = ~pi0307 | ~new_n26965_;
  assign new_n26998_ = ~pi0312 | ~new_n26967_;
  assign new_n26999_ = ~new_n26973_;
  assign new_n27000_ = ~new_n26999_ | ~new_n26992_;
  assign new_n27001_ = ~new_n26973_ | ~new_n26966_;
  assign new_n27002_ = ~pi0308 | ~new_n26964_;
  assign new_n27003_ = ~pi0313 | ~new_n26963_;
  assign new_n27004_ = ~new_n26974_;
  assign new_n27005_ = ~new_n26988_ | ~new_n27004_;
  assign new_n27006_ = ~new_n26974_ | ~new_n26977_;
  assign new_n27007_ = ~pi0309 | ~new_n26962_;
  assign new_n27008_ = ~pi0314 | ~new_n26961_;
  assign new_n27009_ = ~new_n26975_;
  assign new_n27010_ = ~new_n26984_ | ~new_n27009_;
  assign new_n27011_ = ~new_n26975_ | ~new_n26978_;
  assign new_n27012_ = ~pi0310 | ~new_n26960_;
  assign new_n27013_ = ~pi0315 | ~new_n26979_;
  assign new_n27014_ = ~new_n26976_;
  assign new_n27015_ = ~new_n27014_ | ~new_n26980_;
  assign new_n27016_ = ~new_n26976_ | ~new_n26959_;
  assign new_n27017_ = ~new_n3777_;
  assign new_n27018_ = ~new_n27037_ | ~new_n27045_;
  assign new_n27019_ = new_n27035_ & new_n27043_;
  assign new_n27020_ = ~new_n3778_;
  assign new_n27021_ = ~new_n3780_;
  assign new_n27022_ = ~new_n3780_ | ~new_n27037_;
  assign new_n27023_ = ~new_n3781_;
  assign new_n27024_ = ~new_n3781_ | ~new_n27041_;
  assign new_n27025_ = ~new_n3782_;
  assign new_n27026_ = ~new_n3782_ | ~new_n27042_;
  assign new_n27027_ = ~new_n3784_;
  assign new_n27028_ = ~new_n3783_;
  assign new_n27029_ = ~new_n3779_;
  assign new_n27030_ = ~new_n27047_ | ~new_n27046_;
  assign new_n27031_ = ~new_n27049_ | ~new_n27048_;
  assign new_n27032_ = ~new_n27051_ | ~new_n27050_;
  assign new_n27033_ = ~new_n27053_ | ~new_n27052_;
  assign new_n27034_ = ~new_n27057_ | ~new_n27056_;
  assign new_n27035_ = new_n3784_ & new_n3783_;
  assign new_n27036_ = ~new_n3783_ | ~new_n27043_;
  assign new_n27037_ = ~new_n27029_ | ~new_n27039_;
  assign new_n27038_ = new_n27055_ & new_n27054_;
  assign new_n27039_ = ~new_n3778_ | ~new_n3777_;
  assign new_n27040_ = ~new_n27037_;
  assign new_n27041_ = ~new_n27022_;
  assign new_n27042_ = ~new_n27024_;
  assign new_n27043_ = ~new_n27026_;
  assign new_n27044_ = ~new_n27036_;
  assign new_n27045_ = ~new_n3779_ | ~new_n3778_ | ~new_n3777_;
  assign new_n27046_ = ~new_n3784_ | ~new_n27036_;
  assign new_n27047_ = ~new_n27044_ | ~new_n27027_;
  assign new_n27048_ = ~new_n3783_ | ~new_n27026_;
  assign new_n27049_ = ~new_n27043_ | ~new_n27028_;
  assign new_n27050_ = ~new_n3782_ | ~new_n27024_;
  assign new_n27051_ = ~new_n27042_ | ~new_n27025_;
  assign new_n27052_ = ~new_n3781_ | ~new_n27022_;
  assign new_n27053_ = ~new_n27041_ | ~new_n27023_;
  assign new_n27054_ = ~new_n3780_ | ~new_n27037_;
  assign new_n27055_ = ~new_n27040_ | ~new_n27021_;
  assign new_n27056_ = ~new_n3778_ | ~new_n27017_;
  assign new_n27057_ = ~new_n3777_ | ~new_n27020_;
  assign new_n27058_ = ~new_n27097_ | ~new_n27096_;
  assign new_n27059_ = ~new_n27061_ | ~new_n27098_;
  assign new_n27060_ = ~pi0311;
  assign new_n27061_ = ~pi0311 | ~new_n27070_;
  assign new_n27062_ = ~pi0315;
  assign new_n27063_ = ~pi0309;
  assign new_n27064_ = ~pi0314;
  assign new_n27065_ = ~pi0308;
  assign new_n27066_ = ~pi0313;
  assign new_n27067_ = ~pi0312;
  assign new_n27068_ = ~new_n27093_ | ~new_n27092_;
  assign new_n27069_ = ~pi0307;
  assign new_n27070_ = ~pi0316;
  assign new_n27071_ = ~new_n27103_ | ~new_n27102_;
  assign new_n27072_ = ~new_n27108_ | ~new_n27107_;
  assign new_n27073_ = ~new_n27113_ | ~new_n27112_;
  assign new_n27074_ = ~new_n27118_ | ~new_n27117_;
  assign new_n27075_ = ~new_n27100_ | ~new_n27099_;
  assign new_n27076_ = ~new_n27105_ | ~new_n27104_;
  assign new_n27077_ = ~new_n27110_ | ~new_n27109_;
  assign new_n27078_ = ~new_n27115_ | ~new_n27114_;
  assign new_n27079_ = ~new_n27089_ | ~new_n27088_;
  assign new_n27080_ = ~new_n27085_ | ~new_n27084_;
  assign new_n27081_ = ~pi0310;
  assign new_n27082_ = ~new_n27061_;
  assign new_n27083_ = ~new_n27082_ | ~new_n27062_;
  assign new_n27084_ = ~new_n27083_ | ~new_n27081_;
  assign new_n27085_ = ~pi0315 | ~new_n27061_;
  assign new_n27086_ = ~new_n27080_;
  assign new_n27087_ = ~pi0309 | ~new_n27064_;
  assign new_n27088_ = ~new_n27087_ | ~new_n27080_;
  assign new_n27089_ = ~pi0314 | ~new_n27063_;
  assign new_n27090_ = ~new_n27079_;
  assign new_n27091_ = ~pi0308 | ~new_n27066_;
  assign new_n27092_ = ~new_n27091_ | ~new_n27079_;
  assign new_n27093_ = ~pi0313 | ~new_n27065_;
  assign new_n27094_ = ~new_n27068_;
  assign new_n27095_ = ~pi0312 | ~new_n27069_;
  assign new_n27096_ = ~new_n27094_ | ~new_n27095_;
  assign new_n27097_ = ~pi0307 | ~new_n27067_;
  assign new_n27098_ = ~pi0316 | ~new_n27060_;
  assign new_n27099_ = ~pi0307 | ~new_n27067_;
  assign new_n27100_ = ~pi0312 | ~new_n27069_;
  assign new_n27101_ = ~new_n27075_;
  assign new_n27102_ = ~new_n27101_ | ~new_n27094_;
  assign new_n27103_ = ~new_n27075_ | ~new_n27068_;
  assign new_n27104_ = ~pi0308 | ~new_n27066_;
  assign new_n27105_ = ~pi0313 | ~new_n27065_;
  assign new_n27106_ = ~new_n27076_;
  assign new_n27107_ = ~new_n27090_ | ~new_n27106_;
  assign new_n27108_ = ~new_n27076_ | ~new_n27079_;
  assign new_n27109_ = ~pi0309 | ~new_n27064_;
  assign new_n27110_ = ~pi0314 | ~new_n27063_;
  assign new_n27111_ = ~new_n27077_;
  assign new_n27112_ = ~new_n27086_ | ~new_n27111_;
  assign new_n27113_ = ~new_n27077_ | ~new_n27080_;
  assign new_n27114_ = ~pi0310 | ~new_n27062_;
  assign new_n27115_ = ~pi0315 | ~new_n27081_;
  assign new_n27116_ = ~new_n27078_;
  assign new_n27117_ = ~new_n27116_ | ~new_n27082_;
  assign new_n27118_ = ~new_n27078_ | ~new_n27061_;
  assign new_n27119_ = ~new_n3783_;
  assign new_n27120_ = ~new_n3778_;
  assign new_n27121_ = ~new_n3784_;
  assign new_n27122_ = ~new_n3782_;
  assign new_n27123_ = ~new_n3777_;
  assign new_n27124_ = ~new_n3780_;
  assign new_n27125_ = ~new_n3779_;
  assign new_n27126_ = ~new_n3781_;
  assign new_n27127_ = ~pi0310;
  assign new_n27128_ = ~pi0309;
  assign new_n27129_ = ~pi0309 | ~pi0310;
  assign new_n27130_ = ~pi0308;
  assign new_n27131_ = ~new_n27139_ | ~new_n27138_;
  assign new_n27132_ = ~new_n27141_ | ~new_n27140_;
  assign new_n27133_ = ~new_n27143_ | ~new_n27142_;
  assign new_n27134_ = ~pi0307;
  assign new_n27135_ = ~pi0308 | ~new_n27136_;
  assign new_n27136_ = ~new_n27129_;
  assign new_n27137_ = ~new_n27135_;
  assign new_n27138_ = ~pi0307 | ~new_n27135_;
  assign new_n27139_ = ~new_n27137_ | ~new_n27134_;
  assign new_n27140_ = ~pi0308 | ~new_n27129_;
  assign new_n27141_ = ~new_n27136_ | ~new_n27130_;
  assign new_n27142_ = ~pi0309 | ~new_n27127_;
  assign new_n27143_ = ~pi0310 | ~new_n27128_;
  assign new_n27144_ = ~new_n26578_ & ~new_n27145_;
  assign new_n27145_ = ~new_n26589_ & ~new_n26588_ & ~new_n26590_ & ~new_n26591_;
  assign new_n27146_ = ~new_n26898_ & ~new_n27147_;
  assign new_n27147_ = ~new_n26909_ & ~new_n26908_ & ~new_n26910_ & ~new_n26911_;
  assign new_n27148_ = ~pi0318;
  assign new_n27149_ = ~pi0319;
  assign new_n27150_ = ~pi0319 | ~pi0318;
  assign new_n27151_ = ~pi0320;
  assign new_n27152_ = ~pi0320 | ~new_n27238_;
  assign new_n27153_ = ~pi0321;
  assign new_n27154_ = ~pi0321 | ~new_n27239_;
  assign new_n27155_ = ~pi0322;
  assign new_n27156_ = ~pi0322 | ~new_n27240_;
  assign new_n27157_ = ~pi0323;
  assign new_n27158_ = ~pi0323 | ~new_n27241_;
  assign new_n27159_ = ~pi0324;
  assign new_n27160_ = ~pi0324 | ~new_n27242_;
  assign new_n27161_ = ~pi0325;
  assign new_n27162_ = ~pi0326;
  assign new_n27163_ = ~pi0325 | ~new_n27243_;
  assign new_n27164_ = ~new_n27244_ | ~pi0326;
  assign new_n27165_ = ~pi0327;
  assign new_n27166_ = ~pi0327 | ~new_n27245_;
  assign new_n27167_ = ~pi0328;
  assign new_n27168_ = ~pi0328 | ~new_n27246_;
  assign new_n27169_ = ~pi0329;
  assign new_n27170_ = ~pi0329 | ~new_n27247_;
  assign new_n27171_ = ~pi0330;
  assign new_n27172_ = ~pi0330 | ~new_n27248_;
  assign new_n27173_ = ~pi0331;
  assign new_n27174_ = ~pi0331 | ~new_n27249_;
  assign new_n27175_ = ~pi0332;
  assign new_n27176_ = ~pi0332 | ~new_n27250_;
  assign new_n27177_ = ~pi0333;
  assign new_n27178_ = ~pi0333 | ~new_n27251_;
  assign new_n27179_ = ~pi0334;
  assign new_n27180_ = ~pi0334 | ~new_n27252_;
  assign new_n27181_ = ~pi0335;
  assign new_n27182_ = ~pi0335 | ~new_n27253_;
  assign new_n27183_ = ~pi0336;
  assign new_n27184_ = ~pi0336 | ~new_n27254_;
  assign new_n27185_ = ~pi0337;
  assign new_n27186_ = ~pi0337 | ~new_n27255_;
  assign new_n27187_ = ~pi0338;
  assign new_n27188_ = ~pi0338 | ~new_n27256_;
  assign new_n27189_ = ~pi0339;
  assign new_n27190_ = ~pi0339 | ~new_n27257_;
  assign new_n27191_ = ~pi0340;
  assign new_n27192_ = ~pi0340 | ~new_n27258_;
  assign new_n27193_ = ~pi0341;
  assign new_n27194_ = ~pi0341 | ~new_n27259_;
  assign new_n27195_ = ~pi0342;
  assign new_n27196_ = ~pi0342 | ~new_n27260_;
  assign new_n27197_ = ~pi0343;
  assign new_n27198_ = ~pi0343 | ~new_n27261_;
  assign new_n27199_ = ~pi0344;
  assign new_n27200_ = ~pi0344 | ~new_n27262_;
  assign new_n27201_ = ~pi0345;
  assign new_n27202_ = ~pi0345 | ~new_n27263_;
  assign new_n27203_ = ~pi0346;
  assign new_n27204_ = ~pi0346 | ~new_n27264_;
  assign new_n27205_ = ~pi0347;
  assign new_n27206_ = ~new_n27268_ | ~new_n27267_;
  assign new_n27207_ = ~new_n27270_ | ~new_n27269_;
  assign new_n27208_ = ~new_n27272_ | ~new_n27271_;
  assign new_n27209_ = ~new_n27274_ | ~new_n27273_;
  assign new_n27210_ = ~new_n27276_ | ~new_n27275_;
  assign new_n27211_ = ~new_n27278_ | ~new_n27277_;
  assign new_n27212_ = ~new_n27280_ | ~new_n27279_;
  assign new_n27213_ = ~new_n27282_ | ~new_n27281_;
  assign new_n27214_ = ~new_n27284_ | ~new_n27283_;
  assign new_n27215_ = ~new_n27286_ | ~new_n27285_;
  assign new_n27216_ = ~new_n27288_ | ~new_n27287_;
  assign new_n27217_ = ~new_n27290_ | ~new_n27289_;
  assign new_n27218_ = ~new_n27292_ | ~new_n27291_;
  assign new_n27219_ = ~new_n27294_ | ~new_n27293_;
  assign new_n27220_ = ~new_n27296_ | ~new_n27295_;
  assign new_n27221_ = ~new_n27298_ | ~new_n27297_;
  assign new_n27222_ = ~new_n27300_ | ~new_n27299_;
  assign new_n27223_ = ~new_n27302_ | ~new_n27301_;
  assign new_n27224_ = ~new_n27304_ | ~new_n27303_;
  assign new_n27225_ = ~new_n27306_ | ~new_n27305_;
  assign new_n27226_ = ~new_n27308_ | ~new_n27307_;
  assign new_n27227_ = ~new_n27310_ | ~new_n27309_;
  assign new_n27228_ = ~new_n27312_ | ~new_n27311_;
  assign new_n27229_ = ~new_n27314_ | ~new_n27313_;
  assign new_n27230_ = ~new_n27316_ | ~new_n27315_;
  assign new_n27231_ = ~new_n27318_ | ~new_n27317_;
  assign new_n27232_ = ~new_n27320_ | ~new_n27319_;
  assign new_n27233_ = ~new_n27322_ | ~new_n27321_;
  assign new_n27234_ = ~new_n27324_ | ~new_n27323_;
  assign new_n27235_ = ~new_n27326_ | ~new_n27325_;
  assign new_n27236_ = ~pi0348;
  assign new_n27237_ = ~pi0347 | ~new_n27265_;
  assign new_n27238_ = ~new_n27150_;
  assign new_n27239_ = ~new_n27152_;
  assign new_n27240_ = ~new_n27154_;
  assign new_n27241_ = ~new_n27156_;
  assign new_n27242_ = ~new_n27158_;
  assign new_n27243_ = ~new_n27160_;
  assign new_n27244_ = ~new_n27163_;
  assign new_n27245_ = ~new_n27164_;
  assign new_n27246_ = ~new_n27166_;
  assign new_n27247_ = ~new_n27168_;
  assign new_n27248_ = ~new_n27170_;
  assign new_n27249_ = ~new_n27172_;
  assign new_n27250_ = ~new_n27174_;
  assign new_n27251_ = ~new_n27176_;
  assign new_n27252_ = ~new_n27178_;
  assign new_n27253_ = ~new_n27180_;
  assign new_n27254_ = ~new_n27182_;
  assign new_n27255_ = ~new_n27184_;
  assign new_n27256_ = ~new_n27186_;
  assign new_n27257_ = ~new_n27188_;
  assign new_n27258_ = ~new_n27190_;
  assign new_n27259_ = ~new_n27192_;
  assign new_n27260_ = ~new_n27194_;
  assign new_n27261_ = ~new_n27196_;
  assign new_n27262_ = ~new_n27198_;
  assign new_n27263_ = ~new_n27200_;
  assign new_n27264_ = ~new_n27202_;
  assign new_n27265_ = ~new_n27204_;
  assign new_n27266_ = ~new_n27237_;
  assign new_n27267_ = ~pi0326 | ~new_n27163_;
  assign new_n27268_ = ~new_n27244_ | ~new_n27162_;
  assign new_n27269_ = ~pi0325 | ~new_n27160_;
  assign new_n27270_ = ~new_n27243_ | ~new_n27161_;
  assign new_n27271_ = ~pi0324 | ~new_n27158_;
  assign new_n27272_ = ~new_n27242_ | ~new_n27159_;
  assign new_n27273_ = ~pi0323 | ~new_n27156_;
  assign new_n27274_ = ~new_n27241_ | ~new_n27157_;
  assign new_n27275_ = ~pi0322 | ~new_n27154_;
  assign new_n27276_ = ~new_n27240_ | ~new_n27155_;
  assign new_n27277_ = ~pi0321 | ~new_n27152_;
  assign new_n27278_ = ~new_n27239_ | ~new_n27153_;
  assign new_n27279_ = ~pi0320 | ~new_n27150_;
  assign new_n27280_ = ~new_n27238_ | ~new_n27151_;
  assign new_n27281_ = ~pi0348 | ~new_n27237_;
  assign new_n27282_ = ~new_n27266_ | ~new_n27236_;
  assign new_n27283_ = ~pi0347 | ~new_n27204_;
  assign new_n27284_ = ~new_n27265_ | ~new_n27205_;
  assign new_n27285_ = ~pi0319 | ~new_n27148_;
  assign new_n27286_ = ~pi0318 | ~new_n27149_;
  assign new_n27287_ = ~pi0346 | ~new_n27202_;
  assign new_n27288_ = ~new_n27264_ | ~new_n27203_;
  assign new_n27289_ = ~pi0345 | ~new_n27200_;
  assign new_n27290_ = ~new_n27263_ | ~new_n27201_;
  assign new_n27291_ = ~pi0344 | ~new_n27198_;
  assign new_n27292_ = ~new_n27262_ | ~new_n27199_;
  assign new_n27293_ = ~pi0343 | ~new_n27196_;
  assign new_n27294_ = ~new_n27261_ | ~new_n27197_;
  assign new_n27295_ = ~pi0342 | ~new_n27194_;
  assign new_n27296_ = ~new_n27260_ | ~new_n27195_;
  assign new_n27297_ = ~pi0341 | ~new_n27192_;
  assign new_n27298_ = ~new_n27259_ | ~new_n27193_;
  assign new_n27299_ = ~pi0340 | ~new_n27190_;
  assign new_n27300_ = ~new_n27258_ | ~new_n27191_;
  assign new_n27301_ = ~pi0339 | ~new_n27188_;
  assign new_n27302_ = ~new_n27257_ | ~new_n27189_;
  assign new_n27303_ = ~pi0338 | ~new_n27186_;
  assign new_n27304_ = ~new_n27256_ | ~new_n27187_;
  assign new_n27305_ = ~pi0337 | ~new_n27184_;
  assign new_n27306_ = ~new_n27255_ | ~new_n27185_;
  assign new_n27307_ = ~pi0336 | ~new_n27182_;
  assign new_n27308_ = ~new_n27254_ | ~new_n27183_;
  assign new_n27309_ = ~pi0335 | ~new_n27180_;
  assign new_n27310_ = ~new_n27253_ | ~new_n27181_;
  assign new_n27311_ = ~pi0334 | ~new_n27178_;
  assign new_n27312_ = ~new_n27252_ | ~new_n27179_;
  assign new_n27313_ = ~pi0333 | ~new_n27176_;
  assign new_n27314_ = ~new_n27251_ | ~new_n27177_;
  assign new_n27315_ = ~pi0332 | ~new_n27174_;
  assign new_n27316_ = ~new_n27250_ | ~new_n27175_;
  assign new_n27317_ = ~pi0331 | ~new_n27172_;
  assign new_n27318_ = ~new_n27249_ | ~new_n27173_;
  assign new_n27319_ = ~pi0330 | ~new_n27170_;
  assign new_n27320_ = ~new_n27248_ | ~new_n27171_;
  assign new_n27321_ = ~pi0329 | ~new_n27168_;
  assign new_n27322_ = ~new_n27247_ | ~new_n27169_;
  assign new_n27323_ = ~pi0328 | ~new_n27166_;
  assign new_n27324_ = ~new_n27246_ | ~new_n27167_;
  assign new_n27325_ = ~pi0327 | ~new_n27164_;
  assign new_n27326_ = ~new_n27245_ | ~new_n27165_;
  assign new_n27327_ = ~pi0318;
  assign new_n27328_ = ~pi0319;
  assign new_n27329_ = ~pi0319 | ~pi0318;
  assign new_n27330_ = ~pi0320;
  assign new_n27331_ = ~pi0320 | ~new_n27417_;
  assign new_n27332_ = ~pi0321;
  assign new_n27333_ = ~pi0321 | ~new_n27418_;
  assign new_n27334_ = ~pi0322;
  assign new_n27335_ = ~pi0322 | ~new_n27419_;
  assign new_n27336_ = ~pi0323;
  assign new_n27337_ = ~pi0323 | ~new_n27420_;
  assign new_n27338_ = ~pi0324;
  assign new_n27339_ = ~pi0324 | ~new_n27421_;
  assign new_n27340_ = ~pi0325;
  assign new_n27341_ = ~pi0326;
  assign new_n27342_ = ~pi0325 | ~new_n27422_;
  assign new_n27343_ = ~new_n27423_ | ~pi0326;
  assign new_n27344_ = ~pi0327;
  assign new_n27345_ = ~pi0327 | ~new_n27424_;
  assign new_n27346_ = ~pi0328;
  assign new_n27347_ = ~pi0328 | ~new_n27425_;
  assign new_n27348_ = ~pi0329;
  assign new_n27349_ = ~pi0329 | ~new_n27426_;
  assign new_n27350_ = ~pi0330;
  assign new_n27351_ = ~pi0330 | ~new_n27427_;
  assign new_n27352_ = ~pi0331;
  assign new_n27353_ = ~pi0331 | ~new_n27428_;
  assign new_n27354_ = ~pi0332;
  assign new_n27355_ = ~pi0332 | ~new_n27429_;
  assign new_n27356_ = ~pi0333;
  assign new_n27357_ = ~pi0333 | ~new_n27430_;
  assign new_n27358_ = ~pi0334;
  assign new_n27359_ = ~pi0334 | ~new_n27431_;
  assign new_n27360_ = ~pi0335;
  assign new_n27361_ = ~pi0335 | ~new_n27432_;
  assign new_n27362_ = ~pi0336;
  assign new_n27363_ = ~pi0336 | ~new_n27433_;
  assign new_n27364_ = ~pi0337;
  assign new_n27365_ = ~pi0337 | ~new_n27434_;
  assign new_n27366_ = ~pi0338;
  assign new_n27367_ = ~pi0338 | ~new_n27435_;
  assign new_n27368_ = ~pi0339;
  assign new_n27369_ = ~pi0339 | ~new_n27436_;
  assign new_n27370_ = ~pi0340;
  assign new_n27371_ = ~pi0340 | ~new_n27437_;
  assign new_n27372_ = ~pi0341;
  assign new_n27373_ = ~pi0341 | ~new_n27438_;
  assign new_n27374_ = ~pi0342;
  assign new_n27375_ = ~pi0342 | ~new_n27439_;
  assign new_n27376_ = ~pi0343;
  assign new_n27377_ = ~pi0343 | ~new_n27440_;
  assign new_n27378_ = ~pi0344;
  assign new_n27379_ = ~pi0344 | ~new_n27441_;
  assign new_n27380_ = ~pi0345;
  assign new_n27381_ = ~pi0345 | ~new_n27442_;
  assign new_n27382_ = ~pi0346;
  assign new_n27383_ = ~pi0346 | ~new_n27443_;
  assign new_n27384_ = ~pi0347;
  assign new_n27385_ = ~new_n27447_ | ~new_n27446_;
  assign new_n27386_ = ~new_n27449_ | ~new_n27448_;
  assign new_n27387_ = ~new_n27451_ | ~new_n27450_;
  assign new_n27388_ = ~new_n27453_ | ~new_n27452_;
  assign new_n27389_ = ~new_n27455_ | ~new_n27454_;
  assign new_n27390_ = ~new_n27457_ | ~new_n27456_;
  assign new_n27391_ = ~new_n27459_ | ~new_n27458_;
  assign new_n27392_ = ~new_n27461_ | ~new_n27460_;
  assign new_n27393_ = ~new_n27463_ | ~new_n27462_;
  assign new_n27394_ = ~new_n27465_ | ~new_n27464_;
  assign new_n27395_ = ~new_n27467_ | ~new_n27466_;
  assign new_n27396_ = ~new_n27469_ | ~new_n27468_;
  assign new_n27397_ = ~new_n27471_ | ~new_n27470_;
  assign new_n27398_ = ~new_n27473_ | ~new_n27472_;
  assign new_n27399_ = ~new_n27475_ | ~new_n27474_;
  assign new_n27400_ = ~new_n27477_ | ~new_n27476_;
  assign new_n27401_ = ~new_n27479_ | ~new_n27478_;
  assign new_n27402_ = ~new_n27481_ | ~new_n27480_;
  assign new_n27403_ = ~new_n27483_ | ~new_n27482_;
  assign new_n27404_ = ~new_n27485_ | ~new_n27484_;
  assign new_n27405_ = ~new_n27487_ | ~new_n27486_;
  assign new_n27406_ = ~new_n27489_ | ~new_n27488_;
  assign new_n27407_ = ~new_n27491_ | ~new_n27490_;
  assign new_n27408_ = ~new_n27493_ | ~new_n27492_;
  assign new_n27409_ = ~new_n27495_ | ~new_n27494_;
  assign new_n27410_ = ~new_n27497_ | ~new_n27496_;
  assign new_n27411_ = ~new_n27499_ | ~new_n27498_;
  assign new_n27412_ = ~new_n27501_ | ~new_n27500_;
  assign new_n27413_ = ~new_n27503_ | ~new_n27502_;
  assign new_n27414_ = ~new_n27505_ | ~new_n27504_;
  assign new_n27415_ = ~pi0348;
  assign new_n27416_ = ~pi0347 | ~new_n27444_;
  assign new_n27417_ = ~new_n27329_;
  assign new_n27418_ = ~new_n27331_;
  assign new_n27419_ = ~new_n27333_;
  assign new_n27420_ = ~new_n27335_;
  assign new_n27421_ = ~new_n27337_;
  assign new_n27422_ = ~new_n27339_;
  assign new_n27423_ = ~new_n27342_;
  assign new_n27424_ = ~new_n27343_;
  assign new_n27425_ = ~new_n27345_;
  assign new_n27426_ = ~new_n27347_;
  assign new_n27427_ = ~new_n27349_;
  assign new_n27428_ = ~new_n27351_;
  assign new_n27429_ = ~new_n27353_;
  assign new_n27430_ = ~new_n27355_;
  assign new_n27431_ = ~new_n27357_;
  assign new_n27432_ = ~new_n27359_;
  assign new_n27433_ = ~new_n27361_;
  assign new_n27434_ = ~new_n27363_;
  assign new_n27435_ = ~new_n27365_;
  assign new_n27436_ = ~new_n27367_;
  assign new_n27437_ = ~new_n27369_;
  assign new_n27438_ = ~new_n27371_;
  assign new_n27439_ = ~new_n27373_;
  assign new_n27440_ = ~new_n27375_;
  assign new_n27441_ = ~new_n27377_;
  assign new_n27442_ = ~new_n27379_;
  assign new_n27443_ = ~new_n27381_;
  assign new_n27444_ = ~new_n27383_;
  assign new_n27445_ = ~new_n27416_;
  assign new_n27446_ = ~pi0326 | ~new_n27342_;
  assign new_n27447_ = ~new_n27423_ | ~new_n27341_;
  assign new_n27448_ = ~pi0325 | ~new_n27339_;
  assign new_n27449_ = ~new_n27422_ | ~new_n27340_;
  assign new_n27450_ = ~pi0324 | ~new_n27337_;
  assign new_n27451_ = ~new_n27421_ | ~new_n27338_;
  assign new_n27452_ = ~pi0323 | ~new_n27335_;
  assign new_n27453_ = ~new_n27420_ | ~new_n27336_;
  assign new_n27454_ = ~pi0322 | ~new_n27333_;
  assign new_n27455_ = ~new_n27419_ | ~new_n27334_;
  assign new_n27456_ = ~pi0321 | ~new_n27331_;
  assign new_n27457_ = ~new_n27418_ | ~new_n27332_;
  assign new_n27458_ = ~pi0320 | ~new_n27329_;
  assign new_n27459_ = ~new_n27417_ | ~new_n27330_;
  assign new_n27460_ = ~pi0348 | ~new_n27416_;
  assign new_n27461_ = ~new_n27445_ | ~new_n27415_;
  assign new_n27462_ = ~pi0347 | ~new_n27383_;
  assign new_n27463_ = ~new_n27444_ | ~new_n27384_;
  assign new_n27464_ = ~pi0319 | ~new_n27327_;
  assign new_n27465_ = ~pi0318 | ~new_n27328_;
  assign new_n27466_ = ~pi0346 | ~new_n27381_;
  assign new_n27467_ = ~new_n27443_ | ~new_n27382_;
  assign new_n27468_ = ~pi0345 | ~new_n27379_;
  assign new_n27469_ = ~new_n27442_ | ~new_n27380_;
  assign new_n27470_ = ~pi0344 | ~new_n27377_;
  assign new_n27471_ = ~new_n27441_ | ~new_n27378_;
  assign new_n27472_ = ~pi0343 | ~new_n27375_;
  assign new_n27473_ = ~new_n27440_ | ~new_n27376_;
  assign new_n27474_ = ~pi0342 | ~new_n27373_;
  assign new_n27475_ = ~new_n27439_ | ~new_n27374_;
  assign new_n27476_ = ~pi0341 | ~new_n27371_;
  assign new_n27477_ = ~new_n27438_ | ~new_n27372_;
  assign new_n27478_ = ~pi0340 | ~new_n27369_;
  assign new_n27479_ = ~new_n27437_ | ~new_n27370_;
  assign new_n27480_ = ~pi0339 | ~new_n27367_;
  assign new_n27481_ = ~new_n27436_ | ~new_n27368_;
  assign new_n27482_ = ~pi0338 | ~new_n27365_;
  assign new_n27483_ = ~new_n27435_ | ~new_n27366_;
  assign new_n27484_ = ~pi0337 | ~new_n27363_;
  assign new_n27485_ = ~new_n27434_ | ~new_n27364_;
  assign new_n27486_ = ~pi0336 | ~new_n27361_;
  assign new_n27487_ = ~new_n27433_ | ~new_n27362_;
  assign new_n27488_ = ~pi0335 | ~new_n27359_;
  assign new_n27489_ = ~new_n27432_ | ~new_n27360_;
  assign new_n27490_ = ~pi0334 | ~new_n27357_;
  assign new_n27491_ = ~new_n27431_ | ~new_n27358_;
  assign new_n27492_ = ~pi0333 | ~new_n27355_;
  assign new_n27493_ = ~new_n27430_ | ~new_n27356_;
  assign new_n27494_ = ~pi0332 | ~new_n27353_;
  assign new_n27495_ = ~new_n27429_ | ~new_n27354_;
  assign new_n27496_ = ~pi0331 | ~new_n27351_;
  assign new_n27497_ = ~new_n27428_ | ~new_n27352_;
  assign new_n27498_ = ~pi0330 | ~new_n27349_;
  assign new_n27499_ = ~new_n27427_ | ~new_n27350_;
  assign new_n27500_ = ~pi0329 | ~new_n27347_;
  assign new_n27501_ = ~new_n27426_ | ~new_n27348_;
  assign new_n27502_ = ~pi0328 | ~new_n27345_;
  assign new_n27503_ = ~new_n27425_ | ~new_n27346_;
  assign new_n27504_ = ~pi0327 | ~new_n27343_;
  assign new_n27505_ = ~new_n27424_ | ~new_n27344_;
  assign new_n27506_ = ~new_n3769_;
  assign new_n27507_ = ~new_n4225_;
  assign new_n27508_ = ~new_n4225_ | ~new_n3769_;
  assign new_n27509_ = ~new_n3770_;
  assign new_n27510_ = ~new_n3770_ | ~new_n27530_;
  assign new_n27511_ = ~new_n3771_;
  assign new_n27512_ = ~new_n3771_ | ~new_n27531_;
  assign new_n27513_ = ~new_n3772_;
  assign new_n27514_ = ~new_n3772_ | ~new_n27532_;
  assign new_n27515_ = ~new_n3773_;
  assign new_n27516_ = ~new_n3773_ | ~new_n27533_;
  assign new_n27517_ = ~new_n3774_;
  assign new_n27518_ = ~new_n3774_ | ~new_n27534_;
  assign new_n27519_ = ~new_n3775_;
  assign new_n27520_ = ~new_n27538_ | ~new_n27537_;
  assign new_n27521_ = ~new_n27540_ | ~new_n27539_;
  assign new_n27522_ = ~new_n27542_ | ~new_n27541_;
  assign new_n27523_ = ~new_n27544_ | ~new_n27543_;
  assign new_n27524_ = ~new_n27546_ | ~new_n27545_;
  assign new_n27525_ = ~new_n27548_ | ~new_n27547_;
  assign new_n27526_ = ~new_n27550_ | ~new_n27549_;
  assign new_n27527_ = ~new_n27552_ | ~new_n27551_;
  assign new_n27528_ = ~new_n3776_;
  assign new_n27529_ = ~new_n3775_ | ~new_n27535_;
  assign new_n27530_ = ~new_n27508_;
  assign new_n27531_ = ~new_n27510_;
  assign new_n27532_ = ~new_n27512_;
  assign new_n27533_ = ~new_n27514_;
  assign new_n27534_ = ~new_n27516_;
  assign new_n27535_ = ~new_n27518_;
  assign new_n27536_ = ~new_n27529_;
  assign new_n27537_ = ~new_n3776_ | ~new_n27529_;
  assign new_n27538_ = ~new_n27536_ | ~new_n27528_;
  assign new_n27539_ = ~new_n3775_ | ~new_n27518_;
  assign new_n27540_ = ~new_n27535_ | ~new_n27519_;
  assign new_n27541_ = ~new_n3774_ | ~new_n27516_;
  assign new_n27542_ = ~new_n27534_ | ~new_n27517_;
  assign new_n27543_ = ~new_n3773_ | ~new_n27514_;
  assign new_n27544_ = ~new_n27533_ | ~new_n27515_;
  assign new_n27545_ = ~new_n3772_ | ~new_n27512_;
  assign new_n27546_ = ~new_n27532_ | ~new_n27513_;
  assign new_n27547_ = ~new_n3771_ | ~new_n27510_;
  assign new_n27548_ = ~new_n27531_ | ~new_n27511_;
  assign new_n27549_ = ~new_n3770_ | ~new_n27508_;
  assign new_n27550_ = ~new_n27530_ | ~new_n27509_;
  assign new_n27551_ = ~new_n4225_ | ~new_n27506_;
  assign new_n27552_ = ~new_n3769_ | ~new_n27507_;
  assign new_n27553_ = ~new_n27655_ | ~new_n27696_;
  assign new_n27554_ = ~new_n9788_;
  assign new_n27555_ = ~new_n9792_;
  assign new_n27556_ = ~new_n9791_;
  assign new_n27557_ = ~new_n9787_;
  assign new_n27558_ = ~new_n9790_;
  assign new_n27559_ = ~new_n9786_;
  assign new_n27560_ = ~new_n9789_;
  assign new_n27561_ = ~new_n9785_;
  assign new_n27562_ = ~new_n9784_;
  assign new_n27563_ = ~new_n9784_ | ~new_n27645_;
  assign new_n27564_ = ~new_n9783_;
  assign new_n27565_ = ~new_n9783_ | ~new_n27668_;
  assign new_n27566_ = ~new_n9782_;
  assign new_n27567_ = ~new_n9782_ | ~new_n27669_;
  assign new_n27568_ = ~new_n9781_;
  assign new_n27569_ = ~new_n9781_ | ~new_n27670_;
  assign new_n27570_ = ~new_n9780_;
  assign new_n27571_ = ~new_n9779_;
  assign new_n27572_ = ~new_n9780_ | ~new_n27671_;
  assign new_n27573_ = ~new_n27672_ | ~new_n9779_;
  assign new_n27574_ = ~new_n9778_;
  assign new_n27575_ = ~new_n9778_ | ~new_n27673_;
  assign new_n27576_ = ~new_n9777_;
  assign new_n27577_ = ~new_n9777_ | ~new_n27674_;
  assign new_n27578_ = ~new_n9776_;
  assign new_n27579_ = ~new_n9776_ | ~new_n27675_;
  assign new_n27580_ = ~new_n9775_;
  assign new_n27581_ = ~new_n9775_ | ~new_n27676_;
  assign new_n27582_ = ~new_n9774_;
  assign new_n27583_ = ~new_n9774_ | ~new_n27677_;
  assign new_n27584_ = ~new_n9773_;
  assign new_n27585_ = ~new_n9773_ | ~new_n27678_;
  assign new_n27586_ = ~new_n9772_;
  assign new_n27587_ = ~new_n9772_ | ~new_n27679_;
  assign new_n27588_ = ~new_n9771_;
  assign new_n27589_ = ~new_n9771_ | ~new_n27680_;
  assign new_n27590_ = ~new_n9770_;
  assign new_n27591_ = ~new_n9770_ | ~new_n27681_;
  assign new_n27592_ = ~new_n9769_;
  assign new_n27593_ = ~new_n9769_ | ~new_n27682_;
  assign new_n27594_ = ~new_n9768_;
  assign new_n27595_ = ~new_n9768_ | ~new_n27683_;
  assign new_n27596_ = ~new_n9767_;
  assign new_n27597_ = ~new_n9767_ | ~new_n27684_;
  assign new_n27598_ = ~new_n9766_;
  assign new_n27599_ = ~new_n9766_ | ~new_n27685_;
  assign new_n27600_ = ~new_n9765_;
  assign new_n27601_ = ~new_n9765_ | ~new_n27686_;
  assign new_n27602_ = ~new_n9764_;
  assign new_n27603_ = ~new_n9764_ | ~new_n27687_;
  assign new_n27604_ = ~new_n9763_;
  assign new_n27605_ = ~new_n9763_ | ~new_n27688_;
  assign new_n27606_ = ~new_n9762_;
  assign new_n27607_ = ~new_n9762_ | ~new_n27689_;
  assign new_n27608_ = ~new_n9761_;
  assign new_n27609_ = ~new_n9761_ | ~new_n27690_;
  assign new_n27610_ = ~new_n9760_;
  assign new_n27611_ = ~new_n9760_ | ~new_n27691_;
  assign new_n27612_ = ~new_n9759_;
  assign new_n27613_ = ~new_n9759_ | ~new_n27692_;
  assign new_n27614_ = ~new_n9758_;
  assign new_n27615_ = ~new_n27698_ | ~new_n27697_;
  assign new_n27616_ = ~new_n27700_ | ~new_n27699_;
  assign new_n27617_ = ~new_n27702_ | ~new_n27701_;
  assign new_n27618_ = ~new_n27704_ | ~new_n27703_;
  assign new_n27619_ = ~new_n27706_ | ~new_n27705_;
  assign new_n27620_ = ~new_n27717_ | ~new_n27716_;
  assign new_n27621_ = ~new_n27719_ | ~new_n27718_;
  assign new_n27622_ = ~new_n27728_ | ~new_n27727_;
  assign new_n27623_ = ~new_n27730_ | ~new_n27729_;
  assign new_n27624_ = ~new_n27732_ | ~new_n27731_;
  assign new_n27625_ = ~new_n27734_ | ~new_n27733_;
  assign new_n27626_ = ~new_n27736_ | ~new_n27735_;
  assign new_n27627_ = ~new_n27738_ | ~new_n27737_;
  assign new_n27628_ = ~new_n27740_ | ~new_n27739_;
  assign new_n27629_ = ~new_n27742_ | ~new_n27741_;
  assign new_n27630_ = ~new_n27744_ | ~new_n27743_;
  assign new_n27631_ = ~new_n27746_ | ~new_n27745_;
  assign new_n27632_ = ~new_n27753_ | ~new_n27752_;
  assign new_n27633_ = ~new_n27755_ | ~new_n27754_;
  assign new_n27634_ = ~new_n27757_ | ~new_n27756_;
  assign new_n27635_ = ~new_n27759_ | ~new_n27758_;
  assign new_n27636_ = ~new_n27761_ | ~new_n27760_;
  assign new_n27637_ = ~new_n27763_ | ~new_n27762_;
  assign new_n27638_ = ~new_n27765_ | ~new_n27764_;
  assign new_n27639_ = ~new_n27767_ | ~new_n27766_;
  assign new_n27640_ = ~new_n27769_ | ~new_n27768_;
  assign new_n27641_ = ~new_n27771_ | ~new_n27770_;
  assign new_n27642_ = ~new_n27773_ | ~new_n27772_;
  assign new_n27643_ = ~new_n27715_ | ~new_n27714_;
  assign new_n27644_ = ~new_n27726_ | ~new_n27725_;
  assign new_n27645_ = ~new_n27666_ | ~new_n27665_;
  assign new_n27646_ = new_n27708_ & new_n27707_;
  assign new_n27647_ = new_n27710_ & new_n27709_;
  assign new_n27648_ = ~new_n27662_ | ~new_n27661_;
  assign new_n27649_ = ~new_n9757_;
  assign new_n27650_ = ~new_n9758_ | ~new_n27693_;
  assign new_n27651_ = new_n27721_ & new_n27720_;
  assign new_n27652_ = ~new_n27654_ | ~new_n27658_;
  assign new_n27653_ = ~new_n9792_ | ~new_n9788_;
  assign new_n27654_ = ~new_n9792_ | ~new_n9787_ | ~new_n9788_;
  assign new_n27655_ = new_n27751_ & new_n27750_;
  assign new_n27656_ = ~new_n27654_;
  assign new_n27657_ = ~new_n27557_ | ~new_n27653_;
  assign new_n27658_ = ~new_n9791_ | ~new_n27657_;
  assign new_n27659_ = ~new_n27652_;
  assign new_n27660_ = new_n9790_ | new_n9786_;
  assign new_n27661_ = ~new_n27660_ | ~new_n27652_;
  assign new_n27662_ = ~new_n9786_ | ~new_n9790_;
  assign new_n27663_ = ~new_n27648_;
  assign new_n27664_ = new_n9789_ | new_n9785_;
  assign new_n27665_ = ~new_n27664_ | ~new_n27648_;
  assign new_n27666_ = ~new_n9785_ | ~new_n9789_;
  assign new_n27667_ = ~new_n27645_;
  assign new_n27668_ = ~new_n27563_;
  assign new_n27669_ = ~new_n27565_;
  assign new_n27670_ = ~new_n27567_;
  assign new_n27671_ = ~new_n27569_;
  assign new_n27672_ = ~new_n27572_;
  assign new_n27673_ = ~new_n27573_;
  assign new_n27674_ = ~new_n27575_;
  assign new_n27675_ = ~new_n27577_;
  assign new_n27676_ = ~new_n27579_;
  assign new_n27677_ = ~new_n27581_;
  assign new_n27678_ = ~new_n27583_;
  assign new_n27679_ = ~new_n27585_;
  assign new_n27680_ = ~new_n27587_;
  assign new_n27681_ = ~new_n27589_;
  assign new_n27682_ = ~new_n27591_;
  assign new_n27683_ = ~new_n27593_;
  assign new_n27684_ = ~new_n27595_;
  assign new_n27685_ = ~new_n27597_;
  assign new_n27686_ = ~new_n27599_;
  assign new_n27687_ = ~new_n27601_;
  assign new_n27688_ = ~new_n27603_;
  assign new_n27689_ = ~new_n27605_;
  assign new_n27690_ = ~new_n27607_;
  assign new_n27691_ = ~new_n27609_;
  assign new_n27692_ = ~new_n27611_;
  assign new_n27693_ = ~new_n27613_;
  assign new_n27694_ = ~new_n27650_;
  assign new_n27695_ = ~new_n27653_;
  assign new_n27696_ = ~new_n27749_ | ~new_n27557_;
  assign new_n27697_ = ~new_n9779_ | ~new_n27572_;
  assign new_n27698_ = ~new_n27672_ | ~new_n27571_;
  assign new_n27699_ = ~new_n9780_ | ~new_n27569_;
  assign new_n27700_ = ~new_n27671_ | ~new_n27570_;
  assign new_n27701_ = ~new_n9781_ | ~new_n27567_;
  assign new_n27702_ = ~new_n27670_ | ~new_n27568_;
  assign new_n27703_ = ~new_n9782_ | ~new_n27565_;
  assign new_n27704_ = ~new_n27669_ | ~new_n27566_;
  assign new_n27705_ = ~new_n9783_ | ~new_n27563_;
  assign new_n27706_ = ~new_n27668_ | ~new_n27564_;
  assign new_n27707_ = ~new_n9784_ | ~new_n27645_;
  assign new_n27708_ = ~new_n27667_ | ~new_n27562_;
  assign new_n27709_ = ~new_n9785_ | ~new_n27560_;
  assign new_n27710_ = ~new_n9789_ | ~new_n27561_;
  assign new_n27711_ = ~new_n9785_ | ~new_n27560_;
  assign new_n27712_ = ~new_n9789_ | ~new_n27561_;
  assign new_n27713_ = ~new_n27712_ | ~new_n27711_;
  assign new_n27714_ = ~new_n27647_ | ~new_n27648_;
  assign new_n27715_ = ~new_n27663_ | ~new_n27713_;
  assign new_n27716_ = ~new_n9757_ | ~new_n27650_;
  assign new_n27717_ = ~new_n27694_ | ~new_n27649_;
  assign new_n27718_ = ~new_n9758_ | ~new_n27613_;
  assign new_n27719_ = ~new_n27693_ | ~new_n27614_;
  assign new_n27720_ = ~new_n9786_ | ~new_n27558_;
  assign new_n27721_ = ~new_n9790_ | ~new_n27559_;
  assign new_n27722_ = ~new_n9786_ | ~new_n27558_;
  assign new_n27723_ = ~new_n9790_ | ~new_n27559_;
  assign new_n27724_ = ~new_n27723_ | ~new_n27722_;
  assign new_n27725_ = ~new_n27651_ | ~new_n27652_;
  assign new_n27726_ = ~new_n27659_ | ~new_n27724_;
  assign new_n27727_ = ~new_n9759_ | ~new_n27611_;
  assign new_n27728_ = ~new_n27692_ | ~new_n27612_;
  assign new_n27729_ = ~new_n9760_ | ~new_n27609_;
  assign new_n27730_ = ~new_n27691_ | ~new_n27610_;
  assign new_n27731_ = ~new_n9761_ | ~new_n27607_;
  assign new_n27732_ = ~new_n27690_ | ~new_n27608_;
  assign new_n27733_ = ~new_n9762_ | ~new_n27605_;
  assign new_n27734_ = ~new_n27689_ | ~new_n27606_;
  assign new_n27735_ = ~new_n9763_ | ~new_n27603_;
  assign new_n27736_ = ~new_n27688_ | ~new_n27604_;
  assign new_n27737_ = ~new_n9764_ | ~new_n27601_;
  assign new_n27738_ = ~new_n27687_ | ~new_n27602_;
  assign new_n27739_ = ~new_n9765_ | ~new_n27599_;
  assign new_n27740_ = ~new_n27686_ | ~new_n27600_;
  assign new_n27741_ = ~new_n9766_ | ~new_n27597_;
  assign new_n27742_ = ~new_n27685_ | ~new_n27598_;
  assign new_n27743_ = ~new_n9767_ | ~new_n27595_;
  assign new_n27744_ = ~new_n27684_ | ~new_n27596_;
  assign new_n27745_ = ~new_n9768_ | ~new_n27593_;
  assign new_n27746_ = ~new_n27683_ | ~new_n27594_;
  assign new_n27747_ = ~new_n9791_ | ~new_n27653_;
  assign new_n27748_ = ~new_n27695_ | ~new_n27556_;
  assign new_n27749_ = ~new_n27748_ | ~new_n27747_;
  assign new_n27750_ = ~new_n27556_ | ~new_n9787_ | ~new_n27653_;
  assign new_n27751_ = ~new_n27656_ | ~new_n9791_;
  assign new_n27752_ = ~new_n9769_ | ~new_n27591_;
  assign new_n27753_ = ~new_n27682_ | ~new_n27592_;
  assign new_n27754_ = ~new_n9770_ | ~new_n27589_;
  assign new_n27755_ = ~new_n27681_ | ~new_n27590_;
  assign new_n27756_ = ~new_n9771_ | ~new_n27587_;
  assign new_n27757_ = ~new_n27680_ | ~new_n27588_;
  assign new_n27758_ = ~new_n9772_ | ~new_n27585_;
  assign new_n27759_ = ~new_n27679_ | ~new_n27586_;
  assign new_n27760_ = ~new_n9773_ | ~new_n27583_;
  assign new_n27761_ = ~new_n27678_ | ~new_n27584_;
  assign new_n27762_ = ~new_n9774_ | ~new_n27581_;
  assign new_n27763_ = ~new_n27677_ | ~new_n27582_;
  assign new_n27764_ = ~new_n9775_ | ~new_n27579_;
  assign new_n27765_ = ~new_n27676_ | ~new_n27580_;
  assign new_n27766_ = ~new_n9776_ | ~new_n27577_;
  assign new_n27767_ = ~new_n27675_ | ~new_n27578_;
  assign new_n27768_ = ~new_n9777_ | ~new_n27575_;
  assign new_n27769_ = ~new_n27674_ | ~new_n27576_;
  assign new_n27770_ = ~new_n9778_ | ~new_n27573_;
  assign new_n27771_ = ~new_n27673_ | ~new_n27574_;
  assign new_n27772_ = ~new_n9792_ | ~new_n27554_;
  assign new_n27773_ = ~new_n9788_ | ~new_n27555_;
  assign new_n27774_ = new_n28070_ & new_n28068_;
  assign new_n27775_ = new_n28065_ & new_n28063_;
  assign new_n27776_ = new_n28061_ & new_n28059_;
  assign new_n27777_ = new_n28056_ & new_n28052_;
  assign new_n27778_ = new_n27974_ & new_n27972_;
  assign new_n27779_ = new_n27970_ & new_n27968_;
  assign new_n27780_ = new_n27965_ & new_n27961_;
  assign new_n27781_ = ~new_n27913_ | ~new_n28075_;
  assign new_n27782_ = ~new_n28365_;
  assign new_n27783_ = ~new_n29207_;
  assign new_n27784_ = ~new_n28366_;
  assign new_n27785_ = ~new_n29208_;
  assign new_n27786_ = ~new_n28367_;
  assign new_n27787_ = ~new_n29209_;
  assign new_n27788_ = ~new_n29204_;
  assign new_n27789_ = ~new_n28362_;
  assign new_n27790_ = ~new_n28361_;
  assign new_n27791_ = ~new_n28362_ | ~new_n29204_;
  assign new_n27792_ = ~new_n29187_;
  assign new_n27793_ = ~new_n28333_;
  assign new_n27794_ = ~new_n29213_;
  assign new_n27795_ = ~new_n28369_;
  assign new_n27796_ = ~new_n29211_;
  assign new_n27797_ = ~new_n28368_;
  assign new_n27798_ = ~new_n29210_;
  assign new_n27799_ = ~new_n27808_ | ~new_n27949_;
  assign new_n27800_ = ~new_n28364_;
  assign new_n27801_ = ~new_n29206_;
  assign new_n27802_ = ~new_n29205_;
  assign new_n27803_ = ~new_n28363_;
  assign new_n27804_ = ~new_n27959_ | ~new_n27958_;
  assign new_n27805_ = ~new_n27804_ | ~new_n27962_;
  assign new_n27806_ = ~new_n27952_ | ~new_n27953_ | ~new_n27951_;
  assign new_n27807_ = ~new_n27945_ | ~new_n27944_;
  assign new_n27808_ = ~new_n27807_ | ~new_n27947_;
  assign new_n27809_ = ~new_n28384_;
  assign new_n27810_ = ~new_n29228_;
  assign new_n27811_ = ~new_n28385_;
  assign new_n27812_ = ~new_n29229_;
  assign new_n27813_ = ~new_n28386_;
  assign new_n27814_ = ~new_n29230_;
  assign new_n27815_ = ~new_n28388_;
  assign new_n27816_ = ~new_n29232_;
  assign new_n27817_ = ~new_n28389_;
  assign new_n27818_ = ~new_n29233_;
  assign new_n27819_ = ~new_n27805_ | ~new_n27975_;
  assign new_n27820_ = ~new_n28387_;
  assign new_n27821_ = ~new_n29231_;
  assign new_n27822_ = ~new_n27854_ | ~new_n27989_;
  assign new_n27823_ = ~new_n28383_;
  assign new_n27824_ = ~new_n29227_;
  assign new_n27825_ = ~new_n28382_;
  assign new_n27826_ = ~new_n29226_;
  assign new_n27827_ = ~new_n28381_;
  assign new_n27828_ = ~new_n29225_;
  assign new_n27829_ = ~new_n28380_;
  assign new_n27830_ = ~new_n29224_;
  assign new_n27831_ = ~new_n28379_;
  assign new_n27832_ = ~new_n29223_;
  assign new_n27833_ = ~new_n28378_;
  assign new_n27834_ = ~new_n29222_;
  assign new_n27835_ = ~new_n28377_;
  assign new_n27836_ = ~new_n29221_;
  assign new_n27837_ = ~new_n28376_;
  assign new_n27838_ = ~new_n29220_;
  assign new_n27839_ = ~new_n28375_;
  assign new_n27840_ = ~new_n29219_;
  assign new_n27841_ = ~new_n28374_;
  assign new_n27842_ = ~new_n29218_;
  assign new_n27843_ = ~new_n28373_;
  assign new_n27844_ = ~new_n29217_;
  assign new_n27845_ = ~new_n28372_;
  assign new_n27846_ = ~new_n29216_;
  assign new_n27847_ = ~new_n29215_;
  assign new_n27848_ = ~new_n28371_;
  assign new_n27849_ = ~new_n29214_;
  assign new_n27850_ = ~new_n28370_;
  assign new_n27851_ = ~new_n28047_ | ~new_n28046_;
  assign new_n27852_ = ~new_n27992_ | ~new_n27993_ | ~new_n27991_;
  assign new_n27853_ = ~new_n27985_ | ~new_n27984_;
  assign new_n27854_ = ~new_n27853_ | ~new_n27987_;
  assign new_n27855_ = ~new_n27978_ | ~new_n27979_ | ~new_n27977_;
  assign new_n27856_ = ~new_n28247_ | ~new_n28246_;
  assign new_n27857_ = ~new_n28084_ | ~new_n28083_;
  assign new_n27858_ = ~new_n28091_ | ~new_n28090_;
  assign new_n27859_ = ~new_n28100_ | ~new_n28099_;
  assign new_n27860_ = ~new_n28107_ | ~new_n28106_;
  assign new_n27861_ = ~new_n28119_ | ~new_n28118_;
  assign new_n27862_ = ~new_n28126_ | ~new_n28125_;
  assign new_n27863_ = ~new_n28133_ | ~new_n28132_;
  assign new_n27864_ = ~new_n28140_ | ~new_n28139_;
  assign new_n27865_ = ~new_n28147_ | ~new_n28146_;
  assign new_n27866_ = ~new_n28154_ | ~new_n28153_;
  assign new_n27867_ = ~new_n28161_ | ~new_n28160_;
  assign new_n27868_ = ~new_n28168_ | ~new_n28167_;
  assign new_n27869_ = ~new_n28175_ | ~new_n28174_;
  assign new_n27870_ = ~new_n28182_ | ~new_n28181_;
  assign new_n27871_ = ~new_n28189_ | ~new_n28188_;
  assign new_n27872_ = ~new_n28201_ | ~new_n28200_;
  assign new_n27873_ = ~new_n28208_ | ~new_n28207_;
  assign new_n27874_ = ~new_n28215_ | ~new_n28214_;
  assign new_n27875_ = ~new_n28222_ | ~new_n28221_;
  assign new_n27876_ = ~new_n28229_ | ~new_n28228_;
  assign new_n27877_ = ~new_n28238_ | ~new_n28237_;
  assign new_n27878_ = ~new_n28245_ | ~new_n28244_;
  assign new_n27879_ = new_n28077_ & new_n28076_;
  assign new_n27880_ = new_n28079_ & new_n28078_;
  assign new_n27881_ = ~new_n27806_ | ~new_n27955_;
  assign new_n27882_ = new_n28086_ & new_n28085_;
  assign new_n27883_ = new_n28093_ & new_n28092_;
  assign new_n27884_ = new_n28095_ & new_n28094_;
  assign new_n27885_ = ~new_n27941_ | ~new_n27940_;
  assign new_n27886_ = new_n28102_ & new_n28101_;
  assign new_n27887_ = ~new_n27937_ | ~new_n27936_;
  assign new_n27888_ = ~new_n28334_;
  assign new_n27889_ = ~new_n29212_;
  assign new_n27890_ = new_n28109_ & new_n28108_;
  assign new_n27891_ = new_n28114_ & new_n28113_;
  assign new_n27892_ = ~new_n27912_ | ~new_n27933_;
  assign new_n27893_ = new_n28121_ & new_n28120_;
  assign new_n27894_ = new_n28128_ & new_n28127_;
  assign new_n27895_ = ~new_n28043_ | ~new_n28042_;
  assign new_n27896_ = new_n28135_ & new_n28134_;
  assign new_n27897_ = ~new_n28039_ | ~new_n28038_;
  assign new_n27898_ = new_n28142_ & new_n28141_;
  assign new_n27899_ = ~new_n28035_ | ~new_n28034_;
  assign new_n27900_ = new_n28149_ & new_n28148_;
  assign new_n27901_ = ~new_n28031_ | ~new_n28030_;
  assign new_n27902_ = new_n28156_ & new_n28155_;
  assign new_n27903_ = ~new_n28027_ | ~new_n28026_;
  assign new_n27904_ = new_n28163_ & new_n28162_;
  assign new_n27905_ = ~new_n28023_ | ~new_n28022_;
  assign new_n27906_ = new_n28170_ & new_n28169_;
  assign new_n27907_ = ~new_n28019_ | ~new_n28018_;
  assign new_n27908_ = new_n28177_ & new_n28176_;
  assign new_n27909_ = ~new_n28015_ | ~new_n28014_;
  assign new_n27910_ = new_n28184_ & new_n28183_;
  assign new_n27911_ = ~new_n28011_ | ~new_n28010_;
  assign new_n27912_ = ~new_n29187_ | ~new_n27931_;
  assign new_n27913_ = new_n28194_ & new_n28193_;
  assign new_n27914_ = new_n28196_ & new_n28195_;
  assign new_n27915_ = ~new_n28007_ | ~new_n28006_;
  assign new_n27916_ = new_n28203_ & new_n28202_;
  assign new_n27917_ = ~new_n28003_ | ~new_n28002_;
  assign new_n27918_ = new_n28210_ & new_n28209_;
  assign new_n27919_ = ~new_n27999_ | ~new_n27998_;
  assign new_n27920_ = new_n28217_ & new_n28216_;
  assign new_n27921_ = ~new_n27852_ | ~new_n27995_;
  assign new_n27922_ = new_n28224_ & new_n28223_;
  assign new_n27923_ = new_n28231_ & new_n28230_;
  assign new_n27924_ = new_n28233_ & new_n28232_;
  assign new_n27925_ = ~new_n27855_ | ~new_n27981_;
  assign new_n27926_ = new_n28240_ & new_n28239_;
  assign new_n27927_ = ~new_n29233_ | ~new_n28389_;
  assign new_n27928_ = ~new_n29229_ | ~new_n28385_;
  assign new_n27929_ = ~new_n27912_;
  assign new_n27930_ = ~new_n29208_ | ~new_n28366_;
  assign new_n27931_ = ~new_n27791_;
  assign new_n27932_ = ~new_n27792_ | ~new_n27791_;
  assign new_n27933_ = ~new_n28361_ | ~new_n27932_;
  assign new_n27934_ = ~new_n27892_;
  assign new_n27935_ = new_n28333_ | new_n29213_;
  assign new_n27936_ = ~new_n27935_ | ~new_n27892_;
  assign new_n27937_ = ~new_n29213_ | ~new_n28333_;
  assign new_n27938_ = ~new_n27887_;
  assign new_n27939_ = new_n28369_ | new_n29211_;
  assign new_n27940_ = ~new_n27939_ | ~new_n27887_;
  assign new_n27941_ = ~new_n29211_ | ~new_n28369_;
  assign new_n27942_ = ~new_n27885_;
  assign new_n27943_ = new_n28368_ | new_n29210_;
  assign new_n27944_ = ~new_n27943_ | ~new_n27885_;
  assign new_n27945_ = ~new_n29210_ | ~new_n28368_;
  assign new_n27946_ = ~new_n27807_;
  assign new_n27947_ = new_n29209_ | new_n28367_;
  assign new_n27948_ = ~new_n27808_;
  assign new_n27949_ = ~new_n29209_ | ~new_n28367_;
  assign new_n27950_ = ~new_n27799_;
  assign new_n27951_ = ~new_n27950_ | ~new_n27930_;
  assign new_n27952_ = new_n29207_ | new_n28365_;
  assign new_n27953_ = new_n29208_ | new_n28366_;
  assign new_n27954_ = ~new_n27806_;
  assign new_n27955_ = ~new_n29207_ | ~new_n28365_;
  assign new_n27956_ = ~new_n27881_;
  assign new_n27957_ = new_n28364_ | new_n29206_;
  assign new_n27958_ = ~new_n27957_ | ~new_n27881_;
  assign new_n27959_ = ~new_n29206_ | ~new_n28364_;
  assign new_n27960_ = ~new_n27804_;
  assign new_n27961_ = ~new_n27879_ | ~new_n27960_;
  assign new_n27962_ = new_n29205_ | new_n28363_;
  assign new_n27963_ = ~new_n27805_;
  assign new_n27964_ = ~new_n28363_ | ~new_n29205_;
  assign new_n27965_ = ~new_n27963_ | ~new_n27964_;
  assign new_n27966_ = new_n28366_ | new_n29208_;
  assign new_n27967_ = ~new_n27966_ | ~new_n27799_;
  assign new_n27968_ = ~new_n27882_ | ~new_n27967_ | ~new_n27930_;
  assign new_n27969_ = ~new_n29207_ | ~new_n28365_;
  assign new_n27970_ = ~new_n27954_ | ~new_n27969_;
  assign new_n27971_ = new_n29208_ | new_n28366_;
  assign new_n27972_ = ~new_n27883_ | ~new_n27946_;
  assign new_n27973_ = ~new_n29209_ | ~new_n28367_;
  assign new_n27974_ = ~new_n27948_ | ~new_n27973_;
  assign new_n27975_ = ~new_n28363_ | ~new_n29205_;
  assign new_n27976_ = ~new_n27819_;
  assign new_n27977_ = ~new_n27976_ | ~new_n27927_;
  assign new_n27978_ = new_n29232_ | new_n28388_;
  assign new_n27979_ = new_n29233_ | new_n28389_;
  assign new_n27980_ = ~new_n27855_;
  assign new_n27981_ = ~new_n29232_ | ~new_n28388_;
  assign new_n27982_ = ~new_n27925_;
  assign new_n27983_ = new_n28387_ | new_n29231_;
  assign new_n27984_ = ~new_n27983_ | ~new_n27925_;
  assign new_n27985_ = ~new_n29231_ | ~new_n28387_;
  assign new_n27986_ = ~new_n27853_;
  assign new_n27987_ = new_n29230_ | new_n28386_;
  assign new_n27988_ = ~new_n27854_;
  assign new_n27989_ = ~new_n29230_ | ~new_n28386_;
  assign new_n27990_ = ~new_n27822_;
  assign new_n27991_ = ~new_n27990_ | ~new_n27928_;
  assign new_n27992_ = new_n29228_ | new_n28384_;
  assign new_n27993_ = new_n29229_ | new_n28385_;
  assign new_n27994_ = ~new_n27852_;
  assign new_n27995_ = ~new_n29228_ | ~new_n28384_;
  assign new_n27996_ = ~new_n27921_;
  assign new_n27997_ = new_n28383_ | new_n29227_;
  assign new_n27998_ = ~new_n27997_ | ~new_n27921_;
  assign new_n27999_ = ~new_n29227_ | ~new_n28383_;
  assign new_n28000_ = ~new_n27919_;
  assign new_n28001_ = new_n28382_ | new_n29226_;
  assign new_n28002_ = ~new_n28001_ | ~new_n27919_;
  assign new_n28003_ = ~new_n29226_ | ~new_n28382_;
  assign new_n28004_ = ~new_n27917_;
  assign new_n28005_ = new_n28381_ | new_n29225_;
  assign new_n28006_ = ~new_n28005_ | ~new_n27917_;
  assign new_n28007_ = ~new_n29225_ | ~new_n28381_;
  assign new_n28008_ = ~new_n27915_;
  assign new_n28009_ = new_n28380_ | new_n29224_;
  assign new_n28010_ = ~new_n28009_ | ~new_n27915_;
  assign new_n28011_ = ~new_n29224_ | ~new_n28380_;
  assign new_n28012_ = ~new_n27911_;
  assign new_n28013_ = new_n28379_ | new_n29223_;
  assign new_n28014_ = ~new_n28013_ | ~new_n27911_;
  assign new_n28015_ = ~new_n29223_ | ~new_n28379_;
  assign new_n28016_ = ~new_n27909_;
  assign new_n28017_ = new_n28378_ | new_n29222_;
  assign new_n28018_ = ~new_n28017_ | ~new_n27909_;
  assign new_n28019_ = ~new_n29222_ | ~new_n28378_;
  assign new_n28020_ = ~new_n27907_;
  assign new_n28021_ = new_n28377_ | new_n29221_;
  assign new_n28022_ = ~new_n28021_ | ~new_n27907_;
  assign new_n28023_ = ~new_n29221_ | ~new_n28377_;
  assign new_n28024_ = ~new_n27905_;
  assign new_n28025_ = new_n28376_ | new_n29220_;
  assign new_n28026_ = ~new_n28025_ | ~new_n27905_;
  assign new_n28027_ = ~new_n29220_ | ~new_n28376_;
  assign new_n28028_ = ~new_n27903_;
  assign new_n28029_ = new_n28375_ | new_n29219_;
  assign new_n28030_ = ~new_n28029_ | ~new_n27903_;
  assign new_n28031_ = ~new_n29219_ | ~new_n28375_;
  assign new_n28032_ = ~new_n27901_;
  assign new_n28033_ = new_n28374_ | new_n29218_;
  assign new_n28034_ = ~new_n28033_ | ~new_n27901_;
  assign new_n28035_ = ~new_n29218_ | ~new_n28374_;
  assign new_n28036_ = ~new_n27899_;
  assign new_n28037_ = new_n28373_ | new_n29217_;
  assign new_n28038_ = ~new_n28037_ | ~new_n27899_;
  assign new_n28039_ = ~new_n29217_ | ~new_n28373_;
  assign new_n28040_ = ~new_n27897_;
  assign new_n28041_ = new_n28372_ | new_n29216_;
  assign new_n28042_ = ~new_n28041_ | ~new_n27897_;
  assign new_n28043_ = ~new_n29216_ | ~new_n28372_;
  assign new_n28044_ = ~new_n27895_;
  assign new_n28045_ = new_n29215_ | new_n28371_;
  assign new_n28046_ = ~new_n28045_ | ~new_n27895_;
  assign new_n28047_ = ~new_n28371_ | ~new_n29215_;
  assign new_n28048_ = ~new_n27851_;
  assign new_n28049_ = new_n29214_ | new_n28370_;
  assign new_n28050_ = ~new_n28049_ | ~new_n27851_;
  assign new_n28051_ = ~new_n28370_ | ~new_n29214_;
  assign new_n28052_ = ~new_n27890_ | ~new_n28051_ | ~new_n28050_;
  assign new_n28053_ = ~new_n28370_ | ~new_n29214_;
  assign new_n28054_ = ~new_n28048_ | ~new_n28053_;
  assign new_n28055_ = new_n28370_ | new_n29214_;
  assign new_n28056_ = ~new_n28112_ | ~new_n28055_ | ~new_n28054_;
  assign new_n28057_ = new_n28385_ | new_n29229_;
  assign new_n28058_ = ~new_n28057_ | ~new_n27822_;
  assign new_n28059_ = ~new_n27922_ | ~new_n28058_ | ~new_n27928_;
  assign new_n28060_ = ~new_n29228_ | ~new_n28384_;
  assign new_n28061_ = ~new_n27994_ | ~new_n28060_;
  assign new_n28062_ = new_n29229_ | new_n28385_;
  assign new_n28063_ = ~new_n27923_ | ~new_n27986_;
  assign new_n28064_ = ~new_n29230_ | ~new_n28386_;
  assign new_n28065_ = ~new_n27988_ | ~new_n28064_;
  assign new_n28066_ = new_n28389_ | new_n29233_;
  assign new_n28067_ = ~new_n28066_ | ~new_n27819_;
  assign new_n28068_ = ~new_n27926_ | ~new_n28067_ | ~new_n27927_;
  assign new_n28069_ = ~new_n29232_ | ~new_n28388_;
  assign new_n28070_ = ~new_n27980_ | ~new_n28069_;
  assign new_n28071_ = new_n29233_ | new_n28389_;
  assign new_n28072_ = ~new_n27971_ | ~new_n27930_;
  assign new_n28073_ = ~new_n28062_ | ~new_n27928_;
  assign new_n28074_ = ~new_n28071_ | ~new_n27927_;
  assign new_n28075_ = ~new_n28192_ | ~new_n27792_;
  assign new_n28076_ = ~new_n29205_ | ~new_n27803_;
  assign new_n28077_ = ~new_n28363_ | ~new_n27802_;
  assign new_n28078_ = ~new_n29206_ | ~new_n27800_;
  assign new_n28079_ = ~new_n28364_ | ~new_n27801_;
  assign new_n28080_ = ~new_n29206_ | ~new_n27800_;
  assign new_n28081_ = ~new_n28364_ | ~new_n27801_;
  assign new_n28082_ = ~new_n28081_ | ~new_n28080_;
  assign new_n28083_ = ~new_n27880_ | ~new_n27881_;
  assign new_n28084_ = ~new_n27956_ | ~new_n28082_;
  assign new_n28085_ = ~new_n29207_ | ~new_n27782_;
  assign new_n28086_ = ~new_n28365_ | ~new_n27783_;
  assign new_n28087_ = ~new_n29208_ | ~new_n27784_;
  assign new_n28088_ = ~new_n28366_ | ~new_n27785_;
  assign new_n28089_ = ~new_n28088_ | ~new_n28087_;
  assign new_n28090_ = ~new_n28072_ | ~new_n27799_;
  assign new_n28091_ = ~new_n28089_ | ~new_n27950_;
  assign new_n28092_ = ~new_n29209_ | ~new_n27786_;
  assign new_n28093_ = ~new_n28367_ | ~new_n27787_;
  assign new_n28094_ = ~new_n29210_ | ~new_n27797_;
  assign new_n28095_ = ~new_n28368_ | ~new_n27798_;
  assign new_n28096_ = ~new_n29210_ | ~new_n27797_;
  assign new_n28097_ = ~new_n28368_ | ~new_n27798_;
  assign new_n28098_ = ~new_n28097_ | ~new_n28096_;
  assign new_n28099_ = ~new_n27884_ | ~new_n27885_;
  assign new_n28100_ = ~new_n27942_ | ~new_n28098_;
  assign new_n28101_ = ~new_n29211_ | ~new_n27795_;
  assign new_n28102_ = ~new_n28369_ | ~new_n27796_;
  assign new_n28103_ = ~new_n29211_ | ~new_n27795_;
  assign new_n28104_ = ~new_n28369_ | ~new_n27796_;
  assign new_n28105_ = ~new_n28104_ | ~new_n28103_;
  assign new_n28106_ = ~new_n27886_ | ~new_n27887_;
  assign new_n28107_ = ~new_n27938_ | ~new_n28105_;
  assign new_n28108_ = ~new_n28334_ | ~new_n27889_;
  assign new_n28109_ = ~new_n29212_ | ~new_n27888_;
  assign new_n28110_ = ~new_n28334_ | ~new_n27889_;
  assign new_n28111_ = ~new_n29212_ | ~new_n27888_;
  assign new_n28112_ = ~new_n28111_ | ~new_n28110_;
  assign new_n28113_ = ~new_n29213_ | ~new_n27793_;
  assign new_n28114_ = ~new_n28333_ | ~new_n27794_;
  assign new_n28115_ = ~new_n29213_ | ~new_n27793_;
  assign new_n28116_ = ~new_n28333_ | ~new_n27794_;
  assign new_n28117_ = ~new_n28116_ | ~new_n28115_;
  assign new_n28118_ = ~new_n27891_ | ~new_n27892_;
  assign new_n28119_ = ~new_n27934_ | ~new_n28117_;
  assign new_n28120_ = ~new_n28370_ | ~new_n27849_;
  assign new_n28121_ = ~new_n29214_ | ~new_n27850_;
  assign new_n28122_ = ~new_n28370_ | ~new_n27849_;
  assign new_n28123_ = ~new_n29214_ | ~new_n27850_;
  assign new_n28124_ = ~new_n28123_ | ~new_n28122_;
  assign new_n28125_ = ~new_n27893_ | ~new_n27851_;
  assign new_n28126_ = ~new_n28124_ | ~new_n28048_;
  assign new_n28127_ = ~new_n28371_ | ~new_n27847_;
  assign new_n28128_ = ~new_n29215_ | ~new_n27848_;
  assign new_n28129_ = ~new_n28371_ | ~new_n27847_;
  assign new_n28130_ = ~new_n29215_ | ~new_n27848_;
  assign new_n28131_ = ~new_n28130_ | ~new_n28129_;
  assign new_n28132_ = ~new_n27894_ | ~new_n27895_;
  assign new_n28133_ = ~new_n28044_ | ~new_n28131_;
  assign new_n28134_ = ~new_n29216_ | ~new_n27845_;
  assign new_n28135_ = ~new_n28372_ | ~new_n27846_;
  assign new_n28136_ = ~new_n29216_ | ~new_n27845_;
  assign new_n28137_ = ~new_n28372_ | ~new_n27846_;
  assign new_n28138_ = ~new_n28137_ | ~new_n28136_;
  assign new_n28139_ = ~new_n27896_ | ~new_n27897_;
  assign new_n28140_ = ~new_n28040_ | ~new_n28138_;
  assign new_n28141_ = ~new_n29217_ | ~new_n27843_;
  assign new_n28142_ = ~new_n28373_ | ~new_n27844_;
  assign new_n28143_ = ~new_n29217_ | ~new_n27843_;
  assign new_n28144_ = ~new_n28373_ | ~new_n27844_;
  assign new_n28145_ = ~new_n28144_ | ~new_n28143_;
  assign new_n28146_ = ~new_n27898_ | ~new_n27899_;
  assign new_n28147_ = ~new_n28036_ | ~new_n28145_;
  assign new_n28148_ = ~new_n29218_ | ~new_n27841_;
  assign new_n28149_ = ~new_n28374_ | ~new_n27842_;
  assign new_n28150_ = ~new_n29218_ | ~new_n27841_;
  assign new_n28151_ = ~new_n28374_ | ~new_n27842_;
  assign new_n28152_ = ~new_n28151_ | ~new_n28150_;
  assign new_n28153_ = ~new_n27900_ | ~new_n27901_;
  assign new_n28154_ = ~new_n28032_ | ~new_n28152_;
  assign new_n28155_ = ~new_n29219_ | ~new_n27839_;
  assign new_n28156_ = ~new_n28375_ | ~new_n27840_;
  assign new_n28157_ = ~new_n29219_ | ~new_n27839_;
  assign new_n28158_ = ~new_n28375_ | ~new_n27840_;
  assign new_n28159_ = ~new_n28158_ | ~new_n28157_;
  assign new_n28160_ = ~new_n27902_ | ~new_n27903_;
  assign new_n28161_ = ~new_n28028_ | ~new_n28159_;
  assign new_n28162_ = ~new_n29220_ | ~new_n27837_;
  assign new_n28163_ = ~new_n28376_ | ~new_n27838_;
  assign new_n28164_ = ~new_n29220_ | ~new_n27837_;
  assign new_n28165_ = ~new_n28376_ | ~new_n27838_;
  assign new_n28166_ = ~new_n28165_ | ~new_n28164_;
  assign new_n28167_ = ~new_n27904_ | ~new_n27905_;
  assign new_n28168_ = ~new_n28024_ | ~new_n28166_;
  assign new_n28169_ = ~new_n29221_ | ~new_n27835_;
  assign new_n28170_ = ~new_n28377_ | ~new_n27836_;
  assign new_n28171_ = ~new_n29221_ | ~new_n27835_;
  assign new_n28172_ = ~new_n28377_ | ~new_n27836_;
  assign new_n28173_ = ~new_n28172_ | ~new_n28171_;
  assign new_n28174_ = ~new_n27906_ | ~new_n27907_;
  assign new_n28175_ = ~new_n28020_ | ~new_n28173_;
  assign new_n28176_ = ~new_n29222_ | ~new_n27833_;
  assign new_n28177_ = ~new_n28378_ | ~new_n27834_;
  assign new_n28178_ = ~new_n29222_ | ~new_n27833_;
  assign new_n28179_ = ~new_n28378_ | ~new_n27834_;
  assign new_n28180_ = ~new_n28179_ | ~new_n28178_;
  assign new_n28181_ = ~new_n27908_ | ~new_n27909_;
  assign new_n28182_ = ~new_n28016_ | ~new_n28180_;
  assign new_n28183_ = ~new_n29223_ | ~new_n27831_;
  assign new_n28184_ = ~new_n28379_ | ~new_n27832_;
  assign new_n28185_ = ~new_n29223_ | ~new_n27831_;
  assign new_n28186_ = ~new_n28379_ | ~new_n27832_;
  assign new_n28187_ = ~new_n28186_ | ~new_n28185_;
  assign new_n28188_ = ~new_n27910_ | ~new_n27911_;
  assign new_n28189_ = ~new_n28012_ | ~new_n28187_;
  assign new_n28190_ = ~new_n28361_ | ~new_n27791_;
  assign new_n28191_ = ~new_n27931_ | ~new_n27790_;
  assign new_n28192_ = ~new_n28191_ | ~new_n28190_;
  assign new_n28193_ = ~new_n27790_ | ~new_n29187_ | ~new_n27791_;
  assign new_n28194_ = ~new_n27929_ | ~new_n28361_;
  assign new_n28195_ = ~new_n29224_ | ~new_n27829_;
  assign new_n28196_ = ~new_n28380_ | ~new_n27830_;
  assign new_n28197_ = ~new_n29224_ | ~new_n27829_;
  assign new_n28198_ = ~new_n28380_ | ~new_n27830_;
  assign new_n28199_ = ~new_n28198_ | ~new_n28197_;
  assign new_n28200_ = ~new_n27914_ | ~new_n27915_;
  assign new_n28201_ = ~new_n28008_ | ~new_n28199_;
  assign new_n28202_ = ~new_n29225_ | ~new_n27827_;
  assign new_n28203_ = ~new_n28381_ | ~new_n27828_;
  assign new_n28204_ = ~new_n29225_ | ~new_n27827_;
  assign new_n28205_ = ~new_n28381_ | ~new_n27828_;
  assign new_n28206_ = ~new_n28205_ | ~new_n28204_;
  assign new_n28207_ = ~new_n27916_ | ~new_n27917_;
  assign new_n28208_ = ~new_n28004_ | ~new_n28206_;
  assign new_n28209_ = ~new_n29226_ | ~new_n27825_;
  assign new_n28210_ = ~new_n28382_ | ~new_n27826_;
  assign new_n28211_ = ~new_n29226_ | ~new_n27825_;
  assign new_n28212_ = ~new_n28382_ | ~new_n27826_;
  assign new_n28213_ = ~new_n28212_ | ~new_n28211_;
  assign new_n28214_ = ~new_n27918_ | ~new_n27919_;
  assign new_n28215_ = ~new_n28000_ | ~new_n28213_;
  assign new_n28216_ = ~new_n29227_ | ~new_n27823_;
  assign new_n28217_ = ~new_n28383_ | ~new_n27824_;
  assign new_n28218_ = ~new_n29227_ | ~new_n27823_;
  assign new_n28219_ = ~new_n28383_ | ~new_n27824_;
  assign new_n28220_ = ~new_n28219_ | ~new_n28218_;
  assign new_n28221_ = ~new_n27920_ | ~new_n27921_;
  assign new_n28222_ = ~new_n27996_ | ~new_n28220_;
  assign new_n28223_ = ~new_n29228_ | ~new_n27809_;
  assign new_n28224_ = ~new_n28384_ | ~new_n27810_;
  assign new_n28225_ = ~new_n29229_ | ~new_n27811_;
  assign new_n28226_ = ~new_n28385_ | ~new_n27812_;
  assign new_n28227_ = ~new_n28226_ | ~new_n28225_;
  assign new_n28228_ = ~new_n28073_ | ~new_n27822_;
  assign new_n28229_ = ~new_n28227_ | ~new_n27990_;
  assign new_n28230_ = ~new_n29230_ | ~new_n27813_;
  assign new_n28231_ = ~new_n28386_ | ~new_n27814_;
  assign new_n28232_ = ~new_n29231_ | ~new_n27820_;
  assign new_n28233_ = ~new_n28387_ | ~new_n27821_;
  assign new_n28234_ = ~new_n29231_ | ~new_n27820_;
  assign new_n28235_ = ~new_n28387_ | ~new_n27821_;
  assign new_n28236_ = ~new_n28235_ | ~new_n28234_;
  assign new_n28237_ = ~new_n27924_ | ~new_n27925_;
  assign new_n28238_ = ~new_n27982_ | ~new_n28236_;
  assign new_n28239_ = ~new_n29232_ | ~new_n27815_;
  assign new_n28240_ = ~new_n28388_ | ~new_n27816_;
  assign new_n28241_ = ~new_n29233_ | ~new_n27817_;
  assign new_n28242_ = ~new_n28389_ | ~new_n27818_;
  assign new_n28243_ = ~new_n28242_ | ~new_n28241_;
  assign new_n28244_ = ~new_n28074_ | ~new_n27819_;
  assign new_n28245_ = ~new_n28243_ | ~new_n27976_;
  assign new_n28246_ = ~new_n28362_ | ~new_n27788_;
  assign new_n28247_ = ~new_n29204_ | ~new_n27789_;
  assign new_n28248_ = ~new_n9647_;
  assign new_n28249_ = ~new_n9632_;
  assign new_n28250_ = ~new_n9632_ | ~new_n9647_;
  assign new_n28251_ = ~new_n9633_;
  assign new_n28252_ = ~new_n9633_ | ~new_n28272_;
  assign new_n28253_ = ~new_n9634_;
  assign new_n28254_ = ~new_n9634_ | ~new_n28273_;
  assign new_n28255_ = ~new_n9635_;
  assign new_n28256_ = ~new_n9635_ | ~new_n28274_;
  assign new_n28257_ = ~new_n9636_;
  assign new_n28258_ = ~new_n9636_ | ~new_n28275_;
  assign new_n28259_ = ~new_n9637_;
  assign new_n28260_ = ~new_n9637_ | ~new_n28276_;
  assign new_n28261_ = ~new_n9638_;
  assign new_n28262_ = ~new_n28280_ | ~new_n28279_;
  assign new_n28263_ = ~new_n28282_ | ~new_n28281_;
  assign new_n28264_ = ~new_n28284_ | ~new_n28283_;
  assign new_n28265_ = ~new_n28286_ | ~new_n28285_;
  assign new_n28266_ = ~new_n28288_ | ~new_n28287_;
  assign new_n28267_ = ~new_n28290_ | ~new_n28289_;
  assign new_n28268_ = ~new_n28292_ | ~new_n28291_;
  assign new_n28269_ = ~new_n28294_ | ~new_n28293_;
  assign new_n28270_ = ~new_n9639_;
  assign new_n28271_ = ~new_n9638_ | ~new_n28277_;
  assign new_n28272_ = ~new_n28250_;
  assign new_n28273_ = ~new_n28252_;
  assign new_n28274_ = ~new_n28254_;
  assign new_n28275_ = ~new_n28256_;
  assign new_n28276_ = ~new_n28258_;
  assign new_n28277_ = ~new_n28260_;
  assign new_n28278_ = ~new_n28271_;
  assign new_n28279_ = ~new_n9639_ | ~new_n28271_;
  assign new_n28280_ = ~new_n28278_ | ~new_n28270_;
  assign new_n28281_ = ~new_n9638_ | ~new_n28260_;
  assign new_n28282_ = ~new_n28277_ | ~new_n28261_;
  assign new_n28283_ = ~new_n9633_ | ~new_n28250_;
  assign new_n28284_ = ~new_n28272_ | ~new_n28251_;
  assign new_n28285_ = ~new_n9635_ | ~new_n28254_;
  assign new_n28286_ = ~new_n28274_ | ~new_n28255_;
  assign new_n28287_ = ~new_n9636_ | ~new_n28256_;
  assign new_n28288_ = ~new_n28275_ | ~new_n28257_;
  assign new_n28289_ = ~new_n9632_ | ~new_n28248_;
  assign new_n28290_ = ~new_n9647_ | ~new_n28249_;
  assign new_n28291_ = ~new_n9637_ | ~new_n28258_;
  assign new_n28292_ = ~new_n28276_ | ~new_n28259_;
  assign new_n28293_ = ~new_n9634_ | ~new_n28252_;
  assign new_n28294_ = ~new_n28273_ | ~new_n28253_;
  assign new_n28295_ = ~new_n10659_;
  assign new_n28296_ = ~new_n10660_;
  assign new_n28297_ = new_n9712_ & new_n28313_;
  assign new_n28298_ = new_n9711_ & new_n28297_;
  assign new_n28299_ = new_n9710_ & new_n28298_;
  assign new_n28300_ = new_n9731_ & new_n28301_;
  assign new_n28301_ = new_n9732_ & new_n28304_;
  assign new_n28302_ = new_n9716_ & new_n28314_;
  assign new_n28303_ = new_n9715_ & new_n28302_;
  assign new_n28304_ = new_n9733_ & new_n28306_;
  assign new_n28305_ = new_n9735_ & new_n28311_;
  assign new_n28306_ = new_n9734_ & new_n28305_;
  assign new_n28307_ = new_n9709_ & new_n28299_;
  assign new_n28308_ = new_n9708_ & new_n28307_;
  assign new_n28309_ = new_n9707_ & new_n28308_;
  assign new_n28310_ = new_n9737_ & new_n28309_;
  assign new_n28311_ = new_n9736_ & new_n28310_;
  assign new_n28312_ = new_n9714_ & new_n28303_;
  assign new_n28313_ = new_n9713_ & new_n28312_;
  assign new_n28314_ = new_n9717_ & new_n28395_;
  assign new_n28315_ = ~new_n9716_;
  assign new_n28316_ = ~new_n9712_;
  assign new_n28317_ = ~new_n9717_;
  assign new_n28318_ = ~new_n9707_;
  assign new_n28319_ = ~new_n9708_;
  assign new_n28320_ = ~new_n9737_;
  assign new_n28321_ = ~new_n9736_;
  assign new_n28322_ = ~new_n9735_;
  assign new_n28323_ = ~new_n9734_;
  assign new_n28324_ = ~new_n9733_;
  assign new_n28325_ = ~new_n9732_;
  assign new_n28326_ = ~new_n9711_;
  assign new_n28327_ = ~new_n9713_;
  assign new_n28328_ = ~new_n9715_;
  assign new_n28329_ = ~new_n9714_;
  assign new_n28330_ = ~new_n9731_;
  assign new_n28331_ = ~new_n9709_;
  assign new_n28332_ = ~new_n9710_;
  assign new_n28333_ = new_n28485_ & new_n28483_;
  assign new_n28334_ = new_n28479_ & new_n28475_;
  assign new_n28335_ = ~new_n9741_;
  assign new_n28336_ = ~new_n9720_;
  assign new_n28337_ = ~new_n9743_;
  assign new_n28338_ = ~new_n9722_;
  assign new_n28339_ = ~new_n9722_ | ~new_n9743_;
  assign new_n28340_ = ~new_n9721_;
  assign new_n28341_ = ~new_n9740_;
  assign new_n28342_ = ~new_n9719_;
  assign new_n28343_ = ~new_n9739_;
  assign new_n28344_ = ~new_n9718_;
  assign new_n28345_ = ~new_n9730_;
  assign new_n28346_ = ~new_n9706_;
  assign new_n28347_ = ~new_n9729_;
  assign new_n28348_ = ~new_n9705_;
  assign new_n28349_ = ~new_n9728_;
  assign new_n28350_ = ~new_n9704_;
  assign new_n28351_ = ~new_n9727_;
  assign new_n28352_ = ~new_n9703_;
  assign new_n28353_ = ~new_n9726_;
  assign new_n28354_ = ~new_n9702_;
  assign new_n28355_ = ~new_n9725_;
  assign new_n28356_ = ~new_n9701_;
  assign new_n28357_ = ~new_n9724_;
  assign new_n28358_ = ~new_n9700_;
  assign new_n28359_ = ~new_n28470_ | ~new_n28469_;
  assign new_n28360_ = ~new_n9742_;
  assign new_n28361_ = ~new_n28576_ | ~new_n28575_;
  assign new_n28362_ = ~new_n28598_ | ~new_n28597_;
  assign new_n28363_ = ~new_n28487_ | ~new_n28486_;
  assign new_n28364_ = ~new_n28489_ | ~new_n28488_;
  assign new_n28365_ = ~new_n28491_ | ~new_n28490_;
  assign new_n28366_ = ~new_n28493_ | ~new_n28492_;
  assign new_n28367_ = ~new_n28495_ | ~new_n28494_;
  assign new_n28368_ = ~new_n28502_ | ~new_n28501_;
  assign new_n28369_ = ~new_n28509_ | ~new_n28508_;
  assign new_n28370_ = ~new_n28523_ | ~new_n28522_;
  assign new_n28371_ = ~new_n28530_ | ~new_n28529_;
  assign new_n28372_ = ~new_n28537_ | ~new_n28536_;
  assign new_n28373_ = ~new_n28544_ | ~new_n28543_;
  assign new_n28374_ = ~new_n28551_ | ~new_n28550_;
  assign new_n28375_ = ~new_n28558_ | ~new_n28557_;
  assign new_n28376_ = ~new_n28565_ | ~new_n28564_;
  assign new_n28377_ = ~new_n28567_ | ~new_n28566_;
  assign new_n28378_ = ~new_n28569_ | ~new_n28568_;
  assign new_n28379_ = ~new_n28571_ | ~new_n28570_;
  assign new_n28380_ = ~new_n28578_ | ~new_n28577_;
  assign new_n28381_ = ~new_n28580_ | ~new_n28579_;
  assign new_n28382_ = ~new_n28582_ | ~new_n28581_;
  assign new_n28383_ = ~new_n28584_ | ~new_n28583_;
  assign new_n28384_ = ~new_n28586_ | ~new_n28585_;
  assign new_n28385_ = ~new_n28588_ | ~new_n28587_;
  assign new_n28386_ = ~new_n28590_ | ~new_n28589_;
  assign new_n28387_ = ~new_n28592_ | ~new_n28591_;
  assign new_n28388_ = ~new_n28594_ | ~new_n28593_;
  assign new_n28389_ = ~new_n28596_ | ~new_n28595_;
  assign new_n28390_ = new_n28474_ & new_n28511_ & new_n28510_;
  assign new_n28391_ = new_n28478_ & new_n28514_;
  assign new_n28392_ = new_n28482_ & new_n28516_ & new_n28515_;
  assign new_n28393_ = new_n28484_ & new_n28418_;
  assign new_n28394_ = ~new_n28573_ | ~new_n28572_;
  assign new_n28395_ = ~new_n28428_ | ~new_n28427_;
  assign new_n28396_ = new_n28497_ & new_n28496_;
  assign new_n28397_ = ~new_n28424_ | ~new_n28423_;
  assign new_n28398_ = new_n28504_ & new_n28503_;
  assign new_n28399_ = ~new_n28419_ | ~new_n28420_;
  assign new_n28400_ = ~new_n9699_;
  assign new_n28401_ = ~new_n9723_;
  assign new_n28402_ = new_n28518_ & new_n28517_;
  assign new_n28403_ = new_n28525_ & new_n28524_;
  assign new_n28404_ = ~new_n28466_ | ~new_n28465_;
  assign new_n28405_ = new_n28532_ & new_n28531_;
  assign new_n28406_ = ~new_n28462_ | ~new_n28461_;
  assign new_n28407_ = new_n28539_ & new_n28538_;
  assign new_n28408_ = ~new_n28458_ | ~new_n28457_;
  assign new_n28409_ = new_n28546_ & new_n28545_;
  assign new_n28410_ = ~new_n28454_ | ~new_n28453_;
  assign new_n28411_ = new_n28553_ & new_n28552_;
  assign new_n28412_ = ~new_n28450_ | ~new_n28449_;
  assign new_n28413_ = new_n28560_ & new_n28559_;
  assign new_n28414_ = ~new_n28339_;
  assign new_n28415_ = ~new_n9721_ | ~new_n28414_;
  assign new_n28416_ = ~new_n28415_ | ~new_n28360_;
  assign new_n28417_ = new_n9720_ | new_n9741_;
  assign new_n28418_ = ~new_n28339_ | ~new_n28340_;
  assign new_n28419_ = ~new_n28417_ | ~new_n28418_ | ~new_n28416_;
  assign new_n28420_ = ~new_n9720_ | ~new_n9741_;
  assign new_n28421_ = ~new_n28399_;
  assign new_n28422_ = new_n9740_ | new_n9719_;
  assign new_n28423_ = ~new_n28422_ | ~new_n28399_;
  assign new_n28424_ = ~new_n9719_ | ~new_n9740_;
  assign new_n28425_ = ~new_n28397_;
  assign new_n28426_ = new_n9739_ | new_n9718_;
  assign new_n28427_ = ~new_n28426_ | ~new_n28397_;
  assign new_n28428_ = ~new_n9718_ | ~new_n9739_;
  assign new_n28429_ = ~new_n28395_;
  assign new_n28430_ = ~new_n28314_;
  assign new_n28431_ = ~new_n28302_;
  assign new_n28432_ = ~new_n28303_;
  assign new_n28433_ = ~new_n28312_;
  assign new_n28434_ = ~new_n28313_;
  assign new_n28435_ = ~new_n28297_;
  assign new_n28436_ = ~new_n28298_;
  assign new_n28437_ = ~new_n28299_;
  assign new_n28438_ = ~new_n28307_;
  assign new_n28439_ = ~new_n28308_;
  assign new_n28440_ = ~new_n28309_;
  assign new_n28441_ = ~new_n28310_;
  assign new_n28442_ = ~new_n28311_;
  assign new_n28443_ = ~new_n28305_;
  assign new_n28444_ = ~new_n28306_;
  assign new_n28445_ = ~new_n28304_;
  assign new_n28446_ = ~new_n28301_;
  assign new_n28447_ = ~new_n28300_;
  assign new_n28448_ = new_n9730_ | new_n9706_;
  assign new_n28449_ = ~new_n28448_ | ~new_n28300_;
  assign new_n28450_ = ~new_n9706_ | ~new_n9730_;
  assign new_n28451_ = ~new_n28412_;
  assign new_n28452_ = new_n9729_ | new_n9705_;
  assign new_n28453_ = ~new_n28452_ | ~new_n28412_;
  assign new_n28454_ = ~new_n9705_ | ~new_n9729_;
  assign new_n28455_ = ~new_n28410_;
  assign new_n28456_ = new_n9728_ | new_n9704_;
  assign new_n28457_ = ~new_n28456_ | ~new_n28410_;
  assign new_n28458_ = ~new_n9704_ | ~new_n9728_;
  assign new_n28459_ = ~new_n28408_;
  assign new_n28460_ = new_n9727_ | new_n9703_;
  assign new_n28461_ = ~new_n28460_ | ~new_n28408_;
  assign new_n28462_ = ~new_n9703_ | ~new_n9727_;
  assign new_n28463_ = ~new_n28406_;
  assign new_n28464_ = new_n9726_ | new_n9702_;
  assign new_n28465_ = ~new_n28464_ | ~new_n28406_;
  assign new_n28466_ = ~new_n9702_ | ~new_n9726_;
  assign new_n28467_ = ~new_n28404_;
  assign new_n28468_ = new_n9725_ | new_n9701_;
  assign new_n28469_ = ~new_n28468_ | ~new_n28404_;
  assign new_n28470_ = ~new_n9701_ | ~new_n9725_;
  assign new_n28471_ = ~new_n28359_;
  assign new_n28472_ = new_n9724_ | new_n9700_;
  assign new_n28473_ = ~new_n28472_ | ~new_n28359_;
  assign new_n28474_ = ~new_n9700_ | ~new_n9724_;
  assign new_n28475_ = ~new_n28390_ | ~new_n28473_;
  assign new_n28476_ = ~new_n9700_ | ~new_n9724_;
  assign new_n28477_ = ~new_n28471_ | ~new_n28476_;
  assign new_n28478_ = new_n9700_ | new_n9724_;
  assign new_n28479_ = ~new_n28391_ | ~new_n28477_;
  assign new_n28480_ = ~new_n28340_ | ~new_n28339_;
  assign new_n28481_ = ~new_n9742_ | ~new_n28480_;
  assign new_n28482_ = ~new_n9721_ | ~new_n28414_;
  assign new_n28483_ = ~new_n28392_ | ~new_n28481_;
  assign new_n28484_ = ~new_n9720_ | ~new_n9741_;
  assign new_n28485_ = ~new_n28393_ | ~new_n28417_ | ~new_n28416_;
  assign new_n28486_ = ~new_n28327_ | ~new_n28312_;
  assign new_n28487_ = ~new_n28433_ | ~new_n9713_;
  assign new_n28488_ = ~new_n28329_ | ~new_n28303_;
  assign new_n28489_ = ~new_n28432_ | ~new_n9714_;
  assign new_n28490_ = ~new_n28328_ | ~new_n28302_;
  assign new_n28491_ = ~new_n28431_ | ~new_n9715_;
  assign new_n28492_ = ~new_n28315_ | ~new_n28314_;
  assign new_n28493_ = ~new_n28430_ | ~new_n9716_;
  assign new_n28494_ = ~new_n28317_ | ~new_n28395_;
  assign new_n28495_ = ~new_n28429_ | ~new_n9717_;
  assign new_n28496_ = ~new_n9718_ | ~new_n28343_;
  assign new_n28497_ = ~new_n9739_ | ~new_n28344_;
  assign new_n28498_ = ~new_n9718_ | ~new_n28343_;
  assign new_n28499_ = ~new_n9739_ | ~new_n28344_;
  assign new_n28500_ = ~new_n28499_ | ~new_n28498_;
  assign new_n28501_ = ~new_n28396_ | ~new_n28397_;
  assign new_n28502_ = ~new_n28425_ | ~new_n28500_;
  assign new_n28503_ = ~new_n9719_ | ~new_n28341_;
  assign new_n28504_ = ~new_n9740_ | ~new_n28342_;
  assign new_n28505_ = ~new_n9719_ | ~new_n28341_;
  assign new_n28506_ = ~new_n9740_ | ~new_n28342_;
  assign new_n28507_ = ~new_n28506_ | ~new_n28505_;
  assign new_n28508_ = ~new_n28398_ | ~new_n28399_;
  assign new_n28509_ = ~new_n28421_ | ~new_n28507_;
  assign new_n28510_ = ~new_n9699_ | ~new_n28401_;
  assign new_n28511_ = ~new_n9723_ | ~new_n28400_;
  assign new_n28512_ = ~new_n9699_ | ~new_n28401_;
  assign new_n28513_ = ~new_n9723_ | ~new_n28400_;
  assign new_n28514_ = ~new_n28513_ | ~new_n28512_;
  assign new_n28515_ = ~new_n9720_ | ~new_n28335_;
  assign new_n28516_ = ~new_n9741_ | ~new_n28336_;
  assign new_n28517_ = ~new_n9700_ | ~new_n28357_;
  assign new_n28518_ = ~new_n9724_ | ~new_n28358_;
  assign new_n28519_ = ~new_n9700_ | ~new_n28357_;
  assign new_n28520_ = ~new_n9724_ | ~new_n28358_;
  assign new_n28521_ = ~new_n28520_ | ~new_n28519_;
  assign new_n28522_ = ~new_n28402_ | ~new_n28359_;
  assign new_n28523_ = ~new_n28521_ | ~new_n28471_;
  assign new_n28524_ = ~new_n9701_ | ~new_n28355_;
  assign new_n28525_ = ~new_n9725_ | ~new_n28356_;
  assign new_n28526_ = ~new_n9701_ | ~new_n28355_;
  assign new_n28527_ = ~new_n9725_ | ~new_n28356_;
  assign new_n28528_ = ~new_n28527_ | ~new_n28526_;
  assign new_n28529_ = ~new_n28403_ | ~new_n28404_;
  assign new_n28530_ = ~new_n28467_ | ~new_n28528_;
  assign new_n28531_ = ~new_n9702_ | ~new_n28353_;
  assign new_n28532_ = ~new_n9726_ | ~new_n28354_;
  assign new_n28533_ = ~new_n9702_ | ~new_n28353_;
  assign new_n28534_ = ~new_n9726_ | ~new_n28354_;
  assign new_n28535_ = ~new_n28534_ | ~new_n28533_;
  assign new_n28536_ = ~new_n28405_ | ~new_n28406_;
  assign new_n28537_ = ~new_n28463_ | ~new_n28535_;
  assign new_n28538_ = ~new_n9703_ | ~new_n28351_;
  assign new_n28539_ = ~new_n9727_ | ~new_n28352_;
  assign new_n28540_ = ~new_n9703_ | ~new_n28351_;
  assign new_n28541_ = ~new_n9727_ | ~new_n28352_;
  assign new_n28542_ = ~new_n28541_ | ~new_n28540_;
  assign new_n28543_ = ~new_n28407_ | ~new_n28408_;
  assign new_n28544_ = ~new_n28459_ | ~new_n28542_;
  assign new_n28545_ = ~new_n9704_ | ~new_n28349_;
  assign new_n28546_ = ~new_n9728_ | ~new_n28350_;
  assign new_n28547_ = ~new_n9704_ | ~new_n28349_;
  assign new_n28548_ = ~new_n9728_ | ~new_n28350_;
  assign new_n28549_ = ~new_n28548_ | ~new_n28547_;
  assign new_n28550_ = ~new_n28409_ | ~new_n28410_;
  assign new_n28551_ = ~new_n28455_ | ~new_n28549_;
  assign new_n28552_ = ~new_n9705_ | ~new_n28347_;
  assign new_n28553_ = ~new_n9729_ | ~new_n28348_;
  assign new_n28554_ = ~new_n9705_ | ~new_n28347_;
  assign new_n28555_ = ~new_n9729_ | ~new_n28348_;
  assign new_n28556_ = ~new_n28555_ | ~new_n28554_;
  assign new_n28557_ = ~new_n28411_ | ~new_n28412_;
  assign new_n28558_ = ~new_n28451_ | ~new_n28556_;
  assign new_n28559_ = ~new_n9706_ | ~new_n28345_;
  assign new_n28560_ = ~new_n9730_ | ~new_n28346_;
  assign new_n28561_ = ~new_n9706_ | ~new_n28345_;
  assign new_n28562_ = ~new_n9730_ | ~new_n28346_;
  assign new_n28563_ = ~new_n28562_ | ~new_n28561_;
  assign new_n28564_ = ~new_n28413_ | ~new_n28300_;
  assign new_n28565_ = ~new_n28447_ | ~new_n28563_;
  assign new_n28566_ = ~new_n28330_ | ~new_n28301_;
  assign new_n28567_ = ~new_n28446_ | ~new_n9731_;
  assign new_n28568_ = ~new_n28325_ | ~new_n28304_;
  assign new_n28569_ = ~new_n28445_ | ~new_n9732_;
  assign new_n28570_ = ~new_n28324_ | ~new_n28306_;
  assign new_n28571_ = ~new_n28444_ | ~new_n9733_;
  assign new_n28572_ = ~new_n28414_ | ~new_n28340_;
  assign new_n28573_ = ~new_n9721_ | ~new_n28339_;
  assign new_n28574_ = ~new_n28394_;
  assign new_n28575_ = ~new_n28574_ | ~new_n9742_;
  assign new_n28576_ = ~new_n28394_ | ~new_n28360_;
  assign new_n28577_ = ~new_n28323_ | ~new_n28305_;
  assign new_n28578_ = ~new_n28443_ | ~new_n9734_;
  assign new_n28579_ = ~new_n28322_ | ~new_n28311_;
  assign new_n28580_ = ~new_n28442_ | ~new_n9735_;
  assign new_n28581_ = ~new_n28321_ | ~new_n28310_;
  assign new_n28582_ = ~new_n28441_ | ~new_n9736_;
  assign new_n28583_ = ~new_n28320_ | ~new_n28309_;
  assign new_n28584_ = ~new_n28440_ | ~new_n9737_;
  assign new_n28585_ = ~new_n28318_ | ~new_n28308_;
  assign new_n28586_ = ~new_n28439_ | ~new_n9707_;
  assign new_n28587_ = ~new_n28319_ | ~new_n28307_;
  assign new_n28588_ = ~new_n28438_ | ~new_n9708_;
  assign new_n28589_ = ~new_n28331_ | ~new_n28299_;
  assign new_n28590_ = ~new_n28437_ | ~new_n9709_;
  assign new_n28591_ = ~new_n28332_ | ~new_n28298_;
  assign new_n28592_ = ~new_n28436_ | ~new_n9710_;
  assign new_n28593_ = ~new_n28326_ | ~new_n28297_;
  assign new_n28594_ = ~new_n28435_ | ~new_n9711_;
  assign new_n28595_ = ~new_n28316_ | ~new_n28313_;
  assign new_n28596_ = ~new_n28434_ | ~new_n9712_;
  assign new_n28597_ = ~new_n9722_ | ~new_n28337_;
  assign new_n28598_ = ~new_n9743_ | ~new_n28338_;
  assign new_n28599_ = ~new_n28631_ | ~new_n28635_ | ~new_n28634_;
  assign new_n28600_ = ~new_n9747_;
  assign new_n28601_ = ~new_n9754_;
  assign new_n28602_ = ~new_n9753_;
  assign new_n28603_ = ~new_n9746_;
  assign new_n28604_ = ~new_n9745_;
  assign new_n28605_ = ~new_n9752_;
  assign new_n28606_ = ~new_n9751_;
  assign new_n28607_ = ~new_n9744_;
  assign new_n28608_ = ~new_n9402_;
  assign new_n28609_ = ~new_n9750_;
  assign new_n28610_ = ~pi0627;
  assign new_n28611_ = ~new_n9749_;
  assign new_n28612_ = ~new_n9755_ | ~new_n9756_;
  assign new_n28613_ = ~new_n9748_ | ~new_n28612_;
  assign new_n28614_ = new_n9755_ | new_n9756_;
  assign new_n28615_ = ~new_n9747_ | ~new_n28601_;
  assign new_n28616_ = ~new_n28615_ | ~new_n28614_ | ~new_n28613_;
  assign new_n28617_ = ~new_n9754_ | ~new_n28600_;
  assign new_n28618_ = ~new_n9753_ | ~new_n28603_;
  assign new_n28619_ = ~new_n28616_ | ~new_n28617_ | ~new_n28618_;
  assign new_n28620_ = ~new_n9746_ | ~new_n28602_;
  assign new_n28621_ = ~new_n9745_ | ~new_n28605_;
  assign new_n28622_ = ~new_n28619_ | ~new_n28620_ | ~new_n28621_;
  assign new_n28623_ = ~new_n9752_ | ~new_n28604_;
  assign new_n28624_ = ~new_n9751_ | ~new_n28607_;
  assign new_n28625_ = ~new_n28624_ | ~new_n28623_ | ~new_n28622_;
  assign new_n28626_ = ~new_n9744_ | ~new_n28606_;
  assign new_n28627_ = ~new_n9402_ | ~new_n28609_;
  assign new_n28628_ = ~new_n28627_ | ~new_n28626_ | ~new_n28625_;
  assign new_n28629_ = ~new_n9750_ | ~new_n28608_;
  assign new_n28630_ = ~new_n28629_ | ~new_n28628_;
  assign new_n28631_ = ~new_n28630_ | ~new_n28633_ | ~new_n28632_;
  assign new_n28632_ = ~new_n9402_ | ~new_n28611_;
  assign new_n28633_ = ~new_n9749_ | ~new_n28608_;
  assign new_n28634_ = ~new_n28611_ | ~pi0627 | ~new_n9402_;
  assign new_n28635_ = ~new_n9749_ | ~new_n28610_ | ~new_n28608_;
  assign new_n28636_ = ~pi0766;
  assign new_n28637_ = ~pi0767;
  assign new_n28638_ = ~pi0767 | ~pi0766;
  assign new_n28639_ = ~pi0768;
  assign new_n28640_ = ~pi0768 | ~new_n28729_;
  assign new_n28641_ = ~pi0769;
  assign new_n28642_ = ~pi0769 | ~new_n28730_;
  assign new_n28643_ = ~pi0770;
  assign new_n28644_ = ~pi0770 | ~new_n28731_;
  assign new_n28645_ = ~pi0771;
  assign new_n28646_ = ~pi0771 | ~new_n28732_;
  assign new_n28647_ = ~pi0772;
  assign new_n28648_ = ~pi0772 | ~new_n28733_;
  assign new_n28649_ = ~pi0773;
  assign new_n28650_ = ~pi0773 | ~new_n28734_;
  assign new_n28651_ = ~pi0774;
  assign new_n28652_ = ~pi0775;
  assign new_n28653_ = ~pi0774 | ~new_n28735_;
  assign new_n28654_ = ~new_n28736_ | ~pi0775;
  assign new_n28655_ = ~pi0776;
  assign new_n28656_ = ~pi0776 | ~new_n28737_;
  assign new_n28657_ = ~pi0777;
  assign new_n28658_ = ~pi0777 | ~new_n28738_;
  assign new_n28659_ = ~pi0778;
  assign new_n28660_ = ~pi0778 | ~new_n28739_;
  assign new_n28661_ = ~pi0779;
  assign new_n28662_ = ~pi0779 | ~new_n28740_;
  assign new_n28663_ = ~pi0780;
  assign new_n28664_ = ~pi0780 | ~new_n28741_;
  assign new_n28665_ = ~pi0781;
  assign new_n28666_ = ~pi0781 | ~new_n28742_;
  assign new_n28667_ = ~pi0782;
  assign new_n28668_ = ~pi0782 | ~new_n28743_;
  assign new_n28669_ = ~pi0783;
  assign new_n28670_ = ~pi0783 | ~new_n28744_;
  assign new_n28671_ = ~pi0784;
  assign new_n28672_ = ~pi0784 | ~new_n28745_;
  assign new_n28673_ = ~pi0785;
  assign new_n28674_ = ~pi0785 | ~new_n28746_;
  assign new_n28675_ = ~pi0786;
  assign new_n28676_ = ~pi0786 | ~new_n28747_;
  assign new_n28677_ = ~pi0787;
  assign new_n28678_ = ~pi0787 | ~new_n28748_;
  assign new_n28679_ = ~pi0788;
  assign new_n28680_ = ~pi0788 | ~new_n28749_;
  assign new_n28681_ = ~pi0789;
  assign new_n28682_ = ~pi0789 | ~new_n28750_;
  assign new_n28683_ = ~pi0790;
  assign new_n28684_ = ~pi0790 | ~new_n28751_;
  assign new_n28685_ = ~pi0791;
  assign new_n28686_ = ~pi0791 | ~new_n28752_;
  assign new_n28687_ = ~pi0792;
  assign new_n28688_ = ~pi0792 | ~new_n28753_;
  assign new_n28689_ = ~pi0793;
  assign new_n28690_ = ~pi0793 | ~new_n28754_;
  assign new_n28691_ = ~pi0794;
  assign new_n28692_ = ~pi0794 | ~new_n28755_;
  assign new_n28693_ = ~pi0795;
  assign new_n28694_ = ~pi0795 | ~new_n28756_;
  assign new_n28695_ = ~pi0796;
  assign new_n28696_ = ~new_n28760_ | ~new_n28759_;
  assign new_n28697_ = ~new_n28762_ | ~new_n28761_;
  assign new_n28698_ = ~new_n28764_ | ~new_n28763_;
  assign new_n28699_ = ~new_n28766_ | ~new_n28765_;
  assign new_n28700_ = ~new_n28768_ | ~new_n28767_;
  assign new_n28701_ = ~new_n28770_ | ~new_n28769_;
  assign new_n28702_ = ~new_n28772_ | ~new_n28771_;
  assign new_n28703_ = ~new_n28774_ | ~new_n28773_;
  assign new_n28704_ = ~new_n28776_ | ~new_n28775_;
  assign new_n28705_ = ~new_n28778_ | ~new_n28777_;
  assign new_n28706_ = ~new_n28780_ | ~new_n28779_;
  assign new_n28707_ = ~new_n28782_ | ~new_n28781_;
  assign new_n28708_ = ~new_n28784_ | ~new_n28783_;
  assign new_n28709_ = ~new_n28786_ | ~new_n28785_;
  assign new_n28710_ = ~new_n28788_ | ~new_n28787_;
  assign new_n28711_ = ~new_n28790_ | ~new_n28789_;
  assign new_n28712_ = ~new_n28792_ | ~new_n28791_;
  assign new_n28713_ = ~new_n28794_ | ~new_n28793_;
  assign new_n28714_ = ~new_n28796_ | ~new_n28795_;
  assign new_n28715_ = ~new_n28798_ | ~new_n28797_;
  assign new_n28716_ = ~new_n28800_ | ~new_n28799_;
  assign new_n28717_ = ~new_n28802_ | ~new_n28801_;
  assign new_n28718_ = ~new_n28804_ | ~new_n28803_;
  assign new_n28719_ = ~new_n28806_ | ~new_n28805_;
  assign new_n28720_ = ~new_n28808_ | ~new_n28807_;
  assign new_n28721_ = ~new_n28810_ | ~new_n28809_;
  assign new_n28722_ = ~new_n28812_ | ~new_n28811_;
  assign new_n28723_ = ~new_n28814_ | ~new_n28813_;
  assign new_n28724_ = ~new_n28816_ | ~new_n28815_;
  assign new_n28725_ = ~new_n28818_ | ~new_n28817_;
  assign new_n28726_ = ~new_n28820_ | ~new_n28819_;
  assign new_n28727_ = ~pi0797;
  assign new_n28728_ = ~pi0796 | ~new_n28757_;
  assign new_n28729_ = ~new_n28638_;
  assign new_n28730_ = ~new_n28640_;
  assign new_n28731_ = ~new_n28642_;
  assign new_n28732_ = ~new_n28644_;
  assign new_n28733_ = ~new_n28646_;
  assign new_n28734_ = ~new_n28648_;
  assign new_n28735_ = ~new_n28650_;
  assign new_n28736_ = ~new_n28653_;
  assign new_n28737_ = ~new_n28654_;
  assign new_n28738_ = ~new_n28656_;
  assign new_n28739_ = ~new_n28658_;
  assign new_n28740_ = ~new_n28660_;
  assign new_n28741_ = ~new_n28662_;
  assign new_n28742_ = ~new_n28664_;
  assign new_n28743_ = ~new_n28666_;
  assign new_n28744_ = ~new_n28668_;
  assign new_n28745_ = ~new_n28670_;
  assign new_n28746_ = ~new_n28672_;
  assign new_n28747_ = ~new_n28674_;
  assign new_n28748_ = ~new_n28676_;
  assign new_n28749_ = ~new_n28678_;
  assign new_n28750_ = ~new_n28680_;
  assign new_n28751_ = ~new_n28682_;
  assign new_n28752_ = ~new_n28684_;
  assign new_n28753_ = ~new_n28686_;
  assign new_n28754_ = ~new_n28688_;
  assign new_n28755_ = ~new_n28690_;
  assign new_n28756_ = ~new_n28692_;
  assign new_n28757_ = ~new_n28694_;
  assign new_n28758_ = ~new_n28728_;
  assign new_n28759_ = ~pi0775 | ~new_n28653_;
  assign new_n28760_ = ~new_n28736_ | ~new_n28652_;
  assign new_n28761_ = ~pi0774 | ~new_n28650_;
  assign new_n28762_ = ~new_n28735_ | ~new_n28651_;
  assign new_n28763_ = ~pi0773 | ~new_n28648_;
  assign new_n28764_ = ~new_n28734_ | ~new_n28649_;
  assign new_n28765_ = ~pi0772 | ~new_n28646_;
  assign new_n28766_ = ~new_n28733_ | ~new_n28647_;
  assign new_n28767_ = ~pi0771 | ~new_n28644_;
  assign new_n28768_ = ~new_n28732_ | ~new_n28645_;
  assign new_n28769_ = ~pi0770 | ~new_n28642_;
  assign new_n28770_ = ~new_n28731_ | ~new_n28643_;
  assign new_n28771_ = ~pi0769 | ~new_n28640_;
  assign new_n28772_ = ~new_n28730_ | ~new_n28641_;
  assign new_n28773_ = ~pi0797 | ~new_n28728_;
  assign new_n28774_ = ~new_n28758_ | ~new_n28727_;
  assign new_n28775_ = ~pi0796 | ~new_n28694_;
  assign new_n28776_ = ~new_n28757_ | ~new_n28695_;
  assign new_n28777_ = ~pi0768 | ~new_n28638_;
  assign new_n28778_ = ~new_n28729_ | ~new_n28639_;
  assign new_n28779_ = ~pi0795 | ~new_n28692_;
  assign new_n28780_ = ~new_n28756_ | ~new_n28693_;
  assign new_n28781_ = ~pi0794 | ~new_n28690_;
  assign new_n28782_ = ~new_n28755_ | ~new_n28691_;
  assign new_n28783_ = ~pi0793 | ~new_n28688_;
  assign new_n28784_ = ~new_n28754_ | ~new_n28689_;
  assign new_n28785_ = ~pi0792 | ~new_n28686_;
  assign new_n28786_ = ~new_n28753_ | ~new_n28687_;
  assign new_n28787_ = ~pi0791 | ~new_n28684_;
  assign new_n28788_ = ~new_n28752_ | ~new_n28685_;
  assign new_n28789_ = ~pi0790 | ~new_n28682_;
  assign new_n28790_ = ~new_n28751_ | ~new_n28683_;
  assign new_n28791_ = ~pi0789 | ~new_n28680_;
  assign new_n28792_ = ~new_n28750_ | ~new_n28681_;
  assign new_n28793_ = ~pi0788 | ~new_n28678_;
  assign new_n28794_ = ~new_n28749_ | ~new_n28679_;
  assign new_n28795_ = ~pi0787 | ~new_n28676_;
  assign new_n28796_ = ~new_n28748_ | ~new_n28677_;
  assign new_n28797_ = ~pi0786 | ~new_n28674_;
  assign new_n28798_ = ~new_n28747_ | ~new_n28675_;
  assign new_n28799_ = ~pi0767 | ~new_n28636_;
  assign new_n28800_ = ~pi0766 | ~new_n28637_;
  assign new_n28801_ = ~pi0785 | ~new_n28672_;
  assign new_n28802_ = ~new_n28746_ | ~new_n28673_;
  assign new_n28803_ = ~pi0784 | ~new_n28670_;
  assign new_n28804_ = ~new_n28745_ | ~new_n28671_;
  assign new_n28805_ = ~pi0783 | ~new_n28668_;
  assign new_n28806_ = ~new_n28744_ | ~new_n28669_;
  assign new_n28807_ = ~pi0782 | ~new_n28666_;
  assign new_n28808_ = ~new_n28743_ | ~new_n28667_;
  assign new_n28809_ = ~pi0781 | ~new_n28664_;
  assign new_n28810_ = ~new_n28742_ | ~new_n28665_;
  assign new_n28811_ = ~pi0780 | ~new_n28662_;
  assign new_n28812_ = ~new_n28741_ | ~new_n28663_;
  assign new_n28813_ = ~pi0779 | ~new_n28660_;
  assign new_n28814_ = ~new_n28740_ | ~new_n28661_;
  assign new_n28815_ = ~pi0778 | ~new_n28658_;
  assign new_n28816_ = ~new_n28739_ | ~new_n28659_;
  assign new_n28817_ = ~pi0777 | ~new_n28656_;
  assign new_n28818_ = ~new_n28738_ | ~new_n28657_;
  assign new_n28819_ = ~pi0776 | ~new_n28654_;
  assign new_n28820_ = ~new_n28737_ | ~new_n28655_;
  assign new_n28821_ = new_n28822_ | new_n10658_;
  assign new_n28822_ = ~new_n28295_ & ~new_n28296_;
  assign new_n28823_ = ~pi0799;
  assign new_n28824_ = ~pi0801;
  assign new_n28825_ = ~pi0800;
  assign new_n28826_ = ~pi0800 | ~pi0801 | ~pi0799;
  assign new_n28827_ = ~pi0802;
  assign new_n28828_ = ~pi0802 | ~new_n28914_;
  assign new_n28829_ = ~pi0803;
  assign new_n28830_ = ~pi0803 | ~new_n28915_;
  assign new_n28831_ = ~pi0804;
  assign new_n28832_ = ~pi0804 | ~new_n28916_;
  assign new_n28833_ = ~pi0805;
  assign new_n28834_ = ~pi0805 | ~new_n28917_;
  assign new_n28835_ = ~pi0806;
  assign new_n28836_ = ~pi0807;
  assign new_n28837_ = ~pi0806 | ~new_n28918_;
  assign new_n28838_ = ~new_n28919_ | ~pi0807;
  assign new_n28839_ = ~pi0808;
  assign new_n28840_ = ~pi0808 | ~new_n28920_;
  assign new_n28841_ = ~pi0809;
  assign new_n28842_ = ~pi0809 | ~new_n28921_;
  assign new_n28843_ = ~pi0810;
  assign new_n28844_ = ~pi0810 | ~new_n28922_;
  assign new_n28845_ = ~pi0811;
  assign new_n28846_ = ~pi0811 | ~new_n28923_;
  assign new_n28847_ = ~pi0812;
  assign new_n28848_ = ~pi0812 | ~new_n28924_;
  assign new_n28849_ = ~pi0813;
  assign new_n28850_ = ~pi0813 | ~new_n28925_;
  assign new_n28851_ = ~pi0814;
  assign new_n28852_ = ~pi0814 | ~new_n28926_;
  assign new_n28853_ = ~pi0815;
  assign new_n28854_ = ~pi0815 | ~new_n28927_;
  assign new_n28855_ = ~pi0816;
  assign new_n28856_ = ~pi0816 | ~new_n28928_;
  assign new_n28857_ = ~pi0817;
  assign new_n28858_ = ~pi0817 | ~new_n28929_;
  assign new_n28859_ = ~pi0818;
  assign new_n28860_ = ~pi0818 | ~new_n28930_;
  assign new_n28861_ = ~pi0819;
  assign new_n28862_ = ~pi0819 | ~new_n28931_;
  assign new_n28863_ = ~pi0820;
  assign new_n28864_ = ~pi0820 | ~new_n28932_;
  assign new_n28865_ = ~pi0821;
  assign new_n28866_ = ~pi0821 | ~new_n28933_;
  assign new_n28867_ = ~pi0822;
  assign new_n28868_ = ~pi0822 | ~new_n28934_;
  assign new_n28869_ = ~pi0823;
  assign new_n28870_ = ~pi0823 | ~new_n28935_;
  assign new_n28871_ = ~pi0824;
  assign new_n28872_ = ~pi0824 | ~new_n28936_;
  assign new_n28873_ = ~pi0825;
  assign new_n28874_ = ~pi0825 | ~new_n28937_;
  assign new_n28875_ = ~pi0826;
  assign new_n28876_ = ~pi0826 | ~new_n28938_;
  assign new_n28877_ = ~pi0827;
  assign new_n28878_ = ~pi0827 | ~new_n28939_;
  assign new_n28879_ = ~pi0828;
  assign new_n28880_ = ~new_n28943_ | ~new_n28942_;
  assign new_n28881_ = ~new_n28945_ | ~new_n28944_;
  assign new_n28882_ = ~new_n28947_ | ~new_n28946_;
  assign new_n28883_ = ~new_n28949_ | ~new_n28948_;
  assign new_n28884_ = ~new_n28951_ | ~new_n28950_;
  assign new_n28885_ = ~new_n28953_ | ~new_n28952_;
  assign new_n28886_ = ~new_n28955_ | ~new_n28954_;
  assign new_n28887_ = ~new_n28957_ | ~new_n28956_;
  assign new_n28888_ = ~new_n28959_ | ~new_n28958_;
  assign new_n28889_ = ~new_n28961_ | ~new_n28960_;
  assign new_n28890_ = ~new_n28963_ | ~new_n28962_;
  assign new_n28891_ = ~new_n28965_ | ~new_n28964_;
  assign new_n28892_ = ~new_n28967_ | ~new_n28966_;
  assign new_n28893_ = ~new_n28969_ | ~new_n28968_;
  assign new_n28894_ = ~new_n28971_ | ~new_n28970_;
  assign new_n28895_ = ~new_n28973_ | ~new_n28972_;
  assign new_n28896_ = ~new_n28975_ | ~new_n28974_;
  assign new_n28897_ = ~new_n28977_ | ~new_n28976_;
  assign new_n28898_ = ~new_n28979_ | ~new_n28978_;
  assign new_n28899_ = ~new_n28981_ | ~new_n28980_;
  assign new_n28900_ = ~new_n28983_ | ~new_n28982_;
  assign new_n28901_ = ~new_n28985_ | ~new_n28984_;
  assign new_n28902_ = ~new_n28987_ | ~new_n28986_;
  assign new_n28903_ = ~new_n28989_ | ~new_n28988_;
  assign new_n28904_ = ~new_n28991_ | ~new_n28990_;
  assign new_n28905_ = ~new_n28993_ | ~new_n28992_;
  assign new_n28906_ = ~new_n28995_ | ~new_n28994_;
  assign new_n28907_ = ~new_n28997_ | ~new_n28996_;
  assign new_n28908_ = ~new_n28999_ | ~new_n28998_;
  assign new_n28909_ = ~new_n29001_ | ~new_n29000_;
  assign new_n28910_ = ~pi0800 | ~pi0799;
  assign new_n28911_ = ~pi0829;
  assign new_n28912_ = ~pi0828 | ~new_n28940_;
  assign new_n28913_ = ~new_n28910_;
  assign new_n28914_ = ~new_n28826_;
  assign new_n28915_ = ~new_n28828_;
  assign new_n28916_ = ~new_n28830_;
  assign new_n28917_ = ~new_n28832_;
  assign new_n28918_ = ~new_n28834_;
  assign new_n28919_ = ~new_n28837_;
  assign new_n28920_ = ~new_n28838_;
  assign new_n28921_ = ~new_n28840_;
  assign new_n28922_ = ~new_n28842_;
  assign new_n28923_ = ~new_n28844_;
  assign new_n28924_ = ~new_n28846_;
  assign new_n28925_ = ~new_n28848_;
  assign new_n28926_ = ~new_n28850_;
  assign new_n28927_ = ~new_n28852_;
  assign new_n28928_ = ~new_n28854_;
  assign new_n28929_ = ~new_n28856_;
  assign new_n28930_ = ~new_n28858_;
  assign new_n28931_ = ~new_n28860_;
  assign new_n28932_ = ~new_n28862_;
  assign new_n28933_ = ~new_n28864_;
  assign new_n28934_ = ~new_n28866_;
  assign new_n28935_ = ~new_n28868_;
  assign new_n28936_ = ~new_n28870_;
  assign new_n28937_ = ~new_n28872_;
  assign new_n28938_ = ~new_n28874_;
  assign new_n28939_ = ~new_n28876_;
  assign new_n28940_ = ~new_n28878_;
  assign new_n28941_ = ~new_n28912_;
  assign new_n28942_ = ~pi0807 | ~new_n28837_;
  assign new_n28943_ = ~new_n28919_ | ~new_n28836_;
  assign new_n28944_ = ~pi0806 | ~new_n28834_;
  assign new_n28945_ = ~new_n28918_ | ~new_n28835_;
  assign new_n28946_ = ~pi0805 | ~new_n28832_;
  assign new_n28947_ = ~new_n28917_ | ~new_n28833_;
  assign new_n28948_ = ~pi0804 | ~new_n28830_;
  assign new_n28949_ = ~new_n28916_ | ~new_n28831_;
  assign new_n28950_ = ~pi0803 | ~new_n28828_;
  assign new_n28951_ = ~new_n28915_ | ~new_n28829_;
  assign new_n28952_ = ~pi0802 | ~new_n28826_;
  assign new_n28953_ = ~new_n28914_ | ~new_n28827_;
  assign new_n28954_ = ~pi0801 | ~new_n28910_;
  assign new_n28955_ = ~new_n28913_ | ~new_n28824_;
  assign new_n28956_ = ~pi0829 | ~new_n28912_;
  assign new_n28957_ = ~new_n28941_ | ~new_n28911_;
  assign new_n28958_ = ~pi0828 | ~new_n28878_;
  assign new_n28959_ = ~new_n28940_ | ~new_n28879_;
  assign new_n28960_ = ~pi0800 | ~new_n28823_;
  assign new_n28961_ = ~pi0799 | ~new_n28825_;
  assign new_n28962_ = ~pi0827 | ~new_n28876_;
  assign new_n28963_ = ~new_n28939_ | ~new_n28877_;
  assign new_n28964_ = ~pi0826 | ~new_n28874_;
  assign new_n28965_ = ~new_n28938_ | ~new_n28875_;
  assign new_n28966_ = ~pi0825 | ~new_n28872_;
  assign new_n28967_ = ~new_n28937_ | ~new_n28873_;
  assign new_n28968_ = ~pi0824 | ~new_n28870_;
  assign new_n28969_ = ~new_n28936_ | ~new_n28871_;
  assign new_n28970_ = ~pi0823 | ~new_n28868_;
  assign new_n28971_ = ~new_n28935_ | ~new_n28869_;
  assign new_n28972_ = ~pi0822 | ~new_n28866_;
  assign new_n28973_ = ~new_n28934_ | ~new_n28867_;
  assign new_n28974_ = ~pi0821 | ~new_n28864_;
  assign new_n28975_ = ~new_n28933_ | ~new_n28865_;
  assign new_n28976_ = ~pi0820 | ~new_n28862_;
  assign new_n28977_ = ~new_n28932_ | ~new_n28863_;
  assign new_n28978_ = ~pi0819 | ~new_n28860_;
  assign new_n28979_ = ~new_n28931_ | ~new_n28861_;
  assign new_n28980_ = ~pi0818 | ~new_n28858_;
  assign new_n28981_ = ~new_n28930_ | ~new_n28859_;
  assign new_n28982_ = ~pi0817 | ~new_n28856_;
  assign new_n28983_ = ~new_n28929_ | ~new_n28857_;
  assign new_n28984_ = ~pi0816 | ~new_n28854_;
  assign new_n28985_ = ~new_n28928_ | ~new_n28855_;
  assign new_n28986_ = ~pi0815 | ~new_n28852_;
  assign new_n28987_ = ~new_n28927_ | ~new_n28853_;
  assign new_n28988_ = ~pi0814 | ~new_n28850_;
  assign new_n28989_ = ~new_n28926_ | ~new_n28851_;
  assign new_n28990_ = ~pi0813 | ~new_n28848_;
  assign new_n28991_ = ~new_n28925_ | ~new_n28849_;
  assign new_n28992_ = ~pi0812 | ~new_n28846_;
  assign new_n28993_ = ~new_n28924_ | ~new_n28847_;
  assign new_n28994_ = ~pi0811 | ~new_n28844_;
  assign new_n28995_ = ~new_n28923_ | ~new_n28845_;
  assign new_n28996_ = ~pi0810 | ~new_n28842_;
  assign new_n28997_ = ~new_n28922_ | ~new_n28843_;
  assign new_n28998_ = ~pi0809 | ~new_n28840_;
  assign new_n28999_ = ~new_n28921_ | ~new_n28841_;
  assign new_n29000_ = ~pi0808 | ~new_n28838_;
  assign new_n29001_ = ~new_n28920_ | ~new_n28839_;
  assign new_n29002_ = ~pi0759;
  assign new_n29003_ = ~pi0757;
  assign new_n29004_ = ~pi0758;
  assign new_n29005_ = ~new_n29014_ | ~new_n29013_;
  assign new_n29006_ = ~new_n29016_ | ~new_n29015_;
  assign new_n29007_ = ~new_n29018_ | ~new_n29017_;
  assign new_n29008_ = ~new_n9793_;
  assign new_n29009_ = ~pi0758 | ~pi0757 | ~pi0759;
  assign new_n29010_ = ~pi0758 | ~pi0759;
  assign new_n29011_ = ~new_n29009_;
  assign new_n29012_ = ~new_n29010_;
  assign new_n29013_ = ~new_n9793_ | ~new_n29009_;
  assign new_n29014_ = ~new_n29011_ | ~new_n29008_;
  assign new_n29015_ = ~pi0757 | ~new_n29010_;
  assign new_n29016_ = ~new_n29012_ | ~new_n29003_;
  assign new_n29017_ = ~pi0758 | ~new_n29002_;
  assign new_n29018_ = ~pi0759 | ~new_n29004_;
  assign new_n29019_ = new_n29065_ & new_n29061_;
  assign new_n29020_ = new_n29081_ & new_n29079_;
  assign new_n29021_ = ~new_n29058_ | ~new_n29082_;
  assign new_n29022_ = ~new_n11469_;
  assign new_n29023_ = ~new_n9794_;
  assign new_n29024_ = ~new_n9802_;
  assign new_n29025_ = ~new_n9804_;
  assign new_n29026_ = ~new_n9803_;
  assign new_n29027_ = ~new_n9797_;
  assign new_n29028_ = ~new_n9806_;
  assign new_n29029_ = ~new_n9805_;
  assign new_n29030_ = ~new_n9796_;
  assign new_n29031_ = ~new_n9795_;
  assign new_n29032_ = ~new_n29085_ | ~new_n29089_;
  assign new_n29033_ = ~new_n9801_;
  assign new_n29034_ = ~new_n9800_;
  assign new_n29035_ = ~new_n9799_;
  assign new_n29036_ = ~new_n9798_;
  assign new_n29037_ = ~new_n29099_ | ~new_n29098_;
  assign new_n29038_ = ~new_n29104_ | ~new_n29103_;
  assign new_n29039_ = ~new_n29109_ | ~new_n29108_;
  assign new_n29040_ = ~new_n29114_ | ~new_n29113_;
  assign new_n29041_ = ~new_n29119_ | ~new_n29118_;
  assign new_n29042_ = ~new_n29124_ | ~new_n29123_;
  assign new_n29043_ = ~new_n29129_ | ~new_n29128_;
  assign new_n29044_ = new_n29019_ & new_n29068_;
  assign new_n29045_ = ~new_n29096_ | ~new_n29095_;
  assign new_n29046_ = ~new_n29101_ | ~new_n29100_;
  assign new_n29047_ = ~new_n29106_ | ~new_n29105_;
  assign new_n29048_ = ~new_n29111_ | ~new_n29110_;
  assign new_n29049_ = ~new_n29116_ | ~new_n29115_;
  assign new_n29050_ = ~new_n29121_ | ~new_n29120_;
  assign new_n29051_ = ~new_n29126_ | ~new_n29125_;
  assign new_n29052_ = ~new_n29077_ | ~new_n29076_;
  assign new_n29053_ = ~new_n29073_ | ~new_n29072_;
  assign new_n29054_ = ~new_n29087_ | ~new_n29088_ | ~new_n29069_;
  assign new_n29055_ = ~new_n29032_ | ~new_n29084_;
  assign new_n29056_ = ~new_n29063_ | ~new_n29062_;
  assign new_n29057_ = ~new_n29091_ | ~new_n29083_;
  assign new_n29058_ = ~new_n9806_ | ~new_n29036_;
  assign new_n29059_ = ~new_n29058_;
  assign new_n29060_ = ~new_n9805_ | ~new_n29027_;
  assign new_n29061_ = ~new_n9804_ | ~new_n29030_;
  assign new_n29062_ = ~new_n29061_ | ~new_n29094_;
  assign new_n29063_ = ~new_n9796_ | ~new_n29025_;
  assign new_n29064_ = ~new_n29056_;
  assign new_n29065_ = ~new_n9803_ | ~new_n29031_;
  assign new_n29066_ = ~new_n9795_ | ~new_n29026_;
  assign new_n29067_ = ~new_n29055_;
  assign new_n29068_ = ~new_n9802_ | ~new_n29023_;
  assign new_n29069_ = ~new_n9794_ | ~new_n29024_;
  assign new_n29070_ = ~new_n29054_;
  assign new_n29071_ = ~new_n9801_ | ~new_n29022_;
  assign new_n29072_ = ~new_n29071_ | ~new_n29054_;
  assign new_n29073_ = ~new_n11469_ | ~new_n29033_;
  assign new_n29074_ = ~new_n29053_;
  assign new_n29075_ = ~new_n9800_ | ~new_n29022_;
  assign new_n29076_ = ~new_n29075_ | ~new_n29053_;
  assign new_n29077_ = ~new_n11469_ | ~new_n29034_;
  assign new_n29078_ = ~new_n29052_;
  assign new_n29079_ = ~new_n11469_ | ~new_n29035_;
  assign new_n29080_ = ~new_n9799_ | ~new_n29022_;
  assign new_n29081_ = ~new_n29080_ | ~new_n29052_;
  assign new_n29082_ = ~new_n9798_ | ~new_n29028_;
  assign new_n29083_ = ~new_n9797_ | ~new_n29029_;
  assign new_n29084_ = ~new_n29019_ | ~new_n29057_;
  assign new_n29085_ = ~new_n29066_ | ~new_n29063_;
  assign new_n29086_ = ~new_n29032_;
  assign new_n29087_ = ~new_n29044_ | ~new_n29057_;
  assign new_n29088_ = ~new_n29086_ | ~new_n29068_;
  assign new_n29089_ = ~new_n9803_ | ~new_n29031_;
  assign new_n29090_ = ~new_n9805_ | ~new_n29027_;
  assign new_n29091_ = ~new_n29060_ | ~new_n29058_;
  assign new_n29092_ = ~new_n29057_;
  assign new_n29093_ = ~new_n29090_ | ~new_n29058_;
  assign new_n29094_ = ~new_n29093_ | ~new_n29083_;
  assign new_n29095_ = ~new_n9799_ | ~new_n29022_;
  assign new_n29096_ = ~new_n11469_ | ~new_n29035_;
  assign new_n29097_ = ~new_n29045_;
  assign new_n29098_ = ~new_n29078_ | ~new_n29097_;
  assign new_n29099_ = ~new_n29045_ | ~new_n29052_;
  assign new_n29100_ = ~new_n9800_ | ~new_n29022_;
  assign new_n29101_ = ~new_n11469_ | ~new_n29034_;
  assign new_n29102_ = ~new_n29046_;
  assign new_n29103_ = ~new_n29074_ | ~new_n29102_;
  assign new_n29104_ = ~new_n29046_ | ~new_n29053_;
  assign new_n29105_ = ~new_n9801_ | ~new_n29022_;
  assign new_n29106_ = ~new_n11469_ | ~new_n29033_;
  assign new_n29107_ = ~new_n29047_;
  assign new_n29108_ = ~new_n29070_ | ~new_n29107_;
  assign new_n29109_ = ~new_n29047_ | ~new_n29054_;
  assign new_n29110_ = ~new_n9802_ | ~new_n29023_;
  assign new_n29111_ = ~new_n9794_ | ~new_n29024_;
  assign new_n29112_ = ~new_n29048_;
  assign new_n29113_ = ~new_n29067_ | ~new_n29112_;
  assign new_n29114_ = ~new_n29048_ | ~new_n29055_;
  assign new_n29115_ = ~new_n9803_ | ~new_n29031_;
  assign new_n29116_ = ~new_n9795_ | ~new_n29026_;
  assign new_n29117_ = ~new_n29049_;
  assign new_n29118_ = ~new_n29064_ | ~new_n29117_;
  assign new_n29119_ = ~new_n29049_ | ~new_n29056_;
  assign new_n29120_ = ~new_n9804_ | ~new_n29030_;
  assign new_n29121_ = ~new_n9796_ | ~new_n29025_;
  assign new_n29122_ = ~new_n29050_;
  assign new_n29123_ = ~new_n29092_ | ~new_n29122_;
  assign new_n29124_ = ~new_n29050_ | ~new_n29057_;
  assign new_n29125_ = ~new_n9805_ | ~new_n29027_;
  assign new_n29126_ = ~new_n9797_ | ~new_n29029_;
  assign new_n29127_ = ~new_n29051_;
  assign new_n29128_ = ~new_n29059_ | ~new_n29127_;
  assign new_n29129_ = ~new_n29051_ | ~new_n29058_;
  assign new_n29130_ = ~new_n10726_ & ~new_n10727_ & ~new_n10728_ & ~new_n10725_;
  assign new_n29131_ = ~new_n10725_ & ~new_n29133_;
  assign new_n29132_ = ~new_n29131_ | ~new_n29135_;
  assign new_n29133_ = ~new_n10728_ & ~new_n10730_ & ~new_n10725_ & ~new_n10726_ & ~new_n10727_;
  assign new_n29134_ = ~new_n10729_;
  assign new_n29135_ = ~new_n29130_ | ~new_n29134_;
  assign new_n29136_ = ~new_n10655_;
  assign new_n29137_ = ~new_n10656_;
  assign new_n29138_ = ~new_n9854_;
  assign new_n29139_ = ~new_n10654_;
  assign new_n29140_ = new_n9681_ & new_n29159_;
  assign new_n29141_ = new_n9674_ & new_n29154_;
  assign new_n29142_ = new_n9672_ & new_n29161_;
  assign new_n29143_ = new_n9670_ & new_n29152_;
  assign new_n29144_ = new_n9669_ & new_n29143_;
  assign new_n29145_ = new_n9668_ & new_n29144_;
  assign new_n29146_ = new_n9667_ & new_n29145_;
  assign new_n29147_ = new_n9666_ & new_n29146_;
  assign new_n29148_ = new_n9665_ & new_n29147_;
  assign new_n29149_ = new_n9663_ & new_n29151_;
  assign new_n29150_ = new_n9662_ & new_n29149_;
  assign new_n29151_ = new_n9664_ & new_n29148_;
  assign new_n29152_ = new_n9671_ & new_n29142_;
  assign new_n29153_ = new_n9676_ & new_n29157_;
  assign new_n29154_ = new_n9675_ & new_n29153_;
  assign new_n29155_ = new_n9679_ & new_n29160_;
  assign new_n29156_ = new_n9678_ & new_n29155_;
  assign new_n29157_ = new_n9677_ & new_n29156_;
  assign new_n29158_ = new_n9661_ & new_n29150_;
  assign new_n29159_ = new_n9682_ & new_n29235_;
  assign new_n29160_ = new_n9680_ & new_n29140_;
  assign new_n29161_ = new_n9673_ & new_n29141_;
  assign new_n29162_ = ~new_n9672_;
  assign new_n29163_ = ~new_n9679_;
  assign new_n29164_ = ~new_n9681_;
  assign new_n29165_ = ~new_n9659_;
  assign new_n29166_ = ~new_n9660_;
  assign new_n29167_ = ~new_n9676_;
  assign new_n29168_ = ~new_n9677_;
  assign new_n29169_ = ~new_n9678_;
  assign new_n29170_ = ~new_n9674_;
  assign new_n29171_ = ~new_n9675_;
  assign new_n29172_ = ~new_n9670_;
  assign new_n29173_ = ~new_n9682_;
  assign new_n29174_ = ~new_n9663_;
  assign new_n29175_ = ~new_n9668_;
  assign new_n29176_ = ~new_n9661_;
  assign new_n29177_ = ~new_n9662_;
  assign new_n29178_ = ~new_n9664_;
  assign new_n29179_ = ~new_n9665_;
  assign new_n29180_ = ~new_n9666_;
  assign new_n29181_ = ~new_n9667_;
  assign new_n29182_ = ~new_n9669_;
  assign new_n29183_ = ~new_n9671_;
  assign new_n29184_ = ~new_n9673_;
  assign new_n29185_ = ~new_n9680_;
  assign new_n29186_ = new_n29304_ & new_n29303_;
  assign new_n29187_ = ~new_n29250_ | ~new_n29306_;
  assign new_n29188_ = ~new_n9698_;
  assign new_n29189_ = ~new_n9690_;
  assign new_n29190_ = ~new_n9689_;
  assign new_n29191_ = ~new_n9697_;
  assign new_n29192_ = ~new_n9696_;
  assign new_n29193_ = ~new_n9688_;
  assign new_n29194_ = ~new_n9695_;
  assign new_n29195_ = ~new_n9687_;
  assign new_n29196_ = ~new_n9694_;
  assign new_n29197_ = ~new_n9686_;
  assign new_n29198_ = ~new_n9693_;
  assign new_n29199_ = ~new_n9685_;
  assign new_n29200_ = ~new_n9692_;
  assign new_n29201_ = ~new_n9684_;
  assign new_n29202_ = ~new_n9691_;
  assign new_n29203_ = ~new_n9683_;
  assign new_n29204_ = ~new_n29401_ | ~new_n29400_;
  assign new_n29205_ = ~new_n29308_ | ~new_n29307_;
  assign new_n29206_ = ~new_n29310_ | ~new_n29309_;
  assign new_n29207_ = ~new_n29317_ | ~new_n29316_;
  assign new_n29208_ = ~new_n29324_ | ~new_n29323_;
  assign new_n29209_ = ~new_n29331_ | ~new_n29330_;
  assign new_n29210_ = ~new_n29338_ | ~new_n29337_;
  assign new_n29211_ = ~new_n29345_ | ~new_n29344_;
  assign new_n29212_ = ~new_n29347_ | ~new_n29346_;
  assign new_n29213_ = ~new_n29354_ | ~new_n29353_;
  assign new_n29214_ = ~new_n29356_ | ~new_n29355_;
  assign new_n29215_ = ~new_n29358_ | ~new_n29357_;
  assign new_n29216_ = ~new_n29360_ | ~new_n29359_;
  assign new_n29217_ = ~new_n29362_ | ~new_n29361_;
  assign new_n29218_ = ~new_n29364_ | ~new_n29363_;
  assign new_n29219_ = ~new_n29366_ | ~new_n29365_;
  assign new_n29220_ = ~new_n29368_ | ~new_n29367_;
  assign new_n29221_ = ~new_n29370_ | ~new_n29369_;
  assign new_n29222_ = ~new_n29372_ | ~new_n29371_;
  assign new_n29223_ = ~new_n29374_ | ~new_n29373_;
  assign new_n29224_ = ~new_n29381_ | ~new_n29380_;
  assign new_n29225_ = ~new_n29383_ | ~new_n29382_;
  assign new_n29226_ = ~new_n29385_ | ~new_n29384_;
  assign new_n29227_ = ~new_n29387_ | ~new_n29386_;
  assign new_n29228_ = ~new_n29389_ | ~new_n29388_;
  assign new_n29229_ = ~new_n29391_ | ~new_n29390_;
  assign new_n29230_ = ~new_n29393_ | ~new_n29392_;
  assign new_n29231_ = ~new_n29395_ | ~new_n29394_;
  assign new_n29232_ = ~new_n29397_ | ~new_n29396_;
  assign new_n29233_ = ~new_n29399_ | ~new_n29398_;
  assign new_n29234_ = new_n9660_ & new_n9659_;
  assign new_n29235_ = ~new_n29278_ | ~new_n29277_;
  assign new_n29236_ = new_n29312_ & new_n29311_;
  assign new_n29237_ = ~new_n29274_ | ~new_n29273_;
  assign new_n29238_ = new_n29319_ & new_n29318_;
  assign new_n29239_ = ~new_n29270_ | ~new_n29269_;
  assign new_n29240_ = new_n29326_ & new_n29325_;
  assign new_n29241_ = ~new_n29266_ | ~new_n29265_;
  assign new_n29242_ = new_n29333_ & new_n29332_;
  assign new_n29243_ = ~new_n29262_ | ~new_n29261_;
  assign new_n29244_ = new_n29340_ & new_n29339_;
  assign new_n29245_ = ~new_n29258_ | ~new_n29257_;
  assign new_n29246_ = new_n29349_ & new_n29348_;
  assign new_n29247_ = ~new_n29249_ | ~new_n29254_;
  assign new_n29248_ = ~new_n9690_ | ~new_n9698_;
  assign new_n29249_ = ~new_n9697_ | ~new_n9690_ | ~new_n9698_;
  assign new_n29250_ = new_n29379_ & new_n29378_;
  assign new_n29251_ = ~new_n29249_;
  assign new_n29252_ = ~new_n9690_ | ~new_n9698_;
  assign new_n29253_ = ~new_n29191_ | ~new_n29252_;
  assign new_n29254_ = ~new_n9689_ | ~new_n29253_;
  assign new_n29255_ = ~new_n29247_;
  assign new_n29256_ = new_n9696_ | new_n9688_;
  assign new_n29257_ = ~new_n29256_ | ~new_n29247_;
  assign new_n29258_ = ~new_n9688_ | ~new_n9696_;
  assign new_n29259_ = ~new_n29245_;
  assign new_n29260_ = new_n9695_ | new_n9687_;
  assign new_n29261_ = ~new_n29260_ | ~new_n29245_;
  assign new_n29262_ = ~new_n9687_ | ~new_n9695_;
  assign new_n29263_ = ~new_n29243_;
  assign new_n29264_ = new_n9694_ | new_n9686_;
  assign new_n29265_ = ~new_n29264_ | ~new_n29243_;
  assign new_n29266_ = ~new_n9686_ | ~new_n9694_;
  assign new_n29267_ = ~new_n29241_;
  assign new_n29268_ = new_n9693_ | new_n9685_;
  assign new_n29269_ = ~new_n29268_ | ~new_n29241_;
  assign new_n29270_ = ~new_n9685_ | ~new_n9693_;
  assign new_n29271_ = ~new_n29239_;
  assign new_n29272_ = new_n9692_ | new_n9684_;
  assign new_n29273_ = ~new_n29272_ | ~new_n29239_;
  assign new_n29274_ = ~new_n9684_ | ~new_n9692_;
  assign new_n29275_ = ~new_n29237_;
  assign new_n29276_ = new_n9691_ | new_n9683_;
  assign new_n29277_ = ~new_n29276_ | ~new_n29237_;
  assign new_n29278_ = ~new_n9683_ | ~new_n9691_;
  assign new_n29279_ = ~new_n29235_;
  assign new_n29280_ = ~new_n29159_;
  assign new_n29281_ = ~new_n29140_;
  assign new_n29282_ = ~new_n29160_;
  assign new_n29283_ = ~new_n29155_;
  assign new_n29284_ = ~new_n29156_;
  assign new_n29285_ = ~new_n29157_;
  assign new_n29286_ = ~new_n29153_;
  assign new_n29287_ = ~new_n29154_;
  assign new_n29288_ = ~new_n29141_;
  assign new_n29289_ = ~new_n29161_;
  assign new_n29290_ = ~new_n29142_;
  assign new_n29291_ = ~new_n29152_;
  assign new_n29292_ = ~new_n29143_;
  assign new_n29293_ = ~new_n29144_;
  assign new_n29294_ = ~new_n29145_;
  assign new_n29295_ = ~new_n29146_;
  assign new_n29296_ = ~new_n29147_;
  assign new_n29297_ = ~new_n29148_;
  assign new_n29298_ = ~new_n29151_;
  assign new_n29299_ = ~new_n29149_;
  assign new_n29300_ = ~new_n29150_;
  assign new_n29301_ = ~new_n29158_;
  assign new_n29302_ = ~new_n9660_ | ~new_n29158_;
  assign new_n29303_ = ~new_n29165_ | ~new_n29302_;
  assign new_n29304_ = ~new_n29234_ | ~new_n29158_;
  assign new_n29305_ = ~new_n29248_;
  assign new_n29306_ = ~new_n29377_ | ~new_n29191_;
  assign new_n29307_ = ~new_n29164_ | ~new_n29159_;
  assign new_n29308_ = ~new_n29280_ | ~new_n9681_;
  assign new_n29309_ = ~new_n29173_ | ~new_n29235_;
  assign new_n29310_ = ~new_n29279_ | ~new_n9682_;
  assign new_n29311_ = ~new_n9683_ | ~new_n29202_;
  assign new_n29312_ = ~new_n9691_ | ~new_n29203_;
  assign new_n29313_ = ~new_n9683_ | ~new_n29202_;
  assign new_n29314_ = ~new_n9691_ | ~new_n29203_;
  assign new_n29315_ = ~new_n29314_ | ~new_n29313_;
  assign new_n29316_ = ~new_n29236_ | ~new_n29237_;
  assign new_n29317_ = ~new_n29275_ | ~new_n29315_;
  assign new_n29318_ = ~new_n9684_ | ~new_n29200_;
  assign new_n29319_ = ~new_n9692_ | ~new_n29201_;
  assign new_n29320_ = ~new_n9684_ | ~new_n29200_;
  assign new_n29321_ = ~new_n9692_ | ~new_n29201_;
  assign new_n29322_ = ~new_n29321_ | ~new_n29320_;
  assign new_n29323_ = ~new_n29238_ | ~new_n29239_;
  assign new_n29324_ = ~new_n29271_ | ~new_n29322_;
  assign new_n29325_ = ~new_n9685_ | ~new_n29198_;
  assign new_n29326_ = ~new_n9693_ | ~new_n29199_;
  assign new_n29327_ = ~new_n9685_ | ~new_n29198_;
  assign new_n29328_ = ~new_n9693_ | ~new_n29199_;
  assign new_n29329_ = ~new_n29328_ | ~new_n29327_;
  assign new_n29330_ = ~new_n29240_ | ~new_n29241_;
  assign new_n29331_ = ~new_n29267_ | ~new_n29329_;
  assign new_n29332_ = ~new_n9686_ | ~new_n29196_;
  assign new_n29333_ = ~new_n9694_ | ~new_n29197_;
  assign new_n29334_ = ~new_n9686_ | ~new_n29196_;
  assign new_n29335_ = ~new_n9694_ | ~new_n29197_;
  assign new_n29336_ = ~new_n29335_ | ~new_n29334_;
  assign new_n29337_ = ~new_n29242_ | ~new_n29243_;
  assign new_n29338_ = ~new_n29263_ | ~new_n29336_;
  assign new_n29339_ = ~new_n9687_ | ~new_n29194_;
  assign new_n29340_ = ~new_n9695_ | ~new_n29195_;
  assign new_n29341_ = ~new_n9687_ | ~new_n29194_;
  assign new_n29342_ = ~new_n9695_ | ~new_n29195_;
  assign new_n29343_ = ~new_n29342_ | ~new_n29341_;
  assign new_n29344_ = ~new_n29244_ | ~new_n29245_;
  assign new_n29345_ = ~new_n29259_ | ~new_n29343_;
  assign new_n29346_ = ~new_n29166_ | ~new_n29158_;
  assign new_n29347_ = ~new_n9660_ | ~new_n29301_;
  assign new_n29348_ = ~new_n9688_ | ~new_n29192_;
  assign new_n29349_ = ~new_n9696_ | ~new_n29193_;
  assign new_n29350_ = ~new_n9688_ | ~new_n29192_;
  assign new_n29351_ = ~new_n9696_ | ~new_n29193_;
  assign new_n29352_ = ~new_n29351_ | ~new_n29350_;
  assign new_n29353_ = ~new_n29246_ | ~new_n29247_;
  assign new_n29354_ = ~new_n29255_ | ~new_n29352_;
  assign new_n29355_ = ~new_n29176_ | ~new_n29150_;
  assign new_n29356_ = ~new_n29300_ | ~new_n9661_;
  assign new_n29357_ = ~new_n29177_ | ~new_n29149_;
  assign new_n29358_ = ~new_n29299_ | ~new_n9662_;
  assign new_n29359_ = ~new_n29174_ | ~new_n29151_;
  assign new_n29360_ = ~new_n29298_ | ~new_n9663_;
  assign new_n29361_ = ~new_n29178_ | ~new_n29148_;
  assign new_n29362_ = ~new_n29297_ | ~new_n9664_;
  assign new_n29363_ = ~new_n29179_ | ~new_n29147_;
  assign new_n29364_ = ~new_n29296_ | ~new_n9665_;
  assign new_n29365_ = ~new_n29180_ | ~new_n29146_;
  assign new_n29366_ = ~new_n29295_ | ~new_n9666_;
  assign new_n29367_ = ~new_n29181_ | ~new_n29145_;
  assign new_n29368_ = ~new_n29294_ | ~new_n9667_;
  assign new_n29369_ = ~new_n29175_ | ~new_n29144_;
  assign new_n29370_ = ~new_n29293_ | ~new_n9668_;
  assign new_n29371_ = ~new_n29182_ | ~new_n29143_;
  assign new_n29372_ = ~new_n29292_ | ~new_n9669_;
  assign new_n29373_ = ~new_n29172_ | ~new_n29152_;
  assign new_n29374_ = ~new_n29291_ | ~new_n9670_;
  assign new_n29375_ = ~new_n9689_ | ~new_n29248_;
  assign new_n29376_ = ~new_n29305_ | ~new_n29190_;
  assign new_n29377_ = ~new_n29376_ | ~new_n29375_;
  assign new_n29378_ = ~new_n29190_ | ~new_n9697_ | ~new_n29252_;
  assign new_n29379_ = ~new_n29251_ | ~new_n9689_;
  assign new_n29380_ = ~new_n29183_ | ~new_n29142_;
  assign new_n29381_ = ~new_n29290_ | ~new_n9671_;
  assign new_n29382_ = ~new_n29162_ | ~new_n29161_;
  assign new_n29383_ = ~new_n29289_ | ~new_n9672_;
  assign new_n29384_ = ~new_n29184_ | ~new_n29141_;
  assign new_n29385_ = ~new_n29288_ | ~new_n9673_;
  assign new_n29386_ = ~new_n29170_ | ~new_n29154_;
  assign new_n29387_ = ~new_n29287_ | ~new_n9674_;
  assign new_n29388_ = ~new_n29171_ | ~new_n29153_;
  assign new_n29389_ = ~new_n29286_ | ~new_n9675_;
  assign new_n29390_ = ~new_n29167_ | ~new_n29157_;
  assign new_n29391_ = ~new_n29285_ | ~new_n9676_;
  assign new_n29392_ = ~new_n29168_ | ~new_n29156_;
  assign new_n29393_ = ~new_n29284_ | ~new_n9677_;
  assign new_n29394_ = ~new_n29169_ | ~new_n29155_;
  assign new_n29395_ = ~new_n29283_ | ~new_n9678_;
  assign new_n29396_ = ~new_n29163_ | ~new_n29160_;
  assign new_n29397_ = ~new_n29282_ | ~new_n9679_;
  assign new_n29398_ = ~new_n29185_ | ~new_n29140_;
  assign new_n29399_ = ~new_n29281_ | ~new_n9680_;
  assign new_n29400_ = ~new_n9690_ | ~new_n29188_;
  assign new_n29401_ = ~new_n9698_ | ~new_n29189_;
  assign new_n29402_ = ~new_n29038_ & ~new_n29404_;
  assign new_n29403_ = new_n29042_ & new_n29405_;
  assign new_n29404_ = ~new_n29040_ & ~new_n29039_ & ~new_n29403_ & ~new_n29041_;
  assign new_n29405_ = new_n29021_ | new_n29043_;
  assign new_n29406_ = new_n29427_ & new_n29426_;
  assign new_n29407_ = ~new_n10661_;
  assign new_n29408_ = ~pi0764;
  assign new_n29409_ = ~pi0763;
  assign new_n29410_ = ~new_n10660_;
  assign new_n29411_ = ~new_n10659_;
  assign new_n29412_ = ~pi0762;
  assign new_n29413_ = ~pi0761;
  assign new_n29414_ = ~new_n10658_;
  assign new_n29415_ = ~new_n10662_;
  assign new_n29416_ = ~new_n10661_ | ~new_n29408_;
  assign new_n29417_ = ~new_n29416_ | ~pi0765 | ~new_n29415_;
  assign new_n29418_ = ~pi0764 | ~new_n29407_;
  assign new_n29419_ = ~pi0763 | ~new_n29410_;
  assign new_n29420_ = ~new_n29417_ | ~new_n29418_ | ~new_n29419_;
  assign new_n29421_ = ~new_n10660_ | ~new_n29409_;
  assign new_n29422_ = ~new_n10659_ | ~new_n29412_;
  assign new_n29423_ = ~new_n29420_ | ~new_n29421_ | ~new_n29422_;
  assign new_n29424_ = ~pi0762 | ~new_n29411_;
  assign new_n29425_ = ~pi0761 | ~new_n29414_;
  assign new_n29426_ = ~new_n29423_ | ~new_n29424_ | ~new_n29425_;
  assign new_n29427_ = ~new_n10658_ | ~new_n29413_;
  assign new_n29428_ = ~new_n29455_ | ~new_n29470_;
  assign new_n29429_ = new_n29447_ & new_n29467_;
  assign new_n29430_ = ~new_n10670_;
  assign new_n29431_ = ~new_n10669_;
  assign new_n29432_ = ~new_n10668_;
  assign new_n29433_ = ~new_n10667_;
  assign new_n29434_ = ~new_n10667_ | ~new_n29449_;
  assign new_n29435_ = ~new_n10666_;
  assign new_n29436_ = ~new_n10666_ | ~new_n29465_;
  assign new_n29437_ = ~new_n10665_;
  assign new_n29438_ = ~new_n10665_ | ~new_n29466_;
  assign new_n29439_ = ~new_n10663_;
  assign new_n29440_ = ~new_n10664_;
  assign new_n29441_ = ~new_n29472_ | ~new_n29471_;
  assign new_n29442_ = ~new_n29474_ | ~new_n29473_;
  assign new_n29443_ = ~new_n29476_ | ~new_n29475_;
  assign new_n29444_ = ~new_n29478_ | ~new_n29477_;
  assign new_n29445_ = ~new_n29494_ | ~new_n29493_;
  assign new_n29446_ = ~new_n29487_ | ~new_n29486_;
  assign new_n29447_ = new_n10663_ & new_n10664_;
  assign new_n29448_ = ~new_n10664_ | ~new_n29467_;
  assign new_n29449_ = ~new_n29463_ | ~new_n29462_;
  assign new_n29450_ = new_n29480_ & new_n29479_;
  assign new_n29451_ = new_n29482_ & new_n29481_;
  assign new_n29452_ = ~new_n29454_ | ~new_n29459_;
  assign new_n29453_ = ~new_n14914_ | ~new_n10670_;
  assign new_n29454_ = ~new_n10669_ | ~new_n14914_ | ~new_n10670_;
  assign new_n29455_ = new_n29492_ & new_n29491_;
  assign new_n29456_ = ~new_n29454_;
  assign new_n29457_ = ~new_n14914_ | ~new_n10670_;
  assign new_n29458_ = ~new_n29431_ | ~new_n29457_;
  assign new_n29459_ = ~new_n9657_ | ~new_n29458_;
  assign new_n29460_ = ~new_n29452_;
  assign new_n29461_ = new_n10668_ | new_n14914_;
  assign new_n29462_ = ~new_n29461_ | ~new_n29452_;
  assign new_n29463_ = ~new_n14914_ | ~new_n10668_;
  assign new_n29464_ = ~new_n29449_;
  assign new_n29465_ = ~new_n29434_;
  assign new_n29466_ = ~new_n29436_;
  assign new_n29467_ = ~new_n29438_;
  assign new_n29468_ = ~new_n29448_;
  assign new_n29469_ = ~new_n29453_;
  assign new_n29470_ = ~new_n29490_ | ~new_n29431_;
  assign new_n29471_ = ~new_n10663_ | ~new_n29448_;
  assign new_n29472_ = ~new_n29468_ | ~new_n29439_;
  assign new_n29473_ = ~new_n10664_ | ~new_n29438_;
  assign new_n29474_ = ~new_n29467_ | ~new_n29440_;
  assign new_n29475_ = ~new_n10665_ | ~new_n29436_;
  assign new_n29476_ = ~new_n29466_ | ~new_n29437_;
  assign new_n29477_ = ~new_n10666_ | ~new_n29434_;
  assign new_n29478_ = ~new_n29465_ | ~new_n29435_;
  assign new_n29479_ = ~new_n10667_ | ~new_n29449_;
  assign new_n29480_ = ~new_n29464_ | ~new_n29433_;
  assign new_n29481_ = ~new_n14914_ | ~new_n29432_;
  assign new_n29482_ = ~new_n10668_ | ~new_n9657_;
  assign new_n29483_ = ~new_n14914_ | ~new_n29432_;
  assign new_n29484_ = ~new_n10668_ | ~new_n9657_;
  assign new_n29485_ = ~new_n29484_ | ~new_n29483_;
  assign new_n29486_ = ~new_n29451_ | ~new_n29452_;
  assign new_n29487_ = ~new_n29460_ | ~new_n29485_;
  assign new_n29488_ = ~new_n9657_ | ~new_n29453_;
  assign new_n29489_ = ~new_n29469_ | ~new_n14914_;
  assign new_n29490_ = ~new_n29489_ | ~new_n29488_;
  assign new_n29491_ = ~new_n14914_ | ~new_n10669_ | ~new_n29457_;
  assign new_n29492_ = ~new_n29456_ | ~new_n9657_;
  assign new_n29493_ = ~new_n14914_ | ~new_n29430_;
  assign new_n29494_ = ~new_n10670_ | ~new_n9657_;
  assign new_n29495_ = ~new_n29534_ | ~new_n29533_;
  assign new_n29496_ = ~new_n29498_ | ~new_n29535_;
  assign new_n29497_ = ~pi0760;
  assign new_n29498_ = ~pi0760 | ~new_n29507_;
  assign new_n29499_ = ~pi0764;
  assign new_n29500_ = ~pi0758;
  assign new_n29501_ = ~pi0763;
  assign new_n29502_ = ~pi0757;
  assign new_n29503_ = ~pi0762;
  assign new_n29504_ = ~pi0761;
  assign new_n29505_ = ~new_n29530_ | ~new_n29529_;
  assign new_n29506_ = ~pi0756;
  assign new_n29507_ = ~pi0765;
  assign new_n29508_ = ~new_n29540_ | ~new_n29539_;
  assign new_n29509_ = ~new_n29545_ | ~new_n29544_;
  assign new_n29510_ = ~new_n29550_ | ~new_n29549_;
  assign new_n29511_ = ~new_n29555_ | ~new_n29554_;
  assign new_n29512_ = ~new_n29537_ | ~new_n29536_;
  assign new_n29513_ = ~new_n29542_ | ~new_n29541_;
  assign new_n29514_ = ~new_n29547_ | ~new_n29546_;
  assign new_n29515_ = ~new_n29552_ | ~new_n29551_;
  assign new_n29516_ = ~new_n29526_ | ~new_n29525_;
  assign new_n29517_ = ~new_n29522_ | ~new_n29521_;
  assign new_n29518_ = ~pi0759;
  assign new_n29519_ = ~new_n29498_;
  assign new_n29520_ = ~new_n29519_ | ~new_n29499_;
  assign new_n29521_ = ~new_n29520_ | ~new_n29518_;
  assign new_n29522_ = ~pi0764 | ~new_n29498_;
  assign new_n29523_ = ~new_n29517_;
  assign new_n29524_ = ~pi0758 | ~new_n29501_;
  assign new_n29525_ = ~new_n29524_ | ~new_n29517_;
  assign new_n29526_ = ~pi0763 | ~new_n29500_;
  assign new_n29527_ = ~new_n29516_;
  assign new_n29528_ = ~pi0757 | ~new_n29503_;
  assign new_n29529_ = ~new_n29528_ | ~new_n29516_;
  assign new_n29530_ = ~pi0762 | ~new_n29502_;
  assign new_n29531_ = ~new_n29505_;
  assign new_n29532_ = ~pi0761 | ~new_n29506_;
  assign new_n29533_ = ~new_n29531_ | ~new_n29532_;
  assign new_n29534_ = ~pi0756 | ~new_n29504_;
  assign new_n29535_ = ~pi0765 | ~new_n29497_;
  assign new_n29536_ = ~pi0756 | ~new_n29504_;
  assign new_n29537_ = ~pi0761 | ~new_n29506_;
  assign new_n29538_ = ~new_n29512_;
  assign new_n29539_ = ~new_n29538_ | ~new_n29531_;
  assign new_n29540_ = ~new_n29512_ | ~new_n29505_;
  assign new_n29541_ = ~pi0757 | ~new_n29503_;
  assign new_n29542_ = ~pi0762 | ~new_n29502_;
  assign new_n29543_ = ~new_n29513_;
  assign new_n29544_ = ~new_n29527_ | ~new_n29543_;
  assign new_n29545_ = ~new_n29513_ | ~new_n29516_;
  assign new_n29546_ = ~pi0758 | ~new_n29501_;
  assign new_n29547_ = ~pi0763 | ~new_n29500_;
  assign new_n29548_ = ~new_n29514_;
  assign new_n29549_ = ~new_n29523_ | ~new_n29548_;
  assign new_n29550_ = ~new_n29514_ | ~new_n29517_;
  assign new_n29551_ = ~pi0759 | ~new_n29499_;
  assign new_n29552_ = ~pi0764 | ~new_n29518_;
  assign new_n29553_ = ~new_n29515_;
  assign new_n29554_ = ~new_n29553_ | ~new_n29519_;
  assign new_n29555_ = ~new_n29515_ | ~new_n29498_;
  assign new_n29556_ = new_n29676_ & new_n29577_;
  assign new_n29557_ = new_n29674_ & new_n29578_;
  assign new_n29558_ = new_n29672_ & new_n29579_;
  assign new_n29559_ = new_n29670_ & new_n29580_;
  assign new_n29560_ = new_n29668_ & new_n29581_;
  assign new_n29561_ = new_n29666_ & new_n29582_;
  assign new_n29562_ = new_n29664_ & new_n29583_;
  assign new_n29563_ = new_n29662_ & new_n29584_;
  assign new_n29564_ = new_n29660_ & new_n29585_;
  assign new_n29565_ = new_n29658_ & new_n29586_;
  assign new_n29566_ = new_n29656_ & new_n29587_;
  assign new_n29567_ = new_n29655_ & new_n29571_;
  assign new_n29568_ = new_n29642_ & new_n29572_;
  assign new_n29569_ = new_n29640_ & new_n29573_;
  assign new_n29570_ = new_n29638_ & new_n29574_;
  assign new_n29571_ = new_n10724_ | new_n10712_ | new_n10723_;
  assign new_n29572_ = ~new_n29601_ | ~new_n29633_;
  assign new_n29573_ = ~new_n29576_ | ~new_n29634_ | ~new_n29606_;
  assign new_n29574_ = ~new_n29575_ | ~new_n29635_ | ~new_n29604_;
  assign new_n29575_ = ~new_n10695_;
  assign new_n29576_ = ~new_n10697_;
  assign new_n29577_ = ~new_n29598_ | ~new_n29602_ | ~new_n29636_;
  assign new_n29578_ = ~new_n29597_ | ~new_n29643_ | ~new_n29631_;
  assign new_n29579_ = ~new_n29596_ | ~new_n29644_ | ~new_n29629_;
  assign new_n29580_ = ~new_n29595_ | ~new_n29645_ | ~new_n29627_;
  assign new_n29581_ = ~new_n29594_ | ~new_n29646_ | ~new_n29625_;
  assign new_n29582_ = ~new_n29593_ | ~new_n29647_ | ~new_n29623_;
  assign new_n29583_ = ~new_n29592_ | ~new_n29648_ | ~new_n29619_;
  assign new_n29584_ = ~new_n29591_ | ~new_n29649_ | ~new_n29617_;
  assign new_n29585_ = ~new_n29590_ | ~new_n29650_ | ~new_n29615_;
  assign new_n29586_ = ~new_n29589_ | ~new_n29651_ | ~new_n29613_;
  assign new_n29587_ = ~new_n29652_ | ~new_n29588_;
  assign new_n29588_ = ~new_n10702_;
  assign new_n29589_ = ~new_n10703_;
  assign new_n29590_ = ~new_n10705_;
  assign new_n29591_ = ~new_n10707_;
  assign new_n29592_ = ~new_n10709_;
  assign new_n29593_ = ~new_n10711_;
  assign new_n29594_ = ~new_n10714_;
  assign new_n29595_ = ~new_n10716_;
  assign new_n29596_ = ~new_n10718_;
  assign new_n29597_ = ~new_n10720_;
  assign new_n29598_ = ~new_n10722_;
  assign new_n29599_ = ~new_n29699_ | ~new_n29698_;
  assign new_n29600_ = ~new_n29687_ | ~new_n29686_;
  assign new_n29601_ = ~new_n10701_ & ~new_n10699_;
  assign new_n29602_ = ~new_n10694_;
  assign new_n29603_ = new_n29679_ & new_n29678_;
  assign new_n29604_ = ~new_n10696_;
  assign new_n29605_ = new_n29681_ & new_n29680_;
  assign new_n29606_ = ~new_n10698_;
  assign new_n29607_ = new_n29683_ & new_n29682_;
  assign new_n29608_ = ~new_n10701_;
  assign new_n29609_ = new_n29685_ & new_n29684_;
  assign new_n29610_ = ~new_n10688_;
  assign new_n29611_ = ~new_n10700_;
  assign new_n29612_ = new_n29689_ & new_n29688_;
  assign new_n29613_ = ~new_n10704_;
  assign new_n29614_ = new_n29691_ & new_n29690_;
  assign new_n29615_ = ~new_n10706_;
  assign new_n29616_ = new_n29693_ & new_n29692_;
  assign new_n29617_ = ~new_n10708_;
  assign new_n29618_ = new_n29695_ & new_n29694_;
  assign new_n29619_ = ~new_n10710_;
  assign new_n29620_ = new_n29697_ & new_n29696_;
  assign new_n29621_ = ~new_n10723_;
  assign new_n29622_ = ~new_n10724_;
  assign new_n29623_ = ~new_n10713_;
  assign new_n29624_ = new_n29701_ & new_n29700_;
  assign new_n29625_ = ~new_n10715_;
  assign new_n29626_ = new_n29703_ & new_n29702_;
  assign new_n29627_ = ~new_n10717_;
  assign new_n29628_ = new_n29705_ & new_n29704_;
  assign new_n29629_ = ~new_n10719_;
  assign new_n29630_ = new_n29707_ & new_n29706_;
  assign new_n29631_ = ~new_n10721_;
  assign new_n29632_ = new_n29709_ & new_n29708_;
  assign new_n29633_ = ~new_n29571_;
  assign new_n29634_ = ~new_n29572_;
  assign new_n29635_ = ~new_n29573_;
  assign new_n29636_ = ~new_n29574_;
  assign new_n29637_ = ~new_n29635_ | ~new_n29604_;
  assign new_n29638_ = ~new_n10695_ | ~new_n29637_;
  assign new_n29639_ = ~new_n29634_ | ~new_n29606_;
  assign new_n29640_ = ~new_n10697_ | ~new_n29639_;
  assign new_n29641_ = ~new_n29633_ | ~new_n29608_;
  assign new_n29642_ = ~new_n10699_ | ~new_n29641_;
  assign new_n29643_ = ~new_n29577_;
  assign new_n29644_ = ~new_n29578_;
  assign new_n29645_ = ~new_n29579_;
  assign new_n29646_ = ~new_n29580_;
  assign new_n29647_ = ~new_n29581_;
  assign new_n29648_ = ~new_n29582_;
  assign new_n29649_ = ~new_n29583_;
  assign new_n29650_ = ~new_n29584_;
  assign new_n29651_ = ~new_n29585_;
  assign new_n29652_ = ~new_n29586_;
  assign new_n29653_ = ~new_n29587_;
  assign new_n29654_ = new_n10723_ | new_n10724_;
  assign new_n29655_ = ~new_n10712_ | ~new_n29654_;
  assign new_n29656_ = ~new_n10702_ | ~new_n29586_;
  assign new_n29657_ = ~new_n29651_ | ~new_n29613_;
  assign new_n29658_ = ~new_n10703_ | ~new_n29657_;
  assign new_n29659_ = ~new_n29650_ | ~new_n29615_;
  assign new_n29660_ = ~new_n10705_ | ~new_n29659_;
  assign new_n29661_ = ~new_n29649_ | ~new_n29617_;
  assign new_n29662_ = ~new_n10707_ | ~new_n29661_;
  assign new_n29663_ = ~new_n29648_ | ~new_n29619_;
  assign new_n29664_ = ~new_n10709_ | ~new_n29663_;
  assign new_n29665_ = ~new_n29647_ | ~new_n29623_;
  assign new_n29666_ = ~new_n10711_ | ~new_n29665_;
  assign new_n29667_ = ~new_n29646_ | ~new_n29625_;
  assign new_n29668_ = ~new_n10714_ | ~new_n29667_;
  assign new_n29669_ = ~new_n29645_ | ~new_n29627_;
  assign new_n29670_ = ~new_n10716_ | ~new_n29669_;
  assign new_n29671_ = ~new_n29644_ | ~new_n29629_;
  assign new_n29672_ = ~new_n10718_ | ~new_n29671_;
  assign new_n29673_ = ~new_n29643_ | ~new_n29631_;
  assign new_n29674_ = ~new_n10720_ | ~new_n29673_;
  assign new_n29675_ = ~new_n29636_ | ~new_n29602_;
  assign new_n29676_ = ~new_n10722_ | ~new_n29675_;
  assign new_n29677_ = ~new_n29653_ | ~new_n29611_;
  assign new_n29678_ = ~new_n10694_ | ~new_n29574_;
  assign new_n29679_ = ~new_n29636_ | ~new_n29602_;
  assign new_n29680_ = ~new_n10696_ | ~new_n29573_;
  assign new_n29681_ = ~new_n29635_ | ~new_n29604_;
  assign new_n29682_ = ~new_n10698_ | ~new_n29572_;
  assign new_n29683_ = ~new_n29634_ | ~new_n29606_;
  assign new_n29684_ = ~new_n10701_ | ~new_n29571_;
  assign new_n29685_ = ~new_n29633_ | ~new_n29608_;
  assign new_n29686_ = ~new_n29677_ | ~new_n29610_;
  assign new_n29687_ = ~new_n10688_ | ~new_n29653_ | ~new_n29611_;
  assign new_n29688_ = ~new_n10700_ | ~new_n29587_;
  assign new_n29689_ = ~new_n29653_ | ~new_n29611_;
  assign new_n29690_ = ~new_n10704_ | ~new_n29585_;
  assign new_n29691_ = ~new_n29651_ | ~new_n29613_;
  assign new_n29692_ = ~new_n10706_ | ~new_n29584_;
  assign new_n29693_ = ~new_n29650_ | ~new_n29615_;
  assign new_n29694_ = ~new_n10708_ | ~new_n29583_;
  assign new_n29695_ = ~new_n29649_ | ~new_n29617_;
  assign new_n29696_ = ~new_n10710_ | ~new_n29582_;
  assign new_n29697_ = ~new_n29648_ | ~new_n29619_;
  assign new_n29698_ = ~new_n10723_ | ~new_n29622_;
  assign new_n29699_ = ~new_n10724_ | ~new_n29621_;
  assign new_n29700_ = ~new_n10713_ | ~new_n29581_;
  assign new_n29701_ = ~new_n29647_ | ~new_n29623_;
  assign new_n29702_ = ~new_n10715_ | ~new_n29580_;
  assign new_n29703_ = ~new_n29646_ | ~new_n29625_;
  assign new_n29704_ = ~new_n10717_ | ~new_n29579_;
  assign new_n29705_ = ~new_n29645_ | ~new_n29627_;
  assign new_n29706_ = ~new_n10719_ | ~new_n29578_;
  assign new_n29707_ = ~new_n29644_ | ~new_n29629_;
  assign new_n29708_ = ~new_n10721_ | ~new_n29577_;
  assign new_n29709_ = ~new_n29643_ | ~new_n29631_;
  assign new_n29710_ = new_n30105_ & new_n30104_;
  assign new_n29711_ = new_n29912_ & new_n29867_ & new_n30015_;
  assign new_n29712_ = ~new_n30051_ | ~new_n30196_ | ~new_n30195_;
  assign new_n29713_ = ~new_n10672_;
  assign new_n29714_ = ~pi0773;
  assign new_n29715_ = ~new_n10674_;
  assign new_n29716_ = ~pi0771;
  assign new_n29717_ = ~new_n10676_;
  assign new_n29718_ = ~pi0769;
  assign new_n29719_ = ~new_n10679_;
  assign new_n29720_ = ~pi0766;
  assign new_n29721_ = ~pi0766 | ~new_n10679_;
  assign new_n29722_ = ~new_n10678_;
  assign new_n29723_ = ~pi0767;
  assign new_n29724_ = ~new_n10677_;
  assign new_n29725_ = ~pi0768;
  assign new_n29726_ = ~pi0768 | ~new_n10677_;
  assign new_n29727_ = ~new_n10675_;
  assign new_n29728_ = ~pi0770;
  assign new_n29729_ = ~pi0770 | ~new_n10675_;
  assign new_n29730_ = ~new_n10673_;
  assign new_n29731_ = ~pi0772;
  assign new_n29732_ = ~pi0772 | ~new_n10673_;
  assign new_n29733_ = ~new_n10671_;
  assign new_n29734_ = ~pi0774;
  assign new_n29735_ = ~pi0775;
  assign new_n29736_ = ~new_n9853_;
  assign new_n29737_ = ~new_n9834_;
  assign new_n29738_ = ~pi0794;
  assign new_n29739_ = ~new_n9833_;
  assign new_n29740_ = ~pi0795;
  assign new_n29741_ = ~new_n9838_;
  assign new_n29742_ = ~pi0790;
  assign new_n29743_ = ~new_n9840_;
  assign new_n29744_ = ~pi0788;
  assign new_n29745_ = ~new_n9842_;
  assign new_n29746_ = ~pi0786;
  assign new_n29747_ = ~new_n9845_;
  assign new_n29748_ = ~pi0783;
  assign new_n29749_ = ~new_n9847_;
  assign new_n29750_ = ~pi0781;
  assign new_n29751_ = ~new_n9849_;
  assign new_n29752_ = ~pi0779;
  assign new_n29753_ = ~new_n9851_;
  assign new_n29754_ = ~pi0777;
  assign new_n29755_ = ~pi0774 | ~new_n10671_;
  assign new_n29756_ = ~new_n9852_;
  assign new_n29757_ = ~pi0776;
  assign new_n29758_ = ~pi0776 | ~new_n9852_;
  assign new_n29759_ = ~new_n9850_;
  assign new_n29760_ = ~pi0778;
  assign new_n29761_ = ~pi0778 | ~new_n9850_;
  assign new_n29762_ = ~new_n9848_;
  assign new_n29763_ = ~pi0780;
  assign new_n29764_ = ~pi0780 | ~new_n9848_;
  assign new_n29765_ = ~new_n9846_;
  assign new_n29766_ = ~pi0782;
  assign new_n29767_ = ~pi0782 | ~new_n9846_;
  assign new_n29768_ = ~new_n9843_;
  assign new_n29769_ = ~pi0785;
  assign new_n29770_ = ~new_n9844_;
  assign new_n29771_ = ~pi0784;
  assign new_n29772_ = ~new_n9841_;
  assign new_n29773_ = ~pi0787;
  assign new_n29774_ = ~pi0787 | ~new_n9841_;
  assign new_n29775_ = ~new_n9839_;
  assign new_n29776_ = ~pi0789;
  assign new_n29777_ = ~pi0789 | ~new_n9839_;
  assign new_n29778_ = ~new_n9837_;
  assign new_n29779_ = ~pi0791;
  assign new_n29780_ = ~new_n9835_;
  assign new_n29781_ = ~pi0793;
  assign new_n29782_ = ~new_n9836_;
  assign new_n29783_ = ~pi0792;
  assign new_n29784_ = ~pi0792 | ~new_n9836_;
  assign new_n29785_ = ~new_n9832_;
  assign new_n29786_ = ~pi0796;
  assign new_n29787_ = ~new_n30046_ | ~new_n30003_;
  assign new_n29788_ = ~new_n10678_ | ~new_n29914_;
  assign new_n29789_ = ~new_n30268_ | ~new_n30267_;
  assign new_n29790_ = ~new_n30058_ | ~new_n30057_;
  assign new_n29791_ = ~new_n30065_ | ~new_n30064_;
  assign new_n29792_ = ~new_n30072_ | ~new_n30071_;
  assign new_n29793_ = ~new_n30079_ | ~new_n30078_;
  assign new_n29794_ = ~new_n30086_ | ~new_n30085_;
  assign new_n29795_ = ~new_n30093_ | ~new_n30092_;
  assign new_n29796_ = ~new_n30100_ | ~new_n30099_;
  assign new_n29797_ = ~new_n30114_ | ~new_n30113_;
  assign new_n29798_ = ~new_n30121_ | ~new_n30120_;
  assign new_n29799_ = ~new_n30128_ | ~new_n30127_;
  assign new_n29800_ = ~new_n30135_ | ~new_n30134_;
  assign new_n29801_ = ~new_n30142_ | ~new_n30141_;
  assign new_n29802_ = ~new_n30149_ | ~new_n30148_;
  assign new_n29803_ = ~new_n30156_ | ~new_n30155_;
  assign new_n29804_ = ~new_n30163_ | ~new_n30162_;
  assign new_n29805_ = ~new_n30170_ | ~new_n30169_;
  assign new_n29806_ = ~new_n30177_ | ~new_n30176_;
  assign new_n29807_ = ~new_n30184_ | ~new_n30183_;
  assign new_n29808_ = ~new_n30191_ | ~new_n30190_;
  assign new_n29809_ = ~new_n30203_ | ~new_n30202_;
  assign new_n29810_ = ~new_n30210_ | ~new_n30209_;
  assign new_n29811_ = ~new_n30217_ | ~new_n30216_;
  assign new_n29812_ = ~new_n30224_ | ~new_n30223_;
  assign new_n29813_ = ~new_n30231_ | ~new_n30230_;
  assign new_n29814_ = ~new_n30238_ | ~new_n30237_;
  assign new_n29815_ = ~new_n30245_ | ~new_n30244_;
  assign new_n29816_ = ~new_n30252_ | ~new_n30251_;
  assign new_n29817_ = ~new_n30259_ | ~new_n30258_;
  assign new_n29818_ = ~new_n30266_ | ~new_n30265_;
  assign new_n29819_ = new_n29916_ & new_n30020_;
  assign new_n29820_ = new_n30019_ & new_n29921_;
  assign new_n29821_ = new_n29923_ & new_n29927_;
  assign new_n29822_ = new_n30022_ & new_n29928_;
  assign new_n29823_ = new_n29930_ & new_n29934_;
  assign new_n29824_ = new_n30024_ & new_n29935_;
  assign new_n29825_ = new_n29937_ & new_n29941_;
  assign new_n29826_ = new_n30026_ & new_n29942_;
  assign new_n29827_ = new_n29944_ & new_n29948_;
  assign new_n29828_ = new_n30028_ & new_n29949_;
  assign new_n29829_ = new_n29951_ & new_n29955_;
  assign new_n29830_ = new_n30030_ & new_n29956_;
  assign new_n29831_ = new_n29958_ & new_n29962_;
  assign new_n29832_ = new_n30032_ & new_n29963_;
  assign new_n29833_ = new_n29965_ & new_n29969_;
  assign new_n29834_ = new_n30034_ & new_n29970_;
  assign new_n29835_ = new_n29979_ & new_n29976_;
  assign new_n29836_ = new_n30037_ & new_n29979_;
  assign new_n29837_ = new_n30040_ & new_n29980_;
  assign new_n29838_ = new_n29982_ & new_n29986_;
  assign new_n29839_ = new_n30042_ & new_n29987_;
  assign new_n29840_ = new_n29989_ & new_n29993_;
  assign new_n29841_ = new_n30044_ & new_n29994_;
  assign new_n29842_ = new_n29998_ & new_n30005_ & new_n30002_;
  assign new_n29843_ = new_n30010_ & new_n30006_;
  assign new_n29844_ = new_n30013_ & new_n30008_;
  assign new_n29845_ = new_n30103_ & new_n29844_;
  assign new_n29846_ = new_n30049_ & new_n30006_;
  assign new_n29847_ = new_n29710_ & new_n29848_;
  assign new_n29848_ = new_n30010_ & new_n30012_;
  assign new_n29849_ = new_n29998_ & new_n30002_;
  assign new_n29850_ = new_n29972_ & new_n29976_;
  assign new_n29851_ = new_n30053_ & new_n30052_;
  assign new_n29852_ = ~new_n29755_ | ~new_n29938_;
  assign new_n29853_ = new_n30060_ & new_n30059_;
  assign new_n29854_ = ~new_n29824_ | ~new_n30023_;
  assign new_n29855_ = new_n30067_ & new_n30066_;
  assign new_n29856_ = ~new_n29732_ | ~new_n29931_;
  assign new_n29857_ = new_n30074_ & new_n30073_;
  assign new_n29858_ = ~new_n29822_ | ~new_n30021_;
  assign new_n29859_ = new_n30081_ & new_n30080_;
  assign new_n29860_ = ~new_n29729_ | ~new_n29924_;
  assign new_n29861_ = new_n30088_ & new_n30087_;
  assign new_n29862_ = ~new_n29820_ | ~new_n30018_;
  assign new_n29863_ = new_n30095_ & new_n30094_;
  assign new_n29864_ = ~new_n29726_ | ~new_n29917_;
  assign new_n29865_ = ~pi0797;
  assign new_n29866_ = ~new_n9831_;
  assign new_n29867_ = new_n30107_ & new_n30106_;
  assign new_n29868_ = new_n30109_ & new_n30108_;
  assign new_n29869_ = ~new_n30010_ | ~new_n30009_;
  assign new_n29870_ = new_n30116_ & new_n30115_;
  assign new_n29871_ = ~new_n30017_ | ~new_n30016_ | ~new_n29788_;
  assign new_n29872_ = new_n30123_ & new_n30122_;
  assign new_n29873_ = ~new_n29846_ | ~new_n30048_;
  assign new_n29874_ = new_n30130_ & new_n30129_;
  assign new_n29875_ = ~new_n30047_ | ~new_n30045_;
  assign new_n29876_ = new_n30137_ & new_n30136_;
  assign new_n29877_ = ~new_n29784_ | ~new_n29999_;
  assign new_n29878_ = new_n30144_ & new_n30143_;
  assign new_n29879_ = ~new_n30014_ | ~new_n29996_ | ~new_n29911_;
  assign new_n29880_ = ~new_n29841_ | ~new_n30043_;
  assign new_n29881_ = new_n30158_ & new_n30157_;
  assign new_n29882_ = ~new_n29777_ | ~new_n29990_;
  assign new_n29883_ = new_n30165_ & new_n30164_;
  assign new_n29884_ = ~new_n29839_ | ~new_n30041_;
  assign new_n29885_ = new_n30172_ & new_n30171_;
  assign new_n29886_ = ~new_n29774_ | ~new_n29983_;
  assign new_n29887_ = new_n30179_ & new_n30178_;
  assign new_n29888_ = ~new_n29837_ | ~new_n30039_;
  assign new_n29889_ = new_n30186_ & new_n30185_;
  assign new_n29890_ = ~new_n30036_ | ~new_n30035_;
  assign new_n29891_ = new_n30198_ & new_n30197_;
  assign new_n29892_ = ~new_n29974_ | ~new_n29973_;
  assign new_n29893_ = new_n30205_ & new_n30204_;
  assign new_n29894_ = ~new_n29834_ | ~new_n30033_;
  assign new_n29895_ = new_n30212_ & new_n30211_;
  assign new_n29896_ = ~new_n29767_ | ~new_n29966_;
  assign new_n29897_ = new_n30219_ & new_n30218_;
  assign new_n29898_ = ~new_n29832_ | ~new_n30031_;
  assign new_n29899_ = new_n30226_ & new_n30225_;
  assign new_n29900_ = ~new_n29764_ | ~new_n29959_;
  assign new_n29901_ = new_n30233_ & new_n30232_;
  assign new_n29902_ = ~new_n29830_ | ~new_n30029_;
  assign new_n29903_ = new_n30240_ & new_n30239_;
  assign new_n29904_ = ~new_n29761_ | ~new_n29952_;
  assign new_n29905_ = new_n30247_ & new_n30246_;
  assign new_n29906_ = ~new_n29828_ | ~new_n30027_;
  assign new_n29907_ = new_n30254_ & new_n30253_;
  assign new_n29908_ = ~new_n29758_ | ~new_n29945_;
  assign new_n29909_ = new_n30261_ & new_n30260_;
  assign new_n29910_ = ~new_n29826_ | ~new_n30025_;
  assign new_n29911_ = ~new_n9837_ | ~new_n29880_;
  assign new_n29912_ = ~new_n29845_ | ~new_n30050_;
  assign new_n29913_ = ~new_n29788_;
  assign new_n29914_ = ~new_n29721_;
  assign new_n29915_ = ~new_n29871_;
  assign new_n29916_ = new_n10677_ | pi0768;
  assign new_n29917_ = ~new_n29916_ | ~new_n29871_;
  assign new_n29918_ = ~new_n29726_;
  assign new_n29919_ = ~new_n29864_;
  assign new_n29920_ = new_n10676_ | pi0769;
  assign new_n29921_ = ~pi0769 | ~new_n10676_;
  assign new_n29922_ = ~new_n29862_;
  assign new_n29923_ = new_n10675_ | pi0770;
  assign new_n29924_ = ~new_n29923_ | ~new_n29862_;
  assign new_n29925_ = ~new_n29729_;
  assign new_n29926_ = ~new_n29860_;
  assign new_n29927_ = new_n10674_ | pi0771;
  assign new_n29928_ = ~pi0771 | ~new_n10674_;
  assign new_n29929_ = ~new_n29858_;
  assign new_n29930_ = new_n10673_ | pi0772;
  assign new_n29931_ = ~new_n29930_ | ~new_n29858_;
  assign new_n29932_ = ~new_n29732_;
  assign new_n29933_ = ~new_n29856_;
  assign new_n29934_ = new_n10672_ | pi0773;
  assign new_n29935_ = ~pi0773 | ~new_n10672_;
  assign new_n29936_ = ~new_n29854_;
  assign new_n29937_ = new_n10671_ | pi0774;
  assign new_n29938_ = ~new_n29937_ | ~new_n29854_;
  assign new_n29939_ = ~new_n29755_;
  assign new_n29940_ = ~new_n29852_;
  assign new_n29941_ = new_n9853_ | pi0775;
  assign new_n29942_ = ~new_n9853_ | ~pi0775;
  assign new_n29943_ = ~new_n29910_;
  assign new_n29944_ = new_n9852_ | pi0776;
  assign new_n29945_ = ~new_n29944_ | ~new_n29910_;
  assign new_n29946_ = ~new_n29758_;
  assign new_n29947_ = ~new_n29908_;
  assign new_n29948_ = new_n9851_ | pi0777;
  assign new_n29949_ = ~pi0777 | ~new_n9851_;
  assign new_n29950_ = ~new_n29906_;
  assign new_n29951_ = new_n9850_ | pi0778;
  assign new_n29952_ = ~new_n29951_ | ~new_n29906_;
  assign new_n29953_ = ~new_n29761_;
  assign new_n29954_ = ~new_n29904_;
  assign new_n29955_ = new_n9849_ | pi0779;
  assign new_n29956_ = ~pi0779 | ~new_n9849_;
  assign new_n29957_ = ~new_n29902_;
  assign new_n29958_ = new_n9848_ | pi0780;
  assign new_n29959_ = ~new_n29958_ | ~new_n29902_;
  assign new_n29960_ = ~new_n29764_;
  assign new_n29961_ = ~new_n29900_;
  assign new_n29962_ = new_n9847_ | pi0781;
  assign new_n29963_ = ~pi0781 | ~new_n9847_;
  assign new_n29964_ = ~new_n29898_;
  assign new_n29965_ = new_n9846_ | pi0782;
  assign new_n29966_ = ~new_n29965_ | ~new_n29898_;
  assign new_n29967_ = ~new_n29767_;
  assign new_n29968_ = ~new_n29896_;
  assign new_n29969_ = new_n9845_ | pi0783;
  assign new_n29970_ = ~pi0783 | ~new_n9845_;
  assign new_n29971_ = ~new_n29894_;
  assign new_n29972_ = new_n9844_ | pi0784;
  assign new_n29973_ = ~new_n29972_ | ~new_n29894_;
  assign new_n29974_ = ~pi0784 | ~new_n9844_;
  assign new_n29975_ = ~new_n29892_;
  assign new_n29976_ = new_n9843_ | pi0785;
  assign new_n29977_ = ~pi0785 | ~new_n9843_;
  assign new_n29978_ = ~new_n29890_;
  assign new_n29979_ = new_n9842_ | pi0786;
  assign new_n29980_ = ~pi0786 | ~new_n9842_;
  assign new_n29981_ = ~new_n29888_;
  assign new_n29982_ = new_n9841_ | pi0787;
  assign new_n29983_ = ~new_n29982_ | ~new_n29888_;
  assign new_n29984_ = ~new_n29774_;
  assign new_n29985_ = ~new_n29886_;
  assign new_n29986_ = new_n9840_ | pi0788;
  assign new_n29987_ = ~pi0788 | ~new_n9840_;
  assign new_n29988_ = ~new_n29884_;
  assign new_n29989_ = new_n9839_ | pi0789;
  assign new_n29990_ = ~new_n29989_ | ~new_n29884_;
  assign new_n29991_ = ~new_n29777_;
  assign new_n29992_ = ~new_n29882_;
  assign new_n29993_ = new_n9838_ | pi0790;
  assign new_n29994_ = ~pi0790 | ~new_n9838_;
  assign new_n29995_ = ~new_n29880_;
  assign new_n29996_ = ~pi0791 | ~new_n29880_;
  assign new_n29997_ = ~new_n29879_;
  assign new_n29998_ = new_n9836_ | pi0792;
  assign new_n29999_ = ~new_n29998_ | ~new_n29879_;
  assign new_n30000_ = ~new_n29784_;
  assign new_n30001_ = ~new_n29877_;
  assign new_n30002_ = new_n9835_ | pi0793;
  assign new_n30003_ = ~pi0793 | ~new_n9835_;
  assign new_n30004_ = ~new_n29875_;
  assign new_n30005_ = new_n9834_ | pi0794;
  assign new_n30006_ = ~pi0794 | ~new_n9834_;
  assign new_n30007_ = ~new_n29873_;
  assign new_n30008_ = new_n9833_ | pi0795;
  assign new_n30009_ = ~new_n30008_ | ~new_n29873_;
  assign new_n30010_ = ~pi0795 | ~new_n9833_;
  assign new_n30011_ = ~new_n29869_;
  assign new_n30012_ = ~pi0796 | ~new_n9832_;
  assign new_n30013_ = pi0796 | new_n9832_;
  assign new_n30014_ = ~pi0791 | ~new_n9837_;
  assign new_n30015_ = ~new_n30009_ | ~new_n29847_;
  assign new_n30016_ = ~pi0767 | ~new_n29914_;
  assign new_n30017_ = ~pi0767 | ~new_n10678_;
  assign new_n30018_ = ~new_n29819_ | ~new_n29871_;
  assign new_n30019_ = ~new_n29918_ | ~new_n29920_;
  assign new_n30020_ = new_n10676_ | pi0769;
  assign new_n30021_ = ~new_n29821_ | ~new_n29862_;
  assign new_n30022_ = ~new_n29925_ | ~new_n29927_;
  assign new_n30023_ = ~new_n29823_ | ~new_n29858_;
  assign new_n30024_ = ~new_n29932_ | ~new_n29934_;
  assign new_n30025_ = ~new_n29825_ | ~new_n29854_;
  assign new_n30026_ = ~new_n29939_ | ~new_n29941_;
  assign new_n30027_ = ~new_n29827_ | ~new_n29910_;
  assign new_n30028_ = ~new_n29946_ | ~new_n29948_;
  assign new_n30029_ = ~new_n29829_ | ~new_n29906_;
  assign new_n30030_ = ~new_n29953_ | ~new_n29955_;
  assign new_n30031_ = ~new_n29831_ | ~new_n29902_;
  assign new_n30032_ = ~new_n29960_ | ~new_n29962_;
  assign new_n30033_ = ~new_n29833_ | ~new_n29898_;
  assign new_n30034_ = ~new_n29967_ | ~new_n29969_;
  assign new_n30035_ = ~new_n29850_ | ~new_n29894_;
  assign new_n30036_ = ~new_n30037_ | ~new_n30038_;
  assign new_n30037_ = new_n9843_ | pi0785;
  assign new_n30038_ = ~new_n29974_ | ~new_n29977_;
  assign new_n30039_ = ~new_n29835_ | ~new_n29972_ | ~new_n29894_;
  assign new_n30040_ = ~new_n29836_ | ~new_n30038_;
  assign new_n30041_ = ~new_n29838_ | ~new_n29888_;
  assign new_n30042_ = ~new_n29984_ | ~new_n29986_;
  assign new_n30043_ = ~new_n29840_ | ~new_n29884_;
  assign new_n30044_ = ~new_n29991_ | ~new_n29993_;
  assign new_n30045_ = ~new_n29849_ | ~new_n29879_;
  assign new_n30046_ = ~new_n30000_ | ~new_n30002_;
  assign new_n30047_ = ~new_n29787_;
  assign new_n30048_ = ~new_n29879_ | ~new_n29842_;
  assign new_n30049_ = ~new_n29787_ | ~new_n30005_;
  assign new_n30050_ = ~new_n29843_ | ~new_n30049_ | ~new_n30048_;
  assign new_n30051_ = ~new_n29913_ | ~pi0767;
  assign new_n30052_ = ~pi0775 | ~new_n29736_;
  assign new_n30053_ = ~new_n9853_ | ~new_n29735_;
  assign new_n30054_ = ~pi0775 | ~new_n29736_;
  assign new_n30055_ = ~new_n9853_ | ~new_n29735_;
  assign new_n30056_ = ~new_n30055_ | ~new_n30054_;
  assign new_n30057_ = ~new_n29851_ | ~new_n29852_;
  assign new_n30058_ = ~new_n29940_ | ~new_n30056_;
  assign new_n30059_ = ~pi0774 | ~new_n29733_;
  assign new_n30060_ = ~new_n10671_ | ~new_n29734_;
  assign new_n30061_ = ~pi0774 | ~new_n29733_;
  assign new_n30062_ = ~new_n10671_ | ~new_n29734_;
  assign new_n30063_ = ~new_n30062_ | ~new_n30061_;
  assign new_n30064_ = ~new_n29853_ | ~new_n29854_;
  assign new_n30065_ = ~new_n29936_ | ~new_n30063_;
  assign new_n30066_ = ~pi0773 | ~new_n29713_;
  assign new_n30067_ = ~new_n10672_ | ~new_n29714_;
  assign new_n30068_ = ~pi0773 | ~new_n29713_;
  assign new_n30069_ = ~new_n10672_ | ~new_n29714_;
  assign new_n30070_ = ~new_n30069_ | ~new_n30068_;
  assign new_n30071_ = ~new_n29855_ | ~new_n29856_;
  assign new_n30072_ = ~new_n29933_ | ~new_n30070_;
  assign new_n30073_ = ~pi0772 | ~new_n29730_;
  assign new_n30074_ = ~new_n10673_ | ~new_n29731_;
  assign new_n30075_ = ~pi0772 | ~new_n29730_;
  assign new_n30076_ = ~new_n10673_ | ~new_n29731_;
  assign new_n30077_ = ~new_n30076_ | ~new_n30075_;
  assign new_n30078_ = ~new_n29857_ | ~new_n29858_;
  assign new_n30079_ = ~new_n29929_ | ~new_n30077_;
  assign new_n30080_ = ~pi0771 | ~new_n29715_;
  assign new_n30081_ = ~new_n10674_ | ~new_n29716_;
  assign new_n30082_ = ~pi0771 | ~new_n29715_;
  assign new_n30083_ = ~new_n10674_ | ~new_n29716_;
  assign new_n30084_ = ~new_n30083_ | ~new_n30082_;
  assign new_n30085_ = ~new_n29859_ | ~new_n29860_;
  assign new_n30086_ = ~new_n29926_ | ~new_n30084_;
  assign new_n30087_ = ~pi0770 | ~new_n29727_;
  assign new_n30088_ = ~new_n10675_ | ~new_n29728_;
  assign new_n30089_ = ~pi0770 | ~new_n29727_;
  assign new_n30090_ = ~new_n10675_ | ~new_n29728_;
  assign new_n30091_ = ~new_n30090_ | ~new_n30089_;
  assign new_n30092_ = ~new_n29861_ | ~new_n29862_;
  assign new_n30093_ = ~new_n29922_ | ~new_n30091_;
  assign new_n30094_ = ~pi0769 | ~new_n29717_;
  assign new_n30095_ = ~new_n10676_ | ~new_n29718_;
  assign new_n30096_ = ~pi0769 | ~new_n29717_;
  assign new_n30097_ = ~new_n10676_ | ~new_n29718_;
  assign new_n30098_ = ~new_n30097_ | ~new_n30096_;
  assign new_n30099_ = ~new_n29863_ | ~new_n29864_;
  assign new_n30100_ = ~new_n29919_ | ~new_n30098_;
  assign new_n30101_ = ~pi0797 | ~new_n29866_;
  assign new_n30102_ = ~new_n9831_ | ~new_n29865_;
  assign new_n30103_ = ~new_n30102_ | ~new_n30101_;
  assign new_n30104_ = ~pi0797 | ~new_n29866_;
  assign new_n30105_ = ~new_n9831_ | ~new_n29865_;
  assign new_n30106_ = ~new_n29786_ | ~new_n29710_ | ~new_n29785_;
  assign new_n30107_ = ~pi0796 | ~new_n9832_ | ~new_n30103_;
  assign new_n30108_ = ~pi0796 | ~new_n29785_;
  assign new_n30109_ = ~new_n9832_ | ~new_n29786_;
  assign new_n30110_ = ~pi0796 | ~new_n29785_;
  assign new_n30111_ = ~new_n9832_ | ~new_n29786_;
  assign new_n30112_ = ~new_n30111_ | ~new_n30110_;
  assign new_n30113_ = ~new_n29868_ | ~new_n29869_;
  assign new_n30114_ = ~new_n30011_ | ~new_n30112_;
  assign new_n30115_ = ~pi0768 | ~new_n29724_;
  assign new_n30116_ = ~new_n10677_ | ~new_n29725_;
  assign new_n30117_ = ~pi0768 | ~new_n29724_;
  assign new_n30118_ = ~new_n10677_ | ~new_n29725_;
  assign new_n30119_ = ~new_n30118_ | ~new_n30117_;
  assign new_n30120_ = ~new_n29870_ | ~new_n29871_;
  assign new_n30121_ = ~new_n29915_ | ~new_n30119_;
  assign new_n30122_ = ~pi0795 | ~new_n29739_;
  assign new_n30123_ = ~new_n9833_ | ~new_n29740_;
  assign new_n30124_ = ~pi0795 | ~new_n29739_;
  assign new_n30125_ = ~new_n9833_ | ~new_n29740_;
  assign new_n30126_ = ~new_n30125_ | ~new_n30124_;
  assign new_n30127_ = ~new_n29872_ | ~new_n29873_;
  assign new_n30128_ = ~new_n30007_ | ~new_n30126_;
  assign new_n30129_ = ~pi0794 | ~new_n29737_;
  assign new_n30130_ = ~new_n9834_ | ~new_n29738_;
  assign new_n30131_ = ~pi0794 | ~new_n29737_;
  assign new_n30132_ = ~new_n9834_ | ~new_n29738_;
  assign new_n30133_ = ~new_n30132_ | ~new_n30131_;
  assign new_n30134_ = ~new_n29874_ | ~new_n29875_;
  assign new_n30135_ = ~new_n30004_ | ~new_n30133_;
  assign new_n30136_ = ~pi0793 | ~new_n29780_;
  assign new_n30137_ = ~new_n9835_ | ~new_n29781_;
  assign new_n30138_ = ~pi0793 | ~new_n29780_;
  assign new_n30139_ = ~new_n9835_ | ~new_n29781_;
  assign new_n30140_ = ~new_n30139_ | ~new_n30138_;
  assign new_n30141_ = ~new_n29876_ | ~new_n29877_;
  assign new_n30142_ = ~new_n30001_ | ~new_n30140_;
  assign new_n30143_ = ~pi0792 | ~new_n29782_;
  assign new_n30144_ = ~new_n9836_ | ~new_n29783_;
  assign new_n30145_ = ~pi0792 | ~new_n29782_;
  assign new_n30146_ = ~new_n9836_ | ~new_n29783_;
  assign new_n30147_ = ~new_n30146_ | ~new_n30145_;
  assign new_n30148_ = ~new_n29878_ | ~new_n29879_;
  assign new_n30149_ = ~new_n29997_ | ~new_n30147_;
  assign new_n30150_ = ~pi0791 | ~new_n29880_;
  assign new_n30151_ = ~new_n29995_ | ~new_n29779_;
  assign new_n30152_ = ~pi0791 | ~new_n29880_;
  assign new_n30153_ = ~new_n29995_ | ~new_n29779_;
  assign new_n30154_ = ~new_n30153_ | ~new_n30152_;
  assign new_n30155_ = ~new_n29778_ | ~new_n30151_ | ~new_n30150_;
  assign new_n30156_ = ~new_n30154_ | ~new_n9837_;
  assign new_n30157_ = ~pi0790 | ~new_n29741_;
  assign new_n30158_ = ~new_n9838_ | ~new_n29742_;
  assign new_n30159_ = ~pi0790 | ~new_n29741_;
  assign new_n30160_ = ~new_n9838_ | ~new_n29742_;
  assign new_n30161_ = ~new_n30160_ | ~new_n30159_;
  assign new_n30162_ = ~new_n29881_ | ~new_n29882_;
  assign new_n30163_ = ~new_n29992_ | ~new_n30161_;
  assign new_n30164_ = ~pi0789 | ~new_n29775_;
  assign new_n30165_ = ~new_n9839_ | ~new_n29776_;
  assign new_n30166_ = ~pi0789 | ~new_n29775_;
  assign new_n30167_ = ~new_n9839_ | ~new_n29776_;
  assign new_n30168_ = ~new_n30167_ | ~new_n30166_;
  assign new_n30169_ = ~new_n29883_ | ~new_n29884_;
  assign new_n30170_ = ~new_n29988_ | ~new_n30168_;
  assign new_n30171_ = ~pi0788 | ~new_n29743_;
  assign new_n30172_ = ~new_n9840_ | ~new_n29744_;
  assign new_n30173_ = ~pi0788 | ~new_n29743_;
  assign new_n30174_ = ~new_n9840_ | ~new_n29744_;
  assign new_n30175_ = ~new_n30174_ | ~new_n30173_;
  assign new_n30176_ = ~new_n29885_ | ~new_n29886_;
  assign new_n30177_ = ~new_n29985_ | ~new_n30175_;
  assign new_n30178_ = ~pi0787 | ~new_n29772_;
  assign new_n30179_ = ~new_n9841_ | ~new_n29773_;
  assign new_n30180_ = ~pi0787 | ~new_n29772_;
  assign new_n30181_ = ~new_n9841_ | ~new_n29773_;
  assign new_n30182_ = ~new_n30181_ | ~new_n30180_;
  assign new_n30183_ = ~new_n29887_ | ~new_n29888_;
  assign new_n30184_ = ~new_n29981_ | ~new_n30182_;
  assign new_n30185_ = ~pi0786 | ~new_n29745_;
  assign new_n30186_ = ~new_n9842_ | ~new_n29746_;
  assign new_n30187_ = ~pi0786 | ~new_n29745_;
  assign new_n30188_ = ~new_n9842_ | ~new_n29746_;
  assign new_n30189_ = ~new_n30188_ | ~new_n30187_;
  assign new_n30190_ = ~new_n29889_ | ~new_n29890_;
  assign new_n30191_ = ~new_n29978_ | ~new_n30189_;
  assign new_n30192_ = ~pi0767 | ~new_n29721_;
  assign new_n30193_ = ~new_n29914_ | ~new_n29723_;
  assign new_n30194_ = ~new_n30193_ | ~new_n30192_;
  assign new_n30195_ = ~new_n10678_ | ~new_n29721_ | ~new_n29723_;
  assign new_n30196_ = ~new_n30194_ | ~new_n29722_;
  assign new_n30197_ = ~pi0785 | ~new_n29768_;
  assign new_n30198_ = ~new_n9843_ | ~new_n29769_;
  assign new_n30199_ = ~pi0785 | ~new_n29768_;
  assign new_n30200_ = ~new_n9843_ | ~new_n29769_;
  assign new_n30201_ = ~new_n30200_ | ~new_n30199_;
  assign new_n30202_ = ~new_n29891_ | ~new_n29892_;
  assign new_n30203_ = ~new_n29975_ | ~new_n30201_;
  assign new_n30204_ = ~pi0784 | ~new_n29770_;
  assign new_n30205_ = ~new_n9844_ | ~new_n29771_;
  assign new_n30206_ = ~pi0784 | ~new_n29770_;
  assign new_n30207_ = ~new_n9844_ | ~new_n29771_;
  assign new_n30208_ = ~new_n30207_ | ~new_n30206_;
  assign new_n30209_ = ~new_n29893_ | ~new_n29894_;
  assign new_n30210_ = ~new_n29971_ | ~new_n30208_;
  assign new_n30211_ = ~pi0783 | ~new_n29747_;
  assign new_n30212_ = ~new_n9845_ | ~new_n29748_;
  assign new_n30213_ = ~pi0783 | ~new_n29747_;
  assign new_n30214_ = ~new_n9845_ | ~new_n29748_;
  assign new_n30215_ = ~new_n30214_ | ~new_n30213_;
  assign new_n30216_ = ~new_n29895_ | ~new_n29896_;
  assign new_n30217_ = ~new_n29968_ | ~new_n30215_;
  assign new_n30218_ = ~pi0782 | ~new_n29765_;
  assign new_n30219_ = ~new_n9846_ | ~new_n29766_;
  assign new_n30220_ = ~pi0782 | ~new_n29765_;
  assign new_n30221_ = ~new_n9846_ | ~new_n29766_;
  assign new_n30222_ = ~new_n30221_ | ~new_n30220_;
  assign new_n30223_ = ~new_n29897_ | ~new_n29898_;
  assign new_n30224_ = ~new_n29964_ | ~new_n30222_;
  assign new_n30225_ = ~pi0781 | ~new_n29749_;
  assign new_n30226_ = ~new_n9847_ | ~new_n29750_;
  assign new_n30227_ = ~pi0781 | ~new_n29749_;
  assign new_n30228_ = ~new_n9847_ | ~new_n29750_;
  assign new_n30229_ = ~new_n30228_ | ~new_n30227_;
  assign new_n30230_ = ~new_n29899_ | ~new_n29900_;
  assign new_n30231_ = ~new_n29961_ | ~new_n30229_;
  assign new_n30232_ = ~pi0780 | ~new_n29762_;
  assign new_n30233_ = ~new_n9848_ | ~new_n29763_;
  assign new_n30234_ = ~pi0780 | ~new_n29762_;
  assign new_n30235_ = ~new_n9848_ | ~new_n29763_;
  assign new_n30236_ = ~new_n30235_ | ~new_n30234_;
  assign new_n30237_ = ~new_n29901_ | ~new_n29902_;
  assign new_n30238_ = ~new_n29957_ | ~new_n30236_;
  assign new_n30239_ = ~pi0779 | ~new_n29751_;
  assign new_n30240_ = ~new_n9849_ | ~new_n29752_;
  assign new_n30241_ = ~pi0779 | ~new_n29751_;
  assign new_n30242_ = ~new_n9849_ | ~new_n29752_;
  assign new_n30243_ = ~new_n30242_ | ~new_n30241_;
  assign new_n30244_ = ~new_n29903_ | ~new_n29904_;
  assign new_n30245_ = ~new_n29954_ | ~new_n30243_;
  assign new_n30246_ = ~pi0778 | ~new_n29759_;
  assign new_n30247_ = ~new_n9850_ | ~new_n29760_;
  assign new_n30248_ = ~pi0778 | ~new_n29759_;
  assign new_n30249_ = ~new_n9850_ | ~new_n29760_;
  assign new_n30250_ = ~new_n30249_ | ~new_n30248_;
  assign new_n30251_ = ~new_n29905_ | ~new_n29906_;
  assign new_n30252_ = ~new_n29950_ | ~new_n30250_;
  assign new_n30253_ = ~pi0777 | ~new_n29753_;
  assign new_n30254_ = ~new_n9851_ | ~new_n29754_;
  assign new_n30255_ = ~pi0777 | ~new_n29753_;
  assign new_n30256_ = ~new_n9851_ | ~new_n29754_;
  assign new_n30257_ = ~new_n30256_ | ~new_n30255_;
  assign new_n30258_ = ~new_n29907_ | ~new_n29908_;
  assign new_n30259_ = ~new_n29947_ | ~new_n30257_;
  assign new_n30260_ = ~pi0776 | ~new_n29756_;
  assign new_n30261_ = ~new_n9852_ | ~new_n29757_;
  assign new_n30262_ = ~pi0776 | ~new_n29756_;
  assign new_n30263_ = ~new_n9852_ | ~new_n29757_;
  assign new_n30264_ = ~new_n30263_ | ~new_n30262_;
  assign new_n30265_ = ~new_n29909_ | ~new_n29910_;
  assign new_n30266_ = ~new_n29943_ | ~new_n30264_;
  assign new_n30267_ = ~pi0766 | ~new_n29719_;
  assign new_n30268_ = ~new_n10679_ | ~new_n29720_;
  assign new_n30269_ = ~new_n30306_ | ~new_n30305_;
  assign new_n30270_ = ~pi0760 | ~new_n30279_;
  assign new_n30271_ = ~pi0764;
  assign new_n30272_ = ~pi0758;
  assign new_n30273_ = ~pi0763;
  assign new_n30274_ = ~pi0757;
  assign new_n30275_ = ~pi0762;
  assign new_n30276_ = ~pi0761;
  assign new_n30277_ = ~new_n30302_ | ~new_n30301_;
  assign new_n30278_ = ~pi0756;
  assign new_n30279_ = ~pi0765;
  assign new_n30280_ = ~new_n30311_ | ~new_n30310_;
  assign new_n30281_ = ~new_n30316_ | ~new_n30315_;
  assign new_n30282_ = ~new_n30321_ | ~new_n30320_;
  assign new_n30283_ = ~new_n30326_ | ~new_n30325_;
  assign new_n30284_ = ~new_n30308_ | ~new_n30307_;
  assign new_n30285_ = ~new_n30313_ | ~new_n30312_;
  assign new_n30286_ = ~new_n30318_ | ~new_n30317_;
  assign new_n30287_ = ~new_n30323_ | ~new_n30322_;
  assign new_n30288_ = ~new_n30298_ | ~new_n30297_;
  assign new_n30289_ = ~new_n30294_ | ~new_n30293_;
  assign new_n30290_ = ~pi0759;
  assign new_n30291_ = ~new_n30270_;
  assign new_n30292_ = ~new_n30291_ | ~new_n30271_;
  assign new_n30293_ = ~new_n30292_ | ~new_n30290_;
  assign new_n30294_ = ~pi0764 | ~new_n30270_;
  assign new_n30295_ = ~new_n30289_;
  assign new_n30296_ = ~pi0758 | ~new_n30273_;
  assign new_n30297_ = ~new_n30296_ | ~new_n30289_;
  assign new_n30298_ = ~pi0763 | ~new_n30272_;
  assign new_n30299_ = ~new_n30288_;
  assign new_n30300_ = ~pi0757 | ~new_n30275_;
  assign new_n30301_ = ~new_n30300_ | ~new_n30288_;
  assign new_n30302_ = ~pi0762 | ~new_n30274_;
  assign new_n30303_ = ~new_n30277_;
  assign new_n30304_ = ~pi0761 | ~new_n30278_;
  assign new_n30305_ = ~new_n30303_ | ~new_n30304_;
  assign new_n30306_ = ~pi0756 | ~new_n30276_;
  assign new_n30307_ = ~pi0756 | ~new_n30276_;
  assign new_n30308_ = ~pi0761 | ~new_n30278_;
  assign new_n30309_ = ~new_n30284_;
  assign new_n30310_ = ~new_n30309_ | ~new_n30303_;
  assign new_n30311_ = ~new_n30284_ | ~new_n30277_;
  assign new_n30312_ = ~pi0757 | ~new_n30275_;
  assign new_n30313_ = ~pi0762 | ~new_n30274_;
  assign new_n30314_ = ~new_n30285_;
  assign new_n30315_ = ~new_n30299_ | ~new_n30314_;
  assign new_n30316_ = ~new_n30285_ | ~new_n30288_;
  assign new_n30317_ = ~pi0758 | ~new_n30273_;
  assign new_n30318_ = ~pi0763 | ~new_n30272_;
  assign new_n30319_ = ~new_n30286_;
  assign new_n30320_ = ~new_n30295_ | ~new_n30319_;
  assign new_n30321_ = ~new_n30286_ | ~new_n30289_;
  assign new_n30322_ = ~pi0759 | ~new_n30271_;
  assign new_n30323_ = ~pi0764 | ~new_n30290_;
  assign new_n30324_ = ~new_n30287_;
  assign new_n30325_ = ~new_n30324_ | ~new_n30291_;
  assign new_n30326_ = ~new_n30287_ | ~new_n30270_;
  assign new_n30327_ = ~new_n10689_ & ~new_n30328_;
  assign new_n30328_ = ~new_n10690_ & ~new_n10689_ & ~new_n10691_ & ~new_n10692_ & ~new_n10693_;
  assign new_n30329_ = ~pi0766;
  assign new_n30330_ = ~new_n30419_ | ~new_n30450_;
  assign new_n30331_ = ~pi0767;
  assign new_n30332_ = ~pi0769;
  assign new_n30333_ = ~pi0769 | ~new_n30419_;
  assign new_n30334_ = ~pi0770;
  assign new_n30335_ = ~pi0770 | ~new_n30423_;
  assign new_n30336_ = ~pi0771;
  assign new_n30337_ = ~pi0772;
  assign new_n30338_ = ~pi0771 | ~new_n30424_;
  assign new_n30339_ = ~new_n30425_ | ~pi0772;
  assign new_n30340_ = ~pi0773;
  assign new_n30341_ = ~pi0773 | ~new_n30426_;
  assign new_n30342_ = ~pi0774;
  assign new_n30343_ = ~pi0774 | ~new_n30427_;
  assign new_n30344_ = ~pi0775;
  assign new_n30345_ = ~pi0775 | ~new_n30428_;
  assign new_n30346_ = ~pi0776;
  assign new_n30347_ = ~pi0776 | ~new_n30429_;
  assign new_n30348_ = ~pi0777;
  assign new_n30349_ = ~pi0777 | ~new_n30430_;
  assign new_n30350_ = ~pi0778;
  assign new_n30351_ = ~pi0778 | ~new_n30431_;
  assign new_n30352_ = ~pi0779;
  assign new_n30353_ = ~pi0779 | ~new_n30432_;
  assign new_n30354_ = ~pi0780;
  assign new_n30355_ = ~pi0780 | ~new_n30433_;
  assign new_n30356_ = ~pi0781;
  assign new_n30357_ = ~pi0781 | ~new_n30434_;
  assign new_n30358_ = ~pi0782;
  assign new_n30359_ = ~pi0782 | ~new_n30435_;
  assign new_n30360_ = ~pi0783;
  assign new_n30361_ = ~pi0783 | ~new_n30436_;
  assign new_n30362_ = ~pi0784;
  assign new_n30363_ = ~pi0784 | ~new_n30437_;
  assign new_n30364_ = ~pi0785;
  assign new_n30365_ = ~pi0785 | ~new_n30438_;
  assign new_n30366_ = ~pi0786;
  assign new_n30367_ = ~pi0786 | ~new_n30439_;
  assign new_n30368_ = ~pi0787;
  assign new_n30369_ = ~pi0787 | ~new_n30440_;
  assign new_n30370_ = ~pi0788;
  assign new_n30371_ = ~pi0788 | ~new_n30441_;
  assign new_n30372_ = ~pi0789;
  assign new_n30373_ = ~pi0789 | ~new_n30442_;
  assign new_n30374_ = ~pi0790;
  assign new_n30375_ = ~pi0790 | ~new_n30443_;
  assign new_n30376_ = ~pi0791;
  assign new_n30377_ = ~pi0791 | ~new_n30444_;
  assign new_n30378_ = ~pi0792;
  assign new_n30379_ = ~pi0792 | ~new_n30445_;
  assign new_n30380_ = ~pi0793;
  assign new_n30381_ = ~pi0793 | ~new_n30446_;
  assign new_n30382_ = ~pi0794;
  assign new_n30383_ = ~pi0794 | ~new_n30447_;
  assign new_n30384_ = ~pi0795;
  assign new_n30385_ = ~pi0796;
  assign new_n30386_ = ~pi0795 | ~new_n30448_;
  assign new_n30387_ = ~pi0768;
  assign new_n30388_ = ~new_n30453_ | ~new_n30452_;
  assign new_n30389_ = ~new_n30455_ | ~new_n30454_;
  assign new_n30390_ = ~new_n30457_ | ~new_n30456_;
  assign new_n30391_ = ~new_n30459_ | ~new_n30458_;
  assign new_n30392_ = ~new_n30461_ | ~new_n30460_;
  assign new_n30393_ = ~new_n30463_ | ~new_n30462_;
  assign new_n30394_ = ~new_n30465_ | ~new_n30464_;
  assign new_n30395_ = ~new_n30467_ | ~new_n30466_;
  assign new_n30396_ = ~new_n30469_ | ~new_n30468_;
  assign new_n30397_ = ~new_n30471_ | ~new_n30470_;
  assign new_n30398_ = ~new_n30473_ | ~new_n30472_;
  assign new_n30399_ = ~new_n30475_ | ~new_n30474_;
  assign new_n30400_ = ~new_n30477_ | ~new_n30476_;
  assign new_n30401_ = ~new_n30479_ | ~new_n30478_;
  assign new_n30402_ = ~new_n30481_ | ~new_n30480_;
  assign new_n30403_ = ~new_n30483_ | ~new_n30482_;
  assign new_n30404_ = ~new_n30485_ | ~new_n30484_;
  assign new_n30405_ = ~new_n30487_ | ~new_n30486_;
  assign new_n30406_ = ~new_n30489_ | ~new_n30488_;
  assign new_n30407_ = ~new_n30491_ | ~new_n30490_;
  assign new_n30408_ = ~new_n30493_ | ~new_n30492_;
  assign new_n30409_ = ~new_n30495_ | ~new_n30494_;
  assign new_n30410_ = ~new_n30499_ | ~new_n30498_;
  assign new_n30411_ = ~new_n30501_ | ~new_n30500_;
  assign new_n30412_ = ~new_n30503_ | ~new_n30502_;
  assign new_n30413_ = ~new_n30505_ | ~new_n30504_;
  assign new_n30414_ = ~new_n30507_ | ~new_n30506_;
  assign new_n30415_ = ~new_n30509_ | ~new_n30508_;
  assign new_n30416_ = ~new_n30511_ | ~new_n30510_;
  assign new_n30417_ = ~pi0797;
  assign new_n30418_ = ~new_n30449_ | ~pi0796;
  assign new_n30419_ = ~new_n30387_ | ~new_n30421_;
  assign new_n30420_ = new_n30497_ & new_n30496_;
  assign new_n30421_ = ~pi0767 | ~pi0766;
  assign new_n30422_ = ~new_n30419_;
  assign new_n30423_ = ~new_n30333_;
  assign new_n30424_ = ~new_n30335_;
  assign new_n30425_ = ~new_n30338_;
  assign new_n30426_ = ~new_n30339_;
  assign new_n30427_ = ~new_n30341_;
  assign new_n30428_ = ~new_n30343_;
  assign new_n30429_ = ~new_n30345_;
  assign new_n30430_ = ~new_n30347_;
  assign new_n30431_ = ~new_n30349_;
  assign new_n30432_ = ~new_n30351_;
  assign new_n30433_ = ~new_n30353_;
  assign new_n30434_ = ~new_n30355_;
  assign new_n30435_ = ~new_n30357_;
  assign new_n30436_ = ~new_n30359_;
  assign new_n30437_ = ~new_n30361_;
  assign new_n30438_ = ~new_n30363_;
  assign new_n30439_ = ~new_n30365_;
  assign new_n30440_ = ~new_n30367_;
  assign new_n30441_ = ~new_n30369_;
  assign new_n30442_ = ~new_n30371_;
  assign new_n30443_ = ~new_n30373_;
  assign new_n30444_ = ~new_n30375_;
  assign new_n30445_ = ~new_n30377_;
  assign new_n30446_ = ~new_n30379_;
  assign new_n30447_ = ~new_n30381_;
  assign new_n30448_ = ~new_n30383_;
  assign new_n30449_ = ~new_n30386_;
  assign new_n30450_ = ~pi0768 | ~pi0767 | ~pi0766;
  assign new_n30451_ = ~new_n30418_;
  assign new_n30452_ = ~pi0772 | ~new_n30338_;
  assign new_n30453_ = ~new_n30425_ | ~new_n30337_;
  assign new_n30454_ = ~pi0796 | ~new_n30386_;
  assign new_n30455_ = ~new_n30449_ | ~new_n30385_;
  assign new_n30456_ = ~pi0795 | ~new_n30383_;
  assign new_n30457_ = ~new_n30448_ | ~new_n30384_;
  assign new_n30458_ = ~pi0790 | ~new_n30373_;
  assign new_n30459_ = ~new_n30443_ | ~new_n30374_;
  assign new_n30460_ = ~pi0783 | ~new_n30359_;
  assign new_n30461_ = ~new_n30436_ | ~new_n30360_;
  assign new_n30462_ = ~pi0786 | ~new_n30365_;
  assign new_n30463_ = ~new_n30439_ | ~new_n30366_;
  assign new_n30464_ = ~pi0779 | ~new_n30351_;
  assign new_n30465_ = ~new_n30432_ | ~new_n30352_;
  assign new_n30466_ = ~pi0775 | ~new_n30343_;
  assign new_n30467_ = ~new_n30428_ | ~new_n30344_;
  assign new_n30468_ = ~pi0788 | ~new_n30369_;
  assign new_n30469_ = ~new_n30441_ | ~new_n30370_;
  assign new_n30470_ = ~pi0784 | ~new_n30361_;
  assign new_n30471_ = ~new_n30437_ | ~new_n30362_;
  assign new_n30472_ = ~pi0777 | ~new_n30347_;
  assign new_n30473_ = ~new_n30430_ | ~new_n30348_;
  assign new_n30474_ = ~pi0792 | ~new_n30377_;
  assign new_n30475_ = ~new_n30445_ | ~new_n30378_;
  assign new_n30476_ = ~pi0781 | ~new_n30355_;
  assign new_n30477_ = ~new_n30434_ | ~new_n30356_;
  assign new_n30478_ = ~pi0770 | ~new_n30333_;
  assign new_n30479_ = ~new_n30423_ | ~new_n30334_;
  assign new_n30480_ = ~pi0793 | ~new_n30379_;
  assign new_n30481_ = ~new_n30446_ | ~new_n30380_;
  assign new_n30482_ = ~pi0780 | ~new_n30353_;
  assign new_n30483_ = ~new_n30433_ | ~new_n30354_;
  assign new_n30484_ = ~pi0771 | ~new_n30335_;
  assign new_n30485_ = ~new_n30424_ | ~new_n30336_;
  assign new_n30486_ = ~pi0774 | ~new_n30341_;
  assign new_n30487_ = ~new_n30427_ | ~new_n30342_;
  assign new_n30488_ = ~pi0789 | ~new_n30371_;
  assign new_n30489_ = ~new_n30442_ | ~new_n30372_;
  assign new_n30490_ = ~pi0785 | ~new_n30363_;
  assign new_n30491_ = ~new_n30438_ | ~new_n30364_;
  assign new_n30492_ = ~pi0776 | ~new_n30345_;
  assign new_n30493_ = ~new_n30429_ | ~new_n30346_;
  assign new_n30494_ = ~pi0797 | ~new_n30418_;
  assign new_n30495_ = ~new_n30451_ | ~new_n30417_;
  assign new_n30496_ = ~pi0769 | ~new_n30419_;
  assign new_n30497_ = ~new_n30422_ | ~new_n30332_;
  assign new_n30498_ = ~pi0767 | ~new_n30329_;
  assign new_n30499_ = ~pi0766 | ~new_n30331_;
  assign new_n30500_ = ~pi0794 | ~new_n30381_;
  assign new_n30501_ = ~new_n30447_ | ~new_n30382_;
  assign new_n30502_ = ~pi0787 | ~new_n30367_;
  assign new_n30503_ = ~new_n30440_ | ~new_n30368_;
  assign new_n30504_ = ~pi0778 | ~new_n30349_;
  assign new_n30505_ = ~new_n30431_ | ~new_n30350_;
  assign new_n30506_ = ~pi0773 | ~new_n30339_;
  assign new_n30507_ = ~new_n30426_ | ~new_n30340_;
  assign new_n30508_ = ~pi0791 | ~new_n30375_;
  assign new_n30509_ = ~new_n30444_ | ~new_n30376_;
  assign new_n30510_ = ~pi0782 | ~new_n30357_;
  assign new_n30511_ = ~new_n30435_ | ~new_n30358_;
  assign new_n30512_ = new_n30639_ & new_n30537_;
  assign new_n30513_ = new_n30637_ & new_n30538_;
  assign new_n30514_ = new_n30635_ & new_n30539_;
  assign new_n30515_ = new_n30633_ & new_n30540_;
  assign new_n30516_ = new_n30631_ & new_n30541_;
  assign new_n30517_ = new_n30629_ & new_n30542_;
  assign new_n30518_ = new_n30627_ & new_n30543_;
  assign new_n30519_ = new_n30625_ & new_n30544_;
  assign new_n30520_ = new_n30623_ & new_n30545_;
  assign new_n30521_ = new_n30621_ & new_n30546_;
  assign new_n30522_ = new_n30619_ & new_n30568_;
  assign new_n30523_ = new_n30607_ & new_n30530_;
  assign new_n30524_ = new_n30605_ & new_n30531_;
  assign new_n30525_ = new_n30603_ & new_n30532_;
  assign new_n30526_ = new_n30601_ & new_n30536_;
  assign new_n30527_ = ~new_n30583_ | ~new_n30640_;
  assign new_n30528_ = ~new_n10687_;
  assign new_n30529_ = ~new_n30582_ | ~new_n30583_;
  assign new_n30530_ = ~new_n30535_ | ~new_n30595_ | ~new_n30570_;
  assign new_n30531_ = ~new_n30534_ | ~new_n30596_ | ~new_n30565_;
  assign new_n30532_ = ~new_n30533_ | ~new_n30597_ | ~new_n30563_;
  assign new_n30533_ = ~new_n10680_;
  assign new_n30534_ = ~new_n10682_;
  assign new_n30535_ = ~new_n10684_;
  assign new_n30536_ = ~new_n30550_ | ~new_n30598_;
  assign new_n30537_ = ~new_n30551_ | ~new_n30599_;
  assign new_n30538_ = ~new_n30552_ | ~new_n30608_;
  assign new_n30539_ = ~new_n30553_ | ~new_n30609_;
  assign new_n30540_ = ~new_n30554_ | ~new_n30610_;
  assign new_n30541_ = ~new_n30555_ | ~new_n30611_;
  assign new_n30542_ = ~new_n30556_ | ~new_n30612_;
  assign new_n30543_ = ~new_n30557_ | ~new_n30613_;
  assign new_n30544_ = ~new_n30558_ | ~new_n30614_;
  assign new_n30545_ = ~new_n30559_ | ~new_n30615_;
  assign new_n30546_ = ~new_n30560_ | ~new_n30616_;
  assign new_n30547_ = ~new_n9808_;
  assign new_n30548_ = ~new_n9658_;
  assign new_n30549_ = ~new_n30662_ | ~new_n30661_;
  assign new_n30550_ = ~new_n9830_ & ~new_n9829_;
  assign new_n30551_ = ~new_n9828_ & ~new_n9827_;
  assign new_n30552_ = ~new_n9826_ & ~new_n9825_;
  assign new_n30553_ = ~new_n9824_ & ~new_n9823_;
  assign new_n30554_ = ~new_n9822_ & ~new_n9821_;
  assign new_n30555_ = ~new_n9820_ & ~new_n9819_;
  assign new_n30556_ = ~new_n9818_ & ~new_n9817_;
  assign new_n30557_ = ~new_n9816_ & ~new_n9815_;
  assign new_n30558_ = ~new_n9814_ & ~new_n9813_;
  assign new_n30559_ = ~new_n9812_ & ~new_n9811_;
  assign new_n30560_ = ~new_n9810_ & ~new_n9809_;
  assign new_n30561_ = ~new_n9830_;
  assign new_n30562_ = new_n30642_ & new_n30641_;
  assign new_n30563_ = ~new_n10681_;
  assign new_n30564_ = new_n30644_ & new_n30643_;
  assign new_n30565_ = ~new_n10683_;
  assign new_n30566_ = new_n30646_ & new_n30645_;
  assign new_n30567_ = ~new_n9807_;
  assign new_n30568_ = ~new_n30617_ | ~new_n30547_;
  assign new_n30569_ = new_n30648_ & new_n30647_;
  assign new_n30570_ = ~new_n10685_;
  assign new_n30571_ = new_n30650_ & new_n30649_;
  assign new_n30572_ = ~new_n9810_;
  assign new_n30573_ = new_n30652_ & new_n30651_;
  assign new_n30574_ = ~new_n9812_;
  assign new_n30575_ = new_n30654_ & new_n30653_;
  assign new_n30576_ = ~new_n9814_;
  assign new_n30577_ = new_n30656_ & new_n30655_;
  assign new_n30578_ = ~new_n9816_;
  assign new_n30579_ = new_n30658_ & new_n30657_;
  assign new_n30580_ = ~new_n9818_;
  assign new_n30581_ = new_n30660_ & new_n30659_;
  assign new_n30582_ = ~new_n10686_;
  assign new_n30583_ = ~new_n10687_ | ~new_n30548_;
  assign new_n30584_ = ~new_n9820_;
  assign new_n30585_ = new_n30664_ & new_n30663_;
  assign new_n30586_ = ~new_n9822_;
  assign new_n30587_ = new_n30666_ & new_n30665_;
  assign new_n30588_ = ~new_n9824_;
  assign new_n30589_ = new_n30668_ & new_n30667_;
  assign new_n30590_ = ~new_n9826_;
  assign new_n30591_ = new_n30670_ & new_n30669_;
  assign new_n30592_ = ~new_n9828_;
  assign new_n30593_ = new_n30672_ & new_n30671_;
  assign new_n30594_ = ~new_n30583_;
  assign new_n30595_ = ~new_n30529_;
  assign new_n30596_ = ~new_n30530_;
  assign new_n30597_ = ~new_n30531_;
  assign new_n30598_ = ~new_n30532_;
  assign new_n30599_ = ~new_n30536_;
  assign new_n30600_ = ~new_n30598_ | ~new_n30561_;
  assign new_n30601_ = ~new_n9829_ | ~new_n30600_;
  assign new_n30602_ = ~new_n30597_ | ~new_n30563_;
  assign new_n30603_ = ~new_n10680_ | ~new_n30602_;
  assign new_n30604_ = ~new_n30596_ | ~new_n30565_;
  assign new_n30605_ = ~new_n10682_ | ~new_n30604_;
  assign new_n30606_ = ~new_n30595_ | ~new_n30570_;
  assign new_n30607_ = ~new_n10684_ | ~new_n30606_;
  assign new_n30608_ = ~new_n30537_;
  assign new_n30609_ = ~new_n30538_;
  assign new_n30610_ = ~new_n30539_;
  assign new_n30611_ = ~new_n30540_;
  assign new_n30612_ = ~new_n30541_;
  assign new_n30613_ = ~new_n30542_;
  assign new_n30614_ = ~new_n30543_;
  assign new_n30615_ = ~new_n30544_;
  assign new_n30616_ = ~new_n30545_;
  assign new_n30617_ = ~new_n30546_;
  assign new_n30618_ = ~new_n30568_;
  assign new_n30619_ = ~new_n9808_ | ~new_n30546_;
  assign new_n30620_ = ~new_n30616_ | ~new_n30572_;
  assign new_n30621_ = ~new_n9809_ | ~new_n30620_;
  assign new_n30622_ = ~new_n30615_ | ~new_n30574_;
  assign new_n30623_ = ~new_n9811_ | ~new_n30622_;
  assign new_n30624_ = ~new_n30614_ | ~new_n30576_;
  assign new_n30625_ = ~new_n9813_ | ~new_n30624_;
  assign new_n30626_ = ~new_n30613_ | ~new_n30578_;
  assign new_n30627_ = ~new_n9815_ | ~new_n30626_;
  assign new_n30628_ = ~new_n30612_ | ~new_n30580_;
  assign new_n30629_ = ~new_n9817_ | ~new_n30628_;
  assign new_n30630_ = ~new_n30611_ | ~new_n30584_;
  assign new_n30631_ = ~new_n9819_ | ~new_n30630_;
  assign new_n30632_ = ~new_n30610_ | ~new_n30586_;
  assign new_n30633_ = ~new_n9821_ | ~new_n30632_;
  assign new_n30634_ = ~new_n30609_ | ~new_n30588_;
  assign new_n30635_ = ~new_n9823_ | ~new_n30634_;
  assign new_n30636_ = ~new_n30608_ | ~new_n30590_;
  assign new_n30637_ = ~new_n9825_ | ~new_n30636_;
  assign new_n30638_ = ~new_n30599_ | ~new_n30592_;
  assign new_n30639_ = ~new_n9827_ | ~new_n30638_;
  assign new_n30640_ = ~new_n9658_ | ~new_n30528_;
  assign new_n30641_ = ~new_n9830_ | ~new_n30532_;
  assign new_n30642_ = ~new_n30598_ | ~new_n30561_;
  assign new_n30643_ = ~new_n10681_ | ~new_n30531_;
  assign new_n30644_ = ~new_n30597_ | ~new_n30563_;
  assign new_n30645_ = ~new_n10683_ | ~new_n30530_;
  assign new_n30646_ = ~new_n30596_ | ~new_n30565_;
  assign new_n30647_ = ~new_n9807_ | ~new_n30568_;
  assign new_n30648_ = ~new_n30618_ | ~new_n30567_;
  assign new_n30649_ = ~new_n10685_ | ~new_n30529_;
  assign new_n30650_ = ~new_n30595_ | ~new_n30570_;
  assign new_n30651_ = ~new_n9810_ | ~new_n30545_;
  assign new_n30652_ = ~new_n30616_ | ~new_n30572_;
  assign new_n30653_ = ~new_n9812_ | ~new_n30544_;
  assign new_n30654_ = ~new_n30615_ | ~new_n30574_;
  assign new_n30655_ = ~new_n9814_ | ~new_n30543_;
  assign new_n30656_ = ~new_n30614_ | ~new_n30576_;
  assign new_n30657_ = ~new_n9816_ | ~new_n30542_;
  assign new_n30658_ = ~new_n30613_ | ~new_n30578_;
  assign new_n30659_ = ~new_n9818_ | ~new_n30541_;
  assign new_n30660_ = ~new_n30612_ | ~new_n30580_;
  assign new_n30661_ = ~new_n10686_ | ~new_n30583_;
  assign new_n30662_ = ~new_n30594_ | ~new_n30582_;
  assign new_n30663_ = ~new_n9820_ | ~new_n30540_;
  assign new_n30664_ = ~new_n30611_ | ~new_n30584_;
  assign new_n30665_ = ~new_n9822_ | ~new_n30539_;
  assign new_n30666_ = ~new_n30610_ | ~new_n30586_;
  assign new_n30667_ = ~new_n9824_ | ~new_n30538_;
  assign new_n30668_ = ~new_n30609_ | ~new_n30588_;
  assign new_n30669_ = ~new_n9826_ | ~new_n30537_;
  assign new_n30670_ = ~new_n30608_ | ~new_n30590_;
  assign new_n30671_ = ~new_n9828_ | ~new_n30536_;
  assign new_n30672_ = ~new_n30599_ | ~new_n30592_;
  assign new_n30673_ = pi0779 & new_n30679_;
  assign new_n30674_ = pi0776 & pi0775;
  assign new_n30675_ = new_n30758_ & new_n30680_;
  assign new_n30676_ = new_n30679_ & new_n30756_;
  assign new_n30677_ = new_n30678_ & new_n30760_;
  assign new_n30678_ = new_n30675_ & new_n30759_;
  assign new_n30679_ = pi0777 & pi0775 & pi0776 & pi0778;
  assign new_n30680_ = new_n30676_ & new_n30757_;
  assign new_n30681_ = new_n30677_ & new_n30761_;
  assign new_n30682_ = new_n30865_ & new_n30837_;
  assign new_n30683_ = new_n30857_ & new_n30801_;
  assign new_n30684_ = new_n30854_ & new_n30839_;
  assign new_n30685_ = new_n30860_ & new_n30789_;
  assign new_n30686_ = new_n30869_ & new_n30783_;
  assign new_n30687_ = new_n30863_ & new_n30843_;
  assign new_n30688_ = new_n30852_ & new_n30800_;
  assign new_n30689_ = new_n30856_ & new_n30845_;
  assign new_n30690_ = new_n30861_ & new_n30782_;
  assign new_n30691_ = new_n30859_ & new_n30792_;
  assign new_n30692_ = new_n30867_ & new_n30849_;
  assign new_n30693_ = new_n30851_ & new_n30781_;
  assign new_n30694_ = ~new_n30873_ | ~new_n30938_ | ~new_n30937_;
  assign new_n30695_ = ~pi0766;
  assign new_n30696_ = ~new_n29445_;
  assign new_n30697_ = ~pi0767;
  assign new_n30698_ = ~new_n29445_ | ~pi0766;
  assign new_n30699_ = ~new_n29428_;
  assign new_n30700_ = ~new_n29446_;
  assign new_n30701_ = ~pi0768;
  assign new_n30702_ = ~new_n29450_;
  assign new_n30703_ = ~pi0769;
  assign new_n30704_ = ~new_n29444_;
  assign new_n30705_ = ~pi0770;
  assign new_n30706_ = ~new_n29443_;
  assign new_n30707_ = ~pi0771;
  assign new_n30708_ = ~pi0772;
  assign new_n30709_ = ~new_n29442_;
  assign new_n30710_ = ~new_n29429_;
  assign new_n30711_ = ~pi0774;
  assign new_n30712_ = ~new_n29441_;
  assign new_n30713_ = ~pi0773;
  assign new_n30714_ = ~pi0775;
  assign new_n30715_ = ~pi0776;
  assign new_n30716_ = ~pi0777;
  assign new_n30717_ = ~pi0778;
  assign new_n30718_ = ~pi0779;
  assign new_n30719_ = ~pi0780;
  assign new_n30720_ = ~pi0781;
  assign new_n30721_ = ~pi0782;
  assign new_n30722_ = ~pi0784;
  assign new_n30723_ = ~pi0783;
  assign new_n30724_ = ~pi0785;
  assign new_n30725_ = ~pi0786;
  assign new_n30726_ = ~pi0787;
  assign new_n30727_ = ~pi0788;
  assign new_n30728_ = ~pi0789;
  assign new_n30729_ = ~pi0790;
  assign new_n30730_ = ~pi0792;
  assign new_n30731_ = ~pi0791;
  assign new_n30732_ = ~pi0793;
  assign new_n30733_ = ~pi0794;
  assign new_n30734_ = ~pi0795;
  assign new_n30735_ = ~pi0796;
  assign new_n30736_ = ~new_n29428_ | ~new_n30806_;
  assign new_n30737_ = ~new_n30875_ | ~new_n30874_;
  assign new_n30738_ = ~new_n30884_ | ~new_n30883_;
  assign new_n30739_ = ~new_n30886_ | ~new_n30885_;
  assign new_n30740_ = ~new_n30888_ | ~new_n30887_;
  assign new_n30741_ = ~new_n30899_ | ~new_n30898_;
  assign new_n30742_ = ~new_n30901_ | ~new_n30900_;
  assign new_n30743_ = ~new_n30910_ | ~new_n30909_;
  assign new_n30744_ = ~new_n30940_ | ~new_n30939_;
  assign new_n30745_ = ~new_n30942_ | ~new_n30941_;
  assign new_n30746_ = ~new_n30951_ | ~new_n30950_;
  assign new_n30747_ = ~new_n30882_ | ~new_n30881_;
  assign new_n30748_ = ~new_n30895_ | ~new_n30894_;
  assign new_n30749_ = ~new_n30908_ | ~new_n30907_;
  assign new_n30750_ = ~new_n30917_ | ~new_n30916_;
  assign new_n30751_ = ~new_n30924_ | ~new_n30923_;
  assign new_n30752_ = ~new_n30926_ | ~new_n30925_;
  assign new_n30753_ = ~new_n30933_ | ~new_n30932_;
  assign new_n30754_ = ~new_n30949_ | ~new_n30948_;
  assign new_n30755_ = new_n30872_ & new_n30835_;
  assign new_n30756_ = pi0779 & pi0781 & pi0780;
  assign new_n30757_ = pi0782 & pi0783 & pi0784;
  assign new_n30758_ = pi0785 & pi0786;
  assign new_n30759_ = pi0787 & pi0789 & pi0788;
  assign new_n30760_ = pi0790 & pi0791 & pi0792;
  assign new_n30761_ = pi0793 & pi0795 & pi0794;
  assign new_n30762_ = new_n30677_ & new_n30763_;
  assign new_n30763_ = pi0794 & pi0793;
  assign new_n30764_ = new_n30676_ & pi0782;
  assign new_n30765_ = new_n30680_ & pi0785;
  assign new_n30766_ = new_n30675_ & new_n30767_;
  assign new_n30767_ = pi0788 & pi0787;
  assign new_n30768_ = new_n30675_ & pi0787;
  assign new_n30769_ = new_n30676_ & new_n30770_;
  assign new_n30770_ = pi0783 & pi0782;
  assign new_n30771_ = pi0777 & new_n30674_;
  assign new_n30772_ = new_n30678_ & new_n30773_;
  assign new_n30773_ = pi0791 & pi0790;
  assign new_n30774_ = pi0780 & new_n30673_;
  assign new_n30775_ = new_n30681_ & pi0796;
  assign new_n30776_ = new_n30681_ & pi0796;
  assign new_n30777_ = new_n30677_ & pi0793;
  assign new_n30778_ = new_n30678_ & pi0790;
  assign new_n30779_ = new_n30877_ & new_n30876_;
  assign new_n30780_ = ~new_n30824_ | ~new_n30823_;
  assign new_n30781_ = ~new_n30681_ | ~new_n30786_;
  assign new_n30782_ = ~new_n30678_ | ~new_n30786_;
  assign new_n30783_ = ~new_n30764_ | ~new_n30786_;
  assign new_n30784_ = new_n30890_ & new_n30889_;
  assign new_n30785_ = ~new_n30736_ | ~new_n30808_;
  assign new_n30786_ = ~new_n30755_ | ~new_n30871_;
  assign new_n30787_ = new_n30897_ & new_n30896_;
  assign new_n30788_ = ~new_n30786_ | ~new_n30769_;
  assign new_n30789_ = ~new_n30774_ | ~new_n30786_;
  assign new_n30790_ = new_n30903_ & new_n30902_;
  assign new_n30791_ = ~new_n30816_ | ~new_n30815_;
  assign new_n30792_ = ~new_n30677_ | ~new_n30786_;
  assign new_n30793_ = new_n30912_ & new_n30911_;
  assign new_n30794_ = ~new_n30820_ | ~new_n30819_;
  assign new_n30795_ = new_n30919_ & new_n30918_;
  assign new_n30796_ = ~new_n30832_ | ~new_n30831_;
  assign new_n30797_ = ~pi0797;
  assign new_n30798_ = new_n30928_ & new_n30927_;
  assign new_n30799_ = ~new_n30812_ | ~new_n30811_;
  assign new_n30800_ = ~new_n30675_ | ~new_n30786_;
  assign new_n30801_ = ~new_n30771_ | ~new_n30786_;
  assign new_n30802_ = new_n30944_ & new_n30943_;
  assign new_n30803_ = ~new_n30828_ | ~new_n30827_;
  assign new_n30804_ = ~new_n30778_ | ~new_n30786_;
  assign new_n30805_ = ~new_n30736_;
  assign new_n30806_ = ~new_n30698_;
  assign new_n30807_ = ~new_n30699_ | ~new_n30698_;
  assign new_n30808_ = ~pi0767 | ~new_n30807_;
  assign new_n30809_ = ~new_n30785_;
  assign new_n30810_ = new_n29446_ | pi0768;
  assign new_n30811_ = ~new_n30810_ | ~new_n30785_;
  assign new_n30812_ = ~pi0768 | ~new_n29446_;
  assign new_n30813_ = ~new_n30799_;
  assign new_n30814_ = new_n29450_ | pi0769;
  assign new_n30815_ = ~new_n30814_ | ~new_n30799_;
  assign new_n30816_ = ~pi0769 | ~new_n29450_;
  assign new_n30817_ = ~new_n30791_;
  assign new_n30818_ = new_n29444_ | pi0770;
  assign new_n30819_ = ~new_n30818_ | ~new_n30791_;
  assign new_n30820_ = ~pi0770 | ~new_n29444_;
  assign new_n30821_ = ~new_n30794_;
  assign new_n30822_ = new_n29443_ | pi0771;
  assign new_n30823_ = ~new_n30822_ | ~new_n30794_;
  assign new_n30824_ = ~pi0771 | ~new_n29443_;
  assign new_n30825_ = ~new_n30780_;
  assign new_n30826_ = new_n29442_ | pi0772;
  assign new_n30827_ = ~new_n30826_ | ~new_n30780_;
  assign new_n30828_ = ~new_n29442_ | ~pi0772;
  assign new_n30829_ = ~new_n30803_;
  assign new_n30830_ = new_n29441_ | pi0773;
  assign new_n30831_ = ~new_n30830_ | ~new_n30803_;
  assign new_n30832_ = ~pi0773 | ~new_n29441_;
  assign new_n30833_ = ~new_n30796_;
  assign new_n30834_ = new_n29429_ | pi0774;
  assign new_n30835_ = ~pi0774 | ~new_n29429_;
  assign new_n30836_ = ~new_n30786_;
  assign new_n30837_ = ~new_n30674_ | ~new_n30786_;
  assign new_n30838_ = ~new_n30801_;
  assign new_n30839_ = ~new_n30673_ | ~new_n30786_;
  assign new_n30840_ = ~new_n30789_;
  assign new_n30841_ = ~new_n30783_;
  assign new_n30842_ = ~new_n30788_;
  assign new_n30843_ = ~new_n30765_ | ~new_n30786_;
  assign new_n30844_ = ~new_n30800_;
  assign new_n30845_ = ~new_n30786_ | ~new_n30766_;
  assign new_n30846_ = ~new_n30782_;
  assign new_n30847_ = ~new_n30804_;
  assign new_n30848_ = ~new_n30792_;
  assign new_n30849_ = ~new_n30786_ | ~new_n30762_;
  assign new_n30850_ = ~new_n30781_;
  assign new_n30851_ = ~new_n30734_ | ~new_n30849_;
  assign new_n30852_ = ~new_n30725_ | ~new_n30843_;
  assign new_n30853_ = ~new_n30679_ | ~new_n30786_;
  assign new_n30854_ = ~new_n30718_ | ~new_n30853_;
  assign new_n30855_ = ~new_n30768_ | ~new_n30786_;
  assign new_n30856_ = ~new_n30727_ | ~new_n30855_;
  assign new_n30857_ = ~new_n30716_ | ~new_n30837_;
  assign new_n30858_ = ~new_n30786_ | ~new_n30772_;
  assign new_n30859_ = ~new_n30730_ | ~new_n30858_;
  assign new_n30860_ = ~new_n30719_ | ~new_n30839_;
  assign new_n30861_ = ~new_n30728_ | ~new_n30845_;
  assign new_n30862_ = ~new_n30680_ | ~new_n30786_;
  assign new_n30863_ = ~new_n30724_ | ~new_n30862_;
  assign new_n30864_ = ~pi0775 | ~new_n30786_;
  assign new_n30865_ = ~new_n30715_ | ~new_n30864_;
  assign new_n30866_ = ~new_n30777_ | ~new_n30786_;
  assign new_n30867_ = ~new_n30733_ | ~new_n30866_;
  assign new_n30868_ = ~new_n30676_ | ~new_n30786_;
  assign new_n30869_ = ~new_n30721_ | ~new_n30868_;
  assign new_n30870_ = ~new_n30776_ | ~new_n30786_;
  assign new_n30871_ = ~new_n30830_ | ~new_n30834_ | ~new_n30803_;
  assign new_n30872_ = ~new_n29441_ | ~pi0773 | ~new_n30834_;
  assign new_n30873_ = ~new_n30805_ | ~pi0767;
  assign new_n30874_ = ~pi0766 | ~new_n30696_;
  assign new_n30875_ = ~new_n29445_ | ~new_n30695_;
  assign new_n30876_ = ~pi0772 | ~new_n30709_;
  assign new_n30877_ = ~new_n29442_ | ~new_n30708_;
  assign new_n30878_ = ~pi0772 | ~new_n30709_;
  assign new_n30879_ = ~new_n29442_ | ~new_n30708_;
  assign new_n30880_ = ~new_n30879_ | ~new_n30878_;
  assign new_n30881_ = ~new_n30779_ | ~new_n30780_;
  assign new_n30882_ = ~new_n30825_ | ~new_n30880_;
  assign new_n30883_ = ~pi0796 | ~new_n30781_;
  assign new_n30884_ = ~new_n30850_ | ~new_n30735_;
  assign new_n30885_ = ~pi0790 | ~new_n30782_;
  assign new_n30886_ = ~new_n30846_ | ~new_n30729_;
  assign new_n30887_ = ~pi0783 | ~new_n30783_;
  assign new_n30888_ = ~new_n30841_ | ~new_n30723_;
  assign new_n30889_ = ~pi0768 | ~new_n30700_;
  assign new_n30890_ = ~new_n29446_ | ~new_n30701_;
  assign new_n30891_ = ~pi0768 | ~new_n30700_;
  assign new_n30892_ = ~new_n29446_ | ~new_n30701_;
  assign new_n30893_ = ~new_n30892_ | ~new_n30891_;
  assign new_n30894_ = ~new_n30784_ | ~new_n30785_;
  assign new_n30895_ = ~new_n30809_ | ~new_n30893_;
  assign new_n30896_ = ~pi0775 | ~new_n30786_;
  assign new_n30897_ = ~new_n30836_ | ~new_n30714_;
  assign new_n30898_ = ~pi0784 | ~new_n30788_;
  assign new_n30899_ = ~new_n30842_ | ~new_n30722_;
  assign new_n30900_ = ~pi0781 | ~new_n30789_;
  assign new_n30901_ = ~new_n30840_ | ~new_n30720_;
  assign new_n30902_ = ~pi0770 | ~new_n30704_;
  assign new_n30903_ = ~new_n29444_ | ~new_n30705_;
  assign new_n30904_ = ~pi0770 | ~new_n30704_;
  assign new_n30905_ = ~new_n29444_ | ~new_n30705_;
  assign new_n30906_ = ~new_n30905_ | ~new_n30904_;
  assign new_n30907_ = ~new_n30790_ | ~new_n30791_;
  assign new_n30908_ = ~new_n30817_ | ~new_n30906_;
  assign new_n30909_ = ~pi0793 | ~new_n30792_;
  assign new_n30910_ = ~new_n30848_ | ~new_n30732_;
  assign new_n30911_ = ~pi0771 | ~new_n30706_;
  assign new_n30912_ = ~new_n29443_ | ~new_n30707_;
  assign new_n30913_ = ~pi0771 | ~new_n30706_;
  assign new_n30914_ = ~new_n29443_ | ~new_n30707_;
  assign new_n30915_ = ~new_n30914_ | ~new_n30913_;
  assign new_n30916_ = ~new_n30793_ | ~new_n30794_;
  assign new_n30917_ = ~new_n30821_ | ~new_n30915_;
  assign new_n30918_ = ~pi0774 | ~new_n30710_;
  assign new_n30919_ = ~new_n29429_ | ~new_n30711_;
  assign new_n30920_ = ~pi0774 | ~new_n30710_;
  assign new_n30921_ = ~new_n29429_ | ~new_n30711_;
  assign new_n30922_ = ~new_n30921_ | ~new_n30920_;
  assign new_n30923_ = ~new_n30795_ | ~new_n30796_;
  assign new_n30924_ = ~new_n30833_ | ~new_n30922_;
  assign new_n30925_ = ~pi0797 | ~new_n30870_;
  assign new_n30926_ = ~new_n30797_ | ~new_n30775_ | ~new_n30786_;
  assign new_n30927_ = ~pi0769 | ~new_n30702_;
  assign new_n30928_ = ~new_n29450_ | ~new_n30703_;
  assign new_n30929_ = ~pi0769 | ~new_n30702_;
  assign new_n30930_ = ~new_n29450_ | ~new_n30703_;
  assign new_n30931_ = ~new_n30930_ | ~new_n30929_;
  assign new_n30932_ = ~new_n30798_ | ~new_n30799_;
  assign new_n30933_ = ~new_n30813_ | ~new_n30931_;
  assign new_n30934_ = ~pi0767 | ~new_n30698_;
  assign new_n30935_ = ~new_n30806_ | ~new_n30697_;
  assign new_n30936_ = ~new_n30935_ | ~new_n30934_;
  assign new_n30937_ = ~new_n29428_ | ~new_n30698_ | ~new_n30697_;
  assign new_n30938_ = ~new_n30936_ | ~new_n30699_;
  assign new_n30939_ = ~pi0787 | ~new_n30800_;
  assign new_n30940_ = ~new_n30844_ | ~new_n30726_;
  assign new_n30941_ = ~pi0778 | ~new_n30801_;
  assign new_n30942_ = ~new_n30838_ | ~new_n30717_;
  assign new_n30943_ = ~pi0773 | ~new_n30712_;
  assign new_n30944_ = ~new_n29441_ | ~new_n30713_;
  assign new_n30945_ = ~pi0773 | ~new_n30712_;
  assign new_n30946_ = ~new_n29441_ | ~new_n30713_;
  assign new_n30947_ = ~new_n30946_ | ~new_n30945_;
  assign new_n30948_ = ~new_n30802_ | ~new_n30803_;
  assign new_n30949_ = ~new_n30829_ | ~new_n30947_;
  assign new_n30950_ = ~pi0791 | ~new_n30804_;
  assign new_n30951_ = ~new_n30847_ | ~new_n30731_;
  assign new_n30952_ = ~pi1215;
  assign new_n30953_ = ~pi1217;
  assign new_n30954_ = ~pi1216;
  assign new_n30955_ = ~pi1219;
  assign new_n30956_ = ~pi1218;
  assign new_n30957_ = ~pi1216 | ~pi1217 | ~pi1215;
  assign new_n30958_ = ~pi1221;
  assign new_n30959_ = ~pi1220;
  assign new_n30960_ = ~new_n31029_ | ~new_n31058_;
  assign new_n30961_ = ~pi1223;
  assign new_n30962_ = ~pi1222;
  assign new_n30963_ = ~new_n31030_ | ~new_n31059_;
  assign new_n30964_ = ~new_n31031_ | ~new_n31065_;
  assign new_n30965_ = ~pi1224;
  assign new_n30966_ = ~pi1225;
  assign new_n30967_ = ~pi1227;
  assign new_n30968_ = ~pi1226;
  assign new_n30969_ = ~new_n31032_ | ~new_n31067_;
  assign new_n30970_ = ~pi1229;
  assign new_n30971_ = ~pi1228;
  assign new_n30972_ = ~new_n31033_ | ~new_n31060_;
  assign new_n30973_ = ~pi1230;
  assign new_n30974_ = ~new_n31034_ | ~new_n31066_;
  assign new_n30975_ = ~pi1231;
  assign new_n30976_ = ~pi1233;
  assign new_n30977_ = ~pi1232;
  assign new_n30978_ = ~new_n31035_ | ~new_n31071_;
  assign new_n30979_ = ~pi1235;
  assign new_n30980_ = ~pi1234;
  assign new_n30981_ = ~new_n31036_ | ~new_n31064_;
  assign new_n30982_ = ~pi1236;
  assign new_n30983_ = ~new_n31037_ | ~new_n31061_;
  assign new_n30984_ = ~pi1237;
  assign new_n30985_ = ~pi1239;
  assign new_n30986_ = ~pi1238;
  assign new_n30987_ = ~new_n31038_ | ~new_n31068_;
  assign new_n30988_ = ~pi1241;
  assign new_n30989_ = ~pi1240;
  assign new_n30990_ = ~new_n31039_ | ~new_n31062_;
  assign new_n30991_ = ~pi1242;
  assign new_n30992_ = ~pi1243;
  assign new_n30993_ = ~new_n31040_ | ~new_n31063_;
  assign new_n30994_ = ~pi1244;
  assign new_n30995_ = ~new_n31041_ | ~new_n31069_;
  assign new_n30996_ = ~new_n31070_ | ~pi1244;
  assign new_n30997_ = ~pi1245;
  assign new_n30998_ = ~new_n31089_ | ~new_n31088_;
  assign new_n30999_ = ~new_n31091_ | ~new_n31090_;
  assign new_n31000_ = ~new_n31093_ | ~new_n31092_;
  assign new_n31001_ = ~new_n31095_ | ~new_n31094_;
  assign new_n31002_ = ~new_n31097_ | ~new_n31096_;
  assign new_n31003_ = ~new_n31099_ | ~new_n31098_;
  assign new_n31004_ = ~new_n31101_ | ~new_n31100_;
  assign new_n31005_ = ~new_n31103_ | ~new_n31102_;
  assign new_n31006_ = ~new_n31105_ | ~new_n31104_;
  assign new_n31007_ = ~new_n31107_ | ~new_n31106_;
  assign new_n31008_ = ~new_n31109_ | ~new_n31108_;
  assign new_n31009_ = ~new_n31111_ | ~new_n31110_;
  assign new_n31010_ = ~new_n31113_ | ~new_n31112_;
  assign new_n31011_ = ~new_n31115_ | ~new_n31114_;
  assign new_n31012_ = ~new_n31117_ | ~new_n31116_;
  assign new_n31013_ = ~new_n31119_ | ~new_n31118_;
  assign new_n31014_ = ~new_n31121_ | ~new_n31120_;
  assign new_n31015_ = ~new_n31123_ | ~new_n31122_;
  assign new_n31016_ = ~new_n31125_ | ~new_n31124_;
  assign new_n31017_ = ~new_n31127_ | ~new_n31126_;
  assign new_n31018_ = ~new_n31129_ | ~new_n31128_;
  assign new_n31019_ = ~new_n31131_ | ~new_n31130_;
  assign new_n31020_ = ~new_n31133_ | ~new_n31132_;
  assign new_n31021_ = ~new_n31135_ | ~new_n31134_;
  assign new_n31022_ = ~new_n31137_ | ~new_n31136_;
  assign new_n31023_ = ~new_n31139_ | ~new_n31138_;
  assign new_n31024_ = ~new_n31141_ | ~new_n31140_;
  assign new_n31025_ = ~new_n31143_ | ~new_n31142_;
  assign new_n31026_ = ~new_n31145_ | ~new_n31144_;
  assign new_n31027_ = ~new_n31147_ | ~new_n31146_;
  assign new_n31028_ = ~new_n31149_ | ~new_n31148_;
  assign new_n31029_ = pi1218 & pi1219;
  assign new_n31030_ = pi1220 & pi1221;
  assign new_n31031_ = pi1222 & pi1223;
  assign new_n31032_ = pi1224 & pi1225;
  assign new_n31033_ = pi1226 & pi1227;
  assign new_n31034_ = pi1228 & pi1229;
  assign new_n31035_ = pi1231 & pi1230;
  assign new_n31036_ = pi1232 & pi1233;
  assign new_n31037_ = pi1234 & pi1235;
  assign new_n31038_ = pi1237 & pi1236;
  assign new_n31039_ = pi1238 & pi1239;
  assign new_n31040_ = pi1240 & pi1241;
  assign new_n31041_ = pi1243 & pi1242;
  assign new_n31042_ = ~new_n31065_ | ~pi1222;
  assign new_n31043_ = ~new_n31059_ | ~pi1220;
  assign new_n31044_ = ~new_n31058_ | ~pi1218;
  assign new_n31045_ = ~pi1246;
  assign new_n31046_ = ~pi1245 | ~new_n31075_;
  assign new_n31047_ = ~pi1216 | ~pi1215;
  assign new_n31048_ = ~new_n31069_ | ~pi1242;
  assign new_n31049_ = ~new_n31063_ | ~pi1240;
  assign new_n31050_ = ~new_n31062_ | ~pi1238;
  assign new_n31051_ = ~new_n31068_ | ~pi1236;
  assign new_n31052_ = ~new_n31061_ | ~pi1234;
  assign new_n31053_ = ~new_n31064_ | ~pi1232;
  assign new_n31054_ = ~new_n31071_ | ~pi1230;
  assign new_n31055_ = ~new_n31066_ | ~pi1228;
  assign new_n31056_ = ~new_n31060_ | ~pi1226;
  assign new_n31057_ = ~pi1224 | ~new_n31067_;
  assign new_n31058_ = ~new_n30957_;
  assign new_n31059_ = ~new_n30960_;
  assign new_n31060_ = ~new_n30969_;
  assign new_n31061_ = ~new_n30981_;
  assign new_n31062_ = ~new_n30987_;
  assign new_n31063_ = ~new_n30990_;
  assign new_n31064_ = ~new_n30978_;
  assign new_n31065_ = ~new_n30963_;
  assign new_n31066_ = ~new_n30972_;
  assign new_n31067_ = ~new_n30964_;
  assign new_n31068_ = ~new_n30983_;
  assign new_n31069_ = ~new_n30993_;
  assign new_n31070_ = ~new_n30995_;
  assign new_n31071_ = ~new_n30974_;
  assign new_n31072_ = ~new_n31042_;
  assign new_n31073_ = ~new_n31043_;
  assign new_n31074_ = ~new_n31044_;
  assign new_n31075_ = ~new_n30996_;
  assign new_n31076_ = ~new_n31046_;
  assign new_n31077_ = ~new_n31047_;
  assign new_n31078_ = ~new_n31048_;
  assign new_n31079_ = ~new_n31049_;
  assign new_n31080_ = ~new_n31050_;
  assign new_n31081_ = ~new_n31051_;
  assign new_n31082_ = ~new_n31052_;
  assign new_n31083_ = ~new_n31053_;
  assign new_n31084_ = ~new_n31054_;
  assign new_n31085_ = ~new_n31055_;
  assign new_n31086_ = ~new_n31056_;
  assign new_n31087_ = ~new_n31057_;
  assign new_n31088_ = ~new_n31067_ | ~new_n30965_;
  assign new_n31089_ = ~pi1224 | ~new_n30964_;
  assign new_n31090_ = ~pi1223 | ~new_n31042_;
  assign new_n31091_ = ~new_n31072_ | ~new_n30961_;
  assign new_n31092_ = ~new_n31065_ | ~new_n30962_;
  assign new_n31093_ = ~pi1222 | ~new_n30963_;
  assign new_n31094_ = ~pi1221 | ~new_n31043_;
  assign new_n31095_ = ~new_n31073_ | ~new_n30958_;
  assign new_n31096_ = ~new_n31059_ | ~new_n30959_;
  assign new_n31097_ = ~pi1220 | ~new_n30960_;
  assign new_n31098_ = ~pi1219 | ~new_n31044_;
  assign new_n31099_ = ~new_n31074_ | ~new_n30955_;
  assign new_n31100_ = ~new_n31058_ | ~new_n30956_;
  assign new_n31101_ = ~pi1218 | ~new_n30957_;
  assign new_n31102_ = ~pi1246 | ~new_n31046_;
  assign new_n31103_ = ~new_n31076_ | ~new_n31045_;
  assign new_n31104_ = ~pi1245 | ~new_n30996_;
  assign new_n31105_ = ~new_n31075_ | ~new_n30997_;
  assign new_n31106_ = ~pi1217 | ~new_n31047_;
  assign new_n31107_ = ~new_n31077_ | ~new_n30953_;
  assign new_n31108_ = ~new_n31070_ | ~new_n30994_;
  assign new_n31109_ = ~pi1244 | ~new_n30995_;
  assign new_n31110_ = ~pi1243 | ~new_n31048_;
  assign new_n31111_ = ~new_n31078_ | ~new_n30992_;
  assign new_n31112_ = ~new_n31069_ | ~new_n30991_;
  assign new_n31113_ = ~pi1242 | ~new_n30993_;
  assign new_n31114_ = ~pi1241 | ~new_n31049_;
  assign new_n31115_ = ~new_n31079_ | ~new_n30988_;
  assign new_n31116_ = ~new_n31063_ | ~new_n30989_;
  assign new_n31117_ = ~pi1240 | ~new_n30990_;
  assign new_n31118_ = ~pi1239 | ~new_n31050_;
  assign new_n31119_ = ~new_n31080_ | ~new_n30985_;
  assign new_n31120_ = ~new_n31062_ | ~new_n30986_;
  assign new_n31121_ = ~pi1238 | ~new_n30987_;
  assign new_n31122_ = ~pi1237 | ~new_n31051_;
  assign new_n31123_ = ~new_n31081_ | ~new_n30984_;
  assign new_n31124_ = ~new_n31068_ | ~new_n30982_;
  assign new_n31125_ = ~pi1236 | ~new_n30983_;
  assign new_n31126_ = ~pi1235 | ~new_n31052_;
  assign new_n31127_ = ~new_n31082_ | ~new_n30979_;
  assign new_n31128_ = ~pi1215 | ~new_n30954_;
  assign new_n31129_ = ~pi1216 | ~new_n30952_;
  assign new_n31130_ = ~new_n31061_ | ~new_n30980_;
  assign new_n31131_ = ~pi1234 | ~new_n30981_;
  assign new_n31132_ = ~pi1233 | ~new_n31053_;
  assign new_n31133_ = ~new_n31083_ | ~new_n30976_;
  assign new_n31134_ = ~new_n31064_ | ~new_n30977_;
  assign new_n31135_ = ~pi1232 | ~new_n30978_;
  assign new_n31136_ = ~pi1231 | ~new_n31054_;
  assign new_n31137_ = ~new_n31084_ | ~new_n30975_;
  assign new_n31138_ = ~new_n31071_ | ~new_n30973_;
  assign new_n31139_ = ~pi1230 | ~new_n30974_;
  assign new_n31140_ = ~pi1229 | ~new_n31055_;
  assign new_n31141_ = ~new_n31085_ | ~new_n30970_;
  assign new_n31142_ = ~new_n31066_ | ~new_n30971_;
  assign new_n31143_ = ~pi1228 | ~new_n30972_;
  assign new_n31144_ = ~pi1227 | ~new_n31056_;
  assign new_n31145_ = ~new_n31086_ | ~new_n30967_;
  assign new_n31146_ = ~new_n31060_ | ~new_n30968_;
  assign new_n31147_ = ~pi1226 | ~new_n30969_;
  assign new_n31148_ = ~pi1225 | ~new_n31057_;
  assign new_n31149_ = ~new_n31087_ | ~new_n30966_;
  assign new_n31150_ = new_n31192_ & new_n15921_;
  assign new_n31151_ = new_n31205_ & new_n31161_;
  assign new_n31152_ = ~new_n15925_;
  assign new_n31153_ = ~new_n16427_;
  assign new_n31154_ = ~new_n16427_ | ~new_n15925_;
  assign new_n31155_ = ~new_n15923_;
  assign new_n31156_ = ~new_n15922_;
  assign new_n31157_ = ~new_n15921_;
  assign new_n31158_ = ~new_n31180_ | ~new_n31186_;
  assign new_n31159_ = ~new_n15918_;
  assign new_n31160_ = ~new_n15919_;
  assign new_n31161_ = ~new_n15904_ | ~new_n15920_;
  assign new_n31162_ = ~new_n15917_;
  assign new_n31163_ = ~new_n15916_;
  assign new_n31164_ = ~new_n31181_ | ~new_n31194_;
  assign new_n31165_ = ~new_n15915_;
  assign new_n31166_ = ~new_n31182_ | ~new_n31191_;
  assign new_n31167_ = ~new_n31193_ | ~new_n15915_;
  assign new_n31168_ = ~new_n15914_;
  assign new_n31169_ = ~new_n31209_ | ~new_n31208_;
  assign new_n31170_ = ~new_n31211_ | ~new_n31210_;
  assign new_n31171_ = ~new_n31213_ | ~new_n31212_;
  assign new_n31172_ = ~new_n31217_ | ~new_n31216_;
  assign new_n31173_ = ~new_n31219_ | ~new_n31218_;
  assign new_n31174_ = ~new_n31221_ | ~new_n31220_;
  assign new_n31175_ = ~new_n31223_ | ~new_n31222_;
  assign new_n31176_ = ~new_n31225_ | ~new_n31224_;
  assign new_n31177_ = ~new_n31227_ | ~new_n31226_;
  assign new_n31178_ = ~new_n31229_ | ~new_n31228_;
  assign new_n31179_ = ~new_n31231_ | ~new_n31230_;
  assign new_n31180_ = new_n15923_ & new_n15922_;
  assign new_n31181_ = new_n15919_ & new_n15918_;
  assign new_n31182_ = new_n15916_ & new_n15917_;
  assign new_n31183_ = ~new_n15923_ | ~new_n31186_;
  assign new_n31184_ = ~new_n15913_;
  assign new_n31185_ = ~new_n15914_ | ~new_n31201_;
  assign new_n31186_ = ~new_n31197_ | ~new_n31198_;
  assign new_n31187_ = new_n31215_ & new_n31214_;
  assign new_n31188_ = ~new_n31191_ | ~new_n15917_;
  assign new_n31189_ = ~new_n31194_ | ~new_n15919_;
  assign new_n31190_ = ~new_n31196_ | ~new_n31207_;
  assign new_n31191_ = ~new_n31164_;
  assign new_n31192_ = ~new_n31158_;
  assign new_n31193_ = ~new_n31166_;
  assign new_n31194_ = ~new_n31161_;
  assign new_n31195_ = ~new_n31154_;
  assign new_n31196_ = new_n15924_ | new_n15912_;
  assign new_n31197_ = ~new_n15912_ | ~new_n15924_;
  assign new_n31198_ = ~new_n31195_ | ~new_n31196_;
  assign new_n31199_ = ~new_n31186_;
  assign new_n31200_ = ~new_n31183_;
  assign new_n31201_ = ~new_n31167_;
  assign new_n31202_ = ~new_n31185_;
  assign new_n31203_ = ~new_n31188_;
  assign new_n31204_ = ~new_n31189_;
  assign new_n31205_ = new_n15920_ | new_n15904_;
  assign new_n31206_ = ~new_n31190_;
  assign new_n31207_ = ~new_n15912_ | ~new_n15924_;
  assign new_n31208_ = ~new_n31192_ | ~new_n31157_;
  assign new_n31209_ = ~new_n15921_ | ~new_n31158_;
  assign new_n31210_ = ~new_n15922_ | ~new_n31183_;
  assign new_n31211_ = ~new_n31200_ | ~new_n31156_;
  assign new_n31212_ = ~new_n15913_ | ~new_n31185_;
  assign new_n31213_ = ~new_n31202_ | ~new_n31184_;
  assign new_n31214_ = ~new_n15923_ | ~new_n31186_;
  assign new_n31215_ = ~new_n31199_ | ~new_n31155_;
  assign new_n31216_ = ~new_n15914_ | ~new_n31167_;
  assign new_n31217_ = ~new_n31201_ | ~new_n31168_;
  assign new_n31218_ = ~new_n31193_ | ~new_n31165_;
  assign new_n31219_ = ~new_n15915_ | ~new_n31166_;
  assign new_n31220_ = ~new_n15916_ | ~new_n31188_;
  assign new_n31221_ = ~new_n31203_ | ~new_n31163_;
  assign new_n31222_ = ~new_n31191_ | ~new_n31162_;
  assign new_n31223_ = ~new_n15917_ | ~new_n31164_;
  assign new_n31224_ = ~new_n15918_ | ~new_n31189_;
  assign new_n31225_ = ~new_n31204_ | ~new_n31159_;
  assign new_n31226_ = ~new_n31194_ | ~new_n31160_;
  assign new_n31227_ = ~new_n15919_ | ~new_n31161_;
  assign new_n31228_ = ~new_n31195_ | ~new_n31190_;
  assign new_n31229_ = ~new_n31206_ | ~new_n31154_;
  assign new_n31230_ = ~new_n16427_ | ~new_n31152_;
  assign new_n31231_ = ~new_n15925_ | ~new_n31153_;
  assign new_n31232_ = new_n31331_ & new_n31330_;
  assign new_n31233_ = new_n31262_ & new_n31256_ & new_n31254_ & new_n31263_;
  assign new_n31234_ = new_n31331_ & new_n31308_;
  assign new_n31235_ = new_n31365_ & new_n31363_;
  assign new_n31236_ = new_n31355_ & new_n31354_;
  assign new_n31237_ = new_n31309_ & new_n31440_ & new_n31439_;
  assign new_n31238_ = ~new_n31371_ | ~new_n31373_;
  assign new_n31239_ = ~new_n15536_;
  assign new_n31240_ = ~new_n15931_;
  assign new_n31241_ = ~new_n15932_;
  assign new_n31242_ = ~new_n15933_;
  assign new_n31243_ = ~new_n15930_;
  assign new_n31244_ = ~new_n15926_;
  assign new_n31245_ = ~new_n15929_;
  assign new_n31246_ = ~new_n15929_ | ~new_n31405_;
  assign new_n31247_ = ~new_n15928_;
  assign new_n31248_ = ~new_n15928_ | ~new_n31397_;
  assign new_n31249_ = ~new_n15927_;
  assign new_n31250_ = ~new_n15927_ | ~new_n31400_;
  assign new_n31251_ = ~new_n31306_ | ~new_n31290_;
  assign new_n31252_ = ~new_n31233_ | ~new_n31306_;
  assign new_n31253_ = ~new_n31292_ | ~new_n31368_;
  assign new_n31254_ = ~new_n31433_ | ~new_n31432_;
  assign new_n31255_ = ~new_n31413_ | ~new_n31412_;
  assign new_n31256_ = ~new_n31430_ | ~new_n31429_;
  assign new_n31257_ = ~new_n31436_ | ~new_n31435_;
  assign new_n31258_ = ~new_n31451_ | ~new_n31450_;
  assign new_n31259_ = ~new_n31448_ | ~new_n31447_;
  assign new_n31260_ = ~new_n31454_ | ~new_n31453_;
  assign new_n31261_ = ~new_n31457_ | ~new_n31456_;
  assign new_n31262_ = ~new_n31460_ | ~new_n31459_;
  assign new_n31263_ = ~new_n31463_ | ~new_n31462_;
  assign new_n31264_ = ~new_n31475_ | ~new_n31474_;
  assign new_n31265_ = ~new_n31477_ | ~new_n31476_;
  assign new_n31266_ = ~new_n31479_ | ~new_n31478_;
  assign new_n31267_ = ~new_n31481_ | ~new_n31480_;
  assign new_n31268_ = ~new_n31483_ | ~new_n31482_;
  assign new_n31269_ = ~new_n31485_ | ~new_n31484_;
  assign new_n31270_ = ~new_n31487_ | ~new_n31486_;
  assign new_n31271_ = new_n31248_ & new_n31332_;
  assign new_n31272_ = ~new_n31444_ | ~new_n31443_;
  assign new_n31273_ = new_n31246_ & new_n31333_;
  assign new_n31274_ = ~new_n31446_ | ~new_n31445_;
  assign new_n31275_ = new_n31389_ & new_n31336_;
  assign new_n31276_ = ~new_n31466_ | ~new_n31465_;
  assign new_n31277_ = ~new_n31473_ | ~new_n31472_;
  assign new_n31278_ = new_n31337_ & new_n31336_;
  assign new_n31279_ = new_n31333_ & new_n31332_;
  assign new_n31280_ = new_n31234_ & new_n31279_;
  assign new_n31281_ = new_n31378_ & new_n31379_ & new_n31380_ & new_n31330_;
  assign new_n31282_ = new_n31336_ & new_n31333_;
  assign new_n31283_ = new_n31386_ & new_n31246_;
  assign new_n31284_ = new_n31383_ & new_n31248_;
  assign new_n31285_ = new_n31386_ & new_n31246_ & new_n31248_;
  assign new_n31286_ = new_n31232_ & new_n31332_;
  assign new_n31287_ = new_n31353_ & new_n31248_;
  assign new_n31288_ = new_n31250_ & new_n31308_;
  assign new_n31289_ = new_n31338_ & new_n31337_;
  assign new_n31290_ = new_n31233_ & new_n31291_;
  assign new_n31291_ = new_n31260_ & new_n31259_ & new_n31258_ & new_n31261_;
  assign new_n31292_ = new_n31261_ & new_n31260_;
  assign new_n31293_ = new_n31256_ & new_n31263_ & new_n31254_;
  assign new_n31294_ = new_n31256_ & new_n31254_;
  assign new_n31295_ = ~new_n15943_;
  assign new_n31296_ = ~new_n15942_;
  assign new_n31297_ = ~new_n15944_;
  assign new_n31298_ = ~new_n15945_;
  assign new_n31299_ = ~new_n15947_;
  assign new_n31300_ = ~new_n15948_;
  assign new_n31301_ = ~new_n15949_;
  assign new_n31302_ = ~new_n15946_;
  assign new_n31303_ = ~new_n15941_;
  assign new_n31304_ = ~new_n15940_;
  assign new_n31305_ = ~new_n31256_ | ~new_n31306_;
  assign new_n31306_ = ~new_n31326_ | ~new_n31281_;
  assign new_n31307_ = new_n31438_ & new_n31437_;
  assign new_n31308_ = ~new_n31249_ | ~new_n31392_ | ~new_n31391_;
  assign new_n31309_ = new_n31442_ & new_n31441_;
  assign new_n31310_ = ~new_n31283_ | ~new_n31385_;
  assign new_n31311_ = ~new_n31338_ | ~new_n31345_;
  assign new_n31312_ = ~new_n15935_;
  assign new_n31313_ = ~new_n15934_;
  assign new_n31314_ = ~new_n15936_;
  assign new_n31315_ = ~new_n15937_;
  assign new_n31316_ = ~new_n15938_;
  assign new_n31317_ = ~new_n15939_;
  assign new_n31318_ = ~new_n31327_ | ~new_n31359_;
  assign new_n31319_ = new_n31468_ & new_n31467_;
  assign new_n31320_ = ~new_n31356_ | ~new_n31340_;
  assign new_n31321_ = ~new_n31370_ | ~new_n31259_;
  assign new_n31322_ = ~new_n31368_ | ~new_n31261_;
  assign new_n31323_ = ~new_n31306_ | ~new_n31293_;
  assign new_n31324_ = ~new_n31294_ | ~new_n31306_;
  assign new_n31325_ = ~new_n31340_ | ~new_n31339_;
  assign new_n31326_ = ~new_n31280_ | ~new_n31311_;
  assign new_n31327_ = ~new_n15932_ | ~new_n31255_;
  assign new_n31328_ = ~new_n31251_;
  assign new_n31329_ = ~new_n31308_;
  assign new_n31330_ = ~new_n15926_ | ~new_n31408_;
  assign new_n31331_ = ~new_n31244_ | ~new_n31394_ | ~new_n31393_;
  assign new_n31332_ = ~new_n31247_ | ~new_n31402_ | ~new_n31401_;
  assign new_n31333_ = ~new_n31245_ | ~new_n31428_ | ~new_n31427_;
  assign new_n31334_ = ~new_n31248_;
  assign new_n31335_ = ~new_n31250_;
  assign new_n31336_ = ~new_n31240_ | ~new_n31421_ | ~new_n31420_;
  assign new_n31337_ = ~new_n31243_ | ~new_n31423_ | ~new_n31422_;
  assign new_n31338_ = ~new_n15930_ | ~new_n31426_;
  assign new_n31339_ = ~new_n31242_ | ~new_n31416_ | ~new_n31415_;
  assign new_n31340_ = ~new_n15933_ | ~new_n31419_;
  assign new_n31341_ = ~new_n31414_ | ~new_n31241_;
  assign new_n31342_ = ~new_n15536_ | ~new_n31339_;
  assign new_n31343_ = ~new_n15931_ | ~new_n31411_;
  assign new_n31344_ = ~new_n31382_ | ~new_n31384_;
  assign new_n31345_ = ~new_n31278_ | ~new_n31344_;
  assign new_n31346_ = ~new_n31311_;
  assign new_n31347_ = ~new_n31246_;
  assign new_n31348_ = ~new_n31306_;
  assign new_n31349_ = ~new_n31305_;
  assign new_n31350_ = ~new_n31310_;
  assign new_n31351_ = ~new_n31310_ | ~new_n31332_;
  assign new_n31352_ = ~new_n31248_ | ~new_n31351_;
  assign new_n31353_ = ~new_n31250_ | ~new_n31308_;
  assign new_n31354_ = ~new_n31287_ | ~new_n31351_;
  assign new_n31355_ = ~new_n31288_ | ~new_n31352_;
  assign new_n31356_ = ~new_n15536_ | ~new_n31339_;
  assign new_n31357_ = ~new_n31320_;
  assign new_n31358_ = ~new_n31414_ | ~new_n31241_;
  assign new_n31359_ = ~new_n31358_ | ~new_n31320_;
  assign new_n31360_ = ~new_n31318_;
  assign new_n31361_ = ~new_n31318_ | ~new_n31336_;
  assign new_n31362_ = ~new_n31361_ | ~new_n31343_;
  assign new_n31363_ = ~new_n31289_ | ~new_n31362_;
  assign new_n31364_ = ~new_n31388_ | ~new_n31337_;
  assign new_n31365_ = ~new_n31364_ | ~new_n31361_ | ~new_n31343_;
  assign new_n31366_ = ~new_n31324_;
  assign new_n31367_ = ~new_n31323_;
  assign new_n31368_ = ~new_n31252_;
  assign new_n31369_ = ~new_n31322_;
  assign new_n31370_ = ~new_n31253_;
  assign new_n31371_ = ~new_n15536_ | ~new_n31251_;
  assign new_n31372_ = ~new_n31371_;
  assign new_n31373_ = ~new_n31328_ | ~new_n31239_;
  assign new_n31374_ = ~new_n31321_;
  assign new_n31375_ = ~new_n31325_;
  assign new_n31376_ = ~new_n31248_ | ~new_n31332_;
  assign new_n31377_ = ~new_n31246_ | ~new_n31333_;
  assign new_n31378_ = ~new_n31234_ | ~new_n31347_ | ~new_n31332_;
  assign new_n31379_ = ~new_n31334_ | ~new_n31234_;
  assign new_n31380_ = ~new_n31335_ | ~new_n31234_;
  assign new_n31381_ = ~new_n31327_ | ~new_n31340_ | ~new_n31342_;
  assign new_n31382_ = ~new_n31381_ | ~new_n31341_;
  assign new_n31383_ = ~new_n31331_ | ~new_n31330_;
  assign new_n31384_ = ~new_n15931_ | ~new_n31411_;
  assign new_n31385_ = ~new_n31282_ | ~new_n31344_ | ~new_n31337_;
  assign new_n31386_ = ~new_n31426_ | ~new_n15930_ | ~new_n31333_;
  assign new_n31387_ = ~new_n31285_ | ~new_n31385_;
  assign new_n31388_ = ~new_n15930_ | ~new_n31426_;
  assign new_n31389_ = ~new_n15931_ | ~new_n31411_;
  assign new_n31390_ = ~new_n31343_ | ~new_n31336_;
  assign new_n31391_ = ~new_n15536_ | ~new_n31295_;
  assign new_n31392_ = ~new_n15943_ | ~new_n31239_;
  assign new_n31393_ = ~new_n15536_ | ~new_n31296_;
  assign new_n31394_ = ~new_n15942_ | ~new_n31239_;
  assign new_n31395_ = ~new_n15536_ | ~new_n31297_;
  assign new_n31396_ = ~new_n15944_ | ~new_n31239_;
  assign new_n31397_ = ~new_n31396_ | ~new_n31395_;
  assign new_n31398_ = ~new_n15536_ | ~new_n31295_;
  assign new_n31399_ = ~new_n15943_ | ~new_n31239_;
  assign new_n31400_ = ~new_n31399_ | ~new_n31398_;
  assign new_n31401_ = ~new_n15536_ | ~new_n31297_;
  assign new_n31402_ = ~new_n15944_ | ~new_n31239_;
  assign new_n31403_ = ~new_n15536_ | ~new_n31298_;
  assign new_n31404_ = ~new_n15945_ | ~new_n31239_;
  assign new_n31405_ = ~new_n31404_ | ~new_n31403_;
  assign new_n31406_ = ~new_n15536_ | ~new_n31296_;
  assign new_n31407_ = ~new_n15942_ | ~new_n31239_;
  assign new_n31408_ = ~new_n31407_ | ~new_n31406_;
  assign new_n31409_ = ~new_n15536_ | ~new_n31299_;
  assign new_n31410_ = ~new_n15947_ | ~new_n31239_;
  assign new_n31411_ = ~new_n31410_ | ~new_n31409_;
  assign new_n31412_ = ~new_n15536_ | ~new_n31300_;
  assign new_n31413_ = ~new_n15948_ | ~new_n31239_;
  assign new_n31414_ = ~new_n31255_;
  assign new_n31415_ = ~new_n15536_ | ~new_n31301_;
  assign new_n31416_ = ~new_n15949_ | ~new_n31239_;
  assign new_n31417_ = ~new_n15536_ | ~new_n31301_;
  assign new_n31418_ = ~new_n15949_ | ~new_n31239_;
  assign new_n31419_ = ~new_n31418_ | ~new_n31417_;
  assign new_n31420_ = ~new_n15536_ | ~new_n31299_;
  assign new_n31421_ = ~new_n15947_ | ~new_n31239_;
  assign new_n31422_ = ~new_n15536_ | ~new_n31302_;
  assign new_n31423_ = ~new_n15946_ | ~new_n31239_;
  assign new_n31424_ = ~new_n15536_ | ~new_n31302_;
  assign new_n31425_ = ~new_n15946_ | ~new_n31239_;
  assign new_n31426_ = ~new_n31425_ | ~new_n31424_;
  assign new_n31427_ = ~new_n15536_ | ~new_n31298_;
  assign new_n31428_ = ~new_n15945_ | ~new_n31239_;
  assign new_n31429_ = ~new_n15536_ | ~new_n31303_;
  assign new_n31430_ = ~new_n15941_ | ~new_n31239_;
  assign new_n31431_ = ~new_n31256_;
  assign new_n31432_ = ~new_n15536_ | ~new_n31304_;
  assign new_n31433_ = ~new_n15940_ | ~new_n31239_;
  assign new_n31434_ = ~new_n31254_;
  assign new_n31435_ = ~new_n31349_ | ~new_n31434_;
  assign new_n31436_ = ~new_n31254_ | ~new_n31305_;
  assign new_n31437_ = ~new_n31348_ | ~new_n31431_;
  assign new_n31438_ = ~new_n31256_ | ~new_n31306_;
  assign new_n31439_ = ~new_n31250_ | ~new_n31284_ | ~new_n31351_;
  assign new_n31440_ = ~new_n31232_ | ~new_n31335_;
  assign new_n31441_ = ~new_n31329_ | ~new_n31383_;
  assign new_n31442_ = ~new_n31308_ | ~new_n31286_ | ~new_n31387_;
  assign new_n31443_ = ~new_n31376_ | ~new_n31310_;
  assign new_n31444_ = ~new_n31271_ | ~new_n31350_;
  assign new_n31445_ = ~new_n31377_ | ~new_n31311_;
  assign new_n31446_ = ~new_n31273_ | ~new_n31346_;
  assign new_n31447_ = ~new_n15536_ | ~new_n31312_;
  assign new_n31448_ = ~new_n15935_ | ~new_n31239_;
  assign new_n31449_ = ~new_n31259_;
  assign new_n31450_ = ~new_n15536_ | ~new_n31313_;
  assign new_n31451_ = ~new_n15934_ | ~new_n31239_;
  assign new_n31452_ = ~new_n31258_;
  assign new_n31453_ = ~new_n15536_ | ~new_n31314_;
  assign new_n31454_ = ~new_n15936_ | ~new_n31239_;
  assign new_n31455_ = ~new_n31260_;
  assign new_n31456_ = ~new_n15536_ | ~new_n31315_;
  assign new_n31457_ = ~new_n15937_ | ~new_n31239_;
  assign new_n31458_ = ~new_n31261_;
  assign new_n31459_ = ~new_n15536_ | ~new_n31316_;
  assign new_n31460_ = ~new_n15938_ | ~new_n31239_;
  assign new_n31461_ = ~new_n31262_;
  assign new_n31462_ = ~new_n15536_ | ~new_n31317_;
  assign new_n31463_ = ~new_n15939_ | ~new_n31239_;
  assign new_n31464_ = ~new_n31263_;
  assign new_n31465_ = ~new_n31390_ | ~new_n31318_;
  assign new_n31466_ = ~new_n31275_ | ~new_n31360_;
  assign new_n31467_ = ~new_n31414_ | ~new_n15932_;
  assign new_n31468_ = ~new_n31255_ | ~new_n31241_;
  assign new_n31469_ = ~new_n31414_ | ~new_n15932_;
  assign new_n31470_ = ~new_n31255_ | ~new_n31241_;
  assign new_n31471_ = ~new_n31470_ | ~new_n31469_;
  assign new_n31472_ = ~new_n31319_ | ~new_n31320_;
  assign new_n31473_ = ~new_n31357_ | ~new_n31471_;
  assign new_n31474_ = ~new_n31374_ | ~new_n31452_;
  assign new_n31475_ = ~new_n31258_ | ~new_n31321_;
  assign new_n31476_ = ~new_n31449_ | ~new_n31370_;
  assign new_n31477_ = ~new_n31259_ | ~new_n31253_;
  assign new_n31478_ = ~new_n31369_ | ~new_n31455_;
  assign new_n31479_ = ~new_n31260_ | ~new_n31322_;
  assign new_n31480_ = ~new_n31458_ | ~new_n31368_;
  assign new_n31481_ = ~new_n31261_ | ~new_n31252_;
  assign new_n31482_ = ~new_n31367_ | ~new_n31461_;
  assign new_n31483_ = ~new_n31262_ | ~new_n31323_;
  assign new_n31484_ = ~new_n31366_ | ~new_n31464_;
  assign new_n31485_ = ~new_n31263_ | ~new_n31324_;
  assign new_n31486_ = ~new_n15536_ | ~new_n31325_;
  assign new_n31487_ = ~new_n31375_ | ~new_n31239_;
  assign new_n31488_ = new_n31949_ & new_n31810_;
  assign new_n31489_ = new_n31775_ & new_n31771_;
  assign new_n31490_ = new_n31489_ & new_n31778_;
  assign new_n31491_ = new_n31788_ & new_n31785_ & new_n31781_;
  assign new_n31492_ = new_n31491_ & new_n31791_;
  assign new_n31493_ = new_n31798_ & new_n31796_ & new_n31794_;
  assign new_n31494_ = new_n31617_ & new_n31493_;
  assign new_n31495_ = new_n31778_ & new_n31775_;
  assign new_n31496_ = new_n31492_ & new_n31804_;
  assign new_n31497_ = new_n31946_ & new_n31945_;
  assign new_n31498_ = new_n31827_ & new_n31825_;
  assign new_n31499_ = new_n31858_ & new_n31950_ & new_n31951_ & new_n31671_;
  assign new_n31500_ = new_n31755_ & new_n31753_;
  assign new_n31501_ = new_n31751_ & new_n31749_;
  assign new_n31502_ = ~new_n31697_ | ~new_n31912_;
  assign new_n31503_ = new_n31897_ & new_n31818_;
  assign new_n31504_ = ~pi1223;
  assign new_n31505_ = ~new_n15973_;
  assign new_n31506_ = ~pi1222;
  assign new_n31507_ = ~new_n15974_;
  assign new_n31508_ = ~pi1221;
  assign new_n31509_ = ~new_n15975_;
  assign new_n31510_ = ~pi1220;
  assign new_n31511_ = ~new_n15976_;
  assign new_n31512_ = ~new_n15981_;
  assign new_n31513_ = ~pi1215;
  assign new_n31514_ = ~pi1216;
  assign new_n31515_ = ~pi1215 | ~new_n15981_;
  assign new_n31516_ = ~new_n15980_;
  assign new_n31517_ = ~pi1217;
  assign new_n31518_ = ~new_n15979_;
  assign new_n31519_ = ~pi1218;
  assign new_n31520_ = ~new_n15978_;
  assign new_n31521_ = ~pi1219;
  assign new_n31522_ = ~new_n15977_;
  assign new_n31523_ = ~new_n31526_ | ~new_n31733_;
  assign new_n31524_ = ~new_n31736_ | ~new_n31737_ | ~new_n31735_;
  assign new_n31525_ = ~new_n31729_ | ~new_n31728_;
  assign new_n31526_ = ~new_n31525_ | ~new_n31731_;
  assign new_n31527_ = ~pi1240;
  assign new_n31528_ = ~new_n15956_;
  assign new_n31529_ = ~pi1241;
  assign new_n31530_ = ~new_n15955_;
  assign new_n31531_ = ~pi1239;
  assign new_n31532_ = ~new_n15957_;
  assign new_n31533_ = ~pi1238;
  assign new_n31534_ = ~new_n15958_;
  assign new_n31535_ = ~pi1236;
  assign new_n31536_ = ~new_n15960_;
  assign new_n31537_ = ~pi1235;
  assign new_n31538_ = ~new_n15961_;
  assign new_n31539_ = ~pi1234;
  assign new_n31540_ = ~new_n15962_;
  assign new_n31541_ = ~pi1226;
  assign new_n31542_ = ~new_n15970_;
  assign new_n31543_ = ~pi1225;
  assign new_n31544_ = ~new_n15971_;
  assign new_n31545_ = ~pi1230;
  assign new_n31546_ = ~new_n15966_;
  assign new_n31547_ = ~pi1228;
  assign new_n31548_ = ~new_n15968_;
  assign new_n31549_ = ~pi1229;
  assign new_n31550_ = ~new_n15967_;
  assign new_n31551_ = ~new_n15969_ | ~pi1227;
  assign new_n31552_ = ~pi1231;
  assign new_n31553_ = ~new_n15965_;
  assign new_n31554_ = ~pi1232;
  assign new_n31555_ = ~new_n15964_;
  assign new_n31556_ = ~new_n31491_ | ~new_n31791_ | ~new_n31842_ | ~new_n31495_;
  assign new_n31557_ = ~pi1237;
  assign new_n31558_ = ~new_n15959_;
  assign new_n31559_ = ~new_n15959_ | ~pi1237;
  assign new_n31560_ = ~pi1233;
  assign new_n31561_ = ~new_n15963_;
  assign new_n31562_ = ~new_n15963_ | ~pi1233;
  assign new_n31563_ = ~new_n31627_ | ~new_n31491_;
  assign new_n31564_ = ~new_n15953_;
  assign new_n31565_ = ~pi1243;
  assign new_n31566_ = ~pi1242;
  assign new_n31567_ = ~new_n15954_;
  assign new_n31568_ = ~new_n15954_ | ~pi1242;
  assign new_n31569_ = ~new_n31862_ | ~new_n31805_;
  assign new_n31570_ = ~new_n31576_ | ~new_n31875_ | ~new_n31575_;
  assign new_n31571_ = ~new_n15951_;
  assign new_n31572_ = ~pi1245;
  assign new_n31573_ = ~new_n15952_;
  assign new_n31574_ = ~pi1244;
  assign new_n31575_ = ~new_n31626_ | ~new_n31494_;
  assign new_n31576_ = ~new_n31860_ | ~new_n31494_ | ~new_n31804_;
  assign new_n31577_ = ~new_n31615_ | ~new_n31855_;
  assign new_n31578_ = ~new_n31619_ | ~new_n31851_;
  assign new_n31579_ = ~new_n31861_ | ~new_n31494_ | ~new_n31804_;
  assign new_n31580_ = ~new_n31712_ | ~new_n31814_;
  assign new_n31581_ = ~new_n31621_ | ~new_n31837_;
  assign new_n31582_ = ~new_n32093_ | ~new_n32092_;
  assign new_n31583_ = new_n31745_ & new_n31744_;
  assign new_n31584_ = ~new_n31914_ | ~new_n31913_;
  assign new_n31585_ = ~new_n31921_ | ~new_n31920_;
  assign new_n31586_ = ~new_n31928_ | ~new_n31927_;
  assign new_n31587_ = ~new_n31937_ | ~new_n31936_;
  assign new_n31588_ = ~new_n31944_ | ~new_n31943_;
  assign new_n31589_ = ~new_n31960_ | ~new_n31959_;
  assign new_n31590_ = ~new_n31967_ | ~new_n31966_;
  assign new_n31591_ = ~new_n31974_ | ~new_n31973_;
  assign new_n31592_ = ~new_n31981_ | ~new_n31980_;
  assign new_n31593_ = ~new_n31988_ | ~new_n31987_;
  assign new_n31594_ = ~new_n31995_ | ~new_n31994_;
  assign new_n31595_ = ~new_n32002_ | ~new_n32001_;
  assign new_n31596_ = ~new_n32009_ | ~new_n32008_;
  assign new_n31597_ = ~new_n32016_ | ~new_n32015_;
  assign new_n31598_ = ~new_n32023_ | ~new_n32022_;
  assign new_n31599_ = ~new_n32030_ | ~new_n32029_;
  assign new_n31600_ = ~new_n32037_ | ~new_n32036_;
  assign new_n31601_ = ~new_n32049_ | ~new_n32048_;
  assign new_n31602_ = ~new_n32056_ | ~new_n32055_;
  assign new_n31603_ = ~new_n32063_ | ~new_n32062_;
  assign new_n31604_ = ~new_n32070_ | ~new_n32069_;
  assign new_n31605_ = ~new_n32077_ | ~new_n32076_;
  assign new_n31606_ = ~new_n32082_ | ~new_n32081_;
  assign new_n31607_ = new_n31551_ & new_n31764_;
  assign new_n31608_ = ~new_n32084_ | ~new_n32083_;
  assign new_n31609_ = ~new_n32091_ | ~new_n32090_;
  assign new_n31610_ = pi1222 & new_n15974_;
  assign new_n31611_ = new_n31741_ & new_n31737_;
  assign new_n31612_ = new_n31835_ & new_n31742_;
  assign new_n31613_ = pi1238 & new_n15958_;
  assign new_n31614_ = new_n31801_ & new_n31799_;
  assign new_n31615_ = new_n31804_ & new_n31802_ & new_n31800_;
  assign new_n31616_ = pi1234 & new_n15962_;
  assign new_n31617_ = new_n31802_ & new_n31800_;
  assign new_n31618_ = new_n31804_ & new_n31791_;
  assign new_n31619_ = new_n31494_ & new_n31618_;
  assign new_n31620_ = new_n31756_ & new_n31742_ & new_n31711_;
  assign new_n31621_ = new_n31872_ & new_n31759_;
  assign new_n31622_ = new_n31840_ & new_n31623_;
  assign new_n31623_ = new_n31767_ & new_n31764_ & new_n31766_;
  assign new_n31624_ = new_n31769_ & new_n31893_;
  assign new_n31625_ = new_n31490_ & new_n31496_;
  assign new_n31626_ = new_n31792_ & new_n31804_;
  assign new_n31627_ = new_n31779_ & new_n31791_;
  assign new_n31628_ = new_n31578_ & new_n31577_;
  assign new_n31629_ = new_n31884_ & new_n31579_;
  assign new_n31630_ = new_n31807_ & new_n31488_;
  assign new_n31631_ = new_n31804_ & new_n31800_ & new_n31802_ & new_n31807_;
  assign new_n31632_ = new_n31807_ & new_n31804_ & new_n31791_;
  assign new_n31633_ = new_n31494_ & new_n31632_;
  assign new_n31634_ = new_n31769_ & new_n31895_;
  assign new_n31635_ = new_n31494_ & new_n31807_;
  assign new_n31636_ = new_n31490_ & new_n31496_;
  assign new_n31637_ = new_n31807_ & new_n31804_;
  assign new_n31638_ = new_n31877_ & new_n31639_ & new_n31881_ & new_n31878_ & new_n31876_;
  assign new_n31639_ = new_n31882_ & new_n31497_ & new_n31883_;
  assign new_n31640_ = new_n31494_ & new_n31807_;
  assign new_n31641_ = new_n31490_ & new_n31496_;
  assign new_n31642_ = new_n31887_ & new_n31886_ & new_n31670_;
  assign new_n31643_ = new_n31769_ & new_n31900_;
  assign new_n31644_ = new_n31492_ & new_n31490_;
  assign new_n31645_ = new_n31852_ & new_n31559_;
  assign new_n31646_ = new_n31556_ & new_n31563_;
  assign new_n31647_ = new_n31800_ & new_n31493_;
  assign new_n31648_ = new_n31854_ & new_n31799_;
  assign new_n31649_ = new_n31794_ & new_n31796_;
  assign new_n31650_ = new_n31853_ & new_n31797_;
  assign new_n31651_ = new_n31769_ & new_n31898_;
  assign new_n31652_ = new_n31845_ & new_n31562_;
  assign new_n31653_ = new_n31850_ & new_n31789_;
  assign new_n31654_ = new_n31781_ & new_n31785_;
  assign new_n31655_ = new_n31847_ & new_n31786_;
  assign new_n31656_ = new_n31768_ & new_n32072_ & new_n32071_;
  assign new_n31657_ = new_n31820_ & new_n31710_;
  assign new_n31658_ = new_n31711_ & new_n32086_ & new_n32085_;
  assign new_n31659_ = ~new_n31612_ | ~new_n31836_;
  assign new_n31660_ = new_n31916_ & new_n31915_;
  assign new_n31661_ = ~new_n31524_ | ~new_n31739_;
  assign new_n31662_ = new_n31923_ & new_n31922_;
  assign new_n31663_ = new_n31930_ & new_n31929_;
  assign new_n31664_ = new_n31932_ & new_n31931_;
  assign new_n31665_ = ~new_n31725_ | ~new_n31724_;
  assign new_n31666_ = new_n31939_ & new_n31938_;
  assign new_n31667_ = ~new_n31721_ | ~new_n31720_;
  assign new_n31668_ = ~pi1246;
  assign new_n31669_ = ~new_n15950_;
  assign new_n31670_ = ~pi1244 | ~new_n15952_;
  assign new_n31671_ = new_n31953_ & new_n31952_;
  assign new_n31672_ = new_n31955_ & new_n31954_;
  assign new_n31673_ = ~new_n31888_ | ~new_n31642_ | ~new_n31890_ | ~new_n31889_;
  assign new_n31674_ = new_n31962_ & new_n31961_;
  assign new_n31675_ = ~new_n31696_ | ~new_n31717_;
  assign new_n31676_ = new_n31969_ & new_n31968_;
  assign new_n31677_ = ~new_n31629_ | ~new_n31628_ | ~new_n31868_;
  assign new_n31678_ = new_n31976_ & new_n31975_;
  assign new_n31679_ = ~new_n31902_ | ~new_n31892_;
  assign new_n31680_ = new_n31983_ & new_n31982_;
  assign new_n31681_ = ~new_n31908_ | ~new_n31856_;
  assign new_n31682_ = new_n31990_ & new_n31989_;
  assign new_n31683_ = ~new_n31648_ | ~new_n31906_;
  assign new_n31684_ = new_n31997_ & new_n31996_;
  assign new_n31685_ = ~new_n31650_ | ~new_n31910_;
  assign new_n31686_ = new_n32004_ & new_n32003_;
  assign new_n31687_ = ~new_n31904_ | ~new_n31795_;
  assign new_n31688_ = new_n32011_ & new_n32010_;
  assign new_n31689_ = ~new_n31645_ | ~new_n31646_ | ~new_n31859_;
  assign new_n31690_ = new_n32018_ & new_n32017_;
  assign new_n31691_ = ~new_n31653_ | ~new_n31848_;
  assign new_n31692_ = new_n32025_ & new_n32024_;
  assign new_n31693_ = ~new_n31655_ | ~new_n31846_;
  assign new_n31694_ = new_n32032_ & new_n32031_;
  assign new_n31695_ = ~new_n31783_ | ~new_n31782_;
  assign new_n31696_ = ~new_n15980_ | ~new_n31715_;
  assign new_n31697_ = new_n32042_ & new_n32041_;
  assign new_n31698_ = new_n32044_ & new_n32043_;
  assign new_n31699_ = ~new_n31652_ | ~new_n31844_;
  assign new_n31700_ = new_n32051_ & new_n32050_;
  assign new_n31701_ = ~new_n31843_ | ~new_n31841_;
  assign new_n31702_ = new_n32058_ & new_n32057_;
  assign new_n31703_ = ~new_n31773_ | ~new_n31772_;
  assign new_n31704_ = new_n32065_ & new_n32064_;
  assign new_n31705_ = ~new_n31651_ | ~new_n31709_;
  assign new_n31706_ = ~new_n31551_ | ~new_n31811_;
  assign new_n31707_ = ~new_n31581_ | ~new_n31762_;
  assign new_n31708_ = ~new_n31757_ | ~new_n31756_;
  assign new_n31709_ = ~new_n31707_ | ~new_n31622_;
  assign new_n31710_ = ~new_n31839_ | ~new_n31838_;
  assign new_n31711_ = ~new_n15971_ | ~pi1225;
  assign new_n31712_ = ~new_n15968_ | ~pi1228;
  assign new_n31713_ = ~new_n31696_;
  assign new_n31714_ = ~new_n15975_ | ~pi1221;
  assign new_n31715_ = ~new_n31515_;
  assign new_n31716_ = ~new_n31516_ | ~new_n31515_;
  assign new_n31717_ = ~pi1216 | ~new_n31716_;
  assign new_n31718_ = ~new_n31675_;
  assign new_n31719_ = pi1217 | new_n15979_;
  assign new_n31720_ = ~new_n31719_ | ~new_n31675_;
  assign new_n31721_ = ~new_n15979_ | ~pi1217;
  assign new_n31722_ = ~new_n31667_;
  assign new_n31723_ = pi1218 | new_n15978_;
  assign new_n31724_ = ~new_n31723_ | ~new_n31667_;
  assign new_n31725_ = ~new_n15978_ | ~pi1218;
  assign new_n31726_ = ~new_n31665_;
  assign new_n31727_ = pi1219 | new_n15977_;
  assign new_n31728_ = ~new_n31727_ | ~new_n31665_;
  assign new_n31729_ = ~new_n15977_ | ~pi1219;
  assign new_n31730_ = ~new_n31525_;
  assign new_n31731_ = new_n15976_ | pi1220;
  assign new_n31732_ = ~new_n31526_;
  assign new_n31733_ = ~new_n15976_ | ~pi1220;
  assign new_n31734_ = ~new_n31523_;
  assign new_n31735_ = ~new_n31734_ | ~new_n31714_;
  assign new_n31736_ = new_n15974_ | pi1222;
  assign new_n31737_ = new_n15975_ | pi1221;
  assign new_n31738_ = ~new_n31524_;
  assign new_n31739_ = ~new_n15974_ | ~pi1222;
  assign new_n31740_ = ~new_n31661_;
  assign new_n31741_ = pi1223 | new_n15973_;
  assign new_n31742_ = ~new_n15973_ | ~pi1223;
  assign new_n31743_ = ~new_n31659_;
  assign new_n31744_ = pi1224 | new_n15972_;
  assign new_n31745_ = ~new_n15972_ | ~pi1224;
  assign new_n31746_ = ~new_n15972_ | ~pi1224;
  assign new_n31747_ = pi1221 | new_n15975_;
  assign new_n31748_ = ~new_n31747_ | ~new_n31523_;
  assign new_n31749_ = ~new_n31662_ | ~new_n31748_ | ~new_n31714_;
  assign new_n31750_ = ~new_n15974_ | ~pi1222;
  assign new_n31751_ = ~new_n31738_ | ~new_n31750_;
  assign new_n31752_ = new_n15975_ | pi1221;
  assign new_n31753_ = ~new_n31663_ | ~new_n31730_;
  assign new_n31754_ = ~new_n15976_ | ~pi1220;
  assign new_n31755_ = ~new_n31732_ | ~new_n31754_;
  assign new_n31756_ = ~new_n15972_ | ~pi1224;
  assign new_n31757_ = ~new_n31744_ | ~new_n31659_;
  assign new_n31758_ = ~new_n31708_;
  assign new_n31759_ = new_n15970_ | pi1226;
  assign new_n31760_ = new_n15971_ | pi1225;
  assign new_n31761_ = ~new_n31581_;
  assign new_n31762_ = ~new_n15970_ | ~pi1226;
  assign new_n31763_ = ~new_n31707_;
  assign new_n31764_ = pi1227 | new_n15969_;
  assign new_n31765_ = ~new_n31551_;
  assign new_n31766_ = new_n15968_ | pi1228;
  assign new_n31767_ = new_n15967_ | pi1229;
  assign new_n31768_ = ~new_n15967_ | ~pi1229;
  assign new_n31769_ = ~new_n15966_ | ~pi1230;
  assign new_n31770_ = ~new_n31768_ | ~new_n31874_ | ~new_n31712_;
  assign new_n31771_ = pi1231 | new_n15965_;
  assign new_n31772_ = ~new_n31771_ | ~new_n31705_;
  assign new_n31773_ = ~new_n15965_ | ~pi1231;
  assign new_n31774_ = ~new_n31703_;
  assign new_n31775_ = pi1232 | new_n15964_;
  assign new_n31776_ = ~new_n15964_ | ~pi1232;
  assign new_n31777_ = ~new_n31701_;
  assign new_n31778_ = pi1233 | new_n15963_;
  assign new_n31779_ = ~new_n31562_;
  assign new_n31780_ = ~new_n31699_;
  assign new_n31781_ = pi1234 | new_n15962_;
  assign new_n31782_ = ~new_n31781_ | ~new_n31699_;
  assign new_n31783_ = ~new_n15962_ | ~pi1234;
  assign new_n31784_ = ~new_n31695_;
  assign new_n31785_ = pi1235 | new_n15961_;
  assign new_n31786_ = ~new_n15961_ | ~pi1235;
  assign new_n31787_ = ~new_n31693_;
  assign new_n31788_ = pi1236 | new_n15960_;
  assign new_n31789_ = ~new_n15960_ | ~pi1236;
  assign new_n31790_ = ~new_n31691_;
  assign new_n31791_ = pi1237 | new_n15959_;
  assign new_n31792_ = ~new_n31559_;
  assign new_n31793_ = ~new_n31689_;
  assign new_n31794_ = pi1238 | new_n15958_;
  assign new_n31795_ = ~new_n15958_ | ~pi1238;
  assign new_n31796_ = pi1239 | new_n15957_;
  assign new_n31797_ = ~new_n15957_ | ~pi1239;
  assign new_n31798_ = pi1240 | new_n15956_;
  assign new_n31799_ = ~new_n15956_ | ~pi1240;
  assign new_n31800_ = pi1241 | new_n15955_;
  assign new_n31801_ = ~new_n15955_ | ~pi1241;
  assign new_n31802_ = pi1242 | new_n15954_;
  assign new_n31803_ = ~new_n31568_;
  assign new_n31804_ = new_n15953_ | pi1243;
  assign new_n31805_ = ~pi1243 | ~new_n15953_;
  assign new_n31806_ = ~new_n31677_;
  assign new_n31807_ = new_n15952_ | pi1244;
  assign new_n31808_ = ~new_n31670_;
  assign new_n31809_ = ~new_n31673_;
  assign new_n31810_ = pi1245 | new_n15951_;
  assign new_n31811_ = ~new_n31764_ | ~new_n31707_;
  assign new_n31812_ = ~new_n31706_;
  assign new_n31813_ = pi1228 | new_n15968_;
  assign new_n31814_ = ~new_n31813_ | ~new_n31706_;
  assign new_n31815_ = ~new_n31580_;
  assign new_n31816_ = pi1229 | new_n15967_;
  assign new_n31817_ = ~new_n31816_ | ~new_n31580_;
  assign new_n31818_ = ~new_n31656_ | ~new_n31817_;
  assign new_n31819_ = ~new_n31815_ | ~new_n31768_;
  assign new_n31820_ = ~new_n15966_ | ~pi1230;
  assign new_n31821_ = new_n15967_ | pi1229;
  assign new_n31822_ = new_n15968_ | pi1228;
  assign new_n31823_ = pi1225 | new_n15971_;
  assign new_n31824_ = ~new_n31823_ | ~new_n31708_;
  assign new_n31825_ = ~new_n31658_ | ~new_n31824_;
  assign new_n31826_ = ~new_n15970_ | ~pi1226;
  assign new_n31827_ = ~new_n31761_ | ~new_n31826_;
  assign new_n31828_ = new_n15971_ | pi1225;
  assign new_n31829_ = ~new_n31746_ | ~new_n31744_;
  assign new_n31830_ = ~new_n31752_ | ~new_n31714_;
  assign new_n31831_ = ~new_n31821_ | ~new_n31768_;
  assign new_n31832_ = ~new_n31822_ | ~new_n31712_;
  assign new_n31833_ = ~new_n31551_ | ~new_n31764_;
  assign new_n31834_ = ~new_n31828_ | ~new_n31711_;
  assign new_n31835_ = ~new_n31610_ | ~new_n31741_;
  assign new_n31836_ = ~new_n31611_ | ~new_n31736_ | ~new_n31735_;
  assign new_n31837_ = ~new_n31620_ | ~new_n31836_ | ~new_n31835_;
  assign new_n31838_ = ~new_n15966_ | ~new_n31767_;
  assign new_n31839_ = ~pi1230 | ~new_n31767_;
  assign new_n31840_ = ~new_n31839_ | ~new_n31546_;
  assign new_n31841_ = ~new_n31489_ | ~new_n31705_;
  assign new_n31842_ = ~new_n31776_ | ~new_n31773_;
  assign new_n31843_ = ~new_n31842_ | ~new_n31775_;
  assign new_n31844_ = ~new_n31490_ | ~new_n31705_;
  assign new_n31845_ = ~new_n31495_ | ~new_n31842_;
  assign new_n31846_ = ~new_n31654_ | ~new_n31699_;
  assign new_n31847_ = ~new_n31616_ | ~new_n31785_;
  assign new_n31848_ = ~new_n31491_ | ~new_n31699_;
  assign new_n31849_ = ~new_n31847_ | ~new_n31786_;
  assign new_n31850_ = ~new_n31849_ | ~new_n31788_;
  assign new_n31851_ = ~new_n31850_ | ~new_n31789_;
  assign new_n31852_ = ~new_n31851_ | ~new_n31791_;
  assign new_n31853_ = ~new_n31613_ | ~new_n31796_;
  assign new_n31854_ = ~new_n31864_ | ~new_n31798_;
  assign new_n31855_ = ~new_n31614_ | ~new_n31854_;
  assign new_n31856_ = ~new_n31855_ | ~new_n31800_;
  assign new_n31857_ = ~new_n31855_ | ~new_n31800_;
  assign new_n31858_ = ~new_n31630_ | ~new_n31677_;
  assign new_n31859_ = ~new_n31644_ | ~new_n31901_;
  assign new_n31860_ = ~new_n31563_;
  assign new_n31861_ = ~new_n31556_;
  assign new_n31862_ = ~new_n31803_ | ~new_n31804_;
  assign new_n31863_ = ~new_n31577_;
  assign new_n31864_ = ~new_n31853_ | ~new_n31797_;
  assign new_n31865_ = ~new_n31768_ | ~new_n31874_ | ~new_n31712_;
  assign new_n31866_ = ~new_n31575_;
  assign new_n31867_ = ~new_n31578_;
  assign new_n31868_ = ~new_n31625_ | ~new_n31494_ | ~new_n31894_;
  assign new_n31869_ = ~new_n31576_;
  assign new_n31870_ = ~new_n31579_;
  assign new_n31871_ = ~new_n31760_ | ~new_n31744_;
  assign new_n31872_ = ~new_n31871_ | ~new_n31711_;
  assign new_n31873_ = ~new_n31768_ | ~new_n31874_ | ~new_n31712_;
  assign new_n31874_ = ~new_n31765_ | ~new_n31766_;
  assign new_n31875_ = ~new_n31569_;
  assign new_n31876_ = ~pi1245 | ~new_n15951_;
  assign new_n31877_ = ~new_n31631_ | ~new_n31855_;
  assign new_n31878_ = ~new_n31866_ | ~new_n31807_;
  assign new_n31879_ = ~new_n31633_ | ~new_n31851_;
  assign new_n31880_ = ~new_n31636_ | ~new_n31635_ | ~new_n31896_;
  assign new_n31881_ = ~new_n31869_ | ~new_n31807_;
  assign new_n31882_ = ~new_n31861_ | ~new_n31637_ | ~new_n31494_;
  assign new_n31883_ = ~new_n31569_ | ~new_n31807_;
  assign new_n31884_ = ~new_n31570_;
  assign new_n31885_ = ~new_n31768_ | ~new_n31874_ | ~new_n31712_;
  assign new_n31886_ = ~new_n31863_ | ~new_n31807_;
  assign new_n31887_ = ~new_n31867_ | ~new_n31807_;
  assign new_n31888_ = ~new_n31641_ | ~new_n31640_ | ~new_n31894_;
  assign new_n31889_ = ~new_n31870_ | ~new_n31807_;
  assign new_n31890_ = ~new_n31570_ | ~new_n31807_;
  assign new_n31891_ = ~new_n31857_ | ~new_n31568_;
  assign new_n31892_ = ~new_n31891_ | ~new_n31802_;
  assign new_n31893_ = ~new_n31885_ | ~new_n31710_;
  assign new_n31894_ = ~new_n31624_ | ~new_n31709_;
  assign new_n31895_ = ~new_n31873_ | ~new_n31710_;
  assign new_n31896_ = ~new_n31634_ | ~new_n31709_;
  assign new_n31897_ = ~new_n31657_ | ~new_n31819_;
  assign new_n31898_ = ~new_n31770_ | ~new_n31710_;
  assign new_n31899_ = ~new_n31705_;
  assign new_n31900_ = ~new_n31865_ | ~new_n31710_;
  assign new_n31901_ = ~new_n31643_ | ~new_n31709_;
  assign new_n31902_ = ~new_n31494_ | ~new_n31689_;
  assign new_n31903_ = ~new_n31679_;
  assign new_n31904_ = ~new_n31794_ | ~new_n31689_;
  assign new_n31905_ = ~new_n31687_;
  assign new_n31906_ = ~new_n31493_ | ~new_n31689_;
  assign new_n31907_ = ~new_n31683_;
  assign new_n31908_ = ~new_n31647_ | ~new_n31689_;
  assign new_n31909_ = ~new_n31681_;
  assign new_n31910_ = ~new_n31649_ | ~new_n31689_;
  assign new_n31911_ = ~new_n31685_;
  assign new_n31912_ = ~new_n32040_ | ~new_n31516_;
  assign new_n31913_ = ~new_n31829_ | ~new_n31659_;
  assign new_n31914_ = ~new_n31583_ | ~new_n31743_;
  assign new_n31915_ = ~new_n15973_ | ~new_n31504_;
  assign new_n31916_ = ~pi1223 | ~new_n31505_;
  assign new_n31917_ = ~new_n15973_ | ~new_n31504_;
  assign new_n31918_ = ~pi1223 | ~new_n31505_;
  assign new_n31919_ = ~new_n31918_ | ~new_n31917_;
  assign new_n31920_ = ~new_n31660_ | ~new_n31661_;
  assign new_n31921_ = ~new_n31740_ | ~new_n31919_;
  assign new_n31922_ = ~new_n15974_ | ~new_n31506_;
  assign new_n31923_ = ~pi1222 | ~new_n31507_;
  assign new_n31924_ = ~new_n15975_ | ~new_n31508_;
  assign new_n31925_ = ~pi1221 | ~new_n31509_;
  assign new_n31926_ = ~new_n31925_ | ~new_n31924_;
  assign new_n31927_ = ~new_n31830_ | ~new_n31523_;
  assign new_n31928_ = ~new_n31926_ | ~new_n31734_;
  assign new_n31929_ = ~new_n15976_ | ~new_n31510_;
  assign new_n31930_ = ~pi1220 | ~new_n31511_;
  assign new_n31931_ = ~new_n15977_ | ~new_n31521_;
  assign new_n31932_ = ~pi1219 | ~new_n31522_;
  assign new_n31933_ = ~new_n15977_ | ~new_n31521_;
  assign new_n31934_ = ~pi1219 | ~new_n31522_;
  assign new_n31935_ = ~new_n31934_ | ~new_n31933_;
  assign new_n31936_ = ~new_n31664_ | ~new_n31665_;
  assign new_n31937_ = ~new_n31726_ | ~new_n31935_;
  assign new_n31938_ = ~new_n15978_ | ~new_n31519_;
  assign new_n31939_ = ~pi1218 | ~new_n31520_;
  assign new_n31940_ = ~new_n15978_ | ~new_n31519_;
  assign new_n31941_ = ~pi1218 | ~new_n31520_;
  assign new_n31942_ = ~new_n31941_ | ~new_n31940_;
  assign new_n31943_ = ~new_n31666_ | ~new_n31667_;
  assign new_n31944_ = ~new_n31722_ | ~new_n31942_;
  assign new_n31945_ = ~pi1246 | ~new_n31669_;
  assign new_n31946_ = ~new_n15950_ | ~new_n31668_;
  assign new_n31947_ = ~pi1246 | ~new_n31669_;
  assign new_n31948_ = ~new_n15950_ | ~new_n31668_;
  assign new_n31949_ = ~new_n31948_ | ~new_n31947_;
  assign new_n31950_ = ~new_n31879_ | ~new_n31670_ | ~new_n31638_ | ~new_n31880_;
  assign new_n31951_ = ~new_n31808_ | ~new_n31488_;
  assign new_n31952_ = ~new_n31572_ | ~new_n31497_ | ~new_n31571_;
  assign new_n31953_ = ~pi1245 | ~new_n15951_ | ~new_n31949_;
  assign new_n31954_ = ~pi1245 | ~new_n31571_;
  assign new_n31955_ = ~new_n15951_ | ~new_n31572_;
  assign new_n31956_ = ~pi1245 | ~new_n31571_;
  assign new_n31957_ = ~new_n15951_ | ~new_n31572_;
  assign new_n31958_ = ~new_n31957_ | ~new_n31956_;
  assign new_n31959_ = ~new_n31672_ | ~new_n31673_;
  assign new_n31960_ = ~new_n31809_ | ~new_n31958_;
  assign new_n31961_ = ~new_n15979_ | ~new_n31517_;
  assign new_n31962_ = ~pi1217 | ~new_n31518_;
  assign new_n31963_ = ~new_n15979_ | ~new_n31517_;
  assign new_n31964_ = ~pi1217 | ~new_n31518_;
  assign new_n31965_ = ~new_n31964_ | ~new_n31963_;
  assign new_n31966_ = ~new_n31674_ | ~new_n31675_;
  assign new_n31967_ = ~new_n31718_ | ~new_n31965_;
  assign new_n31968_ = ~pi1244 | ~new_n31573_;
  assign new_n31969_ = ~new_n15952_ | ~new_n31574_;
  assign new_n31970_ = ~pi1244 | ~new_n31573_;
  assign new_n31971_ = ~new_n15952_ | ~new_n31574_;
  assign new_n31972_ = ~new_n31971_ | ~new_n31970_;
  assign new_n31973_ = ~new_n31676_ | ~new_n31677_;
  assign new_n31974_ = ~new_n31806_ | ~new_n31972_;
  assign new_n31975_ = ~pi1243 | ~new_n31564_;
  assign new_n31976_ = ~new_n15953_ | ~new_n31565_;
  assign new_n31977_ = ~pi1243 | ~new_n31564_;
  assign new_n31978_ = ~new_n15953_ | ~new_n31565_;
  assign new_n31979_ = ~new_n31978_ | ~new_n31977_;
  assign new_n31980_ = ~new_n31678_ | ~new_n31679_;
  assign new_n31981_ = ~new_n31903_ | ~new_n31979_;
  assign new_n31982_ = ~new_n15954_ | ~new_n31566_;
  assign new_n31983_ = ~pi1242 | ~new_n31567_;
  assign new_n31984_ = ~new_n15954_ | ~new_n31566_;
  assign new_n31985_ = ~pi1242 | ~new_n31567_;
  assign new_n31986_ = ~new_n31985_ | ~new_n31984_;
  assign new_n31987_ = ~new_n31680_ | ~new_n31681_;
  assign new_n31988_ = ~new_n31909_ | ~new_n31986_;
  assign new_n31989_ = ~new_n15955_ | ~new_n31529_;
  assign new_n31990_ = ~pi1241 | ~new_n31530_;
  assign new_n31991_ = ~new_n15955_ | ~new_n31529_;
  assign new_n31992_ = ~pi1241 | ~new_n31530_;
  assign new_n31993_ = ~new_n31992_ | ~new_n31991_;
  assign new_n31994_ = ~new_n31682_ | ~new_n31683_;
  assign new_n31995_ = ~new_n31907_ | ~new_n31993_;
  assign new_n31996_ = ~new_n15956_ | ~new_n31527_;
  assign new_n31997_ = ~pi1240 | ~new_n31528_;
  assign new_n31998_ = ~new_n15956_ | ~new_n31527_;
  assign new_n31999_ = ~pi1240 | ~new_n31528_;
  assign new_n32000_ = ~new_n31999_ | ~new_n31998_;
  assign new_n32001_ = ~new_n31684_ | ~new_n31685_;
  assign new_n32002_ = ~new_n31911_ | ~new_n32000_;
  assign new_n32003_ = ~new_n15957_ | ~new_n31531_;
  assign new_n32004_ = ~pi1239 | ~new_n31532_;
  assign new_n32005_ = ~new_n15957_ | ~new_n31531_;
  assign new_n32006_ = ~pi1239 | ~new_n31532_;
  assign new_n32007_ = ~new_n32006_ | ~new_n32005_;
  assign new_n32008_ = ~new_n31686_ | ~new_n31687_;
  assign new_n32009_ = ~new_n31905_ | ~new_n32007_;
  assign new_n32010_ = ~new_n15958_ | ~new_n31533_;
  assign new_n32011_ = ~pi1238 | ~new_n31534_;
  assign new_n32012_ = ~new_n15958_ | ~new_n31533_;
  assign new_n32013_ = ~pi1238 | ~new_n31534_;
  assign new_n32014_ = ~new_n32013_ | ~new_n32012_;
  assign new_n32015_ = ~new_n31688_ | ~new_n31689_;
  assign new_n32016_ = ~new_n31793_ | ~new_n32014_;
  assign new_n32017_ = ~new_n15959_ | ~new_n31557_;
  assign new_n32018_ = ~pi1237 | ~new_n31558_;
  assign new_n32019_ = ~new_n15959_ | ~new_n31557_;
  assign new_n32020_ = ~pi1237 | ~new_n31558_;
  assign new_n32021_ = ~new_n32020_ | ~new_n32019_;
  assign new_n32022_ = ~new_n31690_ | ~new_n31691_;
  assign new_n32023_ = ~new_n31790_ | ~new_n32021_;
  assign new_n32024_ = ~new_n15960_ | ~new_n31535_;
  assign new_n32025_ = ~pi1236 | ~new_n31536_;
  assign new_n32026_ = ~new_n15960_ | ~new_n31535_;
  assign new_n32027_ = ~pi1236 | ~new_n31536_;
  assign new_n32028_ = ~new_n32027_ | ~new_n32026_;
  assign new_n32029_ = ~new_n31692_ | ~new_n31693_;
  assign new_n32030_ = ~new_n31787_ | ~new_n32028_;
  assign new_n32031_ = ~new_n15961_ | ~new_n31537_;
  assign new_n32032_ = ~pi1235 | ~new_n31538_;
  assign new_n32033_ = ~new_n15961_ | ~new_n31537_;
  assign new_n32034_ = ~pi1235 | ~new_n31538_;
  assign new_n32035_ = ~new_n32034_ | ~new_n32033_;
  assign new_n32036_ = ~new_n31694_ | ~new_n31695_;
  assign new_n32037_ = ~new_n31784_ | ~new_n32035_;
  assign new_n32038_ = ~pi1216 | ~new_n31515_;
  assign new_n32039_ = ~new_n31715_ | ~new_n31514_;
  assign new_n32040_ = ~new_n32039_ | ~new_n32038_;
  assign new_n32041_ = ~new_n31514_ | ~new_n15980_ | ~new_n31515_;
  assign new_n32042_ = ~new_n31713_ | ~pi1216;
  assign new_n32043_ = ~new_n15962_ | ~new_n31539_;
  assign new_n32044_ = ~pi1234 | ~new_n31540_;
  assign new_n32045_ = ~new_n15962_ | ~new_n31539_;
  assign new_n32046_ = ~pi1234 | ~new_n31540_;
  assign new_n32047_ = ~new_n32046_ | ~new_n32045_;
  assign new_n32048_ = ~new_n31698_ | ~new_n31699_;
  assign new_n32049_ = ~new_n31780_ | ~new_n32047_;
  assign new_n32050_ = ~new_n15963_ | ~new_n31560_;
  assign new_n32051_ = ~pi1233 | ~new_n31561_;
  assign new_n32052_ = ~new_n15963_ | ~new_n31560_;
  assign new_n32053_ = ~pi1233 | ~new_n31561_;
  assign new_n32054_ = ~new_n32053_ | ~new_n32052_;
  assign new_n32055_ = ~new_n31700_ | ~new_n31701_;
  assign new_n32056_ = ~new_n31777_ | ~new_n32054_;
  assign new_n32057_ = ~new_n15964_ | ~new_n31554_;
  assign new_n32058_ = ~pi1232 | ~new_n31555_;
  assign new_n32059_ = ~new_n15964_ | ~new_n31554_;
  assign new_n32060_ = ~pi1232 | ~new_n31555_;
  assign new_n32061_ = ~new_n32060_ | ~new_n32059_;
  assign new_n32062_ = ~new_n31702_ | ~new_n31703_;
  assign new_n32063_ = ~new_n31774_ | ~new_n32061_;
  assign new_n32064_ = ~new_n15965_ | ~new_n31552_;
  assign new_n32065_ = ~pi1231 | ~new_n31553_;
  assign new_n32066_ = ~new_n15965_ | ~new_n31552_;
  assign new_n32067_ = ~pi1231 | ~new_n31553_;
  assign new_n32068_ = ~new_n32067_ | ~new_n32066_;
  assign new_n32069_ = ~new_n31704_ | ~new_n31705_;
  assign new_n32070_ = ~new_n31899_ | ~new_n32068_;
  assign new_n32071_ = ~new_n15966_ | ~new_n31545_;
  assign new_n32072_ = ~pi1230 | ~new_n31546_;
  assign new_n32073_ = ~new_n15967_ | ~new_n31549_;
  assign new_n32074_ = ~pi1229 | ~new_n31550_;
  assign new_n32075_ = ~new_n32074_ | ~new_n32073_;
  assign new_n32076_ = ~new_n31831_ | ~new_n31580_;
  assign new_n32077_ = ~new_n32075_ | ~new_n31815_;
  assign new_n32078_ = ~new_n15968_ | ~new_n31547_;
  assign new_n32079_ = ~pi1228 | ~new_n31548_;
  assign new_n32080_ = ~new_n32079_ | ~new_n32078_;
  assign new_n32081_ = ~new_n31832_ | ~new_n31706_;
  assign new_n32082_ = ~new_n31812_ | ~new_n32080_;
  assign new_n32083_ = ~new_n31833_ | ~new_n31707_;
  assign new_n32084_ = ~new_n31607_ | ~new_n31763_;
  assign new_n32085_ = ~new_n15970_ | ~new_n31541_;
  assign new_n32086_ = ~pi1226 | ~new_n31542_;
  assign new_n32087_ = ~new_n15971_ | ~new_n31543_;
  assign new_n32088_ = ~pi1225 | ~new_n31544_;
  assign new_n32089_ = ~new_n32088_ | ~new_n32087_;
  assign new_n32090_ = ~new_n31834_ | ~new_n31708_;
  assign new_n32091_ = ~new_n31758_ | ~new_n32089_;
  assign new_n32092_ = ~pi1215 | ~new_n31512_;
  assign new_n32093_ = ~new_n15981_ | ~new_n31513_;
  assign new_n32094_ = new_n32363_ & new_n32361_;
  assign new_n32095_ = new_n32369_ & new_n32367_;
  assign new_n32096_ = new_n32095_ & new_n32371_;
  assign new_n32097_ = new_n32377_ & new_n32375_;
  assign new_n32098_ = new_n32097_ & new_n32379_;
  assign new_n32099_ = new_n32098_ & new_n32381_;
  assign new_n32100_ = new_n32547_ & new_n32546_;
  assign new_n32101_ = new_n32570_ & new_n32569_;
  assign new_n32102_ = new_n32644_ & new_n32643_;
  assign new_n32103_ = new_n32419_ & new_n32418_;
  assign new_n32104_ = new_n32416_ & new_n32414_;
  assign new_n32105_ = new_n32409_ & new_n32408_;
  assign new_n32106_ = new_n32406_ & new_n32404_;
  assign new_n32107_ = new_n32397_ & new_n32396_;
  assign new_n32108_ = new_n32343_ & new_n32341_;
  assign new_n32109_ = new_n32334_ & new_n32333_;
  assign new_n32110_ = new_n32331_ & new_n32329_;
  assign new_n32111_ = new_n32225_ & new_n32655_ & new_n32654_;
  assign new_n32112_ = ~new_n15533_;
  assign new_n32113_ = ~new_n15824_;
  assign new_n32114_ = ~new_n15825_;
  assign new_n32115_ = ~new_n15826_;
  assign new_n32116_ = ~new_n15827_;
  assign new_n32117_ = ~new_n15827_ | ~new_n32502_;
  assign new_n32118_ = ~new_n15830_;
  assign new_n32119_ = ~new_n15829_;
  assign new_n32120_ = ~new_n15831_;
  assign new_n32121_ = ~new_n15828_;
  assign new_n32122_ = ~new_n15823_;
  assign new_n32123_ = ~new_n15822_;
  assign new_n32124_ = ~new_n32325_ | ~new_n32309_;
  assign new_n32125_ = ~new_n32124_ | ~new_n32307_;
  assign new_n32126_ = ~new_n15804_;
  assign new_n32127_ = ~new_n15805_;
  assign new_n32128_ = ~new_n15806_;
  assign new_n32129_ = ~new_n15807_;
  assign new_n32130_ = ~new_n15808_;
  assign new_n32131_ = ~new_n15808_ | ~new_n32635_;
  assign new_n32132_ = ~new_n15809_;
  assign new_n32133_ = ~new_n15810_;
  assign new_n32134_ = ~new_n15811_;
  assign new_n32135_ = ~new_n15812_;
  assign new_n32136_ = ~new_n15812_ | ~new_n32610_;
  assign new_n32137_ = ~new_n15813_;
  assign new_n32138_ = ~new_n15814_;
  assign new_n32139_ = ~new_n15815_;
  assign new_n32140_ = ~new_n15815_ | ~new_n32590_;
  assign new_n32141_ = ~new_n15820_;
  assign new_n32142_ = ~new_n15821_;
  assign new_n32143_ = ~new_n32123_ | ~new_n32489_ | ~new_n32488_;
  assign new_n32144_ = ~new_n15816_;
  assign new_n32145_ = ~new_n15819_;
  assign new_n32146_ = ~new_n15819_ | ~new_n32560_;
  assign new_n32147_ = ~new_n15818_;
  assign new_n32148_ = ~new_n15818_ | ~new_n32552_;
  assign new_n32149_ = ~new_n15817_;
  assign new_n32150_ = ~new_n15817_ | ~new_n32555_;
  assign new_n32151_ = ~new_n15803_;
  assign new_n32152_ = ~new_n15801_;
  assign new_n32153_ = ~new_n15802_;
  assign new_n32154_ = ~new_n32295_ | ~new_n32337_;
  assign new_n32155_ = ~new_n32154_ | ~new_n32291_;
  assign new_n32156_ = ~new_n32460_ | ~new_n32382_;
  assign new_n32157_ = ~new_n32458_ | ~new_n32380_;
  assign new_n32158_ = ~new_n32453_ | ~new_n32372_;
  assign new_n32159_ = ~new_n32447_ | ~new_n32364_;
  assign new_n32160_ = ~new_n32148_ | ~new_n32400_;
  assign new_n32161_ = ~new_n32160_ | ~new_n32344_;
  assign new_n32162_ = ~new_n32322_ | ~new_n32410_;
  assign new_n32163_ = ~new_n32162_ | ~new_n32351_;
  assign new_n32164_ = ~new_n32646_ | ~new_n32645_;
  assign new_n32165_ = ~new_n32700_ | ~new_n32699_;
  assign new_n32166_ = new_n32322_ & new_n32143_;
  assign new_n32167_ = ~new_n32539_ | ~new_n32538_;
  assign new_n32168_ = new_n32318_ & new_n32317_;
  assign new_n32169_ = ~new_n32541_ | ~new_n32540_;
  assign new_n32170_ = new_n32309_ & new_n32308_;
  assign new_n32171_ = ~new_n32543_ | ~new_n32542_;
  assign new_n32172_ = new_n32314_ & new_n32117_;
  assign new_n32173_ = ~new_n32545_ | ~new_n32544_;
  assign new_n32174_ = ~new_n32664_ | ~new_n32663_;
  assign new_n32175_ = new_n32268_ & new_n32389_;
  assign new_n32176_ = ~new_n32666_ | ~new_n32665_;
  assign new_n32177_ = new_n32386_ & new_n32385_;
  assign new_n32178_ = ~new_n32668_ | ~new_n32667_;
  assign new_n32179_ = new_n32384_ & new_n32383_;
  assign new_n32180_ = ~new_n32670_ | ~new_n32669_;
  assign new_n32181_ = new_n32382_ & new_n32381_;
  assign new_n32182_ = ~new_n32672_ | ~new_n32671_;
  assign new_n32183_ = new_n32380_ & new_n32379_;
  assign new_n32184_ = ~new_n32674_ | ~new_n32673_;
  assign new_n32185_ = new_n32378_ & new_n32377_;
  assign new_n32186_ = ~new_n32676_ | ~new_n32675_;
  assign new_n32187_ = new_n32131_ & new_n32375_;
  assign new_n32188_ = ~new_n32678_ | ~new_n32677_;
  assign new_n32189_ = new_n32374_ & new_n32373_;
  assign new_n32190_ = ~new_n32680_ | ~new_n32679_;
  assign new_n32191_ = new_n32372_ & new_n32371_;
  assign new_n32192_ = ~new_n32682_ | ~new_n32681_;
  assign new_n32193_ = new_n32370_ & new_n32369_;
  assign new_n32194_ = ~new_n32684_ | ~new_n32683_;
  assign new_n32195_ = new_n32295_ & new_n32294_;
  assign new_n32196_ = ~new_n32686_ | ~new_n32685_;
  assign new_n32197_ = new_n32136_ & new_n32367_;
  assign new_n32198_ = ~new_n32688_ | ~new_n32687_;
  assign new_n32199_ = new_n32366_ & new_n32365_;
  assign new_n32200_ = ~new_n32690_ | ~new_n32689_;
  assign new_n32201_ = new_n32364_ & new_n32363_;
  assign new_n32202_ = ~new_n32692_ | ~new_n32691_;
  assign new_n32203_ = new_n32140_ & new_n32361_;
  assign new_n32204_ = ~new_n32694_ | ~new_n32693_;
  assign new_n32205_ = new_n32148_ & new_n32347_;
  assign new_n32206_ = ~new_n32696_ | ~new_n32695_;
  assign new_n32207_ = new_n32146_ & new_n32348_;
  assign new_n32208_ = ~new_n32698_ | ~new_n32697_;
  assign new_n32209_ = new_n32297_ & new_n32294_;
  assign new_n32210_ = new_n32293_ & new_n32291_;
  assign new_n32211_ = new_n32306_ & new_n32305_;
  assign new_n32212_ = new_n32293_ & new_n32292_;
  assign new_n32213_ = new_n32318_ & new_n32143_;
  assign new_n32214_ = new_n32354_ & new_n32351_;
  assign new_n32215_ = new_n32348_ & new_n32445_ & new_n32344_ & new_n32347_;
  assign new_n32216_ = new_n32442_ & new_n32443_ & new_n32444_ & new_n32345_;
  assign new_n32217_ = new_n32365_ & new_n32094_;
  assign new_n32218_ = new_n32450_ & new_n32366_;
  assign new_n32219_ = new_n32096_ & new_n32373_;
  assign new_n32220_ = new_n32455_ & new_n32374_;
  assign new_n32221_ = new_n32099_ & new_n32383_;
  assign new_n32222_ = new_n32462_ & new_n32384_;
  assign new_n32223_ = new_n32650_ & new_n32394_;
  assign new_n32224_ = new_n32393_ & new_n32102_;
  assign new_n32225_ = new_n32269_ & new_n32463_;
  assign new_n32226_ = new_n32456_ & new_n32378_;
  assign new_n32227_ = new_n32451_ & new_n32370_;
  assign new_n32228_ = new_n32346_ & new_n32345_;
  assign new_n32229_ = new_n32405_ & new_n32150_;
  assign new_n32230_ = new_n32354_ & new_n32353_;
  assign new_n32231_ = new_n32415_ & new_n32352_;
  assign new_n32232_ = ~new_n15799_;
  assign new_n32233_ = ~new_n15796_;
  assign new_n32234_ = ~new_n15795_;
  assign new_n32235_ = ~new_n15848_;
  assign new_n32236_ = ~new_n15849_;
  assign new_n32237_ = ~new_n15851_;
  assign new_n32238_ = ~new_n15852_;
  assign new_n32239_ = ~new_n15853_;
  assign new_n32240_ = ~new_n15850_;
  assign new_n32241_ = ~new_n15798_;
  assign new_n32242_ = ~new_n32317_ | ~new_n32319_;
  assign new_n32243_ = ~new_n32313_ | ~new_n32315_ | ~new_n32305_;
  assign new_n32244_ = ~new_n32117_ | ~new_n32323_;
  assign new_n32245_ = ~new_n32292_ | ~new_n32302_;
  assign new_n32246_ = ~new_n15792_;
  assign new_n32247_ = ~new_n15793_;
  assign new_n32248_ = ~new_n15794_;
  assign new_n32249_ = ~new_n15797_;
  assign new_n32250_ = ~new_n15791_;
  assign new_n32251_ = ~new_n15790_;
  assign new_n32252_ = ~new_n15847_;
  assign new_n32253_ = ~new_n15846_;
  assign new_n32254_ = ~new_n15845_;
  assign new_n32255_ = ~new_n15841_;
  assign new_n32256_ = ~new_n15842_;
  assign new_n32257_ = ~new_n15844_;
  assign new_n32258_ = ~new_n15843_;
  assign new_n32259_ = ~new_n15836_;
  assign new_n32260_ = ~new_n15837_;
  assign new_n32261_ = ~new_n15838_;
  assign new_n32262_ = ~new_n15840_;
  assign new_n32263_ = ~new_n15839_;
  assign new_n32264_ = ~new_n15835_;
  assign new_n32265_ = ~new_n15834_;
  assign new_n32266_ = ~new_n15832_;
  assign new_n32267_ = ~new_n15833_;
  assign new_n32268_ = ~new_n15802_ | ~new_n32653_;
  assign new_n32269_ = new_n32657_ & new_n32656_;
  assign new_n32270_ = new_n32659_ & new_n32658_;
  assign new_n32271_ = ~new_n32268_ | ~new_n32391_;
  assign new_n32272_ = ~new_n32386_ | ~new_n32387_;
  assign new_n32273_ = ~new_n32222_ | ~new_n32472_;
  assign new_n32274_ = ~new_n32461_ | ~new_n32470_;
  assign new_n32275_ = ~new_n32459_ | ~new_n32468_;
  assign new_n32276_ = ~new_n32226_ | ~new_n32466_;
  assign new_n32277_ = ~new_n32464_ | ~new_n32131_;
  assign new_n32278_ = ~new_n32220_ | ~new_n32474_;
  assign new_n32279_ = ~new_n32454_ | ~new_n32476_;
  assign new_n32280_ = ~new_n32227_ | ~new_n32478_;
  assign new_n32281_ = ~new_n32480_ | ~new_n32136_;
  assign new_n32282_ = ~new_n32298_ | ~new_n32335_;
  assign new_n32283_ = ~new_n32218_ | ~new_n32482_;
  assign new_n32284_ = ~new_n32448_ | ~new_n32484_;
  assign new_n32285_ = ~new_n32486_ | ~new_n32140_;
  assign new_n32286_ = ~new_n32290_ | ~new_n32216_;
  assign new_n32287_ = ~new_n32146_ | ~new_n32398_;
  assign new_n32288_ = ~new_n32356_ | ~new_n32357_ | ~new_n32353_;
  assign new_n32289_ = ~new_n32298_ | ~new_n32297_;
  assign new_n32290_ = ~new_n32215_ | ~new_n32288_;
  assign new_n32291_ = ~new_n32119_ | ~new_n32525_ | ~new_n32524_;
  assign new_n32292_ = ~new_n15828_ | ~new_n32530_;
  assign new_n32293_ = ~new_n32121_ | ~new_n32527_ | ~new_n32526_;
  assign new_n32294_ = ~new_n32118_ | ~new_n32521_ | ~new_n32520_;
  assign new_n32295_ = ~new_n15830_ | ~new_n32516_;
  assign new_n32296_ = ~new_n15829_ | ~new_n32513_;
  assign new_n32297_ = ~new_n32120_ | ~new_n32523_ | ~new_n32522_;
  assign new_n32298_ = ~new_n15831_ | ~new_n32519_;
  assign new_n32299_ = ~new_n32298_ | ~new_n32112_;
  assign new_n32300_ = ~new_n32209_ | ~new_n32299_;
  assign new_n32301_ = ~new_n32296_ | ~new_n32300_ | ~new_n32295_;
  assign new_n32302_ = ~new_n32210_ | ~new_n32301_;
  assign new_n32303_ = ~new_n32245_;
  assign new_n32304_ = ~new_n15825_ | ~new_n32497_;
  assign new_n32305_ = ~new_n15824_ | ~new_n32510_;
  assign new_n32306_ = ~new_n32113_ | ~new_n32494_ | ~new_n32493_;
  assign new_n32307_ = ~new_n32114_ | ~new_n32507_ | ~new_n32506_;
  assign new_n32308_ = ~new_n32115_ | ~new_n32499_ | ~new_n32498_;
  assign new_n32309_ = ~new_n15826_ | ~new_n32505_;
  assign new_n32310_ = ~new_n32117_;
  assign new_n32311_ = ~new_n32310_ | ~new_n32308_;
  assign new_n32312_ = ~new_n32304_ | ~new_n32309_ | ~new_n32311_;
  assign new_n32313_ = ~new_n32306_ | ~new_n32307_ | ~new_n32312_;
  assign new_n32314_ = ~new_n32116_ | ~new_n32532_ | ~new_n32531_;
  assign new_n32315_ = ~new_n32314_ | ~new_n32306_ | ~new_n32307_ | ~new_n32308_ | ~new_n32245_;
  assign new_n32316_ = ~new_n32243_;
  assign new_n32317_ = ~new_n15823_ | ~new_n32537_;
  assign new_n32318_ = ~new_n32122_ | ~new_n32534_ | ~new_n32533_;
  assign new_n32319_ = ~new_n32318_ | ~new_n32243_;
  assign new_n32320_ = ~new_n32242_;
  assign new_n32321_ = ~new_n32143_;
  assign new_n32322_ = ~new_n15822_ | ~new_n32492_;
  assign new_n32323_ = ~new_n32314_ | ~new_n32245_;
  assign new_n32324_ = ~new_n32244_;
  assign new_n32325_ = ~new_n32244_ | ~new_n32308_;
  assign new_n32326_ = ~new_n32124_;
  assign new_n32327_ = ~new_n32125_;
  assign new_n32328_ = ~new_n32125_ | ~new_n32304_;
  assign new_n32329_ = ~new_n32211_ | ~new_n32328_;
  assign new_n32330_ = ~new_n32306_ | ~new_n32305_;
  assign new_n32331_ = ~new_n32330_ | ~new_n32125_ | ~new_n32304_;
  assign new_n32332_ = ~new_n32307_ | ~new_n32304_;
  assign new_n32333_ = ~new_n32326_ | ~new_n32332_;
  assign new_n32334_ = ~new_n32327_ | ~new_n32304_;
  assign new_n32335_ = ~new_n15533_ | ~new_n32297_;
  assign new_n32336_ = ~new_n32282_;
  assign new_n32337_ = ~new_n32282_ | ~new_n32294_;
  assign new_n32338_ = ~new_n32154_;
  assign new_n32339_ = ~new_n32155_;
  assign new_n32340_ = ~new_n32155_ | ~new_n32296_;
  assign new_n32341_ = ~new_n32212_ | ~new_n32340_;
  assign new_n32342_ = ~new_n32293_ | ~new_n32292_;
  assign new_n32343_ = ~new_n32342_ | ~new_n32155_ | ~new_n32296_;
  assign new_n32344_ = ~new_n32149_ | ~new_n32549_ | ~new_n32548_;
  assign new_n32345_ = ~new_n15816_ | ~new_n32563_;
  assign new_n32346_ = ~new_n32100_ | ~new_n32144_;
  assign new_n32347_ = ~new_n32147_ | ~new_n32557_ | ~new_n32556_;
  assign new_n32348_ = ~new_n32145_ | ~new_n32575_ | ~new_n32574_;
  assign new_n32349_ = ~new_n32148_;
  assign new_n32350_ = ~new_n32150_;
  assign new_n32351_ = ~new_n32142_ | ~new_n32565_ | ~new_n32564_;
  assign new_n32352_ = ~new_n15821_ | ~new_n32568_;
  assign new_n32353_ = ~new_n15820_ | ~new_n32573_;
  assign new_n32354_ = ~new_n32101_ | ~new_n32141_;
  assign new_n32355_ = ~new_n32352_ | ~new_n32322_ | ~new_n32317_;
  assign new_n32356_ = ~new_n32446_ | ~new_n32351_ | ~new_n32355_ | ~new_n32449_;
  assign new_n32357_ = ~new_n32214_ | ~new_n32213_ | ~new_n32243_;
  assign new_n32358_ = ~new_n32288_;
  assign new_n32359_ = ~new_n32146_;
  assign new_n32360_ = ~new_n32286_;
  assign new_n32361_ = ~new_n32139_ | ~new_n32577_ | ~new_n32576_;
  assign new_n32362_ = ~new_n32140_;
  assign new_n32363_ = ~new_n32138_ | ~new_n32579_ | ~new_n32578_;
  assign new_n32364_ = ~new_n15814_ | ~new_n32587_;
  assign new_n32365_ = ~new_n32137_ | ~new_n32581_ | ~new_n32580_;
  assign new_n32366_ = ~new_n15813_ | ~new_n32584_;
  assign new_n32367_ = ~new_n32135_ | ~new_n32596_ | ~new_n32595_;
  assign new_n32368_ = ~new_n32136_;
  assign new_n32369_ = ~new_n32134_ | ~new_n32598_ | ~new_n32597_;
  assign new_n32370_ = ~new_n15811_ | ~new_n32607_;
  assign new_n32371_ = ~new_n32133_ | ~new_n32594_ | ~new_n32593_;
  assign new_n32372_ = ~new_n15810_ | ~new_n32604_;
  assign new_n32373_ = ~new_n32132_ | ~new_n32592_ | ~new_n32591_;
  assign new_n32374_ = ~new_n15809_ | ~new_n32601_;
  assign new_n32375_ = ~new_n32130_ | ~new_n32618_ | ~new_n32617_;
  assign new_n32376_ = ~new_n32131_;
  assign new_n32377_ = ~new_n32129_ | ~new_n32620_ | ~new_n32619_;
  assign new_n32378_ = ~new_n15807_ | ~new_n32632_;
  assign new_n32379_ = ~new_n32128_ | ~new_n32616_ | ~new_n32615_;
  assign new_n32380_ = ~new_n15806_ | ~new_n32629_;
  assign new_n32381_ = ~new_n32127_ | ~new_n32614_ | ~new_n32613_;
  assign new_n32382_ = ~new_n15805_ | ~new_n32626_;
  assign new_n32383_ = ~new_n32126_ | ~new_n32612_ | ~new_n32611_;
  assign new_n32384_ = ~new_n15804_ | ~new_n32623_;
  assign new_n32385_ = ~new_n32151_ | ~new_n32637_ | ~new_n32636_;
  assign new_n32386_ = ~new_n15803_ | ~new_n32640_;
  assign new_n32387_ = ~new_n32385_ | ~new_n32273_;
  assign new_n32388_ = ~new_n32272_;
  assign new_n32389_ = ~new_n32153_ | ~new_n32642_ | ~new_n32641_;
  assign new_n32390_ = ~new_n32268_;
  assign new_n32391_ = ~new_n32389_ | ~new_n32272_;
  assign new_n32392_ = ~new_n32271_;
  assign new_n32393_ = ~new_n15801_ | ~new_n32164_;
  assign new_n32394_ = ~new_n32647_ | ~new_n32152_;
  assign new_n32395_ = ~new_n32296_ | ~new_n32291_;
  assign new_n32396_ = ~new_n32338_ | ~new_n32395_;
  assign new_n32397_ = ~new_n32339_ | ~new_n32296_;
  assign new_n32398_ = ~new_n32288_ | ~new_n32348_;
  assign new_n32399_ = ~new_n32287_;
  assign new_n32400_ = ~new_n32287_ | ~new_n32347_;
  assign new_n32401_ = ~new_n32160_;
  assign new_n32402_ = ~new_n32161_;
  assign new_n32403_ = ~new_n32161_ | ~new_n32150_;
  assign new_n32404_ = ~new_n32228_ | ~new_n32403_;
  assign new_n32405_ = ~new_n32346_ | ~new_n32345_;
  assign new_n32406_ = ~new_n32229_ | ~new_n32161_;
  assign new_n32407_ = ~new_n32150_ | ~new_n32344_;
  assign new_n32408_ = ~new_n32401_ | ~new_n32407_;
  assign new_n32409_ = ~new_n32402_ | ~new_n32150_;
  assign new_n32410_ = ~new_n32143_ | ~new_n32242_;
  assign new_n32411_ = ~new_n32162_;
  assign new_n32412_ = ~new_n32163_;
  assign new_n32413_ = ~new_n32163_ | ~new_n32352_;
  assign new_n32414_ = ~new_n32230_ | ~new_n32413_;
  assign new_n32415_ = ~new_n32354_ | ~new_n32353_;
  assign new_n32416_ = ~new_n32231_ | ~new_n32163_;
  assign new_n32417_ = ~new_n32352_ | ~new_n32351_;
  assign new_n32418_ = ~new_n32411_ | ~new_n32417_;
  assign new_n32419_ = ~new_n32412_ | ~new_n32352_;
  assign new_n32420_ = ~new_n32289_;
  assign new_n32421_ = ~new_n32322_ | ~new_n32143_;
  assign new_n32422_ = ~new_n32318_ | ~new_n32317_;
  assign new_n32423_ = ~new_n32309_ | ~new_n32308_;
  assign new_n32424_ = ~new_n32314_ | ~new_n32117_;
  assign new_n32425_ = ~new_n32268_ | ~new_n32389_;
  assign new_n32426_ = ~new_n32386_ | ~new_n32385_;
  assign new_n32427_ = ~new_n32384_ | ~new_n32383_;
  assign new_n32428_ = ~new_n32382_ | ~new_n32381_;
  assign new_n32429_ = ~new_n32380_ | ~new_n32379_;
  assign new_n32430_ = ~new_n32378_ | ~new_n32377_;
  assign new_n32431_ = ~new_n32131_ | ~new_n32375_;
  assign new_n32432_ = ~new_n32374_ | ~new_n32373_;
  assign new_n32433_ = ~new_n32372_ | ~new_n32371_;
  assign new_n32434_ = ~new_n32370_ | ~new_n32369_;
  assign new_n32435_ = ~new_n32295_ | ~new_n32294_;
  assign new_n32436_ = ~new_n32136_ | ~new_n32367_;
  assign new_n32437_ = ~new_n32366_ | ~new_n32365_;
  assign new_n32438_ = ~new_n32364_ | ~new_n32363_;
  assign new_n32439_ = ~new_n32140_ | ~new_n32361_;
  assign new_n32440_ = ~new_n32148_ | ~new_n32347_;
  assign new_n32441_ = ~new_n32146_ | ~new_n32348_;
  assign new_n32442_ = ~new_n32347_ | ~new_n32346_ | ~new_n32344_ | ~new_n32359_;
  assign new_n32443_ = ~new_n32346_ | ~new_n32349_ | ~new_n32344_;
  assign new_n32444_ = ~new_n32350_ | ~new_n32346_;
  assign new_n32445_ = ~new_n32100_ | ~new_n32144_;
  assign new_n32446_ = ~new_n32321_ | ~new_n32352_;
  assign new_n32447_ = ~new_n32362_ | ~new_n32363_;
  assign new_n32448_ = ~new_n32159_;
  assign new_n32449_ = ~new_n32101_ | ~new_n32141_;
  assign new_n32450_ = ~new_n32159_ | ~new_n32365_;
  assign new_n32451_ = ~new_n32368_ | ~new_n32369_;
  assign new_n32452_ = ~new_n32451_ | ~new_n32370_;
  assign new_n32453_ = ~new_n32452_ | ~new_n32371_;
  assign new_n32454_ = ~new_n32158_;
  assign new_n32455_ = ~new_n32158_ | ~new_n32373_;
  assign new_n32456_ = ~new_n32376_ | ~new_n32377_;
  assign new_n32457_ = ~new_n32456_ | ~new_n32378_;
  assign new_n32458_ = ~new_n32457_ | ~new_n32379_;
  assign new_n32459_ = ~new_n32157_;
  assign new_n32460_ = ~new_n32157_ | ~new_n32381_;
  assign new_n32461_ = ~new_n32156_;
  assign new_n32462_ = ~new_n32156_ | ~new_n32383_;
  assign new_n32463_ = ~new_n32223_ | ~new_n32389_ | ~new_n32272_;
  assign new_n32464_ = ~new_n32375_ | ~new_n32278_;
  assign new_n32465_ = ~new_n32277_;
  assign new_n32466_ = ~new_n32097_ | ~new_n32278_;
  assign new_n32467_ = ~new_n32276_;
  assign new_n32468_ = ~new_n32098_ | ~new_n32278_;
  assign new_n32469_ = ~new_n32275_;
  assign new_n32470_ = ~new_n32099_ | ~new_n32278_;
  assign new_n32471_ = ~new_n32274_;
  assign new_n32472_ = ~new_n32221_ | ~new_n32278_;
  assign new_n32473_ = ~new_n32273_;
  assign new_n32474_ = ~new_n32219_ | ~new_n32283_;
  assign new_n32475_ = ~new_n32278_;
  assign new_n32476_ = ~new_n32096_ | ~new_n32283_;
  assign new_n32477_ = ~new_n32279_;
  assign new_n32478_ = ~new_n32095_ | ~new_n32283_;
  assign new_n32479_ = ~new_n32280_;
  assign new_n32480_ = ~new_n32367_ | ~new_n32283_;
  assign new_n32481_ = ~new_n32281_;
  assign new_n32482_ = ~new_n32217_ | ~new_n32286_;
  assign new_n32483_ = ~new_n32283_;
  assign new_n32484_ = ~new_n32094_ | ~new_n32286_;
  assign new_n32485_ = ~new_n32284_;
  assign new_n32486_ = ~new_n32361_ | ~new_n32286_;
  assign new_n32487_ = ~new_n32285_;
  assign new_n32488_ = ~new_n15533_ | ~new_n32232_;
  assign new_n32489_ = ~new_n15799_ | ~new_n32112_;
  assign new_n32490_ = ~new_n15533_ | ~new_n32232_;
  assign new_n32491_ = ~new_n15799_ | ~new_n32112_;
  assign new_n32492_ = ~new_n32491_ | ~new_n32490_;
  assign new_n32493_ = ~new_n15533_ | ~new_n32233_;
  assign new_n32494_ = ~new_n15796_ | ~new_n32112_;
  assign new_n32495_ = ~new_n15533_ | ~new_n32234_;
  assign new_n32496_ = ~new_n15795_ | ~new_n32112_;
  assign new_n32497_ = ~new_n32496_ | ~new_n32495_;
  assign new_n32498_ = ~new_n15533_ | ~new_n32235_;
  assign new_n32499_ = ~new_n15848_ | ~new_n32112_;
  assign new_n32500_ = ~new_n15533_ | ~new_n32236_;
  assign new_n32501_ = ~new_n15849_ | ~new_n32112_;
  assign new_n32502_ = ~new_n32501_ | ~new_n32500_;
  assign new_n32503_ = ~new_n15533_ | ~new_n32235_;
  assign new_n32504_ = ~new_n15848_ | ~new_n32112_;
  assign new_n32505_ = ~new_n32504_ | ~new_n32503_;
  assign new_n32506_ = ~new_n15533_ | ~new_n32234_;
  assign new_n32507_ = ~new_n15795_ | ~new_n32112_;
  assign new_n32508_ = ~new_n15533_ | ~new_n32233_;
  assign new_n32509_ = ~new_n15796_ | ~new_n32112_;
  assign new_n32510_ = ~new_n32509_ | ~new_n32508_;
  assign new_n32511_ = ~new_n15533_ | ~new_n32237_;
  assign new_n32512_ = ~new_n15851_ | ~new_n32112_;
  assign new_n32513_ = ~new_n32512_ | ~new_n32511_;
  assign new_n32514_ = ~new_n15533_ | ~new_n32238_;
  assign new_n32515_ = ~new_n15852_ | ~new_n32112_;
  assign new_n32516_ = ~new_n32515_ | ~new_n32514_;
  assign new_n32517_ = ~new_n15533_ | ~new_n32239_;
  assign new_n32518_ = ~new_n15853_ | ~new_n32112_;
  assign new_n32519_ = ~new_n32518_ | ~new_n32517_;
  assign new_n32520_ = ~new_n15533_ | ~new_n32238_;
  assign new_n32521_ = ~new_n15852_ | ~new_n32112_;
  assign new_n32522_ = ~new_n15533_ | ~new_n32239_;
  assign new_n32523_ = ~new_n15853_ | ~new_n32112_;
  assign new_n32524_ = ~new_n15533_ | ~new_n32237_;
  assign new_n32525_ = ~new_n15851_ | ~new_n32112_;
  assign new_n32526_ = ~new_n15533_ | ~new_n32240_;
  assign new_n32527_ = ~new_n15850_ | ~new_n32112_;
  assign new_n32528_ = ~new_n15533_ | ~new_n32240_;
  assign new_n32529_ = ~new_n15850_ | ~new_n32112_;
  assign new_n32530_ = ~new_n32529_ | ~new_n32528_;
  assign new_n32531_ = ~new_n15533_ | ~new_n32236_;
  assign new_n32532_ = ~new_n15849_ | ~new_n32112_;
  assign new_n32533_ = ~new_n15533_ | ~new_n32241_;
  assign new_n32534_ = ~new_n15798_ | ~new_n32112_;
  assign new_n32535_ = ~new_n15533_ | ~new_n32241_;
  assign new_n32536_ = ~new_n15798_ | ~new_n32112_;
  assign new_n32537_ = ~new_n32536_ | ~new_n32535_;
  assign new_n32538_ = ~new_n32421_ | ~new_n32242_;
  assign new_n32539_ = ~new_n32166_ | ~new_n32320_;
  assign new_n32540_ = ~new_n32422_ | ~new_n32243_;
  assign new_n32541_ = ~new_n32168_ | ~new_n32316_;
  assign new_n32542_ = ~new_n32423_ | ~new_n32244_;
  assign new_n32543_ = ~new_n32170_ | ~new_n32324_;
  assign new_n32544_ = ~new_n32424_ | ~new_n32245_;
  assign new_n32545_ = ~new_n32172_ | ~new_n32303_;
  assign new_n32546_ = ~new_n15533_ | ~new_n32246_;
  assign new_n32547_ = ~new_n15792_ | ~new_n32112_;
  assign new_n32548_ = ~new_n15533_ | ~new_n32247_;
  assign new_n32549_ = ~new_n15793_ | ~new_n32112_;
  assign new_n32550_ = ~new_n15533_ | ~new_n32248_;
  assign new_n32551_ = ~new_n15794_ | ~new_n32112_;
  assign new_n32552_ = ~new_n32551_ | ~new_n32550_;
  assign new_n32553_ = ~new_n15533_ | ~new_n32247_;
  assign new_n32554_ = ~new_n15793_ | ~new_n32112_;
  assign new_n32555_ = ~new_n32554_ | ~new_n32553_;
  assign new_n32556_ = ~new_n15533_ | ~new_n32248_;
  assign new_n32557_ = ~new_n15794_ | ~new_n32112_;
  assign new_n32558_ = ~new_n15533_ | ~new_n32249_;
  assign new_n32559_ = ~new_n15797_ | ~new_n32112_;
  assign new_n32560_ = ~new_n32559_ | ~new_n32558_;
  assign new_n32561_ = ~new_n15533_ | ~new_n32246_;
  assign new_n32562_ = ~new_n15792_ | ~new_n32112_;
  assign new_n32563_ = ~new_n32562_ | ~new_n32561_;
  assign new_n32564_ = ~new_n15533_ | ~new_n32250_;
  assign new_n32565_ = ~new_n15791_ | ~new_n32112_;
  assign new_n32566_ = ~new_n15533_ | ~new_n32250_;
  assign new_n32567_ = ~new_n15791_ | ~new_n32112_;
  assign new_n32568_ = ~new_n32567_ | ~new_n32566_;
  assign new_n32569_ = ~new_n15533_ | ~new_n32251_;
  assign new_n32570_ = ~new_n15790_ | ~new_n32112_;
  assign new_n32571_ = ~new_n15533_ | ~new_n32251_;
  assign new_n32572_ = ~new_n15790_ | ~new_n32112_;
  assign new_n32573_ = ~new_n32572_ | ~new_n32571_;
  assign new_n32574_ = ~new_n15533_ | ~new_n32249_;
  assign new_n32575_ = ~new_n15797_ | ~new_n32112_;
  assign new_n32576_ = ~new_n15533_ | ~new_n32252_;
  assign new_n32577_ = ~new_n15847_ | ~new_n32112_;
  assign new_n32578_ = ~new_n15533_ | ~new_n32253_;
  assign new_n32579_ = ~new_n15846_ | ~new_n32112_;
  assign new_n32580_ = ~new_n15533_ | ~new_n32254_;
  assign new_n32581_ = ~new_n15845_ | ~new_n32112_;
  assign new_n32582_ = ~new_n15533_ | ~new_n32254_;
  assign new_n32583_ = ~new_n15845_ | ~new_n32112_;
  assign new_n32584_ = ~new_n32583_ | ~new_n32582_;
  assign new_n32585_ = ~new_n15533_ | ~new_n32253_;
  assign new_n32586_ = ~new_n15846_ | ~new_n32112_;
  assign new_n32587_ = ~new_n32586_ | ~new_n32585_;
  assign new_n32588_ = ~new_n15533_ | ~new_n32252_;
  assign new_n32589_ = ~new_n15847_ | ~new_n32112_;
  assign new_n32590_ = ~new_n32589_ | ~new_n32588_;
  assign new_n32591_ = ~new_n15533_ | ~new_n32255_;
  assign new_n32592_ = ~new_n15841_ | ~new_n32112_;
  assign new_n32593_ = ~new_n15533_ | ~new_n32256_;
  assign new_n32594_ = ~new_n15842_ | ~new_n32112_;
  assign new_n32595_ = ~new_n15533_ | ~new_n32257_;
  assign new_n32596_ = ~new_n15844_ | ~new_n32112_;
  assign new_n32597_ = ~new_n15533_ | ~new_n32258_;
  assign new_n32598_ = ~new_n15843_ | ~new_n32112_;
  assign new_n32599_ = ~new_n15533_ | ~new_n32255_;
  assign new_n32600_ = ~new_n15841_ | ~new_n32112_;
  assign new_n32601_ = ~new_n32600_ | ~new_n32599_;
  assign new_n32602_ = ~new_n15533_ | ~new_n32256_;
  assign new_n32603_ = ~new_n15842_ | ~new_n32112_;
  assign new_n32604_ = ~new_n32603_ | ~new_n32602_;
  assign new_n32605_ = ~new_n15533_ | ~new_n32258_;
  assign new_n32606_ = ~new_n15843_ | ~new_n32112_;
  assign new_n32607_ = ~new_n32606_ | ~new_n32605_;
  assign new_n32608_ = ~new_n15533_ | ~new_n32257_;
  assign new_n32609_ = ~new_n15844_ | ~new_n32112_;
  assign new_n32610_ = ~new_n32609_ | ~new_n32608_;
  assign new_n32611_ = ~new_n15533_ | ~new_n32259_;
  assign new_n32612_ = ~new_n15836_ | ~new_n32112_;
  assign new_n32613_ = ~new_n15533_ | ~new_n32260_;
  assign new_n32614_ = ~new_n15837_ | ~new_n32112_;
  assign new_n32615_ = ~new_n15533_ | ~new_n32261_;
  assign new_n32616_ = ~new_n15838_ | ~new_n32112_;
  assign new_n32617_ = ~new_n15533_ | ~new_n32262_;
  assign new_n32618_ = ~new_n15840_ | ~new_n32112_;
  assign new_n32619_ = ~new_n15533_ | ~new_n32263_;
  assign new_n32620_ = ~new_n15839_ | ~new_n32112_;
  assign new_n32621_ = ~new_n15533_ | ~new_n32259_;
  assign new_n32622_ = ~new_n15836_ | ~new_n32112_;
  assign new_n32623_ = ~new_n32622_ | ~new_n32621_;
  assign new_n32624_ = ~new_n15533_ | ~new_n32260_;
  assign new_n32625_ = ~new_n15837_ | ~new_n32112_;
  assign new_n32626_ = ~new_n32625_ | ~new_n32624_;
  assign new_n32627_ = ~new_n15533_ | ~new_n32261_;
  assign new_n32628_ = ~new_n15838_ | ~new_n32112_;
  assign new_n32629_ = ~new_n32628_ | ~new_n32627_;
  assign new_n32630_ = ~new_n15533_ | ~new_n32263_;
  assign new_n32631_ = ~new_n15839_ | ~new_n32112_;
  assign new_n32632_ = ~new_n32631_ | ~new_n32630_;
  assign new_n32633_ = ~new_n15533_ | ~new_n32262_;
  assign new_n32634_ = ~new_n15840_ | ~new_n32112_;
  assign new_n32635_ = ~new_n32634_ | ~new_n32633_;
  assign new_n32636_ = ~new_n15533_ | ~new_n32264_;
  assign new_n32637_ = ~new_n15835_ | ~new_n32112_;
  assign new_n32638_ = ~new_n15533_ | ~new_n32264_;
  assign new_n32639_ = ~new_n15835_ | ~new_n32112_;
  assign new_n32640_ = ~new_n32639_ | ~new_n32638_;
  assign new_n32641_ = ~new_n15533_ | ~new_n32265_;
  assign new_n32642_ = ~new_n15834_ | ~new_n32112_;
  assign new_n32643_ = ~new_n15533_ | ~new_n32266_;
  assign new_n32644_ = ~new_n15832_ | ~new_n32112_;
  assign new_n32645_ = ~new_n15533_ | ~new_n32267_;
  assign new_n32646_ = ~new_n15833_ | ~new_n32112_;
  assign new_n32647_ = ~new_n32164_;
  assign new_n32648_ = ~new_n15533_ | ~new_n32266_;
  assign new_n32649_ = ~new_n15832_ | ~new_n32112_;
  assign new_n32650_ = ~new_n32649_ | ~new_n32648_;
  assign new_n32651_ = ~new_n15533_ | ~new_n32265_;
  assign new_n32652_ = ~new_n15834_ | ~new_n32112_;
  assign new_n32653_ = ~new_n32652_ | ~new_n32651_;
  assign new_n32654_ = ~new_n32268_ | ~new_n32224_ | ~new_n32391_;
  assign new_n32655_ = ~new_n32390_ | ~new_n32650_ | ~new_n32394_;
  assign new_n32656_ = ~new_n32152_ | ~new_n32102_ | ~new_n32647_;
  assign new_n32657_ = ~new_n15801_ | ~new_n32650_ | ~new_n32164_;
  assign new_n32658_ = ~new_n32647_ | ~new_n15801_;
  assign new_n32659_ = ~new_n32164_ | ~new_n32152_;
  assign new_n32660_ = ~new_n32647_ | ~new_n15801_;
  assign new_n32661_ = ~new_n32164_ | ~new_n32152_;
  assign new_n32662_ = ~new_n32661_ | ~new_n32660_;
  assign new_n32663_ = ~new_n32270_ | ~new_n32271_;
  assign new_n32664_ = ~new_n32392_ | ~new_n32662_;
  assign new_n32665_ = ~new_n32425_ | ~new_n32272_;
  assign new_n32666_ = ~new_n32175_ | ~new_n32388_;
  assign new_n32667_ = ~new_n32273_ | ~new_n32426_;
  assign new_n32668_ = ~new_n32177_ | ~new_n32473_;
  assign new_n32669_ = ~new_n32274_ | ~new_n32427_;
  assign new_n32670_ = ~new_n32179_ | ~new_n32471_;
  assign new_n32671_ = ~new_n32275_ | ~new_n32428_;
  assign new_n32672_ = ~new_n32181_ | ~new_n32469_;
  assign new_n32673_ = ~new_n32276_ | ~new_n32429_;
  assign new_n32674_ = ~new_n32183_ | ~new_n32467_;
  assign new_n32675_ = ~new_n32277_ | ~new_n32430_;
  assign new_n32676_ = ~new_n32185_ | ~new_n32465_;
  assign new_n32677_ = ~new_n32278_ | ~new_n32431_;
  assign new_n32678_ = ~new_n32187_ | ~new_n32475_;
  assign new_n32679_ = ~new_n32279_ | ~new_n32432_;
  assign new_n32680_ = ~new_n32189_ | ~new_n32477_;
  assign new_n32681_ = ~new_n32280_ | ~new_n32433_;
  assign new_n32682_ = ~new_n32191_ | ~new_n32479_;
  assign new_n32683_ = ~new_n32281_ | ~new_n32434_;
  assign new_n32684_ = ~new_n32193_ | ~new_n32481_;
  assign new_n32685_ = ~new_n32435_ | ~new_n32282_;
  assign new_n32686_ = ~new_n32195_ | ~new_n32336_;
  assign new_n32687_ = ~new_n32283_ | ~new_n32436_;
  assign new_n32688_ = ~new_n32197_ | ~new_n32483_;
  assign new_n32689_ = ~new_n32284_ | ~new_n32437_;
  assign new_n32690_ = ~new_n32199_ | ~new_n32485_;
  assign new_n32691_ = ~new_n32285_ | ~new_n32438_;
  assign new_n32692_ = ~new_n32201_ | ~new_n32487_;
  assign new_n32693_ = ~new_n32439_ | ~new_n32286_;
  assign new_n32694_ = ~new_n32203_ | ~new_n32360_;
  assign new_n32695_ = ~new_n32440_ | ~new_n32287_;
  assign new_n32696_ = ~new_n32205_ | ~new_n32399_;
  assign new_n32697_ = ~new_n32441_ | ~new_n32288_;
  assign new_n32698_ = ~new_n32207_ | ~new_n32358_;
  assign new_n32699_ = ~new_n15533_ | ~new_n32289_;
  assign new_n32700_ = ~new_n32420_ | ~new_n32112_;
  assign new_n32701_ = new_n32703_ | new_n15854_;
  assign new_n32702_ = new_n32705_ & new_n32704_;
  assign new_n32703_ = ~new_n32707_ & ~new_n32706_ & ~new_n32702_;
  assign new_n32704_ = ~new_n15857_;
  assign new_n32705_ = ~new_n15858_;
  assign new_n32706_ = ~new_n15855_;
  assign new_n32707_ = ~new_n15856_;
  assign new_n32708_ = ~new_n17371_;
  assign new_n32709_ = ~new_n17370_;
  assign new_n32710_ = ~new_n15859_;
  assign new_n32711_ = ~new_n32792_ | ~new_n32841_;
  assign new_n32712_ = ~new_n32793_ | ~new_n32859_;
  assign new_n32713_ = ~new_n32794_ | ~new_n32861_;
  assign new_n32714_ = ~new_n32795_ | ~new_n32863_;
  assign new_n32715_ = ~new_n32796_ | ~new_n32865_;
  assign new_n32716_ = ~new_n32797_ | ~new_n32867_;
  assign new_n32717_ = ~new_n32798_ | ~new_n32869_;
  assign new_n32718_ = ~new_n32799_ | ~new_n32871_;
  assign new_n32719_ = ~new_n32873_ | ~new_n32759_;
  assign new_n32720_ = ~new_n32874_ | ~new_n32758_;
  assign new_n32721_ = ~new_n32875_ | ~new_n32757_;
  assign new_n32722_ = ~new_n32876_ | ~new_n32756_;
  assign new_n32723_ = ~new_n32877_ | ~new_n32755_;
  assign new_n32724_ = ~new_n32878_ | ~new_n32754_;
  assign new_n32725_ = ~new_n32879_ | ~new_n32753_;
  assign new_n32726_ = ~new_n32880_ | ~new_n32752_;
  assign new_n32727_ = ~new_n32881_ | ~new_n32751_;
  assign new_n32728_ = ~new_n32882_ | ~new_n32750_;
  assign new_n32729_ = ~new_n32883_ | ~new_n32749_;
  assign new_n32730_ = ~new_n32914_ | ~new_n32913_;
  assign new_n32731_ = ~new_n32887_ | ~new_n32886_;
  assign new_n32732_ = ~new_n32908_ | ~new_n32907_;
  assign new_n32733_ = ~new_n32911_ | ~new_n32910_;
  assign new_n32734_ = ~new_n32902_ | ~new_n32901_;
  assign new_n32735_ = ~new_n32905_ | ~new_n32904_;
  assign new_n32736_ = ~new_n32890_ | ~new_n32889_;
  assign new_n32737_ = ~new_n32893_ | ~new_n32892_;
  assign new_n32738_ = ~new_n32899_ | ~new_n32898_;
  assign new_n32739_ = ~new_n32896_ | ~new_n32895_;
  assign new_n32740_ = ~new_n32917_ | ~new_n32916_;
  assign new_n32741_ = ~new_n32919_ | ~new_n32918_;
  assign new_n32742_ = ~new_n32921_ | ~new_n32920_;
  assign new_n32743_ = ~new_n32923_ | ~new_n32922_;
  assign new_n32744_ = ~new_n32925_ | ~new_n32924_;
  assign new_n32745_ = ~new_n32927_ | ~new_n32926_;
  assign new_n32746_ = ~new_n32929_ | ~new_n32928_;
  assign new_n32747_ = ~new_n32988_ | ~new_n32987_;
  assign new_n32748_ = ~new_n32991_ | ~new_n32990_;
  assign new_n32749_ = ~new_n32931_ | ~new_n32930_;
  assign new_n32750_ = ~new_n32934_ | ~new_n32933_;
  assign new_n32751_ = ~new_n32937_ | ~new_n32936_;
  assign new_n32752_ = ~new_n32940_ | ~new_n32939_;
  assign new_n32753_ = ~new_n32943_ | ~new_n32942_;
  assign new_n32754_ = ~new_n32946_ | ~new_n32945_;
  assign new_n32755_ = ~new_n32949_ | ~new_n32948_;
  assign new_n32756_ = ~new_n32952_ | ~new_n32951_;
  assign new_n32757_ = ~new_n32955_ | ~new_n32954_;
  assign new_n32758_ = ~new_n32958_ | ~new_n32957_;
  assign new_n32759_ = ~new_n32961_ | ~new_n32960_;
  assign new_n32760_ = ~new_n32982_ | ~new_n32981_;
  assign new_n32761_ = ~new_n32985_ | ~new_n32984_;
  assign new_n32762_ = ~new_n32976_ | ~new_n32975_;
  assign new_n32763_ = ~new_n32979_ | ~new_n32978_;
  assign new_n32764_ = ~new_n32970_ | ~new_n32969_;
  assign new_n32765_ = ~new_n32973_ | ~new_n32972_;
  assign new_n32766_ = ~new_n32964_ | ~new_n32963_;
  assign new_n32767_ = ~new_n32967_ | ~new_n32966_;
  assign new_n32768_ = ~new_n32997_ | ~new_n32996_;
  assign new_n32769_ = ~new_n32999_ | ~new_n32998_;
  assign new_n32770_ = ~new_n33003_ | ~new_n33002_;
  assign new_n32771_ = ~new_n33005_ | ~new_n33004_;
  assign new_n32772_ = ~new_n33007_ | ~new_n33006_;
  assign new_n32773_ = ~new_n33009_ | ~new_n33008_;
  assign new_n32774_ = ~new_n33011_ | ~new_n33010_;
  assign new_n32775_ = ~new_n33013_ | ~new_n33012_;
  assign new_n32776_ = ~new_n33015_ | ~new_n33014_;
  assign new_n32777_ = ~new_n33017_ | ~new_n33016_;
  assign new_n32778_ = ~new_n33019_ | ~new_n33018_;
  assign new_n32779_ = ~new_n33021_ | ~new_n33020_;
  assign new_n32780_ = ~new_n33030_ | ~new_n33029_;
  assign new_n32781_ = ~new_n33032_ | ~new_n33031_;
  assign new_n32782_ = ~new_n33034_ | ~new_n33033_;
  assign new_n32783_ = ~new_n33036_ | ~new_n33035_;
  assign new_n32784_ = ~new_n33038_ | ~new_n33037_;
  assign new_n32785_ = ~new_n33040_ | ~new_n33039_;
  assign new_n32786_ = ~new_n33042_ | ~new_n33041_;
  assign new_n32787_ = ~new_n33044_ | ~new_n33043_;
  assign new_n32788_ = ~new_n33046_ | ~new_n33045_;
  assign new_n32789_ = ~new_n33048_ | ~new_n33047_;
  assign new_n32790_ = ~new_n33053_ | ~new_n33052_;
  assign new_n32791_ = ~new_n33028_ | ~new_n33027_;
  assign new_n32792_ = new_n32738_ & new_n32739_;
  assign new_n32793_ = new_n32735_ & new_n32734_;
  assign new_n32794_ = new_n32733_ & new_n32732_;
  assign new_n32795_ = new_n32730_ & new_n32731_;
  assign new_n32796_ = new_n32767_ & new_n32766_;
  assign new_n32797_ = new_n32765_ & new_n32764_;
  assign new_n32798_ = new_n32763_ & new_n32762_;
  assign new_n32799_ = new_n32761_ & new_n32760_;
  assign new_n32800_ = new_n32748_ & new_n32747_;
  assign new_n32801_ = ~new_n32994_ | ~new_n32993_;
  assign new_n32802_ = ~new_n33050_ | ~new_n33049_;
  assign new_n32803_ = ~new_n15883_;
  assign new_n32804_ = ~new_n15891_;
  assign new_n32805_ = ~new_n15890_;
  assign new_n32806_ = ~new_n15889_;
  assign new_n32807_ = ~new_n15888_;
  assign new_n32808_ = ~new_n15887_;
  assign new_n32809_ = ~new_n15886_;
  assign new_n32810_ = ~new_n15885_;
  assign new_n32811_ = ~new_n15884_;
  assign new_n32812_ = ~new_n15882_;
  assign new_n32813_ = ~new_n32863_ | ~new_n32731_;
  assign new_n32814_ = ~new_n32861_ | ~new_n32732_;
  assign new_n32815_ = ~new_n32859_ | ~new_n32734_;
  assign new_n32816_ = ~new_n32739_ | ~new_n32841_;
  assign new_n32817_ = ~new_n15863_;
  assign new_n32818_ = ~new_n15864_;
  assign new_n32819_ = ~new_n15865_;
  assign new_n32820_ = ~new_n15866_;
  assign new_n32821_ = ~new_n15867_;
  assign new_n32822_ = ~new_n15868_;
  assign new_n32823_ = ~new_n15869_;
  assign new_n32824_ = ~new_n15870_;
  assign new_n32825_ = ~new_n15871_;
  assign new_n32826_ = ~new_n15872_;
  assign new_n32827_ = ~new_n15873_;
  assign new_n32828_ = ~new_n15881_;
  assign new_n32829_ = ~new_n15880_;
  assign new_n32830_ = ~new_n15879_;
  assign new_n32831_ = ~new_n15878_;
  assign new_n32832_ = ~new_n15877_;
  assign new_n32833_ = ~new_n15876_;
  assign new_n32834_ = ~new_n15875_;
  assign new_n32835_ = ~new_n15874_;
  assign new_n32836_ = ~new_n15861_;
  assign new_n32837_ = ~new_n15862_;
  assign new_n32838_ = ~new_n15860_;
  assign new_n32839_ = ~new_n32800_ | ~new_n32884_;
  assign new_n32840_ = ~new_n32884_ | ~new_n32748_;
  assign new_n32841_ = ~new_n32856_ | ~new_n32855_;
  assign new_n32842_ = new_n33001_ & new_n33000_;
  assign new_n32843_ = new_n33023_ & new_n33022_;
  assign new_n32844_ = ~new_n32852_ | ~new_n32851_;
  assign new_n32845_ = ~new_n32871_ | ~new_n32760_;
  assign new_n32846_ = ~new_n32869_ | ~new_n32762_;
  assign new_n32847_ = ~new_n32867_ | ~new_n32764_;
  assign new_n32848_ = ~new_n32865_ | ~new_n32766_;
  assign new_n32849_ = ~new_n32839_;
  assign new_n32850_ = new_n17371_ | new_n17370_;
  assign new_n32851_ = ~new_n32736_ | ~new_n32850_;
  assign new_n32852_ = ~new_n17370_ | ~new_n17371_;
  assign new_n32853_ = ~new_n32844_;
  assign new_n32854_ = ~new_n32894_ | ~new_n32710_;
  assign new_n32855_ = ~new_n32854_ | ~new_n32844_;
  assign new_n32856_ = ~new_n15859_ | ~new_n32737_;
  assign new_n32857_ = ~new_n32841_;
  assign new_n32858_ = ~new_n32816_;
  assign new_n32859_ = ~new_n32711_;
  assign new_n32860_ = ~new_n32815_;
  assign new_n32861_ = ~new_n32712_;
  assign new_n32862_ = ~new_n32814_;
  assign new_n32863_ = ~new_n32713_;
  assign new_n32864_ = ~new_n32813_;
  assign new_n32865_ = ~new_n32714_;
  assign new_n32866_ = ~new_n32848_;
  assign new_n32867_ = ~new_n32715_;
  assign new_n32868_ = ~new_n32847_;
  assign new_n32869_ = ~new_n32716_;
  assign new_n32870_ = ~new_n32846_;
  assign new_n32871_ = ~new_n32717_;
  assign new_n32872_ = ~new_n32845_;
  assign new_n32873_ = ~new_n32718_;
  assign new_n32874_ = ~new_n32719_;
  assign new_n32875_ = ~new_n32720_;
  assign new_n32876_ = ~new_n32721_;
  assign new_n32877_ = ~new_n32722_;
  assign new_n32878_ = ~new_n32723_;
  assign new_n32879_ = ~new_n32724_;
  assign new_n32880_ = ~new_n32725_;
  assign new_n32881_ = ~new_n32726_;
  assign new_n32882_ = ~new_n32727_;
  assign new_n32883_ = ~new_n32728_;
  assign new_n32884_ = ~new_n32729_;
  assign new_n32885_ = ~new_n32840_;
  assign new_n32886_ = ~new_n17371_ | ~new_n32803_;
  assign new_n32887_ = ~new_n15883_ | ~new_n32708_;
  assign new_n32888_ = ~new_n32731_;
  assign new_n32889_ = ~new_n17371_ | ~new_n32804_;
  assign new_n32890_ = ~new_n15891_ | ~new_n32708_;
  assign new_n32891_ = ~new_n32736_;
  assign new_n32892_ = ~new_n17371_ | ~new_n32805_;
  assign new_n32893_ = ~new_n15890_ | ~new_n32708_;
  assign new_n32894_ = ~new_n32737_;
  assign new_n32895_ = ~new_n17371_ | ~new_n32806_;
  assign new_n32896_ = ~new_n15889_ | ~new_n32708_;
  assign new_n32897_ = ~new_n32739_;
  assign new_n32898_ = ~new_n17371_ | ~new_n32807_;
  assign new_n32899_ = ~new_n15888_ | ~new_n32708_;
  assign new_n32900_ = ~new_n32738_;
  assign new_n32901_ = ~new_n17371_ | ~new_n32808_;
  assign new_n32902_ = ~new_n15887_ | ~new_n32708_;
  assign new_n32903_ = ~new_n32734_;
  assign new_n32904_ = ~new_n17371_ | ~new_n32809_;
  assign new_n32905_ = ~new_n15886_ | ~new_n32708_;
  assign new_n32906_ = ~new_n32735_;
  assign new_n32907_ = ~new_n17371_ | ~new_n32810_;
  assign new_n32908_ = ~new_n15885_ | ~new_n32708_;
  assign new_n32909_ = ~new_n32732_;
  assign new_n32910_ = ~new_n17371_ | ~new_n32811_;
  assign new_n32911_ = ~new_n15884_ | ~new_n32708_;
  assign new_n32912_ = ~new_n32733_;
  assign new_n32913_ = ~new_n17371_ | ~new_n32812_;
  assign new_n32914_ = ~new_n15882_ | ~new_n32708_;
  assign new_n32915_ = ~new_n32730_;
  assign new_n32916_ = ~new_n32864_ | ~new_n32915_;
  assign new_n32917_ = ~new_n32730_ | ~new_n32813_;
  assign new_n32918_ = ~new_n32888_ | ~new_n32863_;
  assign new_n32919_ = ~new_n32731_ | ~new_n32713_;
  assign new_n32920_ = ~new_n32862_ | ~new_n32912_;
  assign new_n32921_ = ~new_n32733_ | ~new_n32814_;
  assign new_n32922_ = ~new_n32909_ | ~new_n32861_;
  assign new_n32923_ = ~new_n32732_ | ~new_n32712_;
  assign new_n32924_ = ~new_n32860_ | ~new_n32906_;
  assign new_n32925_ = ~new_n32735_ | ~new_n32815_;
  assign new_n32926_ = ~new_n32903_ | ~new_n32859_;
  assign new_n32927_ = ~new_n32734_ | ~new_n32711_;
  assign new_n32928_ = ~new_n32858_ | ~new_n32900_;
  assign new_n32929_ = ~new_n32738_ | ~new_n32816_;
  assign new_n32930_ = ~new_n17371_ | ~new_n32817_;
  assign new_n32931_ = ~new_n15863_ | ~new_n32708_;
  assign new_n32932_ = ~new_n32749_;
  assign new_n32933_ = ~new_n17371_ | ~new_n32818_;
  assign new_n32934_ = ~new_n15864_ | ~new_n32708_;
  assign new_n32935_ = ~new_n32750_;
  assign new_n32936_ = ~new_n17371_ | ~new_n32819_;
  assign new_n32937_ = ~new_n15865_ | ~new_n32708_;
  assign new_n32938_ = ~new_n32751_;
  assign new_n32939_ = ~new_n17371_ | ~new_n32820_;
  assign new_n32940_ = ~new_n15866_ | ~new_n32708_;
  assign new_n32941_ = ~new_n32752_;
  assign new_n32942_ = ~new_n17371_ | ~new_n32821_;
  assign new_n32943_ = ~new_n15867_ | ~new_n32708_;
  assign new_n32944_ = ~new_n32753_;
  assign new_n32945_ = ~new_n17371_ | ~new_n32822_;
  assign new_n32946_ = ~new_n15868_ | ~new_n32708_;
  assign new_n32947_ = ~new_n32754_;
  assign new_n32948_ = ~new_n17371_ | ~new_n32823_;
  assign new_n32949_ = ~new_n15869_ | ~new_n32708_;
  assign new_n32950_ = ~new_n32755_;
  assign new_n32951_ = ~new_n17371_ | ~new_n32824_;
  assign new_n32952_ = ~new_n15870_ | ~new_n32708_;
  assign new_n32953_ = ~new_n32756_;
  assign new_n32954_ = ~new_n17371_ | ~new_n32825_;
  assign new_n32955_ = ~new_n15871_ | ~new_n32708_;
  assign new_n32956_ = ~new_n32757_;
  assign new_n32957_ = ~new_n17371_ | ~new_n32826_;
  assign new_n32958_ = ~new_n15872_ | ~new_n32708_;
  assign new_n32959_ = ~new_n32758_;
  assign new_n32960_ = ~new_n17371_ | ~new_n32827_;
  assign new_n32961_ = ~new_n15873_ | ~new_n32708_;
  assign new_n32962_ = ~new_n32759_;
  assign new_n32963_ = ~new_n17371_ | ~new_n32828_;
  assign new_n32964_ = ~new_n15881_ | ~new_n32708_;
  assign new_n32965_ = ~new_n32766_;
  assign new_n32966_ = ~new_n17371_ | ~new_n32829_;
  assign new_n32967_ = ~new_n15880_ | ~new_n32708_;
  assign new_n32968_ = ~new_n32767_;
  assign new_n32969_ = ~new_n17371_ | ~new_n32830_;
  assign new_n32970_ = ~new_n15879_ | ~new_n32708_;
  assign new_n32971_ = ~new_n32764_;
  assign new_n32972_ = ~new_n17371_ | ~new_n32831_;
  assign new_n32973_ = ~new_n15878_ | ~new_n32708_;
  assign new_n32974_ = ~new_n32765_;
  assign new_n32975_ = ~new_n17371_ | ~new_n32832_;
  assign new_n32976_ = ~new_n15877_ | ~new_n32708_;
  assign new_n32977_ = ~new_n32762_;
  assign new_n32978_ = ~new_n17371_ | ~new_n32833_;
  assign new_n32979_ = ~new_n15876_ | ~new_n32708_;
  assign new_n32980_ = ~new_n32763_;
  assign new_n32981_ = ~new_n17371_ | ~new_n32834_;
  assign new_n32982_ = ~new_n15875_ | ~new_n32708_;
  assign new_n32983_ = ~new_n32760_;
  assign new_n32984_ = ~new_n17371_ | ~new_n32835_;
  assign new_n32985_ = ~new_n15874_ | ~new_n32708_;
  assign new_n32986_ = ~new_n32761_;
  assign new_n32987_ = ~new_n17371_ | ~new_n32836_;
  assign new_n32988_ = ~new_n15861_ | ~new_n32708_;
  assign new_n32989_ = ~new_n32747_;
  assign new_n32990_ = ~new_n17371_ | ~new_n32837_;
  assign new_n32991_ = ~new_n15862_ | ~new_n32708_;
  assign new_n32992_ = ~new_n32748_;
  assign new_n32993_ = ~new_n17371_ | ~new_n32838_;
  assign new_n32994_ = ~new_n15860_ | ~new_n32708_;
  assign new_n32995_ = ~new_n32801_;
  assign new_n32996_ = ~new_n32849_ | ~new_n32995_;
  assign new_n32997_ = ~new_n32801_ | ~new_n32839_;
  assign new_n32998_ = ~new_n32885_ | ~new_n32989_;
  assign new_n32999_ = ~new_n32747_ | ~new_n32840_;
  assign new_n33000_ = ~new_n32857_ | ~new_n32897_;
  assign new_n33001_ = ~new_n32739_ | ~new_n32841_;
  assign new_n33002_ = ~new_n32992_ | ~new_n32884_;
  assign new_n33003_ = ~new_n32748_ | ~new_n32729_;
  assign new_n33004_ = ~new_n32932_ | ~new_n32883_;
  assign new_n33005_ = ~new_n32749_ | ~new_n32728_;
  assign new_n33006_ = ~new_n32935_ | ~new_n32882_;
  assign new_n33007_ = ~new_n32750_ | ~new_n32727_;
  assign new_n33008_ = ~new_n32938_ | ~new_n32881_;
  assign new_n33009_ = ~new_n32751_ | ~new_n32726_;
  assign new_n33010_ = ~new_n32941_ | ~new_n32880_;
  assign new_n33011_ = ~new_n32752_ | ~new_n32725_;
  assign new_n33012_ = ~new_n32944_ | ~new_n32879_;
  assign new_n33013_ = ~new_n32753_ | ~new_n32724_;
  assign new_n33014_ = ~new_n32947_ | ~new_n32878_;
  assign new_n33015_ = ~new_n32754_ | ~new_n32723_;
  assign new_n33016_ = ~new_n32950_ | ~new_n32877_;
  assign new_n33017_ = ~new_n32755_ | ~new_n32722_;
  assign new_n33018_ = ~new_n32953_ | ~new_n32876_;
  assign new_n33019_ = ~new_n32756_ | ~new_n32721_;
  assign new_n33020_ = ~new_n32956_ | ~new_n32875_;
  assign new_n33021_ = ~new_n32757_ | ~new_n32720_;
  assign new_n33022_ = ~new_n32894_ | ~new_n15859_;
  assign new_n33023_ = ~new_n32737_ | ~new_n32710_;
  assign new_n33024_ = ~new_n32894_ | ~new_n15859_;
  assign new_n33025_ = ~new_n32737_ | ~new_n32710_;
  assign new_n33026_ = ~new_n33025_ | ~new_n33024_;
  assign new_n33027_ = ~new_n32843_ | ~new_n32844_;
  assign new_n33028_ = ~new_n32853_ | ~new_n33026_;
  assign new_n33029_ = ~new_n32959_ | ~new_n32874_;
  assign new_n33030_ = ~new_n32758_ | ~new_n32719_;
  assign new_n33031_ = ~new_n32962_ | ~new_n32873_;
  assign new_n33032_ = ~new_n32759_ | ~new_n32718_;
  assign new_n33033_ = ~new_n32872_ | ~new_n32986_;
  assign new_n33034_ = ~new_n32761_ | ~new_n32845_;
  assign new_n33035_ = ~new_n32983_ | ~new_n32871_;
  assign new_n33036_ = ~new_n32760_ | ~new_n32717_;
  assign new_n33037_ = ~new_n32870_ | ~new_n32980_;
  assign new_n33038_ = ~new_n32763_ | ~new_n32846_;
  assign new_n33039_ = ~new_n32977_ | ~new_n32869_;
  assign new_n33040_ = ~new_n32762_ | ~new_n32716_;
  assign new_n33041_ = ~new_n32868_ | ~new_n32974_;
  assign new_n33042_ = ~new_n32765_ | ~new_n32847_;
  assign new_n33043_ = ~new_n32971_ | ~new_n32867_;
  assign new_n33044_ = ~new_n32764_ | ~new_n32715_;
  assign new_n33045_ = ~new_n32866_ | ~new_n32968_;
  assign new_n33046_ = ~new_n32767_ | ~new_n32848_;
  assign new_n33047_ = ~new_n32965_ | ~new_n32865_;
  assign new_n33048_ = ~new_n32766_ | ~new_n32714_;
  assign new_n33049_ = ~new_n17370_ | ~new_n32708_;
  assign new_n33050_ = ~new_n17371_ | ~new_n32709_;
  assign new_n33051_ = ~new_n32802_;
  assign new_n33052_ = ~new_n32736_ | ~new_n33051_;
  assign new_n33053_ = ~new_n32802_ | ~new_n32891_;
  assign new_n33054_ = ~new_n15897_;
  assign new_n33055_ = ~new_n15895_;
  assign new_n33056_ = ~new_n15901_;
  assign new_n33057_ = ~new_n15900_;
  assign new_n33058_ = ~new_n15894_;
  assign new_n33059_ = ~new_n15893_;
  assign new_n33060_ = ~new_n15899_;
  assign new_n33061_ = ~new_n15898_;
  assign new_n33062_ = ~new_n15892_;
  assign new_n33063_ = ~new_n15537_;
  assign new_n33064_ = ~pi1076;
  assign new_n33065_ = ~new_n33098_ | ~new_n33097_;
  assign new_n33066_ = new_n33077_ & new_n33078_;
  assign new_n33067_ = new_n33080_ & new_n33081_;
  assign new_n33068_ = new_n33083_ & new_n33084_;
  assign new_n33069_ = new_n33086_ & new_n33087_;
  assign new_n33070_ = ~new_n15902_;
  assign new_n33071_ = ~new_n15903_;
  assign new_n33072_ = ~new_n15896_ | ~new_n33071_;
  assign new_n33073_ = ~new_n15896_ | ~new_n33070_;
  assign new_n33074_ = new_n15902_ | new_n15903_;
  assign new_n33075_ = ~new_n15895_ | ~new_n33056_;
  assign new_n33076_ = ~new_n33074_ | ~new_n33072_ | ~new_n33073_ | ~new_n33075_;
  assign new_n33077_ = ~new_n15901_ | ~new_n33055_;
  assign new_n33078_ = ~new_n15900_ | ~new_n33058_;
  assign new_n33079_ = ~new_n33066_ | ~new_n33076_;
  assign new_n33080_ = ~new_n15894_ | ~new_n33057_;
  assign new_n33081_ = ~new_n15893_ | ~new_n33060_;
  assign new_n33082_ = ~new_n33067_ | ~new_n33079_;
  assign new_n33083_ = ~new_n15899_ | ~new_n33059_;
  assign new_n33084_ = ~new_n15898_ | ~new_n33062_;
  assign new_n33085_ = ~new_n33068_ | ~new_n33082_;
  assign new_n33086_ = ~new_n15892_ | ~new_n33061_;
  assign new_n33087_ = ~new_n15537_ | ~new_n33054_;
  assign new_n33088_ = ~new_n33069_ | ~new_n33085_;
  assign new_n33089_ = ~new_n15897_ | ~new_n33063_;
  assign new_n33090_ = ~new_n33088_ | ~new_n33089_;
  assign new_n33091_ = ~new_n15897_ | ~new_n33064_;
  assign new_n33092_ = ~new_n33090_ | ~new_n33054_;
  assign new_n33093_ = ~new_n33092_ | ~new_n33091_;
  assign new_n33094_ = ~pi1076 | ~new_n33054_;
  assign new_n33095_ = ~new_n15897_ | ~new_n33090_;
  assign new_n33096_ = ~new_n33095_ | ~new_n33094_;
  assign new_n33097_ = ~new_n33093_ | ~new_n33063_;
  assign new_n33098_ = ~new_n15537_ | ~new_n33096_;
  assign new_n33099_ = ~pi1248;
  assign new_n33100_ = ~pi1249;
  assign new_n33101_ = ~pi1249 | ~pi1248;
  assign new_n33102_ = ~pi1250;
  assign new_n33103_ = ~pi1250 | ~new_n33189_;
  assign new_n33104_ = ~pi1251;
  assign new_n33105_ = ~pi1251 | ~new_n33190_;
  assign new_n33106_ = ~pi1252;
  assign new_n33107_ = ~pi1252 | ~new_n33191_;
  assign new_n33108_ = ~pi1253;
  assign new_n33109_ = ~pi1253 | ~new_n33192_;
  assign new_n33110_ = ~pi1254;
  assign new_n33111_ = ~pi1254 | ~new_n33193_;
  assign new_n33112_ = ~pi1255;
  assign new_n33113_ = ~pi1256;
  assign new_n33114_ = ~pi1255 | ~new_n33194_;
  assign new_n33115_ = ~new_n33195_ | ~pi1256;
  assign new_n33116_ = ~pi1257;
  assign new_n33117_ = ~pi1257 | ~new_n33196_;
  assign new_n33118_ = ~pi1258;
  assign new_n33119_ = ~pi1258 | ~new_n33197_;
  assign new_n33120_ = ~pi1259;
  assign new_n33121_ = ~pi1259 | ~new_n33198_;
  assign new_n33122_ = ~pi1260;
  assign new_n33123_ = ~pi1260 | ~new_n33199_;
  assign new_n33124_ = ~pi1261;
  assign new_n33125_ = ~pi1261 | ~new_n33200_;
  assign new_n33126_ = ~pi1262;
  assign new_n33127_ = ~pi1262 | ~new_n33201_;
  assign new_n33128_ = ~pi1263;
  assign new_n33129_ = ~pi1263 | ~new_n33202_;
  assign new_n33130_ = ~pi1264;
  assign new_n33131_ = ~pi1264 | ~new_n33203_;
  assign new_n33132_ = ~pi1265;
  assign new_n33133_ = ~pi1265 | ~new_n33204_;
  assign new_n33134_ = ~pi1266;
  assign new_n33135_ = ~pi1266 | ~new_n33205_;
  assign new_n33136_ = ~pi1267;
  assign new_n33137_ = ~pi1267 | ~new_n33206_;
  assign new_n33138_ = ~pi1268;
  assign new_n33139_ = ~pi1268 | ~new_n33207_;
  assign new_n33140_ = ~pi1269;
  assign new_n33141_ = ~pi1269 | ~new_n33208_;
  assign new_n33142_ = ~pi1270;
  assign new_n33143_ = ~pi1270 | ~new_n33209_;
  assign new_n33144_ = ~pi1271;
  assign new_n33145_ = ~pi1271 | ~new_n33210_;
  assign new_n33146_ = ~pi1272;
  assign new_n33147_ = ~pi1272 | ~new_n33211_;
  assign new_n33148_ = ~pi1273;
  assign new_n33149_ = ~pi1273 | ~new_n33212_;
  assign new_n33150_ = ~pi1274;
  assign new_n33151_ = ~pi1274 | ~new_n33213_;
  assign new_n33152_ = ~pi1275;
  assign new_n33153_ = ~pi1275 | ~new_n33214_;
  assign new_n33154_ = ~pi1276;
  assign new_n33155_ = ~pi1276 | ~new_n33215_;
  assign new_n33156_ = ~pi1277;
  assign new_n33157_ = ~new_n33219_ | ~new_n33218_;
  assign new_n33158_ = ~new_n33221_ | ~new_n33220_;
  assign new_n33159_ = ~new_n33223_ | ~new_n33222_;
  assign new_n33160_ = ~new_n33225_ | ~new_n33224_;
  assign new_n33161_ = ~new_n33227_ | ~new_n33226_;
  assign new_n33162_ = ~new_n33229_ | ~new_n33228_;
  assign new_n33163_ = ~new_n33231_ | ~new_n33230_;
  assign new_n33164_ = ~new_n33233_ | ~new_n33232_;
  assign new_n33165_ = ~new_n33235_ | ~new_n33234_;
  assign new_n33166_ = ~new_n33237_ | ~new_n33236_;
  assign new_n33167_ = ~new_n33239_ | ~new_n33238_;
  assign new_n33168_ = ~new_n33241_ | ~new_n33240_;
  assign new_n33169_ = ~new_n33243_ | ~new_n33242_;
  assign new_n33170_ = ~new_n33245_ | ~new_n33244_;
  assign new_n33171_ = ~new_n33247_ | ~new_n33246_;
  assign new_n33172_ = ~new_n33249_ | ~new_n33248_;
  assign new_n33173_ = ~new_n33251_ | ~new_n33250_;
  assign new_n33174_ = ~new_n33253_ | ~new_n33252_;
  assign new_n33175_ = ~new_n33255_ | ~new_n33254_;
  assign new_n33176_ = ~new_n33257_ | ~new_n33256_;
  assign new_n33177_ = ~new_n33259_ | ~new_n33258_;
  assign new_n33178_ = ~new_n33261_ | ~new_n33260_;
  assign new_n33179_ = ~new_n33263_ | ~new_n33262_;
  assign new_n33180_ = ~new_n33265_ | ~new_n33264_;
  assign new_n33181_ = ~new_n33267_ | ~new_n33266_;
  assign new_n33182_ = ~new_n33269_ | ~new_n33268_;
  assign new_n33183_ = ~new_n33271_ | ~new_n33270_;
  assign new_n33184_ = ~new_n33273_ | ~new_n33272_;
  assign new_n33185_ = ~new_n33275_ | ~new_n33274_;
  assign new_n33186_ = ~new_n33277_ | ~new_n33276_;
  assign new_n33187_ = ~pi1278;
  assign new_n33188_ = ~pi1277 | ~new_n33216_;
  assign new_n33189_ = ~new_n33101_;
  assign new_n33190_ = ~new_n33103_;
  assign new_n33191_ = ~new_n33105_;
  assign new_n33192_ = ~new_n33107_;
  assign new_n33193_ = ~new_n33109_;
  assign new_n33194_ = ~new_n33111_;
  assign new_n33195_ = ~new_n33114_;
  assign new_n33196_ = ~new_n33115_;
  assign new_n33197_ = ~new_n33117_;
  assign new_n33198_ = ~new_n33119_;
  assign new_n33199_ = ~new_n33121_;
  assign new_n33200_ = ~new_n33123_;
  assign new_n33201_ = ~new_n33125_;
  assign new_n33202_ = ~new_n33127_;
  assign new_n33203_ = ~new_n33129_;
  assign new_n33204_ = ~new_n33131_;
  assign new_n33205_ = ~new_n33133_;
  assign new_n33206_ = ~new_n33135_;
  assign new_n33207_ = ~new_n33137_;
  assign new_n33208_ = ~new_n33139_;
  assign new_n33209_ = ~new_n33141_;
  assign new_n33210_ = ~new_n33143_;
  assign new_n33211_ = ~new_n33145_;
  assign new_n33212_ = ~new_n33147_;
  assign new_n33213_ = ~new_n33149_;
  assign new_n33214_ = ~new_n33151_;
  assign new_n33215_ = ~new_n33153_;
  assign new_n33216_ = ~new_n33155_;
  assign new_n33217_ = ~new_n33188_;
  assign new_n33218_ = ~pi1256 | ~new_n33114_;
  assign new_n33219_ = ~new_n33195_ | ~new_n33113_;
  assign new_n33220_ = ~pi1255 | ~new_n33111_;
  assign new_n33221_ = ~new_n33194_ | ~new_n33112_;
  assign new_n33222_ = ~pi1254 | ~new_n33109_;
  assign new_n33223_ = ~new_n33193_ | ~new_n33110_;
  assign new_n33224_ = ~pi1253 | ~new_n33107_;
  assign new_n33225_ = ~new_n33192_ | ~new_n33108_;
  assign new_n33226_ = ~pi1252 | ~new_n33105_;
  assign new_n33227_ = ~new_n33191_ | ~new_n33106_;
  assign new_n33228_ = ~pi1251 | ~new_n33103_;
  assign new_n33229_ = ~new_n33190_ | ~new_n33104_;
  assign new_n33230_ = ~pi1250 | ~new_n33101_;
  assign new_n33231_ = ~new_n33189_ | ~new_n33102_;
  assign new_n33232_ = ~pi1278 | ~new_n33188_;
  assign new_n33233_ = ~new_n33217_ | ~new_n33187_;
  assign new_n33234_ = ~pi1277 | ~new_n33155_;
  assign new_n33235_ = ~new_n33216_ | ~new_n33156_;
  assign new_n33236_ = ~pi1249 | ~new_n33099_;
  assign new_n33237_ = ~pi1248 | ~new_n33100_;
  assign new_n33238_ = ~pi1276 | ~new_n33153_;
  assign new_n33239_ = ~new_n33215_ | ~new_n33154_;
  assign new_n33240_ = ~pi1275 | ~new_n33151_;
  assign new_n33241_ = ~new_n33214_ | ~new_n33152_;
  assign new_n33242_ = ~pi1274 | ~new_n33149_;
  assign new_n33243_ = ~new_n33213_ | ~new_n33150_;
  assign new_n33244_ = ~pi1273 | ~new_n33147_;
  assign new_n33245_ = ~new_n33212_ | ~new_n33148_;
  assign new_n33246_ = ~pi1272 | ~new_n33145_;
  assign new_n33247_ = ~new_n33211_ | ~new_n33146_;
  assign new_n33248_ = ~pi1271 | ~new_n33143_;
  assign new_n33249_ = ~new_n33210_ | ~new_n33144_;
  assign new_n33250_ = ~pi1270 | ~new_n33141_;
  assign new_n33251_ = ~new_n33209_ | ~new_n33142_;
  assign new_n33252_ = ~pi1269 | ~new_n33139_;
  assign new_n33253_ = ~new_n33208_ | ~new_n33140_;
  assign new_n33254_ = ~pi1268 | ~new_n33137_;
  assign new_n33255_ = ~new_n33207_ | ~new_n33138_;
  assign new_n33256_ = ~pi1267 | ~new_n33135_;
  assign new_n33257_ = ~new_n33206_ | ~new_n33136_;
  assign new_n33258_ = ~pi1266 | ~new_n33133_;
  assign new_n33259_ = ~new_n33205_ | ~new_n33134_;
  assign new_n33260_ = ~pi1265 | ~new_n33131_;
  assign new_n33261_ = ~new_n33204_ | ~new_n33132_;
  assign new_n33262_ = ~pi1264 | ~new_n33129_;
  assign new_n33263_ = ~new_n33203_ | ~new_n33130_;
  assign new_n33264_ = ~pi1263 | ~new_n33127_;
  assign new_n33265_ = ~new_n33202_ | ~new_n33128_;
  assign new_n33266_ = ~pi1262 | ~new_n33125_;
  assign new_n33267_ = ~new_n33201_ | ~new_n33126_;
  assign new_n33268_ = ~pi1261 | ~new_n33123_;
  assign new_n33269_ = ~new_n33200_ | ~new_n33124_;
  assign new_n33270_ = ~pi1260 | ~new_n33121_;
  assign new_n33271_ = ~new_n33199_ | ~new_n33122_;
  assign new_n33272_ = ~pi1259 | ~new_n33119_;
  assign new_n33273_ = ~new_n33198_ | ~new_n33120_;
  assign new_n33274_ = ~pi1258 | ~new_n33117_;
  assign new_n33275_ = ~new_n33197_ | ~new_n33118_;
  assign new_n33276_ = ~pi1257 | ~new_n33115_;
  assign new_n33277_ = ~new_n33196_ | ~new_n33116_;
  assign new_n33278_ = ~new_n16414_;
  assign new_n33279_ = ~new_n16409_;
  assign new_n33280_ = ~new_n16415_;
  assign new_n33281_ = ~new_n16413_;
  assign new_n33282_ = ~new_n16408_;
  assign new_n33283_ = ~new_n16411_;
  assign new_n33284_ = ~new_n16410_;
  assign new_n33285_ = ~new_n16412_;
  assign new_n33286_ = new_n33289_ & new_n33288_;
  assign new_n33287_ = ~new_n15854_;
  assign new_n33288_ = ~new_n32706_ | ~new_n33287_;
  assign new_n33289_ = ~new_n32707_ | ~new_n33287_;
  assign new_n33290_ = ~new_n33294_ | ~new_n33293_;
  assign new_n33291_ = ~pi1216;
  assign new_n33292_ = ~pi1215;
  assign new_n33293_ = ~pi1216 | ~new_n33292_;
  assign new_n33294_ = ~pi1215 | ~new_n33291_;
  assign new_n33295_ = ~pi1407;
  assign new_n33296_ = ~pi1408;
  assign new_n33297_ = ~pi1408 | ~pi1407;
  assign new_n33298_ = ~pi1409;
  assign new_n33299_ = ~pi1409 | ~new_n33385_;
  assign new_n33300_ = ~pi1410;
  assign new_n33301_ = ~pi1410 | ~new_n33386_;
  assign new_n33302_ = ~pi1411;
  assign new_n33303_ = ~pi1411 | ~new_n33387_;
  assign new_n33304_ = ~pi1412;
  assign new_n33305_ = ~pi1412 | ~new_n33388_;
  assign new_n33306_ = ~pi1413;
  assign new_n33307_ = ~pi1413 | ~new_n33389_;
  assign new_n33308_ = ~pi1414;
  assign new_n33309_ = ~pi1415;
  assign new_n33310_ = ~pi1414 | ~new_n33390_;
  assign new_n33311_ = ~new_n33391_ | ~pi1415;
  assign new_n33312_ = ~pi1416;
  assign new_n33313_ = ~pi1416 | ~new_n33392_;
  assign new_n33314_ = ~pi1417;
  assign new_n33315_ = ~pi1417 | ~new_n33393_;
  assign new_n33316_ = ~pi1418;
  assign new_n33317_ = ~pi1418 | ~new_n33394_;
  assign new_n33318_ = ~pi1419;
  assign new_n33319_ = ~pi1419 | ~new_n33395_;
  assign new_n33320_ = ~pi1420;
  assign new_n33321_ = ~pi1420 | ~new_n33396_;
  assign new_n33322_ = ~pi1421;
  assign new_n33323_ = ~pi1421 | ~new_n33397_;
  assign new_n33324_ = ~pi1422;
  assign new_n33325_ = ~pi1422 | ~new_n33398_;
  assign new_n33326_ = ~pi1423;
  assign new_n33327_ = ~pi1423 | ~new_n33399_;
  assign new_n33328_ = ~pi1424;
  assign new_n33329_ = ~pi1424 | ~new_n33400_;
  assign new_n33330_ = ~pi1425;
  assign new_n33331_ = ~pi1425 | ~new_n33401_;
  assign new_n33332_ = ~pi1426;
  assign new_n33333_ = ~pi1426 | ~new_n33402_;
  assign new_n33334_ = ~pi1427;
  assign new_n33335_ = ~pi1427 | ~new_n33403_;
  assign new_n33336_ = ~pi1428;
  assign new_n33337_ = ~pi1428 | ~new_n33404_;
  assign new_n33338_ = ~pi1429;
  assign new_n33339_ = ~pi1429 | ~new_n33405_;
  assign new_n33340_ = ~pi1430;
  assign new_n33341_ = ~pi1430 | ~new_n33406_;
  assign new_n33342_ = ~pi1431;
  assign new_n33343_ = ~pi1431 | ~new_n33407_;
  assign new_n33344_ = ~pi1432;
  assign new_n33345_ = ~pi1432 | ~new_n33408_;
  assign new_n33346_ = ~pi1433;
  assign new_n33347_ = ~pi1433 | ~new_n33409_;
  assign new_n33348_ = ~pi1434;
  assign new_n33349_ = ~pi1434 | ~new_n33410_;
  assign new_n33350_ = ~pi1435;
  assign new_n33351_ = ~pi1435 | ~new_n33411_;
  assign new_n33352_ = ~pi1436;
  assign new_n33353_ = ~new_n33415_ | ~new_n33414_;
  assign new_n33354_ = ~new_n33417_ | ~new_n33416_;
  assign new_n33355_ = ~new_n33419_ | ~new_n33418_;
  assign new_n33356_ = ~new_n33421_ | ~new_n33420_;
  assign new_n33357_ = ~new_n33423_ | ~new_n33422_;
  assign new_n33358_ = ~new_n33425_ | ~new_n33424_;
  assign new_n33359_ = ~new_n33427_ | ~new_n33426_;
  assign new_n33360_ = ~new_n33429_ | ~new_n33428_;
  assign new_n33361_ = ~new_n33431_ | ~new_n33430_;
  assign new_n33362_ = ~new_n33433_ | ~new_n33432_;
  assign new_n33363_ = ~new_n33435_ | ~new_n33434_;
  assign new_n33364_ = ~new_n33437_ | ~new_n33436_;
  assign new_n33365_ = ~new_n33439_ | ~new_n33438_;
  assign new_n33366_ = ~new_n33441_ | ~new_n33440_;
  assign new_n33367_ = ~new_n33443_ | ~new_n33442_;
  assign new_n33368_ = ~new_n33445_ | ~new_n33444_;
  assign new_n33369_ = ~new_n33447_ | ~new_n33446_;
  assign new_n33370_ = ~new_n33449_ | ~new_n33448_;
  assign new_n33371_ = ~new_n33451_ | ~new_n33450_;
  assign new_n33372_ = ~new_n33453_ | ~new_n33452_;
  assign new_n33373_ = ~new_n33455_ | ~new_n33454_;
  assign new_n33374_ = ~new_n33457_ | ~new_n33456_;
  assign new_n33375_ = ~new_n33459_ | ~new_n33458_;
  assign new_n33376_ = ~new_n33461_ | ~new_n33460_;
  assign new_n33377_ = ~new_n33463_ | ~new_n33462_;
  assign new_n33378_ = ~new_n33465_ | ~new_n33464_;
  assign new_n33379_ = ~new_n33467_ | ~new_n33466_;
  assign new_n33380_ = ~new_n33469_ | ~new_n33468_;
  assign new_n33381_ = ~new_n33471_ | ~new_n33470_;
  assign new_n33382_ = ~new_n33473_ | ~new_n33472_;
  assign new_n33383_ = ~pi1437;
  assign new_n33384_ = ~pi1436 | ~new_n33412_;
  assign new_n33385_ = ~new_n33297_;
  assign new_n33386_ = ~new_n33299_;
  assign new_n33387_ = ~new_n33301_;
  assign new_n33388_ = ~new_n33303_;
  assign new_n33389_ = ~new_n33305_;
  assign new_n33390_ = ~new_n33307_;
  assign new_n33391_ = ~new_n33310_;
  assign new_n33392_ = ~new_n33311_;
  assign new_n33393_ = ~new_n33313_;
  assign new_n33394_ = ~new_n33315_;
  assign new_n33395_ = ~new_n33317_;
  assign new_n33396_ = ~new_n33319_;
  assign new_n33397_ = ~new_n33321_;
  assign new_n33398_ = ~new_n33323_;
  assign new_n33399_ = ~new_n33325_;
  assign new_n33400_ = ~new_n33327_;
  assign new_n33401_ = ~new_n33329_;
  assign new_n33402_ = ~new_n33331_;
  assign new_n33403_ = ~new_n33333_;
  assign new_n33404_ = ~new_n33335_;
  assign new_n33405_ = ~new_n33337_;
  assign new_n33406_ = ~new_n33339_;
  assign new_n33407_ = ~new_n33341_;
  assign new_n33408_ = ~new_n33343_;
  assign new_n33409_ = ~new_n33345_;
  assign new_n33410_ = ~new_n33347_;
  assign new_n33411_ = ~new_n33349_;
  assign new_n33412_ = ~new_n33351_;
  assign new_n33413_ = ~new_n33384_;
  assign new_n33414_ = ~pi1415 | ~new_n33310_;
  assign new_n33415_ = ~new_n33391_ | ~new_n33309_;
  assign new_n33416_ = ~pi1414 | ~new_n33307_;
  assign new_n33417_ = ~new_n33390_ | ~new_n33308_;
  assign new_n33418_ = ~pi1413 | ~new_n33305_;
  assign new_n33419_ = ~new_n33389_ | ~new_n33306_;
  assign new_n33420_ = ~pi1412 | ~new_n33303_;
  assign new_n33421_ = ~new_n33388_ | ~new_n33304_;
  assign new_n33422_ = ~pi1411 | ~new_n33301_;
  assign new_n33423_ = ~new_n33387_ | ~new_n33302_;
  assign new_n33424_ = ~pi1410 | ~new_n33299_;
  assign new_n33425_ = ~new_n33386_ | ~new_n33300_;
  assign new_n33426_ = ~pi1409 | ~new_n33297_;
  assign new_n33427_ = ~new_n33385_ | ~new_n33298_;
  assign new_n33428_ = ~pi1437 | ~new_n33384_;
  assign new_n33429_ = ~new_n33413_ | ~new_n33383_;
  assign new_n33430_ = ~pi1436 | ~new_n33351_;
  assign new_n33431_ = ~new_n33412_ | ~new_n33352_;
  assign new_n33432_ = ~pi1408 | ~new_n33295_;
  assign new_n33433_ = ~pi1407 | ~new_n33296_;
  assign new_n33434_ = ~pi1435 | ~new_n33349_;
  assign new_n33435_ = ~new_n33411_ | ~new_n33350_;
  assign new_n33436_ = ~pi1434 | ~new_n33347_;
  assign new_n33437_ = ~new_n33410_ | ~new_n33348_;
  assign new_n33438_ = ~pi1433 | ~new_n33345_;
  assign new_n33439_ = ~new_n33409_ | ~new_n33346_;
  assign new_n33440_ = ~pi1432 | ~new_n33343_;
  assign new_n33441_ = ~new_n33408_ | ~new_n33344_;
  assign new_n33442_ = ~pi1431 | ~new_n33341_;
  assign new_n33443_ = ~new_n33407_ | ~new_n33342_;
  assign new_n33444_ = ~pi1430 | ~new_n33339_;
  assign new_n33445_ = ~new_n33406_ | ~new_n33340_;
  assign new_n33446_ = ~pi1429 | ~new_n33337_;
  assign new_n33447_ = ~new_n33405_ | ~new_n33338_;
  assign new_n33448_ = ~pi1428 | ~new_n33335_;
  assign new_n33449_ = ~new_n33404_ | ~new_n33336_;
  assign new_n33450_ = ~pi1427 | ~new_n33333_;
  assign new_n33451_ = ~new_n33403_ | ~new_n33334_;
  assign new_n33452_ = ~pi1426 | ~new_n33331_;
  assign new_n33453_ = ~new_n33402_ | ~new_n33332_;
  assign new_n33454_ = ~pi1425 | ~new_n33329_;
  assign new_n33455_ = ~new_n33401_ | ~new_n33330_;
  assign new_n33456_ = ~pi1424 | ~new_n33327_;
  assign new_n33457_ = ~new_n33400_ | ~new_n33328_;
  assign new_n33458_ = ~pi1423 | ~new_n33325_;
  assign new_n33459_ = ~new_n33399_ | ~new_n33326_;
  assign new_n33460_ = ~pi1422 | ~new_n33323_;
  assign new_n33461_ = ~new_n33398_ | ~new_n33324_;
  assign new_n33462_ = ~pi1421 | ~new_n33321_;
  assign new_n33463_ = ~new_n33397_ | ~new_n33322_;
  assign new_n33464_ = ~pi1420 | ~new_n33319_;
  assign new_n33465_ = ~new_n33396_ | ~new_n33320_;
  assign new_n33466_ = ~pi1419 | ~new_n33317_;
  assign new_n33467_ = ~new_n33395_ | ~new_n33318_;
  assign new_n33468_ = ~pi1418 | ~new_n33315_;
  assign new_n33469_ = ~new_n33394_ | ~new_n33316_;
  assign new_n33470_ = ~pi1417 | ~new_n33313_;
  assign new_n33471_ = ~new_n33393_ | ~new_n33314_;
  assign new_n33472_ = ~pi1416 | ~new_n33311_;
  assign new_n33473_ = ~new_n33392_ | ~new_n33312_;
  assign new_n33474_ = new_n33495_ & new_n33494_;
  assign new_n33475_ = ~pi1212;
  assign new_n33476_ = ~new_n16672_;
  assign new_n33477_ = ~new_n16671_;
  assign new_n33478_ = ~pi1211;
  assign new_n33479_ = ~pi1210;
  assign new_n33480_ = ~new_n16670_;
  assign new_n33481_ = new_n33489_ & new_n33490_;
  assign new_n33482_ = new_n33492_ & new_n33493_;
  assign new_n33483_ = ~new_n16673_;
  assign new_n33484_ = ~new_n16674_;
  assign new_n33485_ = ~pi1214 | ~new_n33484_ | ~new_n33483_;
  assign new_n33486_ = ~pi1213 | ~new_n33483_;
  assign new_n33487_ = ~pi1212 | ~new_n33476_;
  assign new_n33488_ = ~new_n33487_ | ~new_n33485_ | ~new_n33486_ | ~new_n33496_;
  assign new_n33489_ = ~new_n16672_ | ~new_n33475_;
  assign new_n33490_ = ~new_n16671_ | ~new_n33478_;
  assign new_n33491_ = ~new_n33481_ | ~new_n33488_;
  assign new_n33492_ = ~pi1211 | ~new_n33477_;
  assign new_n33493_ = ~pi1210 | ~new_n33480_;
  assign new_n33494_ = ~new_n33482_ | ~new_n33491_;
  assign new_n33495_ = ~new_n16670_ | ~new_n33479_;
  assign new_n33496_ = ~new_n33484_ | ~pi1214 | ~pi1213;
  assign new_n33497_ = ~new_n33536_ | ~new_n33535_;
  assign new_n33498_ = ~new_n33500_ | ~new_n33537_;
  assign new_n33499_ = ~pi1209;
  assign new_n33500_ = ~pi1209 | ~new_n33509_;
  assign new_n33501_ = ~pi1213;
  assign new_n33502_ = ~pi1207;
  assign new_n33503_ = ~pi1212;
  assign new_n33504_ = ~pi1206;
  assign new_n33505_ = ~pi1211;
  assign new_n33506_ = ~pi1210;
  assign new_n33507_ = ~new_n33532_ | ~new_n33531_;
  assign new_n33508_ = ~pi1205;
  assign new_n33509_ = ~pi1214;
  assign new_n33510_ = ~new_n33542_ | ~new_n33541_;
  assign new_n33511_ = ~new_n33547_ | ~new_n33546_;
  assign new_n33512_ = ~new_n33552_ | ~new_n33551_;
  assign new_n33513_ = ~new_n33557_ | ~new_n33556_;
  assign new_n33514_ = ~new_n33539_ | ~new_n33538_;
  assign new_n33515_ = ~new_n33544_ | ~new_n33543_;
  assign new_n33516_ = ~new_n33549_ | ~new_n33548_;
  assign new_n33517_ = ~new_n33554_ | ~new_n33553_;
  assign new_n33518_ = ~new_n33528_ | ~new_n33527_;
  assign new_n33519_ = ~new_n33524_ | ~new_n33523_;
  assign new_n33520_ = ~pi1208;
  assign new_n33521_ = ~new_n33500_;
  assign new_n33522_ = ~new_n33521_ | ~new_n33501_;
  assign new_n33523_ = ~new_n33522_ | ~new_n33520_;
  assign new_n33524_ = ~pi1213 | ~new_n33500_;
  assign new_n33525_ = ~new_n33519_;
  assign new_n33526_ = ~pi1207 | ~new_n33503_;
  assign new_n33527_ = ~new_n33526_ | ~new_n33519_;
  assign new_n33528_ = ~pi1212 | ~new_n33502_;
  assign new_n33529_ = ~new_n33518_;
  assign new_n33530_ = ~pi1206 | ~new_n33505_;
  assign new_n33531_ = ~new_n33530_ | ~new_n33518_;
  assign new_n33532_ = ~pi1211 | ~new_n33504_;
  assign new_n33533_ = ~new_n33507_;
  assign new_n33534_ = ~pi1210 | ~new_n33508_;
  assign new_n33535_ = ~new_n33533_ | ~new_n33534_;
  assign new_n33536_ = ~pi1205 | ~new_n33506_;
  assign new_n33537_ = ~pi1214 | ~new_n33499_;
  assign new_n33538_ = ~pi1205 | ~new_n33506_;
  assign new_n33539_ = ~pi1210 | ~new_n33508_;
  assign new_n33540_ = ~new_n33514_;
  assign new_n33541_ = ~new_n33540_ | ~new_n33533_;
  assign new_n33542_ = ~new_n33514_ | ~new_n33507_;
  assign new_n33543_ = ~pi1206 | ~new_n33505_;
  assign new_n33544_ = ~pi1211 | ~new_n33504_;
  assign new_n33545_ = ~new_n33515_;
  assign new_n33546_ = ~new_n33529_ | ~new_n33545_;
  assign new_n33547_ = ~new_n33515_ | ~new_n33518_;
  assign new_n33548_ = ~pi1207 | ~new_n33503_;
  assign new_n33549_ = ~pi1212 | ~new_n33502_;
  assign new_n33550_ = ~new_n33516_;
  assign new_n33551_ = ~new_n33525_ | ~new_n33550_;
  assign new_n33552_ = ~new_n33516_ | ~new_n33519_;
  assign new_n33553_ = ~pi1208 | ~new_n33501_;
  assign new_n33554_ = ~pi1213 | ~new_n33520_;
  assign new_n33555_ = ~new_n33517_;
  assign new_n33556_ = ~new_n33555_ | ~new_n33521_;
  assign new_n33557_ = ~new_n33517_ | ~new_n33500_;
  assign new_n33558_ = ~new_n33597_ | ~new_n33596_;
  assign new_n33559_ = ~new_n33561_ | ~new_n33598_;
  assign new_n33560_ = ~pi1209;
  assign new_n33561_ = ~pi1209 | ~new_n33570_;
  assign new_n33562_ = ~pi1213;
  assign new_n33563_ = ~pi1207;
  assign new_n33564_ = ~pi1212;
  assign new_n33565_ = ~pi1206;
  assign new_n33566_ = ~pi1211;
  assign new_n33567_ = ~pi1210;
  assign new_n33568_ = ~new_n33593_ | ~new_n33592_;
  assign new_n33569_ = ~pi1205;
  assign new_n33570_ = ~pi1214;
  assign new_n33571_ = ~new_n33603_ | ~new_n33602_;
  assign new_n33572_ = ~new_n33608_ | ~new_n33607_;
  assign new_n33573_ = ~new_n33613_ | ~new_n33612_;
  assign new_n33574_ = ~new_n33618_ | ~new_n33617_;
  assign new_n33575_ = ~new_n33600_ | ~new_n33599_;
  assign new_n33576_ = ~new_n33605_ | ~new_n33604_;
  assign new_n33577_ = ~new_n33610_ | ~new_n33609_;
  assign new_n33578_ = ~new_n33615_ | ~new_n33614_;
  assign new_n33579_ = ~new_n33589_ | ~new_n33588_;
  assign new_n33580_ = ~new_n33585_ | ~new_n33584_;
  assign new_n33581_ = ~pi1208;
  assign new_n33582_ = ~new_n33561_;
  assign new_n33583_ = ~new_n33582_ | ~new_n33562_;
  assign new_n33584_ = ~new_n33583_ | ~new_n33581_;
  assign new_n33585_ = ~pi1213 | ~new_n33561_;
  assign new_n33586_ = ~new_n33580_;
  assign new_n33587_ = ~pi1207 | ~new_n33564_;
  assign new_n33588_ = ~new_n33587_ | ~new_n33580_;
  assign new_n33589_ = ~pi1212 | ~new_n33563_;
  assign new_n33590_ = ~new_n33579_;
  assign new_n33591_ = ~pi1206 | ~new_n33566_;
  assign new_n33592_ = ~new_n33591_ | ~new_n33579_;
  assign new_n33593_ = ~pi1211 | ~new_n33565_;
  assign new_n33594_ = ~new_n33568_;
  assign new_n33595_ = ~pi1210 | ~new_n33569_;
  assign new_n33596_ = ~new_n33594_ | ~new_n33595_;
  assign new_n33597_ = ~pi1205 | ~new_n33567_;
  assign new_n33598_ = ~pi1214 | ~new_n33560_;
  assign new_n33599_ = ~pi1205 | ~new_n33567_;
  assign new_n33600_ = ~pi1210 | ~new_n33569_;
  assign new_n33601_ = ~new_n33575_;
  assign new_n33602_ = ~new_n33601_ | ~new_n33594_;
  assign new_n33603_ = ~new_n33575_ | ~new_n33568_;
  assign new_n33604_ = ~pi1206 | ~new_n33566_;
  assign new_n33605_ = ~pi1211 | ~new_n33565_;
  assign new_n33606_ = ~new_n33576_;
  assign new_n33607_ = ~new_n33590_ | ~new_n33606_;
  assign new_n33608_ = ~new_n33576_ | ~new_n33579_;
  assign new_n33609_ = ~pi1207 | ~new_n33564_;
  assign new_n33610_ = ~pi1212 | ~new_n33563_;
  assign new_n33611_ = ~new_n33577_;
  assign new_n33612_ = ~new_n33586_ | ~new_n33611_;
  assign new_n33613_ = ~new_n33577_ | ~new_n33580_;
  assign new_n33614_ = ~pi1208 | ~new_n33562_;
  assign new_n33615_ = ~pi1213 | ~new_n33581_;
  assign new_n33616_ = ~new_n33578_;
  assign new_n33617_ = ~new_n33616_ | ~new_n33582_;
  assign new_n33618_ = ~new_n33578_ | ~new_n33561_;
  assign new_n33619_ = ~new_n16408_;
  assign new_n33620_ = ~new_n33638_ | ~new_n33646_;
  assign new_n33621_ = new_n33637_ & new_n33645_;
  assign new_n33622_ = ~new_n16409_;
  assign new_n33623_ = ~new_n16411_;
  assign new_n33624_ = ~new_n16411_ | ~new_n33638_;
  assign new_n33625_ = ~new_n16412_;
  assign new_n33626_ = ~new_n16412_ | ~new_n33643_;
  assign new_n33627_ = ~new_n16413_;
  assign new_n33628_ = ~new_n16414_;
  assign new_n33629_ = ~new_n16413_ | ~new_n33644_;
  assign new_n33630_ = ~new_n16410_;
  assign new_n33631_ = ~new_n16415_;
  assign new_n33632_ = ~new_n33649_ | ~new_n33648_;
  assign new_n33633_ = ~new_n33651_ | ~new_n33650_;
  assign new_n33634_ = ~new_n33653_ | ~new_n33652_;
  assign new_n33635_ = ~new_n33657_ | ~new_n33656_;
  assign new_n33636_ = ~new_n33659_ | ~new_n33658_;
  assign new_n33637_ = new_n16415_ & new_n16414_;
  assign new_n33638_ = ~new_n33630_ | ~new_n33641_;
  assign new_n33639_ = new_n33655_ & new_n33654_;
  assign new_n33640_ = ~new_n33645_ | ~new_n16414_;
  assign new_n33641_ = ~new_n16409_ | ~new_n16408_;
  assign new_n33642_ = ~new_n33638_;
  assign new_n33643_ = ~new_n33624_;
  assign new_n33644_ = ~new_n33626_;
  assign new_n33645_ = ~new_n33629_;
  assign new_n33646_ = ~new_n16410_ | ~new_n16409_ | ~new_n16408_;
  assign new_n33647_ = ~new_n33640_;
  assign new_n33648_ = ~new_n16414_ | ~new_n33629_;
  assign new_n33649_ = ~new_n33645_ | ~new_n33628_;
  assign new_n33650_ = ~new_n16412_ | ~new_n33624_;
  assign new_n33651_ = ~new_n33643_ | ~new_n33625_;
  assign new_n33652_ = ~new_n16413_ | ~new_n33626_;
  assign new_n33653_ = ~new_n33644_ | ~new_n33627_;
  assign new_n33654_ = ~new_n16411_ | ~new_n33638_;
  assign new_n33655_ = ~new_n33642_ | ~new_n33623_;
  assign new_n33656_ = ~new_n16409_ | ~new_n33619_;
  assign new_n33657_ = ~new_n16408_ | ~new_n33622_;
  assign new_n33658_ = ~new_n16415_ | ~new_n33640_;
  assign new_n33659_ = ~new_n33647_ | ~new_n33631_;
  assign new_n33660_ = ~pi1215;
  assign new_n33661_ = ~new_n20995_ | ~new_n15522_;
  assign new_n33662_ = ~pi1216;
  assign new_n33663_ = ~pi1218;
  assign new_n33664_ = ~pi1218 | ~new_n20995_;
  assign new_n33665_ = ~pi1219;
  assign new_n33666_ = ~pi1219 | ~new_n20991_;
  assign new_n33667_ = ~pi1220;
  assign new_n33668_ = ~pi1221;
  assign new_n33669_ = ~pi1220 | ~new_n20990_;
  assign new_n33670_ = ~new_n20989_ | ~pi1221;
  assign new_n33671_ = ~pi1222;
  assign new_n33672_ = ~pi1222 | ~new_n20988_;
  assign new_n33673_ = ~pi1223;
  assign new_n33674_ = ~pi1223 | ~new_n20987_;
  assign new_n33675_ = ~pi1224;
  assign new_n33676_ = ~pi1224 | ~new_n20986_;
  assign new_n33677_ = ~pi1225;
  assign new_n33678_ = ~pi1225 | ~new_n20985_;
  assign new_n33679_ = ~pi1226;
  assign new_n33680_ = ~pi1226 | ~new_n20984_;
  assign new_n33681_ = ~pi1227;
  assign new_n33682_ = ~pi1227 | ~new_n20983_;
  assign new_n33683_ = ~pi1228;
  assign new_n33684_ = ~pi1228 | ~new_n20982_;
  assign new_n33685_ = ~pi1229;
  assign new_n33686_ = ~pi1229 | ~new_n20981_;
  assign new_n33687_ = ~pi1230;
  assign new_n33688_ = ~pi1230 | ~new_n20980_;
  assign new_n33689_ = ~pi1231;
  assign new_n33690_ = ~pi1231 | ~new_n20979_;
  assign new_n33691_ = ~pi1232;
  assign new_n33692_ = ~pi1232 | ~new_n20978_;
  assign new_n33693_ = ~pi1233;
  assign new_n33694_ = ~pi1233 | ~new_n20977_;
  assign new_n33695_ = ~pi1234;
  assign new_n33696_ = ~pi1234 | ~new_n20976_;
  assign new_n33697_ = ~pi1235;
  assign new_n33698_ = ~pi1235 | ~new_n15800_;
  assign new_n33699_ = ~pi1236;
  assign new_n33700_ = ~pi1236 | ~new_n15532_;
  assign new_n33701_ = ~pi1237;
  assign new_n33702_ = ~pi1237 | ~new_n15531_;
  assign new_n33703_ = ~pi1238;
  assign new_n33704_ = ~pi1238 | ~new_n15530_;
  assign new_n33705_ = ~pi1239;
  assign new_n33706_ = ~pi1239 | ~new_n15529_;
  assign new_n33707_ = ~pi1240;
  assign new_n33708_ = ~pi1240 | ~new_n15528_;
  assign new_n33709_ = ~pi1241;
  assign new_n33710_ = ~pi1241 | ~new_n15527_;
  assign new_n33711_ = ~pi1242;
  assign new_n33712_ = ~pi1242 | ~new_n15526_;
  assign new_n33713_ = ~pi1243;
  assign new_n33714_ = ~pi1243 | ~new_n15525_;
  assign new_n33715_ = ~pi1244;
  assign new_n33716_ = ~pi1245;
  assign new_n33717_ = ~pi1244 | ~new_n15524_;
  assign new_n33718_ = ~pi1217;
  assign new_n33719_ = ~new_n15519_ | ~new_n15520_;
  assign new_n33720_ = ~new_n15517_ | ~new_n15518_;
  assign new_n33721_ = ~new_n15515_ | ~new_n15516_;
  assign new_n33722_ = ~new_n15513_ | ~new_n15514_;
  assign new_n33723_ = ~new_n15511_ | ~new_n15512_;
  assign new_n33724_ = ~new_n15509_ | ~new_n15510_;
  assign new_n33725_ = ~new_n15507_ | ~new_n15508_;
  assign new_n33726_ = ~new_n15505_ | ~new_n15506_;
  assign new_n33727_ = ~new_n15503_ | ~new_n15504_;
  assign new_n33728_ = ~new_n15501_ | ~new_n15502_;
  assign new_n33729_ = ~new_n15499_ | ~new_n15500_;
  assign new_n33730_ = ~new_n15497_ | ~new_n15498_;
  assign new_n33731_ = ~new_n15495_ | ~new_n15496_;
  assign new_n33732_ = ~new_n15493_ | ~new_n15494_;
  assign new_n33733_ = ~new_n15491_ | ~new_n15492_;
  assign new_n33734_ = ~new_n15489_ | ~new_n15490_;
  assign new_n33735_ = ~new_n15487_ | ~new_n15488_;
  assign new_n33736_ = ~new_n15485_ | ~new_n15486_;
  assign new_n33737_ = ~new_n15483_ | ~new_n15484_;
  assign new_n33738_ = ~new_n15481_ | ~new_n15482_;
  assign new_n33739_ = ~new_n15479_ | ~new_n15480_;
  assign new_n33740_ = ~new_n15477_ | ~new_n15478_;
  assign new_n33741_ = ~new_n9391_ | ~new_n9392_;
  assign new_n33742_ = ~new_n9389_ | ~new_n9390_;
  assign po0000 = pi0443;
  assign po0001 = pi0442;
  assign po0002 = pi0441;
  assign po0003 = pi0440;
  assign po0004 = pi0439;
  assign po0005 = pi0438;
  assign po0006 = pi0437;
  assign po0007 = pi0436;
  assign po0008 = pi0435;
  assign po0009 = pi0434;
  assign po0010 = pi0433;
  assign po0011 = pi0432;
  assign po0012 = pi0431;
  assign po0013 = pi0430;
  assign po0014 = pi0429;
  assign po0015 = pi0428;
  assign po0016 = pi0427;
  assign po0017 = pi0426;
  assign po0018 = pi0425;
  assign po0019 = pi0424;
  assign po0020 = pi0423;
  assign po0021 = pi0422;
  assign po0022 = pi0421;
  assign po0023 = pi0420;
  assign po0024 = pi0419;
  assign po0025 = pi0418;
  assign po0026 = pi0417;
  assign po0027 = pi0416;
  assign po0028 = pi0415;
  assign po0029 = pi0414;
  assign po0030 = pi0413;
  assign po0031 = pi0412;
  assign po0032 = pi1008;
  assign po0033 = pi1009;
  assign po0034 = pi1010;
  assign po0035 = pi1011;
  assign po0036 = pi1012;
  assign po0037 = pi1013;
  assign po0038 = pi1014;
  assign po0039 = pi1015;
  assign po0040 = pi1016;
  assign po0041 = pi1017;
  assign po0042 = pi1018;
  assign po0043 = pi1019;
  assign po0044 = pi1020;
  assign po0045 = pi1021;
  assign po0046 = pi1022;
  assign po0047 = pi1023;
  assign po0048 = pi1024;
  assign po0049 = pi1025;
  assign po0050 = pi1026;
  assign po0051 = pi1027;
  assign po0052 = pi1028;
  assign po0053 = pi1029;
  assign po0054 = pi1030;
  assign po0055 = pi1031;
  assign po0056 = pi1032;
  assign po0057 = pi1033;
  assign po0058 = pi1034;
  assign po0059 = pi1035;
  assign po0060 = pi1036;
  assign po0061 = pi1037;
  assign po0092 = pi0544;
  assign po0093 = pi0549;
  assign po0094 = pi0550;
  assign po0095 = pi1450;
  assign po0096 = pi0552;
endmodule



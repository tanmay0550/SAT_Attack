// Benchmark "b21" written by ABC on Sun Apr 23 00:37:27 2023

module b21 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519,
    pi520, pi521, pi522,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518,
    pi519, pi520, pi521, pi522;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511;
  wire new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1138_, new_n1139_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1693_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1794_, new_n1795_, new_n1797_, new_n1798_,
    new_n1800_, new_n1801_, new_n1803_, new_n1804_, new_n1806_, new_n1807_,
    new_n1809_, new_n1810_, new_n1812_, new_n1813_, new_n1815_, new_n1816_,
    new_n1818_, new_n1819_, new_n1821_, new_n1822_, new_n1824_, new_n1825_,
    new_n1827_, new_n1828_, new_n1830_, new_n1831_, new_n1833_, new_n1834_,
    new_n1836_, new_n1837_, new_n1839_, new_n1840_, new_n1842_, new_n1843_,
    new_n1845_, new_n1846_, new_n1848_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_,
    new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_,
    new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_,
    new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_,
    new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_,
    new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_,
    new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_,
    new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_,
    new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_,
    new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_,
    new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_,
    new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_,
    new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_,
    new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_,
    new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_,
    new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_,
    new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_,
    new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_,
    new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_,
    new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_,
    new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_,
    new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_,
    new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_,
    new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_,
    new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5068_, new_n5069_, new_n5071_, new_n5072_, new_n5074_,
    new_n5075_, new_n5077_, new_n5078_, new_n5080_, new_n5081_, new_n5083_,
    new_n5084_, new_n5086_, new_n5087_, new_n5089_, new_n5090_, new_n5092_,
    new_n5093_, new_n5095_, new_n5096_, new_n5098_, new_n5099_, new_n5101_,
    new_n5102_, new_n5104_, new_n5105_, new_n5107_, new_n5108_, new_n5110_,
    new_n5111_, new_n5113_, new_n5114_, new_n5116_, new_n5117_, new_n5119_,
    new_n5120_, new_n5122_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_,
    new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_,
    new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_,
    new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_,
    new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_,
    new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_,
    new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_,
    new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_,
    new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_,
    new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_,
    new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_,
    new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_,
    new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_,
    new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_,
    new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_,
    new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_,
    new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_,
    new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_,
    new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_,
    new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_,
    new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_,
    new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_,
    new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_,
    new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_,
    new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_,
    new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_,
    new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_,
    new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_,
    new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_,
    new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_,
    new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_,
    new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_,
    new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_,
    new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_,
    new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_,
    new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_,
    new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_,
    new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_,
    new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_,
    new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_,
    new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_,
    new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_,
    new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_,
    new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_,
    new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_,
    new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_,
    new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_,
    new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_,
    new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_,
    new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_,
    new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_,
    new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_,
    new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_,
    new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_,
    new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_,
    new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_,
    new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_,
    new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_,
    new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_,
    new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_,
    new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_,
    new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_,
    new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_,
    new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_,
    new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_,
    new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_,
    new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_,
    new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_,
    new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_,
    new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_,
    new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_,
    new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_,
    new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_,
    new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_,
    new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_,
    new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_,
    new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_,
    new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_,
    new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_,
    new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_,
    new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_,
    new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_,
    new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_,
    new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_,
    new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_,
    new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_,
    new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_,
    new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_,
    new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_,
    new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_,
    new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_,
    new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_,
    new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_,
    new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_,
    new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_,
    new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_,
    new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_,
    new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_,
    new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_,
    new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_,
    new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_,
    new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_,
    new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_,
    new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_,
    new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_,
    new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_,
    new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_,
    new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_,
    new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_,
    new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_,
    new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_,
    new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_,
    new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_,
    new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_,
    new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_,
    new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_,
    new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_,
    new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_,
    new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_,
    new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_,
    new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_,
    new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_,
    new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_,
    new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_,
    new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_,
    new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_,
    new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_,
    new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_,
    new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_,
    new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_,
    new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_,
    new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_,
    new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_,
    new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_,
    new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_,
    new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_,
    new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_,
    new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_,
    new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_,
    new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_,
    new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_,
    new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_,
    new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_,
    new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_,
    new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_,
    new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_,
    new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_,
    new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_,
    new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_,
    new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_,
    new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_,
    new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_,
    new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_,
    new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_,
    new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_,
    new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_,
    new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_,
    new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_,
    new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_,
    new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_,
    new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_,
    new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_,
    new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_,
    new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_,
    new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_,
    new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_,
    new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_,
    new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_,
    new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_,
    new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_,
    new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_,
    new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_,
    new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_,
    new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_,
    new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_,
    new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_,
    new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_,
    new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_,
    new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_,
    new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_,
    new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_,
    new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_,
    new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_,
    new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_,
    new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_,
    new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_,
    new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_,
    new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_,
    new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_,
    new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_,
    new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_,
    new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_,
    new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_,
    new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_,
    new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_,
    new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_,
    new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_,
    new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_,
    new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_,
    new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_,
    new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_,
    new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_,
    new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_,
    new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_,
    new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_,
    new_n7905_, new_n7906_, new_n7907_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_,
    new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_,
    new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_,
    new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_,
    new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_,
    new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_,
    new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_,
    new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_,
    new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_,
    new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_,
    new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_,
    new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_,
    new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_,
    new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_,
    new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_,
    new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_,
    new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_,
    new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_,
    new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_,
    new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_,
    new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_,
    new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_,
    new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_,
    new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_,
    new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_,
    new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_,
    new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_,
    new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_,
    new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_,
    new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_,
    new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_,
    new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_,
    new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_,
    new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_,
    new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_,
    new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_,
    new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_,
    new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_,
    new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_,
    new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_,
    new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_,
    new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_,
    new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_,
    new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_,
    new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_,
    new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_,
    new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_,
    new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_,
    new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_,
    new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_,
    new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_,
    new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_,
    new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_,
    new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_,
    new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_,
    new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_,
    new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_,
    new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_,
    new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_,
    new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_,
    new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_,
    new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_,
    new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_,
    new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_,
    new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_,
    new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_,
    new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_,
    new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_,
    new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_,
    new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_,
    new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_,
    new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_,
    new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_,
    new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_,
    new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_,
    new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_,
    new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_,
    new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_,
    new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_,
    new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_,
    new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_,
    new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_,
    new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_,
    new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_,
    new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_,
    new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_,
    new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_,
    new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_,
    new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_,
    new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_,
    new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_,
    new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_,
    new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_,
    new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_,
    new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_,
    new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_,
    new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_,
    new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_,
    new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_,
    new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_,
    new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_,
    new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_,
    new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_,
    new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_,
    new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_,
    new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_,
    new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_,
    new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_,
    new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_,
    new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_,
    new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_,
    new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_,
    new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_,
    new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_,
    new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_,
    new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_,
    new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_,
    new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_,
    new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_,
    new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_,
    new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_,
    new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_,
    new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_,
    new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_,
    new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_,
    new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_,
    new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_,
    new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_,
    new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_,
    new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_,
    new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_,
    new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_,
    new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_,
    new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_,
    new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_,
    new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_,
    new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_,
    new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_,
    new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_,
    new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_,
    new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_,
    new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_,
    new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_,
    new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_,
    new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_,
    new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_,
    new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_,
    new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_,
    new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_,
    new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_,
    new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_,
    new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_,
    new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_,
    new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_,
    new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_,
    new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_,
    new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_,
    new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_,
    new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_,
    new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_,
    new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_,
    new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_,
    new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_,
    new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_,
    new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_,
    new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_,
    new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_,
    new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_,
    new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_,
    new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_,
    new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_,
    new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_,
    new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_,
    new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_,
    new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_,
    new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_,
    new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_,
    new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_,
    new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_,
    new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_,
    new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_,
    new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_,
    new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_,
    new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_,
    new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_,
    new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_,
    new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_,
    new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_,
    new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_,
    new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_,
    new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_,
    new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_,
    new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_,
    new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_,
    new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_,
    new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_,
    new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_,
    new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_,
    new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_,
    new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_,
    new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_,
    new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_,
    new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_,
    new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_,
    new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_,
    new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_,
    new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_,
    new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_,
    new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_,
    new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_,
    new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_,
    new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_,
    new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_,
    new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_,
    new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_,
    new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_,
    new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_,
    new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_,
    new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_,
    new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_,
    new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_,
    new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_,
    new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_,
    new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_,
    new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_,
    new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_,
    new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_,
    new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_,
    new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_,
    new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_,
    new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_,
    new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_,
    new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_,
    new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_,
    new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_,
    new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10914_,
    new_n10915_, new_n10916_, new_n10917_, new_n10918_, new_n10919_,
    new_n10920_, new_n10921_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10934_,
    new_n10935_, new_n10936_, new_n10937_, new_n10938_, new_n10939_,
    new_n10940_, new_n10941_, new_n10942_, new_n10943_, new_n10944_,
    new_n10945_, new_n10946_, new_n10947_, new_n10948_, new_n10949_,
    new_n10950_, new_n10951_, new_n10952_, new_n10953_, new_n10954_,
    new_n10955_, new_n10956_, new_n10957_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11107_, new_n11108_, new_n11109_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11148_, new_n11149_,
    new_n11150_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11373_, new_n11374_,
    new_n11375_, new_n11376_, new_n11377_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11531_, new_n11532_, new_n11533_, new_n11534_,
    new_n11535_, new_n11536_, new_n11537_, new_n11538_, new_n11539_,
    new_n11540_, new_n11541_, new_n11542_, new_n11543_, new_n11544_,
    new_n11545_, new_n11546_, new_n11547_, new_n11548_, new_n11549_,
    new_n11550_, new_n11551_, new_n11552_, new_n11553_, new_n11554_,
    new_n11555_, new_n11556_, new_n11557_, new_n11558_, new_n11559_,
    new_n11560_, new_n11561_, new_n11562_, new_n11563_, new_n11564_,
    new_n11565_, new_n11566_, new_n11567_, new_n11568_, new_n11569_,
    new_n11570_, new_n11571_, new_n11572_, new_n11573_, new_n11574_,
    new_n11575_, new_n11576_, new_n11577_, new_n11578_, new_n11579_,
    new_n11580_, new_n11581_, new_n11582_, new_n11583_, new_n11584_,
    new_n11585_, new_n11586_, new_n11587_, new_n11588_, new_n11589_,
    new_n11590_, new_n11591_, new_n11592_, new_n11593_, new_n11594_,
    new_n11595_, new_n11596_, new_n11597_, new_n11598_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11606_, new_n11607_, new_n11608_, new_n11609_,
    new_n11610_, new_n11611_, new_n11612_, new_n11613_, new_n11614_,
    new_n11615_, new_n11616_, new_n11617_, new_n11618_, new_n11619_,
    new_n11620_, new_n11621_, new_n11622_, new_n11623_, new_n11624_,
    new_n11625_, new_n11626_, new_n11627_, new_n11628_, new_n11629_,
    new_n11630_, new_n11631_, new_n11632_, new_n11633_, new_n11634_,
    new_n11635_, new_n11636_, new_n11637_, new_n11638_, new_n11639_,
    new_n11640_, new_n11641_, new_n11642_, new_n11643_, new_n11644_,
    new_n11645_, new_n11646_, new_n11647_, new_n11648_, new_n11649_,
    new_n11650_, new_n11651_, new_n11652_, new_n11653_, new_n11654_,
    new_n11655_, new_n11656_, new_n11657_, new_n11658_, new_n11659_,
    new_n11660_, new_n11661_, new_n11662_, new_n11663_, new_n11664_,
    new_n11665_, new_n11666_, new_n11667_, new_n11668_, new_n11669_,
    new_n11670_, new_n11671_, new_n11672_, new_n11673_, new_n11674_,
    new_n11675_, new_n11676_, new_n11677_, new_n11678_, new_n11679_,
    new_n11680_, new_n11681_, new_n11682_, new_n11683_, new_n11684_,
    new_n11685_, new_n11686_, new_n11687_, new_n11688_, new_n11689_,
    new_n11690_, new_n11691_, new_n11692_, new_n11693_, new_n11694_,
    new_n11695_, new_n11696_, new_n11697_, new_n11698_, new_n11699_,
    new_n11700_, new_n11701_, new_n11702_, new_n11703_, new_n11704_,
    new_n11705_, new_n11706_, new_n11707_, new_n11708_, new_n11709_,
    new_n11710_, new_n11711_, new_n11712_, new_n11713_, new_n11714_,
    new_n11715_, new_n11716_, new_n11717_, new_n11718_, new_n11719_,
    new_n11720_, new_n11721_, new_n11722_, new_n11723_, new_n11724_,
    new_n11725_, new_n11726_, new_n11727_, new_n11728_, new_n11729_,
    new_n11730_, new_n11731_, new_n11732_, new_n11733_, new_n11734_,
    new_n11735_, new_n11736_, new_n11737_, new_n11738_, new_n11739_,
    new_n11740_, new_n11741_, new_n11742_, new_n11743_, new_n11744_,
    new_n11745_, new_n11746_, new_n11747_, new_n11748_, new_n11749_,
    new_n11750_, new_n11751_, new_n11752_, new_n11753_, new_n11754_,
    new_n11755_, new_n11756_, new_n11757_, new_n11758_, new_n11759_,
    new_n11760_, new_n11761_, new_n11762_, new_n11763_, new_n11764_,
    new_n11765_, new_n11766_, new_n11767_, new_n11768_, new_n11769_,
    new_n11770_, new_n11771_, new_n11772_, new_n11773_, new_n11774_,
    new_n11775_, new_n11776_, new_n11777_, new_n11778_, new_n11779_,
    new_n11780_, new_n11781_, new_n11782_, new_n11783_, new_n11784_,
    new_n11785_, new_n11786_, new_n11787_, new_n11788_, new_n11789_,
    new_n11790_, new_n11791_, new_n11792_, new_n11793_, new_n11794_,
    new_n11795_, new_n11796_, new_n11797_, new_n11798_, new_n11799_,
    new_n11800_, new_n11801_, new_n11802_, new_n11803_, new_n11804_,
    new_n11805_, new_n11806_, new_n11807_, new_n11808_, new_n11809_,
    new_n11810_, new_n11811_, new_n11812_, new_n11813_, new_n11814_,
    new_n11815_, new_n11816_, new_n11817_, new_n11818_, new_n11819_,
    new_n11820_, new_n11821_, new_n11822_, new_n11823_, new_n11824_,
    new_n11825_, new_n11826_, new_n11827_, new_n11828_, new_n11829_,
    new_n11830_, new_n11831_, new_n11832_, new_n11833_, new_n11834_,
    new_n11835_, new_n11836_, new_n11837_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11850_, new_n11851_, new_n11852_, new_n11853_, new_n11854_,
    new_n11855_, new_n11856_, new_n11857_, new_n11858_, new_n11859_,
    new_n11860_, new_n11861_, new_n11862_, new_n11863_, new_n11864_,
    new_n11865_, new_n11866_, new_n11867_, new_n11868_, new_n11869_,
    new_n11870_, new_n11871_, new_n11872_, new_n11873_, new_n11874_,
    new_n11875_, new_n11876_, new_n11877_, new_n11878_, new_n11879_,
    new_n11880_, new_n11881_, new_n11882_, new_n11883_, new_n11884_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11891_, new_n11892_, new_n11893_, new_n11894_,
    new_n11895_, new_n11896_, new_n11897_, new_n11898_, new_n11899_,
    new_n11900_, new_n11901_, new_n11902_, new_n11903_, new_n11904_,
    new_n11905_, new_n11906_, new_n11907_, new_n11908_, new_n11909_,
    new_n11910_, new_n11911_, new_n11912_, new_n11913_, new_n11914_,
    new_n11915_, new_n11916_, new_n11917_, new_n11918_, new_n11919_,
    new_n11920_, new_n11921_, new_n11922_, new_n11923_, new_n11924_,
    new_n11925_, new_n11926_, new_n11927_, new_n11928_, new_n11929_,
    new_n11930_, new_n11931_, new_n11932_, new_n11933_, new_n11934_,
    new_n11935_, new_n11936_, new_n11937_, new_n11938_, new_n11939_,
    new_n11940_, new_n11941_, new_n11942_, new_n11943_, new_n11944_,
    new_n11945_, new_n11946_, new_n11947_, new_n11948_, new_n11949_,
    new_n11950_, new_n11951_, new_n11952_, new_n11953_, new_n11954_,
    new_n11955_, new_n11956_, new_n11957_, new_n11958_, new_n11959_,
    new_n11960_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11965_, new_n11966_, new_n11967_, new_n11968_, new_n11969_,
    new_n11970_, new_n11971_, new_n11972_, new_n11973_, new_n11974_,
    new_n11975_, new_n11976_, new_n11977_, new_n11978_, new_n11979_,
    new_n11980_, new_n11981_, new_n11982_, new_n11983_, new_n11984_,
    new_n11985_, new_n11986_, new_n11987_, new_n11988_, new_n11989_,
    new_n11990_, new_n11991_, new_n11992_, new_n11993_, new_n11994_,
    new_n11995_, new_n11996_, new_n11997_, new_n11998_, new_n11999_,
    new_n12000_, new_n12001_, new_n12002_, new_n12003_, new_n12004_,
    new_n12005_, new_n12006_, new_n12007_, new_n12008_, new_n12009_,
    new_n12010_, new_n12011_, new_n12012_, new_n12013_, new_n12014_,
    new_n12015_, new_n12016_, new_n12017_, new_n12018_, new_n12019_,
    new_n12020_, new_n12021_, new_n12022_, new_n12023_, new_n12024_,
    new_n12025_, new_n12026_, new_n12027_, new_n12028_, new_n12029_,
    new_n12030_, new_n12031_, new_n12032_, new_n12033_, new_n12034_,
    new_n12035_, new_n12036_, new_n12037_, new_n12038_, new_n12039_,
    new_n12040_, new_n12041_, new_n12042_, new_n12043_, new_n12044_,
    new_n12045_, new_n12046_, new_n12047_, new_n12048_, new_n12049_,
    new_n12050_, new_n12051_, new_n12052_, new_n12053_, new_n12054_,
    new_n12055_, new_n12056_, new_n12057_, new_n12058_, new_n12059_,
    new_n12060_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12098_, new_n12099_,
    new_n12100_, new_n12101_, new_n12102_, new_n12103_, new_n12104_,
    new_n12105_, new_n12106_, new_n12107_, new_n12108_, new_n12109_,
    new_n12110_, new_n12111_, new_n12112_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12221_, new_n12222_, new_n12223_, new_n12224_,
    new_n12225_, new_n12226_, new_n12227_, new_n12228_, new_n12229_,
    new_n12230_, new_n12231_, new_n12232_, new_n12233_, new_n12234_,
    new_n12235_, new_n12236_, new_n12237_, new_n12238_, new_n12239_,
    new_n12240_, new_n12241_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12247_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12260_, new_n12261_, new_n12262_, new_n12263_, new_n12264_,
    new_n12265_, new_n12266_, new_n12267_, new_n12268_, new_n12269_,
    new_n12270_, new_n12271_, new_n12272_, new_n12273_, new_n12274_,
    new_n12275_, new_n12276_, new_n12277_, new_n12278_, new_n12279_,
    new_n12280_, new_n12281_, new_n12282_, new_n12283_, new_n12284_,
    new_n12285_, new_n12286_, new_n12287_, new_n12288_, new_n12289_,
    new_n12290_, new_n12291_, new_n12292_, new_n12293_, new_n12294_,
    new_n12295_, new_n12296_, new_n12297_, new_n12298_, new_n12299_,
    new_n12300_, new_n12301_, new_n12302_, new_n12303_, new_n12304_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12561_, new_n12562_, new_n12563_, new_n12564_,
    new_n12565_, new_n12566_, new_n12567_, new_n12568_, new_n12569_,
    new_n12570_, new_n12571_, new_n12572_, new_n12573_, new_n12574_,
    new_n12575_, new_n12576_, new_n12577_, new_n12578_, new_n12579_,
    new_n12580_, new_n12581_, new_n12582_, new_n12583_, new_n12584_,
    new_n12585_, new_n12586_, new_n12587_, new_n12588_, new_n12589_,
    new_n12590_, new_n12591_, new_n12592_, new_n12593_, new_n12594_,
    new_n12595_, new_n12596_, new_n12597_, new_n12598_, new_n12599_,
    new_n12600_, new_n12601_, new_n12602_, new_n12603_, new_n12604_,
    new_n12605_, new_n12606_, new_n12607_, new_n12608_, new_n12609_,
    new_n12610_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12639_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13102_, new_n13103_, new_n13104_,
    new_n13105_, new_n13106_, new_n13107_, new_n13108_, new_n13109_,
    new_n13110_, new_n13111_, new_n13112_, new_n13113_, new_n13114_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13121_, new_n13122_, new_n13123_, new_n13124_,
    new_n13125_, new_n13126_, new_n13127_, new_n13128_, new_n13129_,
    new_n13130_, new_n13131_, new_n13132_, new_n13133_, new_n13134_,
    new_n13135_, new_n13136_, new_n13137_, new_n13138_, new_n13139_,
    new_n13140_, new_n13141_, new_n13142_, new_n13143_, new_n13144_,
    new_n13145_, new_n13146_, new_n13147_, new_n13148_, new_n13149_,
    new_n13150_, new_n13151_, new_n13152_, new_n13153_, new_n13154_,
    new_n13155_, new_n13156_, new_n13157_, new_n13158_, new_n13159_,
    new_n13160_, new_n13161_, new_n13162_, new_n13163_, new_n13164_,
    new_n13165_, new_n13166_, new_n13167_, new_n13168_, new_n13169_,
    new_n13170_, new_n13171_, new_n13172_, new_n13173_, new_n13174_,
    new_n13175_, new_n13176_, new_n13177_, new_n13178_, new_n13179_,
    new_n13180_, new_n13181_, new_n13182_, new_n13183_, new_n13184_,
    new_n13185_, new_n13186_, new_n13187_, new_n13188_, new_n13189_,
    new_n13190_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13200_, new_n13201_, new_n13202_, new_n13203_, new_n13204_,
    new_n13205_, new_n13206_, new_n13207_, new_n13208_, new_n13209_,
    new_n13210_, new_n13211_, new_n13212_, new_n13213_, new_n13214_,
    new_n13215_, new_n13216_, new_n13217_, new_n13218_, new_n13219_,
    new_n13220_, new_n13221_, new_n13222_, new_n13223_, new_n13224_,
    new_n13225_, new_n13226_, new_n13227_, new_n13228_, new_n13229_,
    new_n13230_, new_n13231_, new_n13232_, new_n13233_, new_n13234_,
    new_n13235_, new_n13236_, new_n13237_, new_n13238_, new_n13239_,
    new_n13240_, new_n13241_, new_n13242_, new_n13243_, new_n13244_,
    new_n13245_, new_n13246_, new_n13247_, new_n13248_, new_n13249_,
    new_n13250_, new_n13251_, new_n13252_, new_n13253_, new_n13254_,
    new_n13255_, new_n13256_, new_n13257_, new_n13258_, new_n13259_,
    new_n13260_, new_n13261_, new_n13262_, new_n13263_, new_n13264_,
    new_n13265_, new_n13266_, new_n13267_, new_n13268_, new_n13269_,
    new_n13270_, new_n13271_, new_n13272_, new_n13273_, new_n13274_,
    new_n13275_, new_n13276_, new_n13277_, new_n13278_, new_n13279_,
    new_n13280_, new_n13281_, new_n13282_, new_n13283_, new_n13284_,
    new_n13285_, new_n13286_, new_n13287_, new_n13288_, new_n13289_,
    new_n13290_, new_n13291_, new_n13292_, new_n13293_, new_n13294_,
    new_n13295_, new_n13296_, new_n13297_, new_n13298_, new_n13299_,
    new_n13300_, new_n13301_, new_n13302_, new_n13303_, new_n13304_,
    new_n13305_, new_n13306_, new_n13307_, new_n13308_, new_n13309_,
    new_n13310_, new_n13311_, new_n13312_, new_n13313_, new_n13314_,
    new_n13315_, new_n13316_, new_n13317_, new_n13318_, new_n13319_,
    new_n13320_, new_n13321_, new_n13322_, new_n13323_, new_n13324_,
    new_n13325_, new_n13326_, new_n13327_, new_n13328_, new_n13329_,
    new_n13330_, new_n13331_, new_n13332_, new_n13333_, new_n13334_,
    new_n13335_, new_n13336_, new_n13337_, new_n13338_, new_n13339_,
    new_n13340_, new_n13341_, new_n13342_, new_n13343_, new_n13344_,
    new_n13345_, new_n13346_, new_n13347_, new_n13348_, new_n13349_,
    new_n13350_, new_n13351_, new_n13352_, new_n13353_, new_n13354_,
    new_n13355_, new_n13356_, new_n13357_, new_n13358_, new_n13359_,
    new_n13360_, new_n13361_, new_n13362_, new_n13363_, new_n13364_,
    new_n13365_, new_n13366_, new_n13367_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13375_, new_n13376_, new_n13377_, new_n13378_, new_n13379_,
    new_n13380_, new_n13381_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13407_, new_n13408_, new_n13409_,
    new_n13410_, new_n13411_, new_n13412_, new_n13413_, new_n13414_,
    new_n13415_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13438_, new_n13439_,
    new_n13440_, new_n13441_, new_n13442_, new_n13443_, new_n13444_,
    new_n13445_, new_n13446_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13452_, new_n13453_, new_n13454_,
    new_n13455_, new_n13456_, new_n13457_, new_n13458_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13464_,
    new_n13465_, new_n13466_, new_n13467_, new_n13468_, new_n13469_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13511_, new_n13512_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13539_,
    new_n13540_, new_n13541_, new_n13542_, new_n13543_, new_n13544_,
    new_n13545_, new_n13546_, new_n13547_, new_n13548_, new_n13549_,
    new_n13550_, new_n13551_, new_n13552_, new_n13553_, new_n13554_,
    new_n13555_, new_n13556_, new_n13557_, new_n13558_, new_n13559_,
    new_n13560_, new_n13561_, new_n13562_, new_n13563_, new_n13564_,
    new_n13565_, new_n13566_, new_n13567_, new_n13568_, new_n13569_,
    new_n13570_, new_n13571_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13591_, new_n13592_, new_n13593_, new_n13594_,
    new_n13595_, new_n13596_, new_n13597_, new_n13598_, new_n13599_,
    new_n13600_, new_n13601_, new_n13602_, new_n13603_, new_n13604_,
    new_n13605_, new_n13606_, new_n13607_, new_n13608_, new_n13609_,
    new_n13610_, new_n13611_, new_n13612_, new_n13613_, new_n13614_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13660_, new_n13661_, new_n13662_, new_n13663_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13685_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13690_, new_n13691_, new_n13692_, new_n13693_, new_n13694_,
    new_n13695_, new_n13696_, new_n13697_, new_n13698_, new_n13699_,
    new_n13700_, new_n13701_, new_n13702_, new_n13703_, new_n13704_,
    new_n13705_, new_n13706_, new_n13707_, new_n13708_, new_n13709_,
    new_n13710_, new_n13711_, new_n13712_, new_n13713_, new_n13714_,
    new_n13715_, new_n13716_, new_n13717_, new_n13718_, new_n13719_,
    new_n13720_, new_n13721_, new_n13722_, new_n13723_, new_n13724_,
    new_n13725_, new_n13726_, new_n13727_, new_n13728_, new_n13729_,
    new_n13730_, new_n13731_, new_n13732_, new_n13733_, new_n13734_,
    new_n13735_, new_n13736_, new_n13737_, new_n13738_, new_n13739_,
    new_n13740_, new_n13741_, new_n13742_, new_n13743_, new_n13744_,
    new_n13745_, new_n13746_, new_n13747_, new_n13748_, new_n13749_,
    new_n13750_, new_n13751_, new_n13752_, new_n13753_, new_n13754_,
    new_n13755_, new_n13756_, new_n13757_, new_n13758_, new_n13759_,
    new_n13760_, new_n13761_, new_n13762_, new_n13763_, new_n13764_,
    new_n13765_, new_n13766_, new_n13767_, new_n13768_, new_n13769_,
    new_n13770_, new_n13771_, new_n13772_, new_n13773_, new_n13774_,
    new_n13775_, new_n13776_, new_n13777_, new_n13778_, new_n13779_,
    new_n13780_, new_n13781_, new_n13782_, new_n13783_, new_n13784_,
    new_n13785_, new_n13786_, new_n13787_, new_n13788_, new_n13789_,
    new_n13790_, new_n13791_, new_n13792_, new_n13793_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13800_, new_n13801_, new_n13802_, new_n13803_, new_n13804_,
    new_n13805_, new_n13806_, new_n13807_, new_n13808_, new_n13809_,
    new_n13810_, new_n13811_, new_n13812_, new_n13813_, new_n13814_,
    new_n13815_, new_n13816_, new_n13817_, new_n13818_, new_n13819_,
    new_n13820_, new_n13821_, new_n13822_, new_n13823_, new_n13824_,
    new_n13825_, new_n13826_, new_n13827_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13835_, new_n13836_, new_n13837_, new_n13838_, new_n13839_,
    new_n13840_, new_n13841_, new_n13842_, new_n13843_, new_n13844_,
    new_n13845_, new_n13846_, new_n13847_, new_n13848_, new_n13849_,
    new_n13850_, new_n13851_, new_n13852_, new_n13853_, new_n13854_,
    new_n13855_, new_n13856_, new_n13857_, new_n13858_, new_n13859_,
    new_n13860_, new_n13861_, new_n13862_, new_n13863_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13869_,
    new_n13870_, new_n13871_, new_n13872_, new_n13873_, new_n13874_,
    new_n13875_, new_n13876_, new_n13877_, new_n13878_, new_n13879_,
    new_n13880_, new_n13881_, new_n13882_, new_n13883_, new_n13884_,
    new_n13885_, new_n13886_, new_n13887_, new_n13888_, new_n13889_,
    new_n13890_, new_n13891_, new_n13892_, new_n13893_, new_n13894_,
    new_n13895_, new_n13896_, new_n13897_, new_n13898_, new_n13899_,
    new_n13900_, new_n13901_, new_n13902_, new_n13903_, new_n13904_,
    new_n13905_, new_n13906_, new_n13907_, new_n13908_, new_n13909_,
    new_n13910_, new_n13911_, new_n13912_, new_n13913_, new_n13914_,
    new_n13915_, new_n13916_, new_n13917_, new_n13918_, new_n13919_,
    new_n13920_, new_n13921_, new_n13922_, new_n13923_, new_n13924_,
    new_n13925_, new_n13926_, new_n13927_, new_n13928_, new_n13929_,
    new_n13930_, new_n13931_, new_n13932_, new_n13933_, new_n13934_,
    new_n13935_, new_n13936_, new_n13937_, new_n13938_, new_n13939_,
    new_n13940_, new_n13941_, new_n13942_, new_n13943_, new_n13944_,
    new_n13945_, new_n13946_, new_n13947_, new_n13948_, new_n13949_,
    new_n13950_, new_n13951_, new_n13952_, new_n13953_, new_n13954_,
    new_n13955_, new_n13956_, new_n13957_, new_n13958_, new_n13959_,
    new_n13960_, new_n13961_, new_n13962_, new_n13963_, new_n13964_,
    new_n13965_, new_n13966_, new_n13967_, new_n13968_, new_n13969_,
    new_n13970_, new_n13971_, new_n13972_, new_n13973_, new_n13974_,
    new_n13975_, new_n13976_, new_n13977_, new_n13978_, new_n13979_,
    new_n13980_, new_n13981_, new_n13982_, new_n13983_, new_n13984_,
    new_n13985_, new_n13986_, new_n13987_, new_n13988_, new_n13989_,
    new_n13990_, new_n13991_, new_n13992_, new_n13993_, new_n13994_,
    new_n13995_, new_n13996_, new_n13997_, new_n13998_, new_n13999_,
    new_n14000_, new_n14001_, new_n14002_, new_n14003_, new_n14004_,
    new_n14005_, new_n14006_, new_n14007_, new_n14008_, new_n14009_,
    new_n14010_, new_n14011_, new_n14012_, new_n14013_, new_n14014_,
    new_n14015_, new_n14016_, new_n14017_, new_n14018_, new_n14019_,
    new_n14020_, new_n14021_, new_n14022_, new_n14023_, new_n14024_,
    new_n14025_, new_n14026_, new_n14027_, new_n14028_, new_n14029_,
    new_n14030_, new_n14031_, new_n14032_, new_n14033_, new_n14034_,
    new_n14035_, new_n14036_, new_n14037_, new_n14038_, new_n14039_,
    new_n14040_, new_n14041_, new_n14042_, new_n14043_, new_n14044_,
    new_n14045_, new_n14046_, new_n14047_, new_n14048_, new_n14049_,
    new_n14050_, new_n14051_, new_n14052_, new_n14053_, new_n14054_,
    new_n14055_, new_n14056_, new_n14057_, new_n14058_, new_n14059_,
    new_n14060_, new_n14061_, new_n14062_, new_n14063_, new_n14064_,
    new_n14065_, new_n14066_, new_n14067_, new_n14068_, new_n14069_,
    new_n14070_, new_n14071_, new_n14072_, new_n14073_, new_n14074_,
    new_n14075_, new_n14076_, new_n14077_, new_n14078_, new_n14079_,
    new_n14080_, new_n14081_, new_n14082_, new_n14083_, new_n14084_,
    new_n14085_, new_n14086_, new_n14087_, new_n14088_, new_n14089_,
    new_n14090_, new_n14091_, new_n14092_, new_n14093_, new_n14094_,
    new_n14095_, new_n14096_, new_n14097_, new_n14098_, new_n14099_,
    new_n14100_, new_n14101_, new_n14102_, new_n14103_, new_n14104_,
    new_n14105_, new_n14106_, new_n14107_, new_n14108_, new_n14109_,
    new_n14110_, new_n14111_, new_n14112_, new_n14113_, new_n14114_,
    new_n14115_, new_n14116_, new_n14117_, new_n14118_, new_n14119_,
    new_n14120_, new_n14121_, new_n14122_, new_n14123_, new_n14124_,
    new_n14125_, new_n14126_, new_n14127_, new_n14128_, new_n14129_,
    new_n14130_, new_n14131_, new_n14132_, new_n14133_, new_n14134_,
    new_n14135_, new_n14136_, new_n14137_, new_n14138_, new_n14139_,
    new_n14140_, new_n14141_, new_n14142_, new_n14143_, new_n14144_,
    new_n14145_, new_n14146_, new_n14147_, new_n14148_, new_n14149_,
    new_n14150_, new_n14151_, new_n14152_, new_n14153_, new_n14154_,
    new_n14155_, new_n14156_, new_n14157_, new_n14158_, new_n14159_,
    new_n14160_, new_n14161_, new_n14162_, new_n14163_, new_n14164_,
    new_n14165_, new_n14166_, new_n14167_, new_n14168_, new_n14169_,
    new_n14170_, new_n14171_, new_n14172_, new_n14173_, new_n14174_,
    new_n14175_, new_n14176_, new_n14177_, new_n14178_, new_n14179_,
    new_n14180_, new_n14181_, new_n14182_, new_n14183_, new_n14184_,
    new_n14185_, new_n14186_, new_n14187_, new_n14188_, new_n14189_,
    new_n14190_, new_n14191_, new_n14192_, new_n14193_, new_n14194_,
    new_n14195_, new_n14196_, new_n14197_, new_n14198_, new_n14199_,
    new_n14200_, new_n14201_, new_n14202_, new_n14203_, new_n14204_,
    new_n14205_, new_n14206_, new_n14207_, new_n14208_, new_n14209_,
    new_n14210_, new_n14211_, new_n14212_, new_n14213_, new_n14214_,
    new_n14215_, new_n14216_, new_n14217_, new_n14218_, new_n14219_,
    new_n14220_, new_n14221_, new_n14222_, new_n14223_, new_n14224_,
    new_n14225_, new_n14226_, new_n14227_, new_n14228_, new_n14229_,
    new_n14230_, new_n14231_, new_n14232_, new_n14233_, new_n14234_,
    new_n14235_, new_n14236_, new_n14237_, new_n14238_, new_n14239_,
    new_n14240_, new_n14241_, new_n14242_, new_n14243_, new_n14244_,
    new_n14245_, new_n14246_, new_n14247_, new_n14248_, new_n14249_,
    new_n14250_, new_n14251_, new_n14252_, new_n14253_, new_n14254_,
    new_n14255_, new_n14256_, new_n14257_, new_n14258_, new_n14259_,
    new_n14260_, new_n14261_, new_n14262_, new_n14263_, new_n14264_,
    new_n14265_, new_n14266_, new_n14267_, new_n14268_, new_n14269_,
    new_n14270_, new_n14271_, new_n14272_, new_n14273_, new_n14274_,
    new_n14275_, new_n14276_, new_n14277_, new_n14278_, new_n14279_,
    new_n14280_, new_n14281_, new_n14282_, new_n14283_, new_n14284_,
    new_n14285_, new_n14286_, new_n14287_, new_n14288_, new_n14289_,
    new_n14290_, new_n14291_, new_n14292_, new_n14293_, new_n14294_,
    new_n14295_, new_n14296_, new_n14297_, new_n14298_, new_n14299_,
    new_n14300_, new_n14301_, new_n14302_, new_n14303_, new_n14304_,
    new_n14305_, new_n14306_, new_n14307_, new_n14308_, new_n14309_,
    new_n14310_, new_n14311_, new_n14312_, new_n14313_, new_n14314_,
    new_n14315_, new_n14316_, new_n14317_, new_n14318_, new_n14319_,
    new_n14320_, new_n14321_, new_n14322_, new_n14323_, new_n14324_,
    new_n14325_, new_n14326_, new_n14327_, new_n14328_, new_n14329_,
    new_n14330_, new_n14331_, new_n14332_, new_n14333_, new_n14334_,
    new_n14335_, new_n14336_, new_n14337_, new_n14338_, new_n14339_,
    new_n14340_, new_n14341_, new_n14342_, new_n14343_, new_n14344_,
    new_n14345_, new_n14346_, new_n14347_, new_n14348_, new_n14349_,
    new_n14350_, new_n14351_, new_n14352_, new_n14353_, new_n14354_,
    new_n14355_, new_n14356_, new_n14357_, new_n14358_, new_n14359_,
    new_n14360_, new_n14361_, new_n14362_, new_n14363_, new_n14364_,
    new_n14365_, new_n14366_, new_n14367_, new_n14368_, new_n14369_,
    new_n14370_, new_n14371_, new_n14372_, new_n14373_, new_n14374_,
    new_n14375_, new_n14376_, new_n14377_, new_n14378_, new_n14379_,
    new_n14380_, new_n14381_, new_n14382_, new_n14383_, new_n14384_,
    new_n14385_, new_n14386_, new_n14387_, new_n14388_, new_n14389_,
    new_n14390_, new_n14391_, new_n14392_, new_n14393_, new_n14394_,
    new_n14395_, new_n14396_, new_n14397_, new_n14398_, new_n14399_,
    new_n14400_, new_n14401_, new_n14402_, new_n14403_, new_n14404_,
    new_n14405_, new_n14406_, new_n14407_, new_n14408_, new_n14409_,
    new_n14410_, new_n14411_, new_n14412_, new_n14413_, new_n14414_,
    new_n14415_, new_n14416_, new_n14417_, new_n14418_, new_n14419_,
    new_n14420_, new_n14421_, new_n14422_, new_n14423_, new_n14424_,
    new_n14425_, new_n14426_, new_n14427_, new_n14428_, new_n14429_,
    new_n14430_, new_n14431_, new_n14432_, new_n14433_, new_n14434_,
    new_n14435_, new_n14436_, new_n14437_, new_n14438_, new_n14439_,
    new_n14440_, new_n14441_, new_n14442_, new_n14443_, new_n14444_,
    new_n14445_, new_n14446_, new_n14447_, new_n14448_, new_n14449_,
    new_n14450_, new_n14451_, new_n14452_, new_n14453_, new_n14454_,
    new_n14455_, new_n14456_, new_n14457_, new_n14458_, new_n14459_,
    new_n14460_, new_n14461_, new_n14462_, new_n14463_, new_n14464_,
    new_n14465_, new_n14466_, new_n14467_, new_n14468_, new_n14469_,
    new_n14470_, new_n14471_, new_n14472_, new_n14473_, new_n14474_,
    new_n14475_, new_n14476_, new_n14477_, new_n14478_, new_n14479_,
    new_n14480_, new_n14481_, new_n14482_, new_n14483_, new_n14484_,
    new_n14485_, new_n14486_, new_n14487_, new_n14488_, new_n14489_,
    new_n14490_, new_n14491_, new_n14492_, new_n14493_, new_n14494_,
    new_n14495_, new_n14496_, new_n14497_, new_n14498_, new_n14499_,
    new_n14500_, new_n14501_, new_n14502_, new_n14503_, new_n14504_,
    new_n14505_, new_n14506_, new_n14507_, new_n14508_, new_n14509_,
    new_n14510_, new_n14511_, new_n14512_, new_n14513_, new_n14514_,
    new_n14515_, new_n14516_, new_n14517_, new_n14518_, new_n14519_,
    new_n14520_, new_n14521_, new_n14522_, new_n14523_, new_n14524_,
    new_n14525_, new_n14526_, new_n14527_, new_n14528_, new_n14529_,
    new_n14530_, new_n14531_, new_n14532_, new_n14533_, new_n14534_,
    new_n14535_, new_n14536_, new_n14537_, new_n14538_, new_n14539_,
    new_n14540_, new_n14541_, new_n14542_, new_n14543_, new_n14544_,
    new_n14545_, new_n14546_, new_n14547_, new_n14548_, new_n14549_,
    new_n14550_, new_n14551_, new_n14552_, new_n14553_, new_n14554_,
    new_n14555_, new_n14556_, new_n14557_, new_n14558_, new_n14559_,
    new_n14560_, new_n14561_, new_n14562_, new_n14563_, new_n14564_,
    new_n14565_, new_n14566_, new_n14567_, new_n14568_, new_n14569_,
    new_n14570_, new_n14571_, new_n14572_, new_n14573_, new_n14574_,
    new_n14575_, new_n14576_, new_n14577_, new_n14578_, new_n14579_,
    new_n14580_, new_n14581_, new_n14582_, new_n14583_, new_n14584_,
    new_n14585_, new_n14586_, new_n14587_, new_n14588_, new_n14589_,
    new_n14590_, new_n14591_, new_n14592_, new_n14593_, new_n14594_,
    new_n14595_, new_n14596_, new_n14597_, new_n14598_, new_n14599_,
    new_n14600_, new_n14601_, new_n14602_, new_n14603_, new_n14604_,
    new_n14605_, new_n14606_, new_n14607_, new_n14608_, new_n14609_,
    new_n14610_, new_n14611_, new_n14612_, new_n14613_, new_n14614_,
    new_n14615_, new_n14616_, new_n14617_, new_n14618_, new_n14619_,
    new_n14620_, new_n14621_, new_n14622_, new_n14623_, new_n14624_,
    new_n14625_, new_n14626_, new_n14627_, new_n14628_, new_n14629_,
    new_n14630_, new_n14631_, new_n14632_, new_n14633_, new_n14634_,
    new_n14635_, new_n14636_, new_n14637_, new_n14638_, new_n14639_,
    new_n14640_, new_n14641_, new_n14642_, new_n14643_, new_n14644_,
    new_n14645_, new_n14646_, new_n14647_, new_n14648_, new_n14649_,
    new_n14650_, new_n14651_, new_n14652_, new_n14653_, new_n14654_,
    new_n14655_, new_n14656_, new_n14657_, new_n14658_, new_n14659_,
    new_n14660_, new_n14661_, new_n14662_, new_n14663_, new_n14664_,
    new_n14665_, new_n14666_, new_n14667_, new_n14668_, new_n14669_,
    new_n14670_, new_n14671_, new_n14672_, new_n14673_, new_n14674_,
    new_n14675_, new_n14676_, new_n14677_, new_n14678_, new_n14679_,
    new_n14680_, new_n14681_, new_n14682_, new_n14683_, new_n14684_,
    new_n14685_, new_n14686_, new_n14687_, new_n14688_, new_n14689_,
    new_n14690_, new_n14691_, new_n14692_, new_n14693_, new_n14694_,
    new_n14695_, new_n14696_, new_n14697_, new_n14698_, new_n14699_,
    new_n14700_, new_n14701_, new_n14702_, new_n14703_, new_n14704_,
    new_n14705_, new_n14706_, new_n14707_, new_n14708_, new_n14709_,
    new_n14710_, new_n14711_, new_n14712_, new_n14713_, new_n14714_,
    new_n14715_, new_n14716_, new_n14717_, new_n14718_, new_n14719_,
    new_n14720_, new_n14721_, new_n14722_, new_n14723_, new_n14724_,
    new_n14725_, new_n14726_, new_n14727_, new_n14728_, new_n14729_,
    new_n14730_, new_n14731_, new_n14732_, new_n14733_, new_n14734_,
    new_n14735_, new_n14736_, new_n14737_, new_n14738_, new_n14739_,
    new_n14740_, new_n14741_, new_n14742_, new_n14743_, new_n14744_,
    new_n14745_, new_n14746_, new_n14747_, new_n14748_, new_n14749_,
    new_n14750_, new_n14751_, new_n14752_, new_n14753_, new_n14754_,
    new_n14755_, new_n14756_, new_n14757_, new_n14758_, new_n14759_,
    new_n14760_, new_n14761_, new_n14762_, new_n14763_, new_n14764_,
    new_n14765_, new_n14766_, new_n14767_, new_n14768_, new_n14769_,
    new_n14770_, new_n14771_, new_n14772_, new_n14773_, new_n14774_,
    new_n14775_, new_n14776_, new_n14777_, new_n14778_, new_n14779_,
    new_n14780_, new_n14781_, new_n14782_, new_n14783_, new_n14784_,
    new_n14785_, new_n14786_, new_n14787_, new_n14788_, new_n14789_,
    new_n14790_, new_n14791_, new_n14792_, new_n14793_, new_n14794_,
    new_n14795_, new_n14796_, new_n14797_, new_n14798_, new_n14799_,
    new_n14800_, new_n14801_, new_n14802_, new_n14803_, new_n14804_,
    new_n14805_, new_n14806_, new_n14807_, new_n14808_, new_n14809_,
    new_n14810_, new_n14811_, new_n14812_, new_n14813_, new_n14814_,
    new_n14815_, new_n14816_, new_n14817_, new_n14818_, new_n14819_,
    new_n14820_, new_n14821_, new_n14822_, new_n14823_, new_n14824_,
    new_n14825_, new_n14826_, new_n14827_, new_n14828_, new_n14829_,
    new_n14830_, new_n14831_, new_n14832_, new_n14833_, new_n14834_,
    new_n14835_, new_n14836_, new_n14837_, new_n14838_, new_n14839_,
    new_n14840_, new_n14841_, new_n14842_, new_n14843_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14908_, new_n14909_,
    new_n14910_, new_n14911_, new_n14912_, new_n14913_, new_n14914_,
    new_n14915_, new_n14916_, new_n14917_, new_n14918_, new_n14919_,
    new_n14920_, new_n14921_, new_n14922_, new_n14923_, new_n14924_,
    new_n14925_, new_n14926_, new_n14927_, new_n14928_, new_n14929_,
    new_n14930_, new_n14931_, new_n14932_, new_n14933_, new_n14934_,
    new_n14935_, new_n14936_, new_n14937_, new_n14938_, new_n14939_,
    new_n14940_, new_n14941_, new_n14942_, new_n14943_, new_n14944_,
    new_n14945_, new_n14946_, new_n14947_, new_n14948_, new_n14949_,
    new_n14950_, new_n14951_, new_n14952_, new_n14953_, new_n14954_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14963_, new_n14964_,
    new_n14965_, new_n14966_, new_n14967_, new_n14968_, new_n14969_,
    new_n14970_, new_n14971_, new_n14972_, new_n14973_, new_n14974_,
    new_n14975_, new_n14976_, new_n14977_, new_n14978_, new_n14979_,
    new_n14980_, new_n14981_, new_n14982_, new_n14983_, new_n14984_,
    new_n14985_, new_n14986_, new_n14987_, new_n14988_, new_n14989_,
    new_n14990_, new_n14991_, new_n14992_, new_n14993_, new_n14994_,
    new_n14995_, new_n14996_, new_n14997_, new_n14998_, new_n14999_,
    new_n15000_, new_n15001_, new_n15002_, new_n15003_, new_n15004_,
    new_n15005_, new_n15006_, new_n15007_, new_n15008_, new_n15009_,
    new_n15010_, new_n15011_, new_n15012_, new_n15013_, new_n15014_,
    new_n15015_, new_n15016_, new_n15017_, new_n15018_, new_n15019_,
    new_n15020_, new_n15021_, new_n15022_, new_n15023_, new_n15024_,
    new_n15025_, new_n15026_, new_n15027_, new_n15028_, new_n15029_,
    new_n15030_, new_n15031_, new_n15032_, new_n15033_, new_n15034_,
    new_n15035_, new_n15036_, new_n15037_, new_n15038_, new_n15039_,
    new_n15040_, new_n15041_, new_n15042_, new_n15043_, new_n15044_,
    new_n15045_, new_n15046_, new_n15047_, new_n15048_, new_n15049_,
    new_n15050_, new_n15051_, new_n15052_, new_n15053_, new_n15054_,
    new_n15055_, new_n15056_, new_n15057_, new_n15058_, new_n15059_,
    new_n15060_, new_n15061_, new_n15062_, new_n15063_, new_n15064_,
    new_n15065_, new_n15066_, new_n15067_, new_n15068_, new_n15069_,
    new_n15070_, new_n15071_, new_n15072_, new_n15073_, new_n15074_,
    new_n15075_, new_n15076_, new_n15077_, new_n15078_, new_n15079_,
    new_n15080_, new_n15081_, new_n15082_, new_n15083_, new_n15084_,
    new_n15085_, new_n15086_, new_n15087_, new_n15088_, new_n15089_,
    new_n15090_, new_n15091_, new_n15092_, new_n15093_, new_n15094_,
    new_n15095_, new_n15096_, new_n15097_, new_n15098_, new_n15099_,
    new_n15100_, new_n15101_, new_n15102_, new_n15103_, new_n15104_,
    new_n15105_, new_n15106_, new_n15107_, new_n15108_, new_n15109_,
    new_n15110_, new_n15111_, new_n15112_, new_n15113_, new_n15114_,
    new_n15115_, new_n15116_, new_n15117_, new_n15118_, new_n15119_,
    new_n15120_, new_n15121_, new_n15122_, new_n15123_, new_n15124_,
    new_n15125_, new_n15126_, new_n15127_, new_n15128_, new_n15129_,
    new_n15130_, new_n15131_, new_n15132_, new_n15133_, new_n15134_,
    new_n15135_, new_n15136_, new_n15137_, new_n15138_, new_n15139_,
    new_n15140_, new_n15141_, new_n15142_, new_n15143_, new_n15144_,
    new_n15145_, new_n15146_, new_n15147_, new_n15148_, new_n15149_,
    new_n15150_, new_n15151_, new_n15152_, new_n15153_, new_n15154_,
    new_n15155_, new_n15156_, new_n15157_, new_n15158_, new_n15159_,
    new_n15160_, new_n15161_, new_n15162_, new_n15163_, new_n15164_,
    new_n15165_, new_n15166_, new_n15167_, new_n15168_, new_n15169_,
    new_n15170_, new_n15171_, new_n15172_, new_n15173_, new_n15174_,
    new_n15175_, new_n15176_, new_n15177_, new_n15178_, new_n15179_,
    new_n15180_, new_n15181_, new_n15182_, new_n15183_, new_n15184_,
    new_n15185_, new_n15186_, new_n15187_, new_n15188_, new_n15189_,
    new_n15190_, new_n15191_, new_n15192_, new_n15193_, new_n15194_,
    new_n15195_, new_n15196_, new_n15197_, new_n15198_, new_n15199_,
    new_n15200_, new_n15201_, new_n15202_, new_n15203_, new_n15204_,
    new_n15205_, new_n15206_, new_n15207_, new_n15208_, new_n15209_,
    new_n15210_, new_n15211_, new_n15212_, new_n15213_, new_n15214_,
    new_n15215_, new_n15216_, new_n15217_, new_n15218_, new_n15219_,
    new_n15220_, new_n15221_, new_n15222_, new_n15223_, new_n15224_,
    new_n15225_, new_n15226_, new_n15227_, new_n15228_, new_n15229_,
    new_n15230_, new_n15231_, new_n15232_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15383_, new_n15384_,
    new_n15385_, new_n15386_, new_n15387_, new_n15388_, new_n15389_,
    new_n15390_, new_n15391_, new_n15392_, new_n15393_, new_n15394_,
    new_n15395_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15403_, new_n15404_,
    new_n15405_, new_n15406_, new_n15407_, new_n15408_, new_n15409_,
    new_n15410_, new_n15411_, new_n15412_, new_n15413_, new_n15414_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15633_, new_n15634_,
    new_n15635_, new_n15636_, new_n15637_, new_n15638_, new_n15639_,
    new_n15640_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15690_, new_n15691_, new_n15692_, new_n15693_, new_n15694_,
    new_n15695_, new_n15696_, new_n15697_, new_n15698_, new_n15699_,
    new_n15700_, new_n15701_, new_n15702_, new_n15703_, new_n15704_,
    new_n15705_, new_n15706_, new_n15707_, new_n15708_, new_n15709_,
    new_n15710_, new_n15711_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15808_, new_n15809_,
    new_n15810_, new_n15811_, new_n15812_, new_n15813_, new_n15814_,
    new_n15815_, new_n15816_, new_n15817_, new_n15818_, new_n15819_,
    new_n15820_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15865_, new_n15866_, new_n15867_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15897_, new_n15898_, new_n15899_,
    new_n15900_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15910_, new_n15911_, new_n15912_, new_n15913_, new_n15914_,
    new_n15915_, new_n15916_, new_n15917_, new_n15918_, new_n15919_,
    new_n15920_, new_n15921_, new_n15922_, new_n15923_, new_n15924_,
    new_n15925_, new_n15926_, new_n15927_, new_n15928_, new_n15929_,
    new_n15930_, new_n15931_, new_n15932_, new_n15933_, new_n15934_,
    new_n15935_, new_n15936_, new_n15937_, new_n15938_, new_n15939_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15945_, new_n15946_, new_n15947_, new_n15948_, new_n15949_,
    new_n15950_, new_n15951_, new_n15952_, new_n15953_, new_n15954_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16001_, new_n16002_, new_n16003_, new_n16004_,
    new_n16005_, new_n16006_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16067_, new_n16068_, new_n16069_,
    new_n16070_, new_n16071_, new_n16072_, new_n16073_, new_n16074_,
    new_n16075_, new_n16076_, new_n16077_, new_n16078_, new_n16079_,
    new_n16080_, new_n16081_, new_n16082_, new_n16083_, new_n16084_,
    new_n16085_, new_n16086_, new_n16087_, new_n16088_, new_n16089_,
    new_n16090_, new_n16091_, new_n16092_, new_n16093_, new_n16094_,
    new_n16095_, new_n16096_, new_n16097_, new_n16098_, new_n16099_,
    new_n16100_, new_n16101_, new_n16102_, new_n16103_, new_n16104_,
    new_n16105_, new_n16106_, new_n16107_, new_n16108_, new_n16109_,
    new_n16110_, new_n16111_, new_n16112_, new_n16113_, new_n16114_,
    new_n16115_, new_n16116_, new_n16117_, new_n16118_, new_n16119_,
    new_n16120_, new_n16121_, new_n16122_, new_n16123_, new_n16124_,
    new_n16125_, new_n16126_, new_n16127_, new_n16128_, new_n16129_,
    new_n16130_, new_n16131_, new_n16132_, new_n16133_, new_n16134_,
    new_n16135_, new_n16136_, new_n16137_, new_n16138_, new_n16139_,
    new_n16140_, new_n16141_, new_n16142_, new_n16143_, new_n16144_,
    new_n16145_, new_n16146_, new_n16147_, new_n16148_, new_n16149_,
    new_n16150_, new_n16151_, new_n16152_, new_n16153_, new_n16154_,
    new_n16155_, new_n16156_, new_n16157_, new_n16158_, new_n16159_,
    new_n16160_, new_n16161_, new_n16162_, new_n16163_, new_n16164_,
    new_n16165_, new_n16166_, new_n16167_, new_n16168_, new_n16169_,
    new_n16170_, new_n16171_, new_n16172_, new_n16173_, new_n16174_,
    new_n16175_, new_n16176_, new_n16177_, new_n16178_, new_n16179_,
    new_n16180_, new_n16181_, new_n16182_, new_n16183_, new_n16184_,
    new_n16185_, new_n16186_, new_n16187_, new_n16188_, new_n16189_,
    new_n16190_, new_n16191_, new_n16192_, new_n16193_, new_n16194_,
    new_n16195_, new_n16196_, new_n16197_, new_n16198_, new_n16199_,
    new_n16200_, new_n16201_, new_n16202_, new_n16203_, new_n16204_,
    new_n16205_, new_n16206_, new_n16207_, new_n16208_, new_n16209_,
    new_n16210_, new_n16211_, new_n16212_, new_n16213_, new_n16214_,
    new_n16215_, new_n16216_, new_n16217_, new_n16218_, new_n16219_,
    new_n16220_, new_n16221_, new_n16222_, new_n16223_, new_n16224_,
    new_n16225_, new_n16226_, new_n16227_, new_n16228_, new_n16229_,
    new_n16230_, new_n16231_, new_n16232_, new_n16233_, new_n16234_,
    new_n16235_, new_n16236_, new_n16237_, new_n16238_, new_n16239_,
    new_n16240_, new_n16241_, new_n16242_, new_n16243_, new_n16244_,
    new_n16245_, new_n16246_, new_n16247_, new_n16248_, new_n16249_,
    new_n16250_, new_n16251_, new_n16252_, new_n16253_, new_n16254_,
    new_n16255_, new_n16256_, new_n16257_, new_n16258_, new_n16259_,
    new_n16260_, new_n16261_, new_n16262_, new_n16263_, new_n16264_,
    new_n16265_, new_n16266_, new_n16267_, new_n16268_, new_n16269_,
    new_n16270_, new_n16271_, new_n16272_, new_n16273_, new_n16274_,
    new_n16275_, new_n16276_, new_n16277_, new_n16278_, new_n16279_,
    new_n16280_, new_n16281_, new_n16282_, new_n16283_, new_n16284_,
    new_n16285_, new_n16286_, new_n16287_, new_n16288_, new_n16289_,
    new_n16290_, new_n16291_, new_n16292_, new_n16293_, new_n16294_,
    new_n16295_, new_n16296_, new_n16297_, new_n16298_, new_n16299_,
    new_n16300_, new_n16301_, new_n16302_, new_n16303_, new_n16304_,
    new_n16305_, new_n16306_, new_n16307_, new_n16308_, new_n16309_,
    new_n16310_, new_n16311_, new_n16312_, new_n16313_, new_n16314_,
    new_n16315_, new_n16316_, new_n16317_, new_n16318_, new_n16319_,
    new_n16320_, new_n16321_, new_n16322_, new_n16323_, new_n16324_,
    new_n16325_, new_n16326_, new_n16327_, new_n16328_, new_n16329_,
    new_n16330_, new_n16331_, new_n16332_, new_n16333_, new_n16334_,
    new_n16335_, new_n16336_, new_n16337_, new_n16338_, new_n16339_,
    new_n16340_, new_n16341_, new_n16342_, new_n16343_, new_n16344_,
    new_n16345_, new_n16346_, new_n16347_, new_n16348_, new_n16349_,
    new_n16350_, new_n16351_, new_n16352_, new_n16353_, new_n16354_,
    new_n16355_, new_n16356_, new_n16357_, new_n16358_, new_n16359_,
    new_n16360_, new_n16361_, new_n16362_, new_n16363_, new_n16364_,
    new_n16365_, new_n16366_, new_n16367_, new_n16368_, new_n16369_,
    new_n16370_, new_n16371_, new_n16372_, new_n16373_, new_n16374_,
    new_n16375_, new_n16376_, new_n16377_, new_n16378_, new_n16379_,
    new_n16380_, new_n16381_, new_n16382_, new_n16383_, new_n16384_,
    new_n16385_, new_n16386_, new_n16387_, new_n16388_, new_n16389_,
    new_n16390_, new_n16391_, new_n16392_, new_n16393_, new_n16394_,
    new_n16395_, new_n16396_, new_n16397_, new_n16398_, new_n16399_,
    new_n16400_, new_n16401_, new_n16402_, new_n16403_, new_n16404_,
    new_n16405_, new_n16406_, new_n16407_, new_n16408_, new_n16409_,
    new_n16410_, new_n16411_, new_n16412_, new_n16413_, new_n16414_,
    new_n16415_, new_n16416_, new_n16417_, new_n16418_, new_n16419_,
    new_n16420_, new_n16421_, new_n16422_, new_n16423_, new_n16424_,
    new_n16425_, new_n16426_, new_n16427_, new_n16428_, new_n16429_,
    new_n16430_, new_n16431_, new_n16432_, new_n16433_, new_n16434_,
    new_n16435_, new_n16436_, new_n16437_, new_n16438_, new_n16439_,
    new_n16440_, new_n16441_, new_n16442_, new_n16443_, new_n16444_,
    new_n16445_, new_n16446_, new_n16447_, new_n16448_, new_n16449_,
    new_n16450_, new_n16451_, new_n16452_, new_n16453_, new_n16454_,
    new_n16455_, new_n16456_, new_n16457_, new_n16458_, new_n16459_,
    new_n16460_, new_n16461_, new_n16462_, new_n16463_, new_n16464_,
    new_n16465_, new_n16466_, new_n16467_, new_n16468_, new_n16469_,
    new_n16470_, new_n16471_, new_n16472_, new_n16473_, new_n16474_,
    new_n16475_, new_n16476_, new_n16477_, new_n16478_, new_n16479_,
    new_n16480_, new_n16481_, new_n16482_, new_n16483_, new_n16484_,
    new_n16485_, new_n16486_, new_n16487_, new_n16488_, new_n16489_,
    new_n16490_, new_n16491_, new_n16492_, new_n16493_, new_n16494_,
    new_n16495_, new_n16496_, new_n16497_, new_n16498_, new_n16499_,
    new_n16500_, new_n16501_, new_n16502_, new_n16503_, new_n16504_,
    new_n16505_, new_n16506_, new_n16507_, new_n16508_, new_n16509_,
    new_n16510_, new_n16511_, new_n16512_, new_n16513_, new_n16514_,
    new_n16515_, new_n16516_, new_n16517_, new_n16518_, new_n16519_,
    new_n16520_, new_n16521_, new_n16522_, new_n16523_, new_n16524_,
    new_n16525_, new_n16526_, new_n16527_, new_n16528_, new_n16529_,
    new_n16530_, new_n16531_, new_n16532_, new_n16533_, new_n16534_,
    new_n16535_, new_n16536_, new_n16537_, new_n16538_, new_n16539_,
    new_n16540_, new_n16541_, new_n16542_, new_n16543_, new_n16544_,
    new_n16545_, new_n16546_, new_n16547_, new_n16548_, new_n16549_,
    new_n16550_, new_n16551_, new_n16552_, new_n16553_, new_n16554_,
    new_n16555_, new_n16556_, new_n16557_, new_n16558_, new_n16559_,
    new_n16560_, new_n16561_, new_n16562_, new_n16563_, new_n16564_,
    new_n16565_, new_n16566_, new_n16567_, new_n16568_, new_n16569_,
    new_n16570_, new_n16571_, new_n16572_, new_n16573_, new_n16574_,
    new_n16575_, new_n16576_, new_n16577_, new_n16578_, new_n16579_,
    new_n16580_, new_n16581_, new_n16582_, new_n16583_, new_n16584_,
    new_n16585_, new_n16586_, new_n16587_, new_n16588_, new_n16589_,
    new_n16590_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16619_,
    new_n16620_, new_n16621_, new_n16622_, new_n16623_, new_n16624_,
    new_n16625_, new_n16626_, new_n16627_, new_n16628_, new_n16629_,
    new_n16630_, new_n16631_, new_n16632_, new_n16633_, new_n16634_,
    new_n16635_, new_n16636_, new_n16637_, new_n16638_, new_n16639_,
    new_n16640_, new_n16641_, new_n16642_, new_n16643_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16666_, new_n16667_, new_n16668_, new_n16669_,
    new_n16670_, new_n16671_, new_n16672_, new_n16673_, new_n16674_,
    new_n16675_, new_n16676_, new_n16677_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16683_, new_n16684_,
    new_n16685_, new_n16686_, new_n16687_, new_n16688_, new_n16689_,
    new_n16690_, new_n16691_, new_n16692_, new_n16693_, new_n16694_,
    new_n16695_, new_n16696_, new_n16697_, new_n16698_, new_n16699_,
    new_n16700_, new_n16701_, new_n16702_, new_n16703_, new_n16704_,
    new_n16705_, new_n16706_, new_n16707_, new_n16708_, new_n16709_,
    new_n16710_, new_n16711_, new_n16712_, new_n16713_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16727_, new_n16728_, new_n16729_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16736_, new_n16737_, new_n16738_, new_n16739_,
    new_n16740_, new_n16741_, new_n16742_, new_n16743_, new_n16744_,
    new_n16745_, new_n16746_, new_n16747_, new_n16748_, new_n16749_,
    new_n16750_, new_n16751_, new_n16752_, new_n16753_, new_n16754_,
    new_n16755_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16765_, new_n16766_, new_n16767_, new_n16768_, new_n16769_,
    new_n16770_, new_n16771_, new_n16772_, new_n16773_, new_n16774_,
    new_n16775_, new_n16776_, new_n16777_, new_n16778_, new_n16779_,
    new_n16780_, new_n16781_, new_n16782_, new_n16783_, new_n16784_,
    new_n16785_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16820_, new_n16821_, new_n16822_, new_n16823_, new_n16824_,
    new_n16825_, new_n16826_, new_n16827_, new_n16828_, new_n16829_,
    new_n16830_, new_n16831_, new_n16832_, new_n16833_, new_n16834_,
    new_n16835_, new_n16836_, new_n16837_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16852_, new_n16853_, new_n16854_,
    new_n16855_, new_n16856_, new_n16857_, new_n16858_, new_n16859_,
    new_n16860_, new_n16861_, new_n16862_, new_n16863_, new_n16864_,
    new_n16865_, new_n16866_, new_n16867_, new_n16868_, new_n16869_,
    new_n16870_, new_n16871_, new_n16872_, new_n16873_, new_n16874_,
    new_n16875_, new_n16876_, new_n16877_, new_n16878_, new_n16879_,
    new_n16880_, new_n16881_, new_n16882_, new_n16883_, new_n16884_,
    new_n16885_, new_n16886_, new_n16887_, new_n16888_, new_n16889_,
    new_n16890_, new_n16891_, new_n16892_, new_n16893_, new_n16894_,
    new_n16895_, new_n16896_, new_n16897_, new_n16898_, new_n16899_,
    new_n16900_, new_n16901_, new_n16902_, new_n16903_, new_n16904_,
    new_n16905_, new_n16906_, new_n16907_, new_n16908_, new_n16909_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16914_,
    new_n16915_, new_n16916_, new_n16917_, new_n16918_, new_n16919_,
    new_n16920_, new_n16921_, new_n16922_, new_n16923_, new_n16924_,
    new_n16925_, new_n16926_, new_n16927_, new_n16928_, new_n16929_,
    new_n16930_, new_n16931_, new_n16932_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16938_, new_n16939_,
    new_n16940_, new_n16941_, new_n16942_, new_n16943_, new_n16944_,
    new_n16945_, new_n16946_, new_n16947_, new_n16948_, new_n16949_,
    new_n16950_, new_n16951_, new_n16952_, new_n16953_, new_n16954_,
    new_n16955_, new_n16956_, new_n16957_, new_n16958_, new_n16959_,
    new_n16960_, new_n16961_, new_n16962_, new_n16963_, new_n16964_,
    new_n16965_, new_n16966_, new_n16967_, new_n16968_, new_n16969_,
    new_n16970_, new_n16971_, new_n16972_, new_n16973_, new_n16974_,
    new_n16975_, new_n16976_, new_n16977_, new_n16978_, new_n16979_,
    new_n16980_, new_n16981_, new_n16982_, new_n16983_, new_n16984_,
    new_n16985_, new_n16986_, new_n16987_, new_n16988_, new_n16989_,
    new_n16990_, new_n16991_, new_n16992_, new_n16993_, new_n16994_,
    new_n16995_, new_n16996_, new_n16997_, new_n16998_, new_n16999_,
    new_n17000_, new_n17001_, new_n17002_, new_n17003_, new_n17004_,
    new_n17005_, new_n17006_, new_n17007_, new_n17008_, new_n17009_,
    new_n17010_, new_n17011_, new_n17012_, new_n17013_, new_n17014_,
    new_n17015_, new_n17016_, new_n17017_, new_n17018_, new_n17019_,
    new_n17020_, new_n17021_, new_n17022_, new_n17023_, new_n17024_,
    new_n17025_, new_n17026_, new_n17027_, new_n17028_, new_n17029_,
    new_n17030_, new_n17031_, new_n17032_, new_n17033_, new_n17034_,
    new_n17035_, new_n17036_, new_n17037_, new_n17038_, new_n17039_,
    new_n17040_, new_n17041_, new_n17042_, new_n17043_, new_n17044_,
    new_n17045_, new_n17046_, new_n17047_, new_n17048_, new_n17049_,
    new_n17050_, new_n17051_, new_n17052_, new_n17053_, new_n17054_,
    new_n17055_, new_n17056_, new_n17057_, new_n17058_, new_n17059_,
    new_n17060_, new_n17061_, new_n17062_, new_n17063_, new_n17064_,
    new_n17065_, new_n17066_, new_n17067_, new_n17068_, new_n17069_,
    new_n17070_, new_n17071_, new_n17072_, new_n17073_, new_n17074_,
    new_n17075_, new_n17076_, new_n17077_, new_n17078_, new_n17079_,
    new_n17080_, new_n17081_, new_n17082_, new_n17083_, new_n17084_,
    new_n17085_, new_n17086_, new_n17087_, new_n17088_, new_n17089_,
    new_n17090_, new_n17091_, new_n17092_, new_n17093_, new_n17094_,
    new_n17095_, new_n17096_, new_n17097_, new_n17098_, new_n17099_,
    new_n17100_, new_n17101_, new_n17102_, new_n17103_, new_n17104_,
    new_n17105_, new_n17106_, new_n17107_, new_n17108_, new_n17109_,
    new_n17110_, new_n17111_, new_n17112_, new_n17113_, new_n17114_,
    new_n17115_, new_n17116_, new_n17117_, new_n17118_, new_n17119_,
    new_n17120_, new_n17121_, new_n17122_, new_n17123_, new_n17124_,
    new_n17125_, new_n17126_, new_n17127_, new_n17128_, new_n17129_,
    new_n17130_, new_n17131_, new_n17132_, new_n17133_, new_n17134_,
    new_n17135_, new_n17136_, new_n17137_, new_n17138_, new_n17139_,
    new_n17140_, new_n17141_, new_n17142_, new_n17143_, new_n17144_,
    new_n17145_, new_n17146_, new_n17147_, new_n17148_, new_n17149_,
    new_n17150_, new_n17151_, new_n17152_, new_n17153_, new_n17154_,
    new_n17155_, new_n17156_, new_n17157_, new_n17158_, new_n17159_,
    new_n17160_, new_n17161_, new_n17162_, new_n17163_, new_n17164_,
    new_n17165_, new_n17166_, new_n17167_, new_n17168_, new_n17169_,
    new_n17170_, new_n17171_, new_n17172_, new_n17173_, new_n17174_,
    new_n17175_, new_n17176_, new_n17177_, new_n17178_, new_n17179_,
    new_n17180_, new_n17181_, new_n17182_, new_n17183_, new_n17184_,
    new_n17185_, new_n17186_, new_n17187_, new_n17188_, new_n17189_,
    new_n17190_, new_n17191_, new_n17192_, new_n17193_, new_n17194_,
    new_n17195_, new_n17196_, new_n17197_, new_n17198_, new_n17199_,
    new_n17200_, new_n17201_, new_n17202_, new_n17203_, new_n17204_,
    new_n17205_, new_n17206_, new_n17207_, new_n17208_, new_n17209_,
    new_n17210_, new_n17211_, new_n17212_, new_n17213_, new_n17214_,
    new_n17215_, new_n17216_, new_n17217_, new_n17218_, new_n17219_,
    new_n17220_, new_n17221_, new_n17222_, new_n17223_, new_n17224_,
    new_n17225_, new_n17226_, new_n17227_, new_n17228_, new_n17229_,
    new_n17230_, new_n17231_, new_n17232_, new_n17233_, new_n17234_,
    new_n17235_, new_n17236_, new_n17237_, new_n17238_, new_n17239_,
    new_n17240_, new_n17241_, new_n17242_, new_n17243_, new_n17244_,
    new_n17245_, new_n17246_, new_n17247_, new_n17248_, new_n17249_,
    new_n17250_, new_n17251_, new_n17252_, new_n17253_, new_n17254_,
    new_n17255_, new_n17256_, new_n17257_, new_n17258_, new_n17259_,
    new_n17260_, new_n17261_, new_n17262_, new_n17263_, new_n17264_,
    new_n17265_, new_n17266_, new_n17267_, new_n17268_, new_n17269_,
    new_n17270_, new_n17271_, new_n17272_, new_n17273_, new_n17274_,
    new_n17275_, new_n17276_, new_n17277_, new_n17278_, new_n17279_,
    new_n17280_, new_n17281_, new_n17282_, new_n17283_, new_n17284_,
    new_n17285_, new_n17286_, new_n17287_, new_n17288_, new_n17289_,
    new_n17290_, new_n17291_, new_n17292_, new_n17293_, new_n17294_,
    new_n17295_, new_n17296_, new_n17297_, new_n17298_, new_n17299_,
    new_n17300_, new_n17301_, new_n17302_, new_n17303_, new_n17304_,
    new_n17305_, new_n17306_, new_n17307_, new_n17308_, new_n17309_,
    new_n17310_, new_n17311_, new_n17312_, new_n17313_, new_n17314_,
    new_n17315_, new_n17316_, new_n17317_, new_n17318_, new_n17319_,
    new_n17320_, new_n17321_, new_n17322_, new_n17323_, new_n17324_,
    new_n17325_, new_n17326_, new_n17327_, new_n17328_, new_n17329_,
    new_n17330_, new_n17331_, new_n17332_, new_n17333_, new_n17334_,
    new_n17335_, new_n17336_, new_n17337_, new_n17338_, new_n17339_,
    new_n17340_, new_n17341_, new_n17342_, new_n17343_, new_n17344_,
    new_n17345_, new_n17346_, new_n17347_, new_n17348_, new_n17349_,
    new_n17350_, new_n17351_, new_n17352_, new_n17353_, new_n17354_,
    new_n17355_, new_n17356_, new_n17357_, new_n17358_, new_n17359_,
    new_n17360_, new_n17361_, new_n17362_, new_n17363_, new_n17364_,
    new_n17365_, new_n17366_, new_n17367_, new_n17368_, new_n17369_,
    new_n17370_, new_n17371_, new_n17372_, new_n17373_, new_n17374_,
    new_n17375_, new_n17376_, new_n17377_, new_n17378_, new_n17379_,
    new_n17380_, new_n17381_, new_n17382_, new_n17383_, new_n17384_,
    new_n17385_, new_n17386_, new_n17387_, new_n17388_, new_n17389_,
    new_n17390_, new_n17391_, new_n17392_, new_n17393_, new_n17394_,
    new_n17395_, new_n17396_, new_n17397_, new_n17398_, new_n17399_,
    new_n17400_, new_n17401_, new_n17402_, new_n17403_, new_n17404_,
    new_n17405_, new_n17406_, new_n17407_, new_n17408_, new_n17409_,
    new_n17410_, new_n17411_, new_n17412_, new_n17413_, new_n17414_,
    new_n17415_, new_n17416_, new_n17417_, new_n17418_, new_n17419_,
    new_n17420_, new_n17421_, new_n17422_, new_n17423_, new_n17424_,
    new_n17425_, new_n17426_, new_n17427_, new_n17428_, new_n17429_,
    new_n17430_, new_n17431_, new_n17432_, new_n17433_, new_n17434_,
    new_n17435_, new_n17436_, new_n17437_, new_n17438_, new_n17439_,
    new_n17440_, new_n17441_, new_n17442_, new_n17443_, new_n17444_,
    new_n17445_, new_n17446_, new_n17447_, new_n17448_, new_n17449_,
    new_n17450_, new_n17451_, new_n17452_, new_n17453_, new_n17454_,
    new_n17455_, new_n17456_, new_n17457_, new_n17458_, new_n17459_,
    new_n17460_, new_n17461_, new_n17462_, new_n17463_, new_n17464_,
    new_n17465_, new_n17466_, new_n17467_, new_n17468_, new_n17469_,
    new_n17470_, new_n17471_, new_n17472_, new_n17473_, new_n17474_,
    new_n17475_, new_n17476_, new_n17477_, new_n17478_, new_n17479_,
    new_n17480_, new_n17481_, new_n17482_, new_n17483_, new_n17484_,
    new_n17485_, new_n17486_, new_n17487_, new_n17488_, new_n17489_,
    new_n17490_, new_n17491_, new_n17492_, new_n17493_, new_n17494_,
    new_n17495_, new_n17496_, new_n17497_, new_n17498_, new_n17499_,
    new_n17500_, new_n17501_, new_n17502_, new_n17503_, new_n17504_,
    new_n17505_, new_n17506_, new_n17507_, new_n17508_, new_n17509_,
    new_n17510_, new_n17511_, new_n17512_, new_n17513_, new_n17514_,
    new_n17515_, new_n17516_, new_n17517_, new_n17518_, new_n17519_,
    new_n17520_, new_n17521_, new_n17522_, new_n17523_, new_n17524_,
    new_n17525_, new_n17526_, new_n17527_, new_n17528_, new_n17529_,
    new_n17530_, new_n17531_, new_n17532_, new_n17533_, new_n17534_,
    new_n17535_, new_n17536_, new_n17537_, new_n17538_, new_n17539_,
    new_n17540_, new_n17541_, new_n17542_, new_n17543_, new_n17544_,
    new_n17545_, new_n17546_, new_n17547_, new_n17548_, new_n17549_,
    new_n17550_, new_n17551_, new_n17552_, new_n17553_, new_n17554_,
    new_n17555_, new_n17556_, new_n17557_, new_n17558_, new_n17559_,
    new_n17560_, new_n17561_, new_n17562_, new_n17563_, new_n17564_,
    new_n17565_, new_n17566_, new_n17567_, new_n17568_, new_n17569_,
    new_n17570_, new_n17571_, new_n17572_, new_n17573_, new_n17574_,
    new_n17575_, new_n17576_, new_n17577_, new_n17578_, new_n17579_,
    new_n17580_, new_n17581_, new_n17582_, new_n17583_, new_n17584_,
    new_n17585_, new_n17586_, new_n17587_, new_n17588_, new_n17589_,
    new_n17590_, new_n17591_, new_n17592_, new_n17593_, new_n17594_,
    new_n17595_, new_n17596_, new_n17597_, new_n17598_, new_n17599_,
    new_n17600_, new_n17601_, new_n17602_, new_n17603_, new_n17604_,
    new_n17605_, new_n17606_, new_n17607_, new_n17608_, new_n17609_,
    new_n17610_, new_n17611_, new_n17612_, new_n17613_, new_n17614_,
    new_n17615_, new_n17616_, new_n17617_, new_n17618_, new_n17619_,
    new_n17620_, new_n17621_, new_n17622_, new_n17623_, new_n17624_,
    new_n17625_, new_n17626_, new_n17627_, new_n17628_, new_n17629_,
    new_n17630_, new_n17631_, new_n17632_, new_n17633_, new_n17634_,
    new_n17635_, new_n17636_, new_n17637_, new_n17638_, new_n17639_,
    new_n17640_, new_n17641_, new_n17642_, new_n17643_, new_n17644_,
    new_n17645_, new_n17646_, new_n17647_, new_n17648_, new_n17649_,
    new_n17650_, new_n17651_, new_n17652_, new_n17653_, new_n17654_,
    new_n17655_, new_n17656_, new_n17657_, new_n17658_, new_n17659_,
    new_n17660_, new_n17661_, new_n17662_, new_n17663_, new_n17664_,
    new_n17665_, new_n17666_, new_n17667_, new_n17668_, new_n17669_,
    new_n17670_, new_n17671_, new_n17672_, new_n17673_, new_n17674_,
    new_n17675_, new_n17676_, new_n17677_, new_n17678_, new_n17679_,
    new_n17680_, new_n17681_, new_n17682_, new_n17683_, new_n17684_,
    new_n17685_, new_n17686_, new_n17687_, new_n17688_, new_n17689_,
    new_n17690_, new_n17691_, new_n17692_, new_n17693_, new_n17694_,
    new_n17695_, new_n17696_, new_n17697_, new_n17698_, new_n17699_,
    new_n17700_, new_n17701_, new_n17702_, new_n17703_, new_n17704_,
    new_n17705_, new_n17706_, new_n17707_, new_n17708_, new_n17709_,
    new_n17710_, new_n17711_, new_n17712_, new_n17713_, new_n17714_,
    new_n17715_, new_n17716_, new_n17717_, new_n17718_, new_n17719_,
    new_n17720_, new_n17721_, new_n17722_, new_n17723_, new_n17724_,
    new_n17725_, new_n17726_, new_n17727_, new_n17728_, new_n17729_,
    new_n17730_, new_n17731_, new_n17732_, new_n17733_, new_n17734_,
    new_n17735_, new_n17736_, new_n17737_, new_n17738_, new_n17739_,
    new_n17740_, new_n17741_, new_n17742_, new_n17743_, new_n17744_,
    new_n17745_, new_n17746_, new_n17747_, new_n17748_, new_n17749_,
    new_n17750_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17762_, new_n17763_, new_n17764_,
    new_n17765_, new_n17766_, new_n17767_, new_n17768_, new_n17769_,
    new_n17770_, new_n17771_, new_n17772_, new_n17773_, new_n17774_,
    new_n17775_, new_n17776_, new_n17777_, new_n17778_, new_n17779_,
    new_n17780_, new_n17781_, new_n17782_, new_n17783_, new_n17784_,
    new_n17785_, new_n17786_, new_n17787_, new_n17788_, new_n17789_,
    new_n17790_, new_n17791_, new_n17792_, new_n17793_, new_n17794_,
    new_n17795_, new_n17796_, new_n17797_, new_n17798_, new_n17799_,
    new_n17800_, new_n17801_, new_n17802_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17810_, new_n17811_, new_n17812_, new_n17813_, new_n17814_,
    new_n17815_, new_n17816_, new_n17817_, new_n17818_, new_n17819_,
    new_n17820_, new_n17821_, new_n17822_, new_n17823_, new_n17824_,
    new_n17825_, new_n17826_, new_n17827_, new_n17828_, new_n17829_,
    new_n17830_, new_n17831_, new_n17832_, new_n17833_, new_n17834_,
    new_n17835_, new_n17836_, new_n17837_, new_n17838_, new_n17839_,
    new_n17840_, new_n17841_, new_n17842_, new_n17843_, new_n17844_,
    new_n17845_, new_n17846_, new_n17847_, new_n17848_, new_n17849_,
    new_n17850_, new_n17851_, new_n17852_, new_n17853_, new_n17854_,
    new_n17855_, new_n17856_, new_n17857_, new_n17858_, new_n17859_,
    new_n17860_, new_n17861_, new_n17862_, new_n17863_, new_n17864_,
    new_n17865_, new_n17866_, new_n17867_, new_n17868_, new_n17869_,
    new_n17870_, new_n17871_, new_n17872_, new_n17873_, new_n17874_,
    new_n17875_, new_n17876_, new_n17877_, new_n17878_, new_n17879_,
    new_n17880_, new_n17881_, new_n17882_, new_n17883_, new_n17884_,
    new_n17885_, new_n17886_, new_n17887_, new_n17888_, new_n17889_,
    new_n17890_, new_n17891_, new_n17892_, new_n17893_, new_n17894_,
    new_n17895_, new_n17896_, new_n17897_, new_n17898_, new_n17899_,
    new_n17900_, new_n17901_, new_n17902_, new_n17903_, new_n17904_,
    new_n17905_, new_n17906_, new_n17907_, new_n17908_, new_n17909_,
    new_n17910_, new_n17911_, new_n17912_, new_n17913_, new_n17914_,
    new_n17915_, new_n17916_, new_n17917_, new_n17918_, new_n17919_,
    new_n17920_, new_n17921_, new_n17922_, new_n17923_, new_n17924_,
    new_n17925_, new_n17926_, new_n17927_, new_n17928_, new_n17929_,
    new_n17930_, new_n17931_, new_n17932_, new_n17933_, new_n17934_,
    new_n17935_, new_n17936_, new_n17937_, new_n17938_, new_n17939_,
    new_n17940_, new_n17941_, new_n17942_, new_n17943_, new_n17944_,
    new_n17945_, new_n17946_, new_n17947_, new_n17948_, new_n17949_,
    new_n17950_, new_n17951_, new_n17952_, new_n17953_, new_n17954_,
    new_n17955_, new_n17956_, new_n17957_, new_n17958_, new_n17959_,
    new_n17960_, new_n17961_, new_n17962_, new_n17963_, new_n17964_,
    new_n17965_, new_n17966_, new_n17967_, new_n17968_, new_n17969_,
    new_n17970_, new_n17971_, new_n17972_, new_n17973_, new_n17974_,
    new_n17975_, new_n17976_, new_n17977_, new_n17978_, new_n17979_,
    new_n17980_, new_n17981_, new_n17982_, new_n17983_, new_n17984_,
    new_n17985_, new_n17986_, new_n17987_, new_n17988_, new_n17989_,
    new_n17990_, new_n17991_, new_n17992_, new_n17993_, new_n17994_,
    new_n17995_, new_n17996_, new_n17997_, new_n17998_, new_n17999_,
    new_n18000_, new_n18001_, new_n18002_, new_n18003_, new_n18004_,
    new_n18005_, new_n18006_, new_n18007_, new_n18008_, new_n18009_,
    new_n18010_, new_n18011_, new_n18012_, new_n18013_, new_n18014_,
    new_n18015_, new_n18016_, new_n18017_, new_n18018_, new_n18019_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18025_, new_n18026_, new_n18027_, new_n18028_, new_n18029_,
    new_n18030_, new_n18031_, new_n18032_, new_n18033_, new_n18034_,
    new_n18035_, new_n18036_, new_n18037_, new_n18038_, new_n18039_,
    new_n18040_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18108_, new_n18109_,
    new_n18110_, new_n18111_, new_n18112_, new_n18113_, new_n18114_,
    new_n18115_, new_n18116_, new_n18117_, new_n18118_, new_n18119_,
    new_n18120_, new_n18121_, new_n18122_, new_n18123_, new_n18124_,
    new_n18125_, new_n18126_, new_n18127_, new_n18128_, new_n18129_,
    new_n18130_, new_n18131_, new_n18132_, new_n18133_, new_n18134_,
    new_n18135_, new_n18136_, new_n18137_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18169_,
    new_n18170_, new_n18171_, new_n18172_, new_n18173_, new_n18174_,
    new_n18175_, new_n18176_, new_n18177_, new_n18178_, new_n18179_,
    new_n18180_, new_n18181_, new_n18182_, new_n18183_, new_n18184_,
    new_n18185_, new_n18186_, new_n18187_, new_n18188_, new_n18189_,
    new_n18190_, new_n18191_, new_n18192_, new_n18193_, new_n18194_,
    new_n18195_, new_n18196_, new_n18197_, new_n18198_, new_n18199_,
    new_n18200_, new_n18201_, new_n18202_, new_n18203_, new_n18204_,
    new_n18205_, new_n18206_, new_n18207_, new_n18208_, new_n18209_,
    new_n18210_, new_n18211_, new_n18212_, new_n18213_, new_n18214_,
    new_n18215_, new_n18216_, new_n18217_, new_n18218_, new_n18219_,
    new_n18220_, new_n18221_, new_n18222_, new_n18223_, new_n18224_,
    new_n18225_, new_n18226_, new_n18227_, new_n18228_, new_n18229_,
    new_n18230_, new_n18231_, new_n18232_, new_n18233_, new_n18234_,
    new_n18235_, new_n18236_, new_n18237_, new_n18238_, new_n18239_,
    new_n18240_, new_n18241_, new_n18242_, new_n18243_, new_n18244_,
    new_n18245_, new_n18246_, new_n18247_, new_n18248_, new_n18249_,
    new_n18250_, new_n18251_, new_n18252_, new_n18253_, new_n18254_,
    new_n18255_, new_n18256_, new_n18257_, new_n18258_, new_n18259_,
    new_n18260_, new_n18261_, new_n18262_, new_n18263_, new_n18264_,
    new_n18265_, new_n18266_, new_n18267_, new_n18268_, new_n18269_,
    new_n18270_, new_n18271_, new_n18272_, new_n18273_, new_n18274_,
    new_n18275_, new_n18276_, new_n18277_, new_n18278_, new_n18279_,
    new_n18280_, new_n18281_, new_n18282_, new_n18283_, new_n18284_,
    new_n18285_, new_n18286_, new_n18287_, new_n18288_, new_n18289_,
    new_n18290_, new_n18291_, new_n18292_, new_n18293_, new_n18294_,
    new_n18295_, new_n18296_, new_n18297_, new_n18298_, new_n18299_,
    new_n18300_, new_n18301_, new_n18302_, new_n18303_, new_n18304_,
    new_n18305_, new_n18306_, new_n18307_, new_n18308_, new_n18309_,
    new_n18310_, new_n18311_, new_n18312_, new_n18313_, new_n18314_,
    new_n18315_, new_n18316_, new_n18317_, new_n18318_, new_n18319_,
    new_n18320_, new_n18321_, new_n18322_, new_n18323_, new_n18324_,
    new_n18325_, new_n18326_, new_n18327_, new_n18328_, new_n18329_,
    new_n18330_, new_n18331_, new_n18332_, new_n18333_, new_n18334_,
    new_n18335_, new_n18336_, new_n18337_, new_n18338_, new_n18339_,
    new_n18340_, new_n18341_, new_n18342_, new_n18343_, new_n18344_,
    new_n18345_, new_n18346_, new_n18347_, new_n18348_, new_n18349_,
    new_n18350_, new_n18351_, new_n18352_, new_n18353_, new_n18354_,
    new_n18355_, new_n18356_, new_n18357_, new_n18358_, new_n18359_,
    new_n18360_, new_n18361_, new_n18362_, new_n18363_, new_n18364_,
    new_n18365_, new_n18366_, new_n18367_, new_n18368_, new_n18369_,
    new_n18370_, new_n18371_, new_n18372_, new_n18373_, new_n18374_,
    new_n18375_, new_n18376_, new_n18377_, new_n18378_, new_n18379_,
    new_n18380_, new_n18381_, new_n18382_, new_n18383_, new_n18384_,
    new_n18385_, new_n18386_, new_n18387_, new_n18388_, new_n18389_,
    new_n18390_, new_n18391_, new_n18392_, new_n18393_, new_n18394_,
    new_n18395_, new_n18396_, new_n18397_, new_n18398_, new_n18399_,
    new_n18400_, new_n18401_, new_n18402_, new_n18403_, new_n18404_,
    new_n18405_, new_n18406_, new_n18407_, new_n18408_, new_n18409_,
    new_n18410_, new_n18411_, new_n18412_, new_n18413_, new_n18414_,
    new_n18415_, new_n18416_, new_n18417_, new_n18418_, new_n18419_,
    new_n18420_, new_n18421_, new_n18422_, new_n18423_, new_n18424_,
    new_n18425_, new_n18426_, new_n18427_, new_n18428_, new_n18429_,
    new_n18430_, new_n18431_, new_n18432_, new_n18433_, new_n18434_,
    new_n18435_, new_n18436_, new_n18437_, new_n18438_, new_n18439_,
    new_n18440_, new_n18441_, new_n18442_, new_n18443_, new_n18444_,
    new_n18445_, new_n18446_, new_n18447_, new_n18448_, new_n18449_,
    new_n18450_, new_n18451_, new_n18452_, new_n18453_, new_n18454_,
    new_n18455_, new_n18456_, new_n18457_, new_n18458_, new_n18459_,
    new_n18460_, new_n18461_, new_n18462_, new_n18463_, new_n18464_,
    new_n18465_, new_n18466_, new_n18467_, new_n18468_, new_n18469_,
    new_n18470_, new_n18471_, new_n18472_, new_n18473_, new_n18474_,
    new_n18475_, new_n18476_, new_n18477_, new_n18478_, new_n18479_,
    new_n18480_, new_n18481_, new_n18482_, new_n18483_, new_n18484_,
    new_n18485_, new_n18486_, new_n18487_, new_n18488_, new_n18489_,
    new_n18490_, new_n18491_, new_n18492_, new_n18493_, new_n18494_,
    new_n18495_, new_n18496_, new_n18497_, new_n18498_, new_n18499_,
    new_n18500_, new_n18501_, new_n18502_, new_n18503_, new_n18504_,
    new_n18505_, new_n18506_, new_n18507_, new_n18508_, new_n18509_,
    new_n18510_, new_n18511_, new_n18512_, new_n18513_, new_n18514_,
    new_n18515_, new_n18516_, new_n18517_, new_n18518_, new_n18519_,
    new_n18520_, new_n18521_, new_n18522_, new_n18523_, new_n18524_,
    new_n18525_, new_n18526_, new_n18527_, new_n18528_, new_n18529_,
    new_n18530_, new_n18531_, new_n18532_, new_n18533_, new_n18534_,
    new_n18535_, new_n18536_, new_n18537_, new_n18538_, new_n18539_,
    new_n18540_, new_n18541_, new_n18542_, new_n18543_, new_n18544_,
    new_n18545_, new_n18546_, new_n18547_, new_n18548_, new_n18549_,
    new_n18550_, new_n18551_, new_n18552_, new_n18553_, new_n18554_,
    new_n18555_, new_n18556_, new_n18557_, new_n18558_, new_n18559_,
    new_n18560_, new_n18561_, new_n18562_, new_n18563_, new_n18564_,
    new_n18565_, new_n18566_, new_n18567_, new_n18568_, new_n18569_,
    new_n18570_, new_n18571_, new_n18572_, new_n18573_, new_n18574_,
    new_n18575_, new_n18576_, new_n18577_, new_n18578_, new_n18579_,
    new_n18580_, new_n18581_, new_n18582_, new_n18583_, new_n18584_,
    new_n18585_, new_n18586_, new_n18587_, new_n18588_, new_n18589_,
    new_n18590_, new_n18591_, new_n18592_, new_n18593_, new_n18594_,
    new_n18595_, new_n18596_, new_n18597_, new_n18598_, new_n18599_,
    new_n18600_, new_n18601_, new_n18602_, new_n18603_, new_n18604_,
    new_n18605_, new_n18606_, new_n18607_, new_n18608_, new_n18609_,
    new_n18610_, new_n18611_, new_n18612_, new_n18613_, new_n18614_,
    new_n18615_, new_n18616_, new_n18617_, new_n18618_, new_n18619_,
    new_n18620_, new_n18621_, new_n18622_, new_n18623_, new_n18624_,
    new_n18625_, new_n18626_, new_n18627_, new_n18628_, new_n18629_,
    new_n18630_, new_n18631_, new_n18632_, new_n18633_, new_n18634_,
    new_n18635_, new_n18636_, new_n18637_, new_n18638_, new_n18639_,
    new_n18640_, new_n18641_, new_n18642_, new_n18643_, new_n18644_,
    new_n18645_, new_n18646_, new_n18647_, new_n18648_, new_n18649_,
    new_n18650_, new_n18651_, new_n18652_, new_n18653_, new_n18654_,
    new_n18655_, new_n18656_, new_n18657_, new_n18658_, new_n18659_,
    new_n18660_, new_n18661_, new_n18662_, new_n18663_, new_n18664_,
    new_n18665_, new_n18666_, new_n18667_, new_n18668_, new_n18669_,
    new_n18670_, new_n18671_, new_n18672_, new_n18673_, new_n18674_,
    new_n18675_, new_n18676_, new_n18677_, new_n18678_, new_n18679_,
    new_n18680_, new_n18681_, new_n18682_, new_n18683_, new_n18684_,
    new_n18685_, new_n18686_, new_n18687_, new_n18688_, new_n18689_,
    new_n18690_, new_n18691_, new_n18692_, new_n18693_, new_n18694_,
    new_n18695_, new_n18696_, new_n18697_, new_n18698_, new_n18699_,
    new_n18700_, new_n18701_, new_n18702_, new_n18703_, new_n18704_,
    new_n18705_, new_n18706_, new_n18707_, new_n18708_, new_n18709_,
    new_n18710_, new_n18711_, new_n18712_, new_n18713_, new_n18714_,
    new_n18715_, new_n18716_, new_n18717_, new_n18718_, new_n18719_,
    new_n18720_, new_n18721_, new_n18722_, new_n18723_, new_n18724_,
    new_n18725_, new_n18726_, new_n18727_, new_n18728_, new_n18729_,
    new_n18730_, new_n18731_, new_n18732_, new_n18733_, new_n18734_,
    new_n18735_, new_n18736_, new_n18737_, new_n18738_, new_n18739_,
    new_n18740_, new_n18741_, new_n18742_, new_n18743_, new_n18744_,
    new_n18745_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18752_, new_n18753_, new_n18754_,
    new_n18755_, new_n18756_, new_n18757_, new_n18758_, new_n18759_,
    new_n18760_, new_n18761_, new_n18762_, new_n18763_, new_n18764_,
    new_n18765_, new_n18766_, new_n18767_, new_n18768_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18773_, new_n18774_,
    new_n18775_, new_n18776_, new_n18777_, new_n18778_, new_n18779_,
    new_n18780_, new_n18781_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18794_,
    new_n18795_, new_n18796_, new_n18797_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18951_, new_n18952_, new_n18953_, new_n18954_,
    new_n18955_, new_n18956_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18962_, new_n18963_, new_n18964_,
    new_n18965_, new_n18966_, new_n18967_, new_n18968_, new_n18969_,
    new_n18970_, new_n18971_, new_n18972_, new_n18973_, new_n18974_,
    new_n18975_, new_n18976_, new_n18977_, new_n18978_, new_n18979_,
    new_n18980_, new_n18981_, new_n18982_, new_n18983_, new_n18984_,
    new_n18985_, new_n18986_, new_n18987_, new_n18988_, new_n18989_,
    new_n18990_, new_n18991_, new_n18992_, new_n18993_, new_n18994_,
    new_n18995_, new_n18996_, new_n18997_, new_n18998_, new_n18999_,
    new_n19000_, new_n19001_, new_n19002_, new_n19003_, new_n19004_,
    new_n19005_, new_n19006_, new_n19007_, new_n19008_, new_n19009_,
    new_n19010_, new_n19011_, new_n19012_, new_n19013_, new_n19014_,
    new_n19015_, new_n19016_, new_n19017_, new_n19018_, new_n19019_,
    new_n19020_, new_n19021_, new_n19022_, new_n19023_, new_n19024_,
    new_n19025_, new_n19026_, new_n19027_, new_n19028_, new_n19029_,
    new_n19030_, new_n19031_, new_n19032_, new_n19033_, new_n19034_,
    new_n19035_, new_n19036_, new_n19037_, new_n19038_, new_n19039_,
    new_n19040_, new_n19041_, new_n19042_, new_n19043_, new_n19044_,
    new_n19045_, new_n19046_, new_n19047_, new_n19048_, new_n19049_,
    new_n19050_, new_n19051_, new_n19052_, new_n19053_, new_n19054_,
    new_n19055_, new_n19056_, new_n19057_, new_n19058_, new_n19059_,
    new_n19060_, new_n19061_, new_n19062_, new_n19063_, new_n19064_,
    new_n19065_, new_n19066_, new_n19067_, new_n19068_, new_n19069_,
    new_n19070_, new_n19071_, new_n19072_, new_n19073_, new_n19074_,
    new_n19075_, new_n19076_, new_n19077_, new_n19078_, new_n19079_,
    new_n19080_, new_n19081_, new_n19082_, new_n19083_, new_n19084_,
    new_n19085_, new_n19086_, new_n19087_, new_n19088_, new_n19089_,
    new_n19090_, new_n19091_, new_n19092_, new_n19093_, new_n19094_,
    new_n19095_, new_n19096_, new_n19097_, new_n19098_, new_n19099_,
    new_n19100_, new_n19101_, new_n19102_, new_n19103_, new_n19104_,
    new_n19105_, new_n19106_, new_n19107_, new_n19108_, new_n19109_,
    new_n19110_, new_n19111_, new_n19112_, new_n19113_, new_n19114_,
    new_n19115_, new_n19116_, new_n19117_, new_n19118_, new_n19119_,
    new_n19120_, new_n19121_, new_n19122_, new_n19123_, new_n19124_,
    new_n19125_, new_n19126_, new_n19127_, new_n19128_, new_n19129_,
    new_n19130_, new_n19131_, new_n19132_, new_n19133_, new_n19134_,
    new_n19135_, new_n19136_, new_n19137_, new_n19138_, new_n19139_,
    new_n19140_, new_n19141_, new_n19142_, new_n19143_, new_n19144_,
    new_n19145_, new_n19146_, new_n19147_, new_n19148_, new_n19149_,
    new_n19150_, new_n19151_, new_n19152_, new_n19153_, new_n19154_,
    new_n19155_, new_n19156_, new_n19157_, new_n19158_, new_n19159_,
    new_n19160_, new_n19161_, new_n19162_, new_n19163_, new_n19164_,
    new_n19165_, new_n19166_, new_n19167_, new_n19168_, new_n19169_,
    new_n19170_, new_n19171_, new_n19172_, new_n19173_, new_n19174_,
    new_n19175_, new_n19176_, new_n19177_, new_n19178_, new_n19179_,
    new_n19180_, new_n19181_, new_n19182_, new_n19183_, new_n19184_,
    new_n19185_, new_n19186_, new_n19187_, new_n19188_, new_n19189_,
    new_n19190_, new_n19191_, new_n19192_, new_n19193_, new_n19194_,
    new_n19195_, new_n19196_, new_n19197_, new_n19198_, new_n19199_,
    new_n19200_, new_n19201_, new_n19202_, new_n19203_, new_n19204_,
    new_n19205_, new_n19206_, new_n19207_, new_n19208_, new_n19209_,
    new_n19210_, new_n19211_, new_n19212_, new_n19213_, new_n19214_,
    new_n19215_, new_n19216_, new_n19217_, new_n19218_, new_n19219_,
    new_n19220_, new_n19221_, new_n19222_, new_n19223_, new_n19224_,
    new_n19225_, new_n19226_, new_n19227_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19233_, new_n19234_,
    new_n19235_, new_n19236_, new_n19237_, new_n19238_, new_n19239_,
    new_n19240_, new_n19241_, new_n19242_, new_n19243_, new_n19244_,
    new_n19245_, new_n19246_, new_n19247_, new_n19248_, new_n19249_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19277_, new_n19278_, new_n19279_,
    new_n19280_, new_n19281_, new_n19282_, new_n19283_, new_n19284_,
    new_n19285_, new_n19286_, new_n19287_, new_n19288_, new_n19289_,
    new_n19290_, new_n19291_, new_n19292_, new_n19293_, new_n19294_,
    new_n19295_, new_n19296_, new_n19297_, new_n19298_, new_n19299_,
    new_n19300_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19346_, new_n19347_, new_n19348_, new_n19349_,
    new_n19350_, new_n19351_, new_n19352_, new_n19353_, new_n19354_,
    new_n19355_, new_n19356_, new_n19357_, new_n19358_, new_n19359_,
    new_n19360_, new_n19361_, new_n19362_, new_n19363_, new_n19364_,
    new_n19365_, new_n19366_, new_n19367_, new_n19368_, new_n19369_,
    new_n19370_, new_n19371_, new_n19372_, new_n19373_, new_n19374_,
    new_n19375_, new_n19376_, new_n19377_, new_n19378_, new_n19379_,
    new_n19380_, new_n19381_, new_n19382_, new_n19383_, new_n19384_,
    new_n19385_, new_n19386_, new_n19387_, new_n19388_, new_n19389_,
    new_n19390_, new_n19391_, new_n19392_, new_n19393_, new_n19394_,
    new_n19395_, new_n19396_, new_n19397_, new_n19398_, new_n19399_,
    new_n19400_, new_n19401_, new_n19402_, new_n19403_, new_n19404_,
    new_n19405_, new_n19406_, new_n19407_, new_n19408_, new_n19409_,
    new_n19410_, new_n19411_, new_n19412_, new_n19413_, new_n19414_,
    new_n19415_, new_n19416_, new_n19417_, new_n19418_, new_n19419_,
    new_n19420_, new_n19421_, new_n19422_, new_n19423_, new_n19424_,
    new_n19425_, new_n19426_, new_n19427_, new_n19428_, new_n19429_,
    new_n19430_, new_n19431_, new_n19432_, new_n19433_, new_n19434_,
    new_n19435_, new_n19436_, new_n19437_, new_n19438_, new_n19439_,
    new_n19440_, new_n19441_, new_n19442_, new_n19443_, new_n19444_,
    new_n19445_, new_n19446_, new_n19447_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19456_, new_n19457_, new_n19458_, new_n19459_,
    new_n19460_, new_n19461_, new_n19462_, new_n19463_, new_n19464_,
    new_n19465_, new_n19466_, new_n19467_, new_n19468_, new_n19469_,
    new_n19470_, new_n19471_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19531_, new_n19532_, new_n19533_, new_n19534_,
    new_n19535_, new_n19536_, new_n19537_, new_n19538_, new_n19539_,
    new_n19540_, new_n19541_, new_n19542_, new_n19543_, new_n19544_,
    new_n19545_, new_n19546_, new_n19547_, new_n19548_, new_n19549_,
    new_n19550_, new_n19551_, new_n19552_, new_n19553_, new_n19554_,
    new_n19555_, new_n19556_, new_n19557_, new_n19558_, new_n19559_,
    new_n19560_, new_n19561_, new_n19562_, new_n19563_, new_n19564_,
    new_n19565_, new_n19566_, new_n19567_, new_n19568_, new_n19569_,
    new_n19570_, new_n19571_, new_n19572_, new_n19573_, new_n19574_,
    new_n19575_, new_n19576_, new_n19577_, new_n19578_, new_n19579_,
    new_n19580_, new_n19581_, new_n19582_, new_n19583_, new_n19584_,
    new_n19585_, new_n19586_, new_n19587_, new_n19588_, new_n19589_,
    new_n19590_, new_n19591_, new_n19592_, new_n19593_, new_n19594_,
    new_n19595_, new_n19596_, new_n19597_, new_n19598_, new_n19599_,
    new_n19600_, new_n19601_, new_n19602_, new_n19603_, new_n19604_,
    new_n19605_, new_n19606_, new_n19607_, new_n19608_, new_n19609_,
    new_n19610_, new_n19611_, new_n19612_, new_n19613_, new_n19614_,
    new_n19615_, new_n19616_, new_n19617_, new_n19618_, new_n19619_,
    new_n19620_, new_n19621_, new_n19622_, new_n19623_, new_n19624_,
    new_n19625_, new_n19626_, new_n19627_, new_n19628_, new_n19629_,
    new_n19630_, new_n19631_, new_n19632_, new_n19633_, new_n19634_,
    new_n19635_, new_n19636_, new_n19637_, new_n19638_, new_n19639_,
    new_n19640_, new_n19641_, new_n19642_, new_n19643_, new_n19644_,
    new_n19645_, new_n19646_, new_n19647_, new_n19648_, new_n19649_,
    new_n19650_, new_n19651_, new_n19652_, new_n19653_, new_n19654_,
    new_n19655_, new_n19656_, new_n19657_, new_n19658_, new_n19659_,
    new_n19660_, new_n19661_, new_n19662_, new_n19663_, new_n19664_,
    new_n19665_, new_n19666_, new_n19667_, new_n19668_, new_n19669_,
    new_n19670_, new_n19671_, new_n19672_, new_n19673_, new_n19674_,
    new_n19675_, new_n19676_, new_n19677_, new_n19678_, new_n19679_,
    new_n19680_, new_n19681_, new_n19682_, new_n19683_, new_n19684_,
    new_n19685_, new_n19686_, new_n19687_, new_n19688_, new_n19689_,
    new_n19690_, new_n19691_, new_n19692_, new_n19693_, new_n19694_,
    new_n19695_, new_n19696_, new_n19697_, new_n19698_, new_n19699_,
    new_n19700_, new_n19701_, new_n19702_, new_n19703_, new_n19704_,
    new_n19705_, new_n19706_, new_n19707_, new_n19708_, new_n19709_,
    new_n19710_, new_n19711_, new_n19712_, new_n19713_, new_n19714_,
    new_n19715_, new_n19716_, new_n19717_, new_n19718_, new_n19719_,
    new_n19720_, new_n19721_, new_n19722_, new_n19723_, new_n19724_,
    new_n19725_, new_n19726_, new_n19727_, new_n19728_, new_n19729_,
    new_n19730_, new_n19731_, new_n19732_, new_n19733_, new_n19734_,
    new_n19735_, new_n19736_, new_n19737_, new_n19738_, new_n19739_,
    new_n19740_, new_n19741_, new_n19742_, new_n19743_, new_n19744_,
    new_n19745_, new_n19746_, new_n19747_, new_n19748_, new_n19749_,
    new_n19750_, new_n19751_, new_n19752_, new_n19753_, new_n19754_,
    new_n19755_, new_n19756_, new_n19757_, new_n19758_, new_n19759_,
    new_n19760_, new_n19761_, new_n19762_, new_n19763_, new_n19764_,
    new_n19765_, new_n19766_, new_n19767_, new_n19768_, new_n19769_,
    new_n19770_, new_n19771_, new_n19772_, new_n19773_, new_n19774_,
    new_n19775_, new_n19776_, new_n19777_, new_n19778_, new_n19779_,
    new_n19780_, new_n19781_, new_n19782_, new_n19783_, new_n19784_,
    new_n19785_, new_n19786_, new_n19787_, new_n19788_, new_n19789_,
    new_n19790_, new_n19791_, new_n19792_, new_n19793_, new_n19794_,
    new_n19795_, new_n19796_, new_n19797_, new_n19798_, new_n19799_,
    new_n19800_, new_n19801_, new_n19802_, new_n19803_, new_n19804_,
    new_n19805_, new_n19806_, new_n19807_, new_n19808_, new_n19809_,
    new_n19810_, new_n19811_, new_n19812_, new_n19813_, new_n19814_,
    new_n19815_, new_n19816_, new_n19817_, new_n19818_, new_n19819_,
    new_n19820_, new_n19821_, new_n19822_, new_n19823_, new_n19824_,
    new_n19825_, new_n19826_, new_n19827_, new_n19828_, new_n19829_,
    new_n19830_, new_n19831_, new_n19832_, new_n19833_, new_n19834_,
    new_n19835_, new_n19836_, new_n19837_, new_n19838_, new_n19839_,
    new_n19840_, new_n19841_, new_n19842_, new_n19843_, new_n19844_,
    new_n19845_, new_n19846_, new_n19847_, new_n19848_, new_n19849_,
    new_n19850_, new_n19851_, new_n19852_, new_n19853_, new_n19854_,
    new_n19855_, new_n19856_, new_n19857_, new_n19858_, new_n19859_,
    new_n19860_, new_n19861_, new_n19862_, new_n19863_, new_n19864_,
    new_n19865_, new_n19866_, new_n19867_, new_n19868_, new_n19869_,
    new_n19870_, new_n19871_, new_n19872_, new_n19873_, new_n19874_,
    new_n19875_, new_n19876_, new_n19877_, new_n19878_, new_n19879_,
    new_n19880_, new_n19881_, new_n19882_, new_n19883_, new_n19884_,
    new_n19885_, new_n19886_, new_n19887_, new_n19888_, new_n19889_,
    new_n19890_, new_n19891_, new_n19892_, new_n19893_, new_n19894_,
    new_n19895_, new_n19896_, new_n19897_, new_n19898_, new_n19899_,
    new_n19900_, new_n19901_, new_n19902_, new_n19903_, new_n19904_,
    new_n19905_, new_n19906_, new_n19907_, new_n19908_, new_n19909_,
    new_n19910_, new_n19911_, new_n19912_, new_n19913_, new_n19914_,
    new_n19915_, new_n19916_, new_n19917_, new_n19918_, new_n19919_,
    new_n19920_, new_n19921_, new_n19922_, new_n19923_, new_n19924_,
    new_n19925_, new_n19926_, new_n19927_, new_n19928_, new_n19929_,
    new_n19930_, new_n19931_, new_n19932_, new_n19933_, new_n19934_,
    new_n19935_, new_n19936_, new_n19937_, new_n19938_, new_n19939_,
    new_n19940_, new_n19941_, new_n19942_, new_n19943_, new_n19944_,
    new_n19945_, new_n19946_, new_n19947_, new_n19948_, new_n19949_,
    new_n19950_, new_n19951_, new_n19952_, new_n19953_, new_n19954_,
    new_n19955_, new_n19956_, new_n19957_, new_n19958_, new_n19959_,
    new_n19960_, new_n19961_, new_n19962_, new_n19963_, new_n19964_,
    new_n19965_, new_n19966_, new_n19967_, new_n19968_, new_n19969_,
    new_n19970_, new_n19971_, new_n19972_, new_n19973_, new_n19974_,
    new_n19975_, new_n19976_, new_n19977_, new_n19978_, new_n19979_,
    new_n19980_, new_n19981_, new_n19982_, new_n19983_, new_n19984_,
    new_n19985_, new_n19986_, new_n19987_, new_n19988_, new_n19989_,
    new_n19990_, new_n19991_, new_n19992_, new_n19993_, new_n19994_,
    new_n19995_, new_n19996_, new_n19997_, new_n19998_, new_n19999_,
    new_n20000_, new_n20001_, new_n20002_, new_n20003_, new_n20004_,
    new_n20005_, new_n20006_, new_n20007_, new_n20008_, new_n20009_,
    new_n20010_, new_n20011_, new_n20012_, new_n20013_, new_n20014_,
    new_n20015_, new_n20016_, new_n20017_, new_n20018_, new_n20019_,
    new_n20020_, new_n20021_, new_n20022_, new_n20023_, new_n20024_,
    new_n20025_, new_n20026_, new_n20027_, new_n20028_, new_n20029_,
    new_n20030_, new_n20031_, new_n20032_, new_n20033_, new_n20034_,
    new_n20035_, new_n20036_, new_n20037_, new_n20038_, new_n20039_,
    new_n20040_, new_n20041_, new_n20042_, new_n20043_, new_n20044_,
    new_n20045_, new_n20046_, new_n20047_, new_n20048_, new_n20049_,
    new_n20050_, new_n20051_, new_n20052_, new_n20053_, new_n20054_,
    new_n20055_, new_n20056_, new_n20057_, new_n20058_, new_n20059_,
    new_n20060_, new_n20061_, new_n20062_, new_n20063_, new_n20064_,
    new_n20065_, new_n20066_, new_n20067_, new_n20068_, new_n20069_,
    new_n20070_, new_n20071_, new_n20072_, new_n20073_, new_n20074_,
    new_n20075_, new_n20076_, new_n20077_, new_n20078_, new_n20079_,
    new_n20080_, new_n20081_, new_n20082_, new_n20083_, new_n20084_,
    new_n20085_, new_n20086_, new_n20087_, new_n20088_, new_n20089_,
    new_n20090_, new_n20091_, new_n20092_, new_n20093_, new_n20094_,
    new_n20095_, new_n20096_, new_n20097_, new_n20098_, new_n20099_,
    new_n20100_, new_n20101_, new_n20102_, new_n20103_, new_n20104_,
    new_n20105_, new_n20106_, new_n20107_, new_n20108_, new_n20109_,
    new_n20110_, new_n20111_, new_n20112_, new_n20113_, new_n20114_,
    new_n20115_, new_n20116_, new_n20117_, new_n20118_, new_n20119_,
    new_n20120_, new_n20121_, new_n20122_, new_n20123_, new_n20124_,
    new_n20125_, new_n20126_, new_n20127_, new_n20128_, new_n20129_,
    new_n20130_, new_n20131_, new_n20132_, new_n20133_, new_n20134_,
    new_n20135_, new_n20136_, new_n20137_, new_n20138_, new_n20139_,
    new_n20140_, new_n20141_, new_n20142_, new_n20143_, new_n20144_,
    new_n20145_, new_n20146_, new_n20147_, new_n20148_, new_n20149_,
    new_n20150_, new_n20151_, new_n20152_, new_n20153_, new_n20154_,
    new_n20155_, new_n20156_, new_n20157_, new_n20158_, new_n20159_,
    new_n20160_, new_n20161_, new_n20162_, new_n20163_, new_n20164_,
    new_n20165_, new_n20166_, new_n20167_, new_n20168_, new_n20169_,
    new_n20170_, new_n20171_, new_n20172_, new_n20173_, new_n20174_,
    new_n20175_, new_n20176_, new_n20177_, new_n20178_, new_n20179_,
    new_n20180_, new_n20181_, new_n20182_, new_n20183_, new_n20184_,
    new_n20185_, new_n20186_, new_n20187_, new_n20188_, new_n20189_,
    new_n20190_, new_n20191_, new_n20192_, new_n20193_, new_n20194_,
    new_n20195_, new_n20196_, new_n20197_, new_n20198_, new_n20199_,
    new_n20200_, new_n20201_, new_n20202_, new_n20203_, new_n20204_,
    new_n20205_, new_n20206_, new_n20207_, new_n20208_, new_n20209_,
    new_n20210_, new_n20211_, new_n20212_, new_n20213_, new_n20214_,
    new_n20215_, new_n20216_, new_n20217_, new_n20218_, new_n20219_,
    new_n20220_, new_n20221_, new_n20222_, new_n20223_, new_n20224_,
    new_n20225_, new_n20226_, new_n20227_, new_n20228_, new_n20229_,
    new_n20230_, new_n20231_, new_n20232_, new_n20233_, new_n20234_,
    new_n20235_, new_n20236_, new_n20237_, new_n20238_, new_n20239_,
    new_n20240_, new_n20241_, new_n20242_, new_n20243_, new_n20244_,
    new_n20245_, new_n20246_, new_n20247_, new_n20248_, new_n20249_,
    new_n20250_, new_n20251_, new_n20252_, new_n20253_, new_n20254_,
    new_n20255_, new_n20256_, new_n20257_, new_n20258_, new_n20259_,
    new_n20260_, new_n20261_, new_n20262_, new_n20263_, new_n20264_,
    new_n20265_, new_n20266_, new_n20267_, new_n20268_, new_n20269_,
    new_n20270_, new_n20271_, new_n20272_, new_n20273_, new_n20274_,
    new_n20275_, new_n20276_, new_n20277_, new_n20278_, new_n20279_,
    new_n20280_, new_n20281_, new_n20282_, new_n20283_, new_n20284_,
    new_n20285_, new_n20286_, new_n20287_, new_n20288_, new_n20289_,
    new_n20290_, new_n20291_, new_n20292_, new_n20293_, new_n20294_,
    new_n20295_, new_n20296_, new_n20297_, new_n20298_, new_n20299_,
    new_n20300_, new_n20301_, new_n20302_, new_n20303_, new_n20304_,
    new_n20305_, new_n20306_, new_n20307_, new_n20308_, new_n20309_,
    new_n20310_, new_n20311_, new_n20312_, new_n20313_, new_n20314_,
    new_n20315_, new_n20316_, new_n20317_, new_n20318_, new_n20319_,
    new_n20320_, new_n20321_, new_n20322_, new_n20323_, new_n20324_,
    new_n20325_, new_n20326_, new_n20327_, new_n20328_, new_n20329_,
    new_n20330_, new_n20331_, new_n20332_, new_n20333_, new_n20334_,
    new_n20335_, new_n20336_, new_n20337_, new_n20338_, new_n20339_,
    new_n20340_, new_n20341_, new_n20342_, new_n20343_, new_n20344_,
    new_n20345_, new_n20346_, new_n20347_, new_n20348_, new_n20349_,
    new_n20350_, new_n20351_, new_n20352_, new_n20353_, new_n20354_,
    new_n20355_, new_n20356_, new_n20357_, new_n20358_, new_n20359_,
    new_n20360_, new_n20361_, new_n20362_, new_n20363_, new_n20364_,
    new_n20365_, new_n20366_, new_n20367_, new_n20368_, new_n20369_,
    new_n20370_, new_n20371_, new_n20372_, new_n20373_, new_n20374_,
    new_n20375_, new_n20376_, new_n20377_, new_n20378_, new_n20379_,
    new_n20380_, new_n20381_, new_n20382_, new_n20383_, new_n20384_,
    new_n20385_, new_n20386_, new_n20387_, new_n20388_, new_n20389_,
    new_n20390_, new_n20391_, new_n20392_, new_n20393_, new_n20394_,
    new_n20395_, new_n20396_, new_n20397_, new_n20398_, new_n20399_,
    new_n20400_, new_n20401_, new_n20402_, new_n20403_, new_n20404_,
    new_n20405_, new_n20406_, new_n20407_, new_n20408_, new_n20409_,
    new_n20410_, new_n20411_, new_n20412_, new_n20413_, new_n20414_,
    new_n20415_, new_n20416_, new_n20417_, new_n20418_, new_n20419_,
    new_n20420_, new_n20421_, new_n20422_, new_n20423_, new_n20424_,
    new_n20425_, new_n20426_, new_n20427_, new_n20428_, new_n20429_,
    new_n20430_, new_n20431_, new_n20432_, new_n20433_, new_n20434_,
    new_n20435_, new_n20436_, new_n20437_, new_n20438_, new_n20439_,
    new_n20440_, new_n20441_, new_n20442_, new_n20443_, new_n20444_,
    new_n20445_, new_n20446_, new_n20447_, new_n20448_, new_n20449_,
    new_n20450_, new_n20451_, new_n20452_, new_n20453_, new_n20454_,
    new_n20455_, new_n20456_, new_n20457_, new_n20458_, new_n20459_,
    new_n20460_, new_n20461_, new_n20462_, new_n20463_, new_n20464_,
    new_n20465_, new_n20466_, new_n20467_, new_n20468_, new_n20469_,
    new_n20470_, new_n20471_, new_n20472_, new_n20473_, new_n20474_,
    new_n20475_, new_n20476_, new_n20477_, new_n20478_, new_n20479_,
    new_n20480_, new_n20481_, new_n20482_, new_n20483_, new_n20484_,
    new_n20485_, new_n20486_, new_n20487_, new_n20488_, new_n20489_,
    new_n20490_, new_n20491_, new_n20492_, new_n20493_, new_n20494_,
    new_n20495_, new_n20496_, new_n20497_, new_n20498_, new_n20499_,
    new_n20500_, new_n20501_, new_n20502_, new_n20503_, new_n20504_,
    new_n20505_, new_n20506_, new_n20507_, new_n20508_, new_n20509_,
    new_n20510_, new_n20511_, new_n20512_, new_n20513_, new_n20514_,
    new_n20515_, new_n20516_, new_n20517_, new_n20518_, new_n20519_,
    new_n20520_, new_n20521_, new_n20522_, new_n20523_, new_n20524_,
    new_n20525_, new_n20526_, new_n20527_, new_n20528_, new_n20529_,
    new_n20530_, new_n20531_, new_n20532_, new_n20533_, new_n20534_,
    new_n20535_, new_n20536_, new_n20537_, new_n20538_, new_n20539_,
    new_n20540_, new_n20541_, new_n20542_, new_n20543_, new_n20544_,
    new_n20545_, new_n20546_, new_n20547_, new_n20548_, new_n20549_,
    new_n20550_, new_n20551_, new_n20552_, new_n20553_, new_n20554_,
    new_n20555_, new_n20556_, new_n20557_, new_n20558_, new_n20559_,
    new_n20560_, new_n20561_, new_n20562_, new_n20563_, new_n20564_,
    new_n20565_, new_n20566_, new_n20567_, new_n20568_, new_n20569_,
    new_n20570_, new_n20571_, new_n20572_, new_n20573_, new_n20574_,
    new_n20575_, new_n20576_, new_n20577_, new_n20578_, new_n20579_,
    new_n20580_, new_n20581_, new_n20582_, new_n20583_, new_n20584_,
    new_n20585_, new_n20586_, new_n20587_, new_n20588_, new_n20589_,
    new_n20590_, new_n20591_, new_n20592_, new_n20593_, new_n20594_,
    new_n20595_, new_n20596_, new_n20597_, new_n20598_, new_n20599_,
    new_n20600_, new_n20601_, new_n20602_, new_n20603_, new_n20604_,
    new_n20605_, new_n20606_, new_n20607_, new_n20608_, new_n20609_,
    new_n20610_, new_n20611_, new_n20612_, new_n20613_, new_n20614_,
    new_n20615_, new_n20616_, new_n20617_, new_n20618_, new_n20619_,
    new_n20620_, new_n20621_, new_n20622_, new_n20623_, new_n20624_,
    new_n20625_, new_n20626_, new_n20627_, new_n20628_, new_n20629_,
    new_n20630_, new_n20631_, new_n20632_, new_n20633_, new_n20634_,
    new_n20635_, new_n20636_, new_n20637_, new_n20638_, new_n20639_,
    new_n20640_, new_n20641_, new_n20642_, new_n20643_, new_n20644_,
    new_n20645_, new_n20646_, new_n20647_, new_n20648_, new_n20649_,
    new_n20650_, new_n20651_, new_n20652_, new_n20653_, new_n20654_,
    new_n20655_, new_n20656_, new_n20657_, new_n20658_, new_n20659_,
    new_n20660_, new_n20661_, new_n20662_, new_n20663_, new_n20664_,
    new_n20665_, new_n20666_, new_n20667_, new_n20668_, new_n20669_,
    new_n20670_, new_n20671_, new_n20672_, new_n20673_, new_n20674_,
    new_n20675_, new_n20676_, new_n20677_, new_n20678_, new_n20679_,
    new_n20680_, new_n20681_, new_n20682_, new_n20683_, new_n20684_,
    new_n20685_, new_n20686_, new_n20687_, new_n20688_, new_n20689_,
    new_n20690_, new_n20691_, new_n20692_, new_n20693_, new_n20694_,
    new_n20695_, new_n20696_, new_n20697_, new_n20698_, new_n20699_,
    new_n20700_, new_n20701_, new_n20702_, new_n20703_, new_n20704_,
    new_n20705_, new_n20706_, new_n20707_, new_n20708_, new_n20709_,
    new_n20710_, new_n20711_, new_n20712_, new_n20713_, new_n20714_,
    new_n20715_, new_n20716_, new_n20717_, new_n20718_, new_n20719_,
    new_n20720_, new_n20721_, new_n20722_, new_n20723_, new_n20724_,
    new_n20725_, new_n20726_, new_n20727_, new_n20728_, new_n20729_,
    new_n20730_, new_n20731_, new_n20732_, new_n20733_, new_n20734_,
    new_n20735_, new_n20736_, new_n20737_, new_n20738_, new_n20739_,
    new_n20740_, new_n20741_, new_n20742_, new_n20743_, new_n20744_,
    new_n20745_, new_n20746_, new_n20747_, new_n20748_, new_n20749_,
    new_n20750_, new_n20751_, new_n20752_, new_n20753_, new_n20754_,
    new_n20755_, new_n20756_, new_n20757_, new_n20758_, new_n20759_,
    new_n20760_, new_n20761_, new_n20762_, new_n20763_, new_n20764_,
    new_n20765_, new_n20766_, new_n20767_, new_n20768_, new_n20769_,
    new_n20770_, new_n20771_, new_n20772_, new_n20773_, new_n20774_,
    new_n20775_, new_n20776_, new_n20777_, new_n20778_, new_n20779_,
    new_n20780_, new_n20781_, new_n20782_, new_n20783_, new_n20784_,
    new_n20785_, new_n20786_, new_n20787_, new_n20788_, new_n20789_,
    new_n20790_, new_n20791_, new_n20792_, new_n20793_, new_n20794_,
    new_n20795_, new_n20796_, new_n20797_, new_n20798_, new_n20799_,
    new_n20800_, new_n20801_, new_n20802_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20836_, new_n20837_, new_n20838_, new_n20839_,
    new_n20840_, new_n20841_, new_n20842_, new_n20843_, new_n20844_,
    new_n20845_, new_n20846_, new_n20847_, new_n20848_, new_n20849_,
    new_n20850_, new_n20851_, new_n20852_, new_n20853_, new_n20854_,
    new_n20855_, new_n20856_, new_n20857_, new_n20858_, new_n20859_,
    new_n20860_, new_n20861_, new_n20862_, new_n20863_, new_n20864_,
    new_n20865_, new_n20866_, new_n20867_, new_n20868_, new_n20869_,
    new_n20870_, new_n20871_, new_n20872_, new_n20873_, new_n20874_,
    new_n20875_, new_n20876_, new_n20877_, new_n20878_, new_n20879_,
    new_n20880_, new_n20881_, new_n20882_, new_n20883_, new_n20884_,
    new_n20885_, new_n20886_, new_n20887_, new_n20888_, new_n20889_,
    new_n20890_, new_n20891_, new_n20892_, new_n20893_, new_n20894_,
    new_n20895_, new_n20896_, new_n20897_, new_n20898_, new_n20899_,
    new_n20900_, new_n20901_, new_n20902_, new_n20903_, new_n20904_,
    new_n20905_, new_n20906_, new_n20907_, new_n20908_, new_n20909_,
    new_n20910_, new_n20911_, new_n20912_, new_n20913_, new_n20914_,
    new_n20915_, new_n20916_, new_n20917_, new_n20918_, new_n20919_,
    new_n20920_, new_n20921_, new_n20922_, new_n20923_, new_n20924_,
    new_n20925_, new_n20926_, new_n20927_, new_n20928_, new_n20929_,
    new_n20930_, new_n20931_, new_n20932_, new_n20933_, new_n20934_,
    new_n20935_, new_n20936_, new_n20937_, new_n20938_, new_n20939_,
    new_n20940_, new_n20941_, new_n20942_, new_n20943_, new_n20944_,
    new_n20945_, new_n20946_, new_n20947_, new_n20948_, new_n20949_,
    new_n20950_, new_n20951_, new_n20952_, new_n20953_, new_n20954_,
    new_n20955_, new_n20956_, new_n20957_, new_n20958_, new_n20959_,
    new_n20960_, new_n20961_, new_n20962_, new_n20963_, new_n20964_,
    new_n20965_, new_n20966_, new_n20967_, new_n20968_, new_n20969_,
    new_n20970_, new_n20971_, new_n20972_, new_n20973_, new_n20974_,
    new_n20975_, new_n20976_, new_n20977_, new_n20978_, new_n20979_,
    new_n20980_, new_n20981_, new_n20982_, new_n20983_, new_n20984_,
    new_n20985_, new_n20986_, new_n20987_, new_n20988_, new_n20989_,
    new_n20990_, new_n20991_, new_n20992_, new_n20993_, new_n20994_,
    new_n20995_, new_n20996_, new_n20997_, new_n20998_, new_n20999_,
    new_n21000_, new_n21001_, new_n21002_, new_n21003_, new_n21004_,
    new_n21005_, new_n21006_, new_n21007_, new_n21008_, new_n21009_,
    new_n21010_, new_n21011_, new_n21012_, new_n21013_, new_n21014_,
    new_n21015_, new_n21016_, new_n21017_, new_n21018_, new_n21019_,
    new_n21020_, new_n21021_, new_n21022_, new_n21023_, new_n21024_,
    new_n21025_, new_n21026_, new_n21027_, new_n21028_, new_n21029_,
    new_n21030_, new_n21031_, new_n21032_, new_n21033_, new_n21034_,
    new_n21035_, new_n21036_, new_n21037_, new_n21038_, new_n21039_,
    new_n21040_, new_n21041_, new_n21042_, new_n21043_, new_n21044_,
    new_n21045_, new_n21046_, new_n21047_, new_n21048_, new_n21049_,
    new_n21050_, new_n21051_, new_n21052_, new_n21053_, new_n21054_,
    new_n21055_, new_n21056_, new_n21057_, new_n21058_, new_n21059_,
    new_n21060_, new_n21061_, new_n21062_;
  assign new_n1036_ = ~new_n20820_ | ~new_n20981_;
  assign new_n1037_ = ~new_n20989_ | ~new_n20732_;
  assign new_n1038_ = ~new_n4678_ | ~new_n20691_;
  assign new_n1039_ = ~new_n1150_ | ~new_n1149_;
  assign new_n1040_ = ~new_n1152_ | ~new_n1151_;
  assign new_n1041_ = ~new_n1154_ | ~new_n1153_;
  assign new_n1042_ = ~new_n1156_ | ~new_n1155_;
  assign new_n1043_ = ~new_n1158_ | ~new_n1157_;
  assign new_n1044_ = ~new_n1160_ | ~new_n1159_;
  assign new_n1045_ = ~new_n1162_ | ~new_n1161_;
  assign new_n1046_ = ~new_n1164_ | ~new_n1163_;
  assign new_n1047_ = ~new_n1166_ | ~new_n1165_;
  assign new_n1048_ = ~new_n1168_ | ~new_n1167_;
  assign new_n1049_ = ~new_n1170_ | ~new_n1169_;
  assign new_n1050_ = ~new_n1172_ | ~new_n1171_;
  assign new_n1051_ = ~new_n1174_ | ~new_n1173_;
  assign new_n1052_ = ~new_n1176_ | ~new_n1175_;
  assign new_n1053_ = ~new_n1178_ | ~new_n1177_;
  assign new_n1054_ = ~new_n1180_ | ~new_n1179_;
  assign new_n1055_ = ~new_n1182_ | ~new_n1181_;
  assign new_n1056_ = ~new_n1184_ | ~new_n1183_;
  assign new_n1057_ = ~new_n1186_ | ~new_n1185_;
  assign new_n1058_ = ~new_n1188_ | ~new_n1187_;
  assign new_n1059_ = ~new_n1190_ | ~new_n1189_;
  assign new_n1060_ = ~new_n1192_ | ~new_n1191_;
  assign new_n1061_ = ~new_n1194_ | ~new_n1193_;
  assign new_n1062_ = ~new_n1196_ | ~new_n1195_;
  assign new_n1063_ = ~new_n1198_ | ~new_n1197_;
  assign new_n1064_ = ~new_n1200_ | ~new_n1199_;
  assign new_n1065_ = ~new_n1202_ | ~new_n1201_;
  assign new_n1066_ = ~new_n1204_ | ~new_n1203_;
  assign new_n1067_ = ~new_n1206_ | ~new_n1205_;
  assign new_n1068_ = ~new_n1208_ | ~new_n1207_;
  assign new_n1069_ = ~new_n1210_ | ~new_n1209_;
  assign new_n1070_ = ~new_n1212_ | ~new_n1211_;
  assign new_n1071_ = ~new_n1214_ | ~new_n1213_;
  assign new_n1072_ = ~new_n1216_ | ~new_n1215_;
  assign new_n1073_ = ~new_n1218_ | ~new_n1217_;
  assign new_n1074_ = ~new_n1220_ | ~new_n1219_;
  assign new_n1075_ = ~new_n1222_ | ~new_n1221_;
  assign new_n1076_ = ~new_n1224_ | ~new_n1223_;
  assign new_n1077_ = ~new_n1226_ | ~new_n1225_;
  assign new_n1078_ = ~new_n1228_ | ~new_n1227_;
  assign new_n1079_ = ~new_n1230_ | ~new_n1229_;
  assign new_n1080_ = ~new_n1232_ | ~new_n1231_;
  assign new_n1081_ = ~new_n1234_ | ~new_n1233_;
  assign new_n1082_ = ~new_n1236_ | ~new_n1235_;
  assign new_n1083_ = ~new_n1238_ | ~new_n1237_;
  assign new_n1084_ = ~new_n1240_ | ~new_n1239_;
  assign new_n1085_ = ~new_n1242_ | ~new_n1241_;
  assign new_n1086_ = ~new_n1244_ | ~new_n1243_;
  assign new_n1087_ = ~new_n1246_ | ~new_n1245_;
  assign new_n1088_ = ~new_n1248_ | ~new_n1247_;
  assign new_n1089_ = ~new_n1250_ | ~new_n1249_;
  assign new_n1090_ = ~new_n1252_ | ~new_n1251_;
  assign new_n1091_ = ~new_n1254_ | ~new_n1253_;
  assign new_n1092_ = ~new_n1256_ | ~new_n1255_;
  assign new_n1093_ = ~new_n1258_ | ~new_n1257_;
  assign new_n1094_ = ~new_n1260_ | ~new_n1259_;
  assign new_n1095_ = ~new_n1262_ | ~new_n1261_;
  assign new_n1096_ = ~new_n1264_ | ~new_n1263_;
  assign new_n1097_ = ~new_n1266_ | ~new_n1265_;
  assign new_n1098_ = ~new_n1268_ | ~new_n1267_;
  assign new_n1099_ = ~new_n1270_ | ~new_n1269_;
  assign new_n1100_ = ~new_n1272_ | ~new_n1271_;
  assign new_n1101_ = ~new_n1274_ | ~new_n1273_;
  assign new_n1102_ = ~new_n1276_ | ~new_n1275_;
  assign new_n1103_ = ~new_n1278_ | ~new_n1277_;
  assign new_n1104_ = ~new_n1280_ | ~new_n1279_;
  assign new_n1105_ = ~new_n1282_ | ~new_n1281_;
  assign new_n1106_ = ~new_n1284_ | ~new_n1283_;
  assign new_n1107_ = ~new_n1286_ | ~new_n1285_;
  assign new_n1108_ = ~new_n1288_ | ~new_n1287_;
  assign new_n1109_ = ~new_n1290_ | ~new_n1289_;
  assign new_n1110_ = ~new_n1292_ | ~new_n1291_;
  assign new_n1111_ = ~new_n1294_ | ~new_n1293_;
  assign new_n1112_ = ~new_n1296_ | ~new_n1295_;
  assign new_n1113_ = ~new_n1298_ | ~new_n1297_;
  assign new_n1114_ = ~new_n1300_ | ~new_n1299_;
  assign new_n1115_ = ~new_n1302_ | ~new_n1301_;
  assign new_n1116_ = ~new_n1304_ | ~new_n1303_;
  assign new_n1117_ = ~new_n1306_ | ~new_n1305_;
  assign new_n1118_ = ~new_n1308_ | ~new_n1307_;
  assign new_n1119_ = ~new_n1310_ | ~new_n1309_;
  assign new_n1120_ = ~new_n1312_ | ~new_n1311_;
  assign new_n1121_ = ~new_n1314_ | ~new_n1313_;
  assign new_n1122_ = ~new_n1316_ | ~new_n1315_;
  assign new_n1123_ = ~new_n1318_ | ~new_n1317_;
  assign new_n1124_ = ~new_n1320_ | ~new_n1319_;
  assign new_n1125_ = ~new_n1322_ | ~new_n1321_;
  assign new_n1126_ = ~new_n1324_ | ~new_n1323_;
  assign new_n1127_ = ~new_n1326_ | ~new_n1325_;
  assign new_n1128_ = ~new_n1328_ | ~new_n1327_;
  assign new_n1129_ = ~new_n1330_ | ~new_n1329_;
  assign new_n1130_ = ~new_n1332_ | ~new_n1331_;
  assign new_n1131_ = ~new_n1334_ | ~new_n1333_;
  assign new_n1132_ = ~new_n1336_ | ~new_n1335_;
  assign new_n1133_ = ~new_n1338_ | ~new_n1337_;
  assign new_n1134_ = ~new_n1340_ | ~new_n1339_;
  assign new_n1135_ = ~pi522;
  assign new_n1136_ = ~pi277;
  assign po021 = new_n1146_ & new_n1145_;
  assign new_n1138_ = ~pi521;
  assign new_n1139_ = ~pi276;
  assign po020 = new_n1148_ & new_n1147_;
  assign new_n1141_ = ~new_n1143_ | ~new_n1142_;
  assign new_n1142_ = ~new_n8734_ | ~new_n7907_ | ~new_n1139_;
  assign new_n1143_ = ~pi438 | ~pi193 | ~new_n1138_;
  assign new_n1144_ = ~new_n1141_;
  assign new_n1145_ = ~pi522 | ~new_n1136_;
  assign new_n1146_ = ~pi277 | ~new_n1135_;
  assign new_n1147_ = ~pi521 | ~new_n1139_;
  assign new_n1148_ = ~pi276 | ~new_n1138_;
  assign new_n1149_ = ~pi222 | ~new_n1141_;
  assign new_n1150_ = ~new_n8276_ | ~new_n1144_;
  assign new_n1151_ = ~pi221 | ~new_n1141_;
  assign new_n1152_ = ~new_n8277_ | ~new_n1144_;
  assign new_n1153_ = ~pi220 | ~new_n1141_;
  assign new_n1154_ = ~new_n8278_ | ~new_n1144_;
  assign new_n1155_ = ~pi219 | ~new_n1141_;
  assign new_n1156_ = ~new_n8279_ | ~new_n1144_;
  assign new_n1157_ = ~pi218 | ~new_n1141_;
  assign new_n1158_ = ~new_n8280_ | ~new_n1144_;
  assign new_n1159_ = ~pi217 | ~new_n1141_;
  assign new_n1160_ = ~new_n8281_ | ~new_n1144_;
  assign new_n1161_ = ~pi216 | ~new_n1141_;
  assign new_n1162_ = ~new_n8282_ | ~new_n1144_;
  assign new_n1163_ = ~pi244 | ~new_n1141_;
  assign new_n1164_ = ~new_n8203_ | ~new_n1144_;
  assign new_n1165_ = ~pi243 | ~new_n1141_;
  assign new_n1166_ = ~new_n8283_ | ~new_n1144_;
  assign new_n1167_ = ~pi215 | ~new_n1141_;
  assign new_n1168_ = ~new_n8284_ | ~new_n1144_;
  assign new_n1169_ = ~pi242 | ~new_n1141_;
  assign new_n1170_ = ~new_n8285_ | ~new_n1144_;
  assign new_n1171_ = ~pi241 | ~new_n1141_;
  assign new_n1172_ = ~new_n8286_ | ~new_n1144_;
  assign new_n1173_ = ~pi240 | ~new_n1141_;
  assign new_n1174_ = ~new_n8287_ | ~new_n1144_;
  assign new_n1175_ = ~pi239 | ~new_n1141_;
  assign new_n1176_ = ~new_n8288_ | ~new_n1144_;
  assign new_n1177_ = ~pi238 | ~new_n1141_;
  assign new_n1178_ = ~new_n8289_ | ~new_n1144_;
  assign new_n1179_ = ~pi237 | ~new_n1141_;
  assign new_n1180_ = ~new_n8290_ | ~new_n1144_;
  assign new_n1181_ = ~pi236 | ~new_n1141_;
  assign new_n1182_ = ~new_n8291_ | ~new_n1144_;
  assign new_n1183_ = ~pi235 | ~new_n1141_;
  assign new_n1184_ = ~new_n8292_ | ~new_n1144_;
  assign new_n1185_ = ~pi234 | ~new_n1141_;
  assign new_n1186_ = ~new_n8293_ | ~new_n1144_;
  assign new_n1187_ = ~pi233 | ~new_n1141_;
  assign new_n1188_ = ~new_n8294_ | ~new_n1144_;
  assign new_n1189_ = ~pi214 | ~new_n1141_;
  assign new_n1190_ = ~new_n8202_ | ~new_n1144_;
  assign new_n1191_ = ~pi232 | ~new_n1141_;
  assign new_n1192_ = ~new_n8295_ | ~new_n1144_;
  assign new_n1193_ = ~pi231 | ~new_n1141_;
  assign new_n1194_ = ~new_n8296_ | ~new_n1144_;
  assign new_n1195_ = ~pi230 | ~new_n1141_;
  assign new_n1196_ = ~new_n8297_ | ~new_n1144_;
  assign new_n1197_ = ~pi229 | ~new_n1141_;
  assign new_n1198_ = ~new_n8298_ | ~new_n1144_;
  assign new_n1199_ = ~pi228 | ~new_n1141_;
  assign new_n1200_ = ~new_n8299_ | ~new_n1144_;
  assign new_n1201_ = ~pi227 | ~new_n1141_;
  assign new_n1202_ = ~new_n8300_ | ~new_n1144_;
  assign new_n1203_ = ~pi226 | ~new_n1141_;
  assign new_n1204_ = ~new_n8301_ | ~new_n1144_;
  assign new_n1205_ = ~pi225 | ~new_n1141_;
  assign new_n1206_ = ~new_n8302_ | ~new_n1144_;
  assign new_n1207_ = ~pi224 | ~new_n1141_;
  assign new_n1208_ = ~new_n8303_ | ~new_n1144_;
  assign new_n1209_ = ~pi223 | ~new_n1141_;
  assign new_n1210_ = ~new_n8304_ | ~new_n1144_;
  assign new_n1211_ = ~pi213 | ~new_n1141_;
  assign new_n1212_ = ~new_n8275_ | ~new_n1144_;
  assign new_n1213_ = ~new_n8276_ | ~new_n1141_;
  assign new_n1214_ = ~pi467 | ~new_n1144_;
  assign new_n1215_ = ~new_n8277_ | ~new_n1141_;
  assign new_n1216_ = ~pi466 | ~new_n1144_;
  assign new_n1217_ = ~new_n8278_ | ~new_n1141_;
  assign new_n1218_ = ~pi465 | ~new_n1144_;
  assign new_n1219_ = ~new_n8279_ | ~new_n1141_;
  assign new_n1220_ = ~pi464 | ~new_n1144_;
  assign new_n1221_ = ~new_n8280_ | ~new_n1141_;
  assign new_n1222_ = ~pi463 | ~new_n1144_;
  assign new_n1223_ = ~new_n8281_ | ~new_n1141_;
  assign new_n1224_ = ~pi462 | ~new_n1144_;
  assign new_n1225_ = ~new_n8282_ | ~new_n1141_;
  assign new_n1226_ = ~pi461 | ~new_n1144_;
  assign new_n1227_ = ~new_n8203_ | ~new_n1141_;
  assign new_n1228_ = ~pi489 | ~new_n1144_;
  assign new_n1229_ = ~new_n8283_ | ~new_n1141_;
  assign new_n1230_ = ~pi488 | ~new_n1144_;
  assign new_n1231_ = ~new_n8284_ | ~new_n1141_;
  assign new_n1232_ = ~pi460 | ~new_n1144_;
  assign new_n1233_ = ~new_n8285_ | ~new_n1141_;
  assign new_n1234_ = ~pi487 | ~new_n1144_;
  assign new_n1235_ = ~new_n8286_ | ~new_n1141_;
  assign new_n1236_ = ~pi486 | ~new_n1144_;
  assign new_n1237_ = ~new_n8287_ | ~new_n1141_;
  assign new_n1238_ = ~pi485 | ~new_n1144_;
  assign new_n1239_ = ~new_n8288_ | ~new_n1141_;
  assign new_n1240_ = ~pi484 | ~new_n1144_;
  assign new_n1241_ = ~new_n8289_ | ~new_n1141_;
  assign new_n1242_ = ~pi483 | ~new_n1144_;
  assign new_n1243_ = ~new_n8290_ | ~new_n1141_;
  assign new_n1244_ = ~pi482 | ~new_n1144_;
  assign new_n1245_ = ~new_n8291_ | ~new_n1141_;
  assign new_n1246_ = ~pi481 | ~new_n1144_;
  assign new_n1247_ = ~new_n8292_ | ~new_n1141_;
  assign new_n1248_ = ~pi480 | ~new_n1144_;
  assign new_n1249_ = ~new_n8293_ | ~new_n1141_;
  assign new_n1250_ = ~pi479 | ~new_n1144_;
  assign new_n1251_ = ~new_n8294_ | ~new_n1141_;
  assign new_n1252_ = ~pi478 | ~new_n1144_;
  assign new_n1253_ = ~new_n8202_ | ~new_n1141_;
  assign new_n1254_ = ~pi459 | ~new_n1144_;
  assign new_n1255_ = ~new_n8295_ | ~new_n1141_;
  assign new_n1256_ = ~pi477 | ~new_n1144_;
  assign new_n1257_ = ~new_n8296_ | ~new_n1141_;
  assign new_n1258_ = ~pi476 | ~new_n1144_;
  assign new_n1259_ = ~new_n8297_ | ~new_n1141_;
  assign new_n1260_ = ~pi475 | ~new_n1144_;
  assign new_n1261_ = ~new_n8298_ | ~new_n1141_;
  assign new_n1262_ = ~pi474 | ~new_n1144_;
  assign new_n1263_ = ~new_n8299_ | ~new_n1141_;
  assign new_n1264_ = ~pi473 | ~new_n1144_;
  assign new_n1265_ = ~new_n8300_ | ~new_n1141_;
  assign new_n1266_ = ~pi472 | ~new_n1144_;
  assign new_n1267_ = ~new_n8301_ | ~new_n1141_;
  assign new_n1268_ = ~pi471 | ~new_n1144_;
  assign new_n1269_ = ~new_n8302_ | ~new_n1141_;
  assign new_n1270_ = ~pi470 | ~new_n1144_;
  assign new_n1271_ = ~new_n8303_ | ~new_n1141_;
  assign new_n1272_ = ~pi469 | ~new_n1144_;
  assign new_n1273_ = ~new_n8304_ | ~new_n1141_;
  assign new_n1274_ = ~pi468 | ~new_n1144_;
  assign new_n1275_ = ~new_n8275_ | ~new_n1141_;
  assign new_n1276_ = ~pi458 | ~new_n1144_;
  assign new_n1277_ = ~pi467 | ~new_n1141_;
  assign new_n1278_ = ~new_n1144_ | ~pi222;
  assign new_n1279_ = ~pi466 | ~new_n1141_;
  assign new_n1280_ = ~pi221 | ~new_n1144_;
  assign new_n1281_ = ~pi465 | ~new_n1141_;
  assign new_n1282_ = ~pi220 | ~new_n1144_;
  assign new_n1283_ = ~pi464 | ~new_n1141_;
  assign new_n1284_ = ~pi219 | ~new_n1144_;
  assign new_n1285_ = ~pi463 | ~new_n1141_;
  assign new_n1286_ = ~pi218 | ~new_n1144_;
  assign new_n1287_ = ~pi462 | ~new_n1141_;
  assign new_n1288_ = ~pi217 | ~new_n1144_;
  assign new_n1289_ = ~pi489 | ~new_n1141_;
  assign new_n1290_ = ~pi244 | ~new_n1144_;
  assign new_n1291_ = ~pi488 | ~new_n1141_;
  assign new_n1292_ = ~pi243 | ~new_n1144_;
  assign new_n1293_ = ~pi461 | ~new_n1141_;
  assign new_n1294_ = ~pi216 | ~new_n1144_;
  assign new_n1295_ = ~pi487 | ~new_n1141_;
  assign new_n1296_ = ~pi242 | ~new_n1144_;
  assign new_n1297_ = ~pi486 | ~new_n1141_;
  assign new_n1298_ = ~pi241 | ~new_n1144_;
  assign new_n1299_ = ~pi485 | ~new_n1141_;
  assign new_n1300_ = ~pi240 | ~new_n1144_;
  assign new_n1301_ = ~pi484 | ~new_n1141_;
  assign new_n1302_ = ~pi239 | ~new_n1144_;
  assign new_n1303_ = ~pi483 | ~new_n1141_;
  assign new_n1304_ = ~pi238 | ~new_n1144_;
  assign new_n1305_ = ~pi482 | ~new_n1141_;
  assign new_n1306_ = ~pi237 | ~new_n1144_;
  assign new_n1307_ = ~pi481 | ~new_n1141_;
  assign new_n1308_ = ~pi236 | ~new_n1144_;
  assign new_n1309_ = ~pi480 | ~new_n1141_;
  assign new_n1310_ = ~pi235 | ~new_n1144_;
  assign new_n1311_ = ~pi479 | ~new_n1141_;
  assign new_n1312_ = ~pi234 | ~new_n1144_;
  assign new_n1313_ = ~pi478 | ~new_n1141_;
  assign new_n1314_ = ~pi233 | ~new_n1144_;
  assign new_n1315_ = ~pi460 | ~new_n1141_;
  assign new_n1316_ = ~pi215 | ~new_n1144_;
  assign new_n1317_ = ~pi477 | ~new_n1141_;
  assign new_n1318_ = ~pi232 | ~new_n1144_;
  assign new_n1319_ = ~pi476 | ~new_n1141_;
  assign new_n1320_ = ~pi231 | ~new_n1144_;
  assign new_n1321_ = ~pi475 | ~new_n1141_;
  assign new_n1322_ = ~pi230 | ~new_n1144_;
  assign new_n1323_ = ~pi474 | ~new_n1141_;
  assign new_n1324_ = ~pi229 | ~new_n1144_;
  assign new_n1325_ = ~pi473 | ~new_n1141_;
  assign new_n1326_ = ~pi228 | ~new_n1144_;
  assign new_n1327_ = ~pi472 | ~new_n1141_;
  assign new_n1328_ = ~pi227 | ~new_n1144_;
  assign new_n1329_ = ~pi471 | ~new_n1141_;
  assign new_n1330_ = ~pi226 | ~new_n1144_;
  assign new_n1331_ = ~pi470 | ~new_n1141_;
  assign new_n1332_ = ~pi225 | ~new_n1144_;
  assign new_n1333_ = ~pi469 | ~new_n1141_;
  assign new_n1334_ = ~pi224 | ~new_n1144_;
  assign new_n1335_ = ~pi468 | ~new_n1141_;
  assign new_n1336_ = ~pi223 | ~new_n1144_;
  assign new_n1337_ = ~pi459 | ~new_n1141_;
  assign new_n1338_ = ~pi214 | ~new_n1144_;
  assign new_n1339_ = ~pi458 | ~new_n1141_;
  assign new_n1340_ = ~pi213 | ~new_n1144_;
  assign new_n1341_ = ~new_n5096_ | ~new_n20694_;
  assign new_n1342_ = ~new_n1343_ | ~new_n1344_;
  assign new_n1343_ = ~new_n4679_ | ~new_n20692_;
  assign new_n1344_ = ~new_n5099_ | ~new_n20693_;
  assign new_n1345_ = ~new_n20788_ | ~new_n20819_;
  assign new_n1346_ = ~new_n20894_ | ~new_n1347_;
  assign new_n1347_ = ~new_n20788_;
  assign new_n1348_ = ~new_n4688_ | ~new_n20696_;
  assign new_n1349_ = ~new_n5102_ | ~new_n20697_;
  assign new_n1350_ = ~new_n20787_ | ~new_n20818_;
  assign new_n1351_ = ~new_n20898_ | ~new_n1352_;
  assign new_n1352_ = ~new_n20787_;
  assign new_n1353_ = new_n2328_ & new_n1783_;
  assign new_n1354_ = new_n1789_ & new_n1786_;
  assign new_n1355_ = new_n1971_ & new_n1966_;
  assign new_n1356_ = new_n1784_ & new_n1785_;
  assign new_n1357_ = new_n4064_ & new_n1784_;
  assign new_n1358_ = new_n4061_ & new_n1785_;
  assign new_n1359_ = new_n4061_ & new_n4064_;
  assign new_n1360_ = new_n3739_ & new_n1760_;
  assign new_n1361_ = new_n1385_ & pi275;
  assign new_n1362_ = new_n1388_ & new_n4055_;
  assign new_n1363_ = new_n2156_ & new_n1762_;
  assign new_n1364_ = new_n2359_ & new_n4067_;
  assign new_n1365_ = new_n2325_ & new_n4055_;
  assign new_n1366_ = new_n2219_ & new_n2344_;
  assign new_n1367_ = new_n1695_ & pi275;
  assign new_n1368_ = new_n2336_ & new_n2361_;
  assign new_n1369_ = new_n2361_ & new_n1761_;
  assign new_n1370_ = new_n2329_ & new_n2361_;
  assign new_n1371_ = new_n2337_ & new_n2361_;
  assign new_n1372_ = new_n2359_ & new_n1786_;
  assign new_n1373_ = new_n2344_ & new_n4067_;
  assign new_n1374_ = new_n2361_ & new_n1364_;
  assign new_n1375_ = new_n2344_ & new_n1786_;
  assign new_n1376_ = new_n4073_ & new_n3252_;
  assign new_n1377_ = new_n1363_ & new_n4073_;
  assign new_n1378_ = new_n4067_ & new_n3252_;
  assign new_n1379_ = new_n1363_ & new_n4067_;
  assign new_n1380_ = new_n1354_ & new_n3252_;
  assign new_n1381_ = new_n1363_ & new_n1354_;
  assign new_n1382_ = new_n1361_ & new_n1762_;
  assign new_n1383_ = new_n3484_ & pi275;
  assign new_n1384_ = new_n1361_ & new_n3486_;
  assign new_n1385_ = new_n4042_ & new_n1760_;
  assign new_n1386_ = new_n1972_ & new_n1355_;
  assign new_n1387_ = new_n4055_ & new_n1782_;
  assign new_n1388_ = new_n4049_ & new_n4058_;
  assign new_n1389_ = new_n1775_ & new_n1777_;
  assign new_n1390_ = ~new_n3011_ | ~new_n3008_ | ~new_n3009_ | ~new_n3010_;
  assign new_n1391_ = ~new_n3030_ | ~new_n3027_ | ~new_n3028_ | ~new_n3029_;
  assign new_n1392_ = ~new_n3046_ | ~new_n3047_ | ~new_n3049_ | ~new_n3048_;
  assign new_n1393_ = ~new_n3085_ | ~new_n3086_ | ~new_n3087_;
  assign new_n1394_ = ~new_n2992_ | ~new_n2989_ | ~new_n2990_ | ~new_n2991_;
  assign new_n1395_ = ~new_n2973_ | ~new_n2970_ | ~new_n2971_ | ~new_n2972_;
  assign new_n1396_ = ~new_n3065_ | ~new_n3066_ | ~new_n3067_;
  assign new_n1397_ = ~new_n2571_ | ~new_n2572_ | ~new_n2574_ | ~new_n2573_;
  assign new_n1398_ = ~new_n2916_ | ~new_n2913_ | ~new_n2914_ | ~new_n2915_;
  assign new_n1399_ = ~new_n2688_ | ~new_n2685_ | ~new_n2686_ | ~new_n2687_;
  assign new_n1400_ = ~new_n2707_ | ~new_n2704_ | ~new_n2705_ | ~new_n2706_;
  assign new_n1401_ = ~new_n2552_ | ~new_n2553_ | ~new_n2555_ | ~new_n2554_;
  assign new_n1402_ = ~new_n2954_ | ~new_n2951_ | ~new_n2952_ | ~new_n2953_;
  assign new_n1403_ = ~new_n2935_ | ~new_n2932_ | ~new_n2933_ | ~new_n2934_;
  assign new_n1404_ = ~new_n2590_ | ~new_n2591_ | ~new_n2593_ | ~new_n2592_;
  assign new_n1405_ = ~new_n2528_ | ~new_n2529_ | ~new_n2531_ | ~new_n2530_;
  assign new_n1406_ = ~new_n2821_ | ~new_n2818_ | ~new_n2819_ | ~new_n2820_;
  assign new_n1407_ = ~new_n2628_ | ~new_n2629_ | ~new_n2631_ | ~new_n2630_;
  assign new_n1408_ = ~new_n2609_ | ~new_n2610_ | ~new_n2612_ | ~new_n2611_;
  assign new_n1409_ = ~new_n2726_ | ~new_n2723_ | ~new_n2724_ | ~new_n2725_;
  assign new_n1410_ = ~new_n2802_ | ~new_n2799_ | ~new_n2800_ | ~new_n2801_;
  assign new_n1411_ = ~new_n2783_ | ~new_n2780_ | ~new_n2781_ | ~new_n2782_;
  assign new_n1412_ = ~new_n2897_ | ~new_n2894_ | ~new_n2895_ | ~new_n2896_;
  assign new_n1413_ = ~new_n2878_ | ~new_n2875_ | ~new_n2876_ | ~new_n2877_;
  assign new_n1414_ = ~new_n2533_ | ~new_n2534_ | ~new_n2536_ | ~new_n2535_;
  assign new_n1415_ = ~new_n2509_ | ~new_n2510_ | ~new_n2512_ | ~new_n2511_;
  assign new_n1416_ = ~new_n2764_ | ~new_n2761_ | ~new_n2762_ | ~new_n2763_;
  assign new_n1417_ = ~new_n2745_ | ~new_n2742_ | ~new_n2743_ | ~new_n2744_;
  assign new_n1418_ = ~new_n2859_ | ~new_n2856_ | ~new_n2857_ | ~new_n2858_;
  assign new_n1419_ = ~new_n2840_ | ~new_n2837_ | ~new_n2838_ | ~new_n2839_;
  assign new_n1420_ = ~new_n2669_ | ~new_n2666_ | ~new_n2667_ | ~new_n2668_;
  assign new_n1421_ = ~new_n2647_ | ~new_n2648_ | ~new_n2650_ | ~new_n2649_;
  assign po265 = ~new_n3259_ | ~pi275;
  assign po264 = ~pi275;
  assign new_n1424_ = ~new_n3947_ | ~new_n3946_;
  assign new_n1425_ = ~new_n3949_ | ~new_n3948_;
  assign new_n1426_ = ~new_n3955_ | ~new_n3954_ | ~new_n3953_;
  assign new_n1427_ = ~new_n2262_ | ~new_n3957_;
  assign new_n1428_ = ~new_n2263_ | ~new_n3960_;
  assign new_n1429_ = ~new_n2264_ | ~new_n3963_;
  assign new_n1430_ = ~new_n2265_ | ~new_n3966_;
  assign new_n1431_ = ~new_n2266_ | ~new_n3969_;
  assign new_n1432_ = ~new_n2267_ | ~new_n3972_;
  assign new_n1433_ = ~new_n2268_ | ~new_n3975_;
  assign new_n1434_ = ~new_n2269_ | ~new_n3978_;
  assign new_n1435_ = ~new_n2270_ | ~new_n3981_;
  assign new_n1436_ = ~new_n2272_ | ~new_n3987_;
  assign new_n1437_ = ~new_n2273_ | ~new_n3990_;
  assign new_n1438_ = ~new_n2274_ | ~new_n3993_;
  assign new_n1439_ = ~new_n2275_ | ~new_n3996_;
  assign new_n1440_ = ~new_n2276_ | ~new_n3999_;
  assign new_n1441_ = ~new_n2277_ | ~new_n4002_;
  assign new_n1442_ = ~new_n2278_ | ~new_n4005_;
  assign new_n1443_ = ~new_n2279_ | ~new_n4008_;
  assign new_n1444_ = ~new_n2280_ | ~new_n4011_;
  assign new_n1445_ = ~new_n2281_ | ~new_n4014_;
  assign new_n1446_ = ~new_n3928_ | ~new_n3929_ | ~new_n3930_;
  assign new_n1447_ = ~new_n3931_ | ~new_n3932_ | ~new_n3933_;
  assign new_n1448_ = ~new_n3934_ | ~new_n3935_ | ~new_n3936_;
  assign new_n1449_ = ~new_n3937_ | ~new_n3938_ | ~new_n3939_;
  assign new_n1450_ = ~new_n3940_ | ~new_n3941_ | ~new_n3942_;
  assign new_n1451_ = ~new_n2260_ | ~new_n3944_;
  assign new_n1452_ = ~new_n2261_ | ~new_n3951_;
  assign new_n1453_ = ~new_n2271_ | ~new_n3984_;
  assign new_n1454_ = ~new_n2282_ | ~new_n4017_;
  assign new_n1455_ = ~new_n4020_ | ~new_n4019_;
  assign new_n1456_ = ~new_n3877_ | ~new_n3876_;
  assign new_n1457_ = ~new_n3879_ | ~new_n3878_;
  assign new_n1458_ = ~new_n2237_ | ~new_n3882_;
  assign new_n1459_ = ~new_n2238_ | ~new_n3884_;
  assign new_n1460_ = ~new_n2239_ | ~new_n3886_;
  assign new_n1461_ = ~new_n2240_ | ~new_n3888_;
  assign new_n1462_ = ~new_n2241_ | ~new_n3890_;
  assign new_n1463_ = ~new_n2242_ | ~new_n3892_;
  assign new_n1464_ = ~new_n2243_ | ~new_n3894_;
  assign new_n1465_ = ~new_n2244_ | ~new_n3896_;
  assign new_n1466_ = ~new_n2245_ | ~new_n3898_;
  assign new_n1467_ = ~new_n2246_ | ~new_n3900_;
  assign new_n1468_ = ~new_n2248_ | ~new_n3905_;
  assign new_n1469_ = ~new_n2249_ | ~new_n3907_;
  assign new_n1470_ = ~new_n2250_ | ~new_n3909_;
  assign new_n1471_ = ~new_n2251_ | ~new_n3911_;
  assign new_n1472_ = ~new_n2252_ | ~new_n3913_;
  assign new_n1473_ = ~new_n2253_ | ~new_n3915_;
  assign new_n1474_ = ~new_n2254_ | ~new_n3917_;
  assign new_n1475_ = ~new_n2255_ | ~new_n3919_;
  assign new_n1476_ = ~new_n2256_ | ~new_n3921_;
  assign new_n1477_ = ~new_n2257_ | ~new_n3923_;
  assign new_n1478_ = ~new_n3864_ | ~new_n3865_ | ~new_n1778_;
  assign new_n1479_ = ~new_n3866_ | ~new_n3867_ | ~new_n1778_;
  assign new_n1480_ = ~new_n3868_ | ~new_n3869_ | ~new_n1778_;
  assign new_n1481_ = ~new_n3870_ | ~new_n3871_ | ~new_n1778_;
  assign new_n1482_ = ~new_n3872_ | ~new_n3873_ | ~new_n1778_;
  assign new_n1483_ = ~new_n2235_ | ~new_n3875_;
  assign new_n1484_ = ~new_n2236_ | ~new_n3881_;
  assign new_n1485_ = ~new_n2247_ | ~new_n3903_;
  assign new_n1486_ = ~new_n2258_ | ~new_n3925_;
  assign new_n1487_ = ~new_n2259_ | ~new_n3927_;
  assign new_n1488_ = ~new_n2325_ | ~new_n1778_;
  assign new_n1489_ = ~new_n4042_ | ~new_n1710_;
  assign new_n1490_ = ~new_n3819_ | ~new_n3818_;
  assign new_n1491_ = ~new_n3821_ | ~new_n3820_;
  assign new_n1492_ = ~new_n3823_ | ~new_n3822_;
  assign new_n1493_ = ~new_n3825_ | ~new_n3824_;
  assign new_n1494_ = ~new_n3827_ | ~new_n3826_;
  assign new_n1495_ = ~new_n3829_ | ~new_n3828_;
  assign new_n1496_ = ~new_n3831_ | ~new_n3830_;
  assign new_n1497_ = ~new_n3833_ | ~new_n3832_;
  assign new_n1498_ = ~new_n3835_ | ~new_n3834_;
  assign new_n1499_ = ~new_n3839_ | ~new_n3838_;
  assign new_n1500_ = ~new_n3841_ | ~new_n3840_;
  assign new_n1501_ = ~new_n3843_ | ~new_n3842_;
  assign new_n1502_ = ~new_n3845_ | ~new_n3844_;
  assign new_n1503_ = ~new_n3847_ | ~new_n3846_;
  assign new_n1504_ = ~new_n3849_ | ~new_n3848_;
  assign new_n1505_ = ~new_n3851_ | ~new_n3850_;
  assign new_n1506_ = ~new_n3853_ | ~new_n3852_;
  assign new_n1507_ = ~new_n3855_ | ~new_n3854_;
  assign new_n1508_ = ~new_n3857_ | ~new_n3856_;
  assign new_n1509_ = ~new_n3805_ | ~new_n3804_;
  assign new_n1510_ = ~new_n3807_ | ~new_n3806_;
  assign new_n1511_ = ~new_n3809_ | ~new_n3808_;
  assign new_n1512_ = ~new_n3811_ | ~new_n3810_;
  assign new_n1513_ = ~new_n3813_ | ~new_n3812_;
  assign new_n1514_ = ~new_n3815_ | ~new_n3814_;
  assign new_n1515_ = ~new_n3817_ | ~new_n3816_;
  assign new_n1516_ = ~new_n3837_ | ~new_n3836_;
  assign new_n1517_ = ~new_n3859_ | ~new_n3858_;
  assign new_n1518_ = ~new_n2234_ | ~new_n3861_;
  assign new_n1519_ = ~new_n3760_ | ~new_n3759_;
  assign new_n1520_ = ~new_n3762_ | ~new_n3761_;
  assign new_n1521_ = ~new_n3764_ | ~new_n3763_;
  assign new_n1522_ = ~new_n3766_ | ~new_n3765_;
  assign new_n1523_ = ~new_n3768_ | ~new_n3767_;
  assign new_n1524_ = ~new_n3770_ | ~new_n3769_;
  assign new_n1525_ = ~new_n3772_ | ~new_n3771_;
  assign new_n1526_ = ~new_n3774_ | ~new_n3773_;
  assign new_n1527_ = ~new_n3776_ | ~new_n3775_;
  assign new_n1528_ = ~new_n3780_ | ~new_n3779_;
  assign new_n1529_ = ~new_n3782_ | ~new_n3781_;
  assign new_n1530_ = ~new_n3784_ | ~new_n3783_;
  assign new_n1531_ = ~new_n3786_ | ~new_n3785_;
  assign new_n1532_ = ~new_n3788_ | ~new_n3787_;
  assign new_n1533_ = ~new_n3790_ | ~new_n3789_;
  assign new_n1534_ = ~new_n3792_ | ~new_n3791_;
  assign new_n1535_ = ~new_n3794_ | ~new_n3793_;
  assign new_n1536_ = ~new_n3796_ | ~new_n3795_;
  assign new_n1537_ = ~new_n3798_ | ~new_n3797_;
  assign new_n1538_ = ~new_n3746_ | ~new_n3745_;
  assign new_n1539_ = ~new_n3748_ | ~new_n3747_;
  assign new_n1540_ = ~new_n3750_ | ~new_n3749_;
  assign new_n1541_ = ~new_n3752_ | ~new_n3751_;
  assign new_n1542_ = ~new_n3754_ | ~new_n3753_;
  assign new_n1543_ = ~new_n3756_ | ~new_n3755_;
  assign new_n1544_ = ~new_n3758_ | ~new_n3757_;
  assign new_n1545_ = ~new_n3778_ | ~new_n3777_;
  assign new_n1546_ = ~new_n3800_ | ~new_n3799_;
  assign new_n1547_ = ~new_n2233_ | ~new_n3801_;
  assign new_n1548_ = new_n3738_ & new_n1760_;
  assign new_n1549_ = ~new_n3736_ | ~new_n4605_ | ~new_n4604_;
  assign po263 = ~new_n3732_ | ~new_n3731_ | ~new_n3733_ | ~new_n3730_ | ~new_n3729_;
  assign po262 = ~new_n3723_ | ~new_n3722_ | ~new_n3724_ | ~new_n3721_ | ~new_n3720_;
  assign po261 = ~new_n3714_ | ~new_n3713_ | ~new_n3715_ | ~new_n3712_ | ~new_n3711_;
  assign po260 = ~new_n3705_ | ~new_n3704_ | ~new_n3706_ | ~new_n3703_ | ~new_n3702_;
  assign po259 = ~new_n3696_ | ~new_n3695_ | ~new_n3697_ | ~new_n3694_ | ~new_n3693_;
  assign po258 = ~new_n3686_ | ~new_n2230_ | ~new_n3685_;
  assign po257 = ~new_n3678_ | ~new_n3677_ | ~new_n3679_ | ~new_n3676_ | ~new_n3675_;
  assign po256 = ~new_n3669_ | ~new_n3668_ | ~new_n3670_ | ~new_n3667_ | ~new_n3666_;
  assign po255 = ~new_n3660_ | ~new_n3659_ | ~new_n3661_ | ~new_n3658_ | ~new_n3657_;
  assign po254 = ~new_n3650_ | ~new_n2228_ | ~new_n3649_;
  assign po253 = ~new_n3642_ | ~new_n3641_ | ~new_n3643_ | ~new_n3640_ | ~new_n3639_;
  assign po252 = ~new_n3633_ | ~new_n3632_ | ~new_n3634_ | ~new_n3631_ | ~new_n3630_;
  assign po251 = ~new_n3624_ | ~new_n3623_ | ~new_n3625_ | ~new_n3622_ | ~new_n3621_;
  assign po250 = ~new_n3615_ | ~new_n3614_ | ~new_n3616_ | ~new_n3613_ | ~new_n3612_;
  assign po249 = ~new_n2227_ | ~new_n3605_ | ~new_n3604_ | ~new_n3603_;
  assign po248 = ~new_n3597_ | ~new_n3596_ | ~new_n3598_ | ~new_n3595_ | ~new_n3594_;
  assign po247 = ~new_n3588_ | ~new_n3587_ | ~new_n3589_ | ~new_n3586_ | ~new_n3585_;
  assign po246 = ~new_n3578_ | ~new_n2225_ | ~new_n3577_;
  assign po245 = ~new_n3570_ | ~new_n3569_ | ~new_n3571_ | ~new_n3568_ | ~new_n3567_;
  assign po244 = ~new_n2223_ | ~new_n2224_ | ~new_n3560_;
  assign po243 = ~new_n3553_ | ~new_n3552_ | ~new_n3554_ | ~new_n3551_ | ~new_n3550_;
  assign po242 = ~new_n3544_ | ~new_n3543_ | ~new_n3545_ | ~new_n3542_ | ~new_n3541_;
  assign po241 = ~new_n3535_ | ~new_n3534_ | ~new_n3536_ | ~new_n3533_ | ~new_n3532_;
  assign po240 = ~new_n3526_ | ~new_n3525_ | ~new_n3527_ | ~new_n3524_ | ~new_n3523_;
  assign po239 = ~new_n3516_ | ~new_n2220_ | ~new_n3515_;
  assign po238 = ~new_n3508_ | ~new_n3507_ | ~new_n3509_ | ~new_n3506_ | ~new_n3505_;
  assign po237 = ~new_n3499_ | ~new_n3498_ | ~new_n3500_ | ~new_n3497_ | ~new_n3496_;
  assign po236 = ~new_n3490_ | ~new_n3489_ | ~new_n3491_ | ~new_n3488_ | ~new_n3487_;
  assign po235 = ~new_n3477_ | ~new_n3476_ | ~new_n3478_ | ~new_n3475_ | ~new_n3474_;
  assign po234 = new_n3459_ & new_n4021_;
  assign po201 = ~new_n2198_ | ~new_n2197_;
  assign po200 = ~new_n2196_ | ~new_n2195_;
  assign po199 = ~new_n2194_ | ~new_n2193_;
  assign po198 = ~new_n2191_ | ~new_n2190_;
  assign po197 = ~new_n2189_ | ~new_n2188_;
  assign po196 = ~new_n2186_ | ~new_n2185_;
  assign po195 = ~new_n2184_ | ~new_n2183_;
  assign po194 = ~new_n3382_ | ~new_n2181_ | ~new_n2182_;
  assign po193 = ~new_n3372_ | ~new_n2179_ | ~new_n2180_;
  assign po192 = ~new_n3362_ | ~new_n2177_ | ~new_n2178_;
  assign po191 = ~new_n3352_ | ~new_n2175_ | ~new_n2176_;
  assign po190 = ~new_n3342_ | ~new_n2173_ | ~new_n2174_;
  assign po189 = ~new_n3332_ | ~new_n2171_ | ~new_n2172_;
  assign po188 = ~new_n3322_ | ~new_n2169_ | ~new_n2170_;
  assign po187 = ~new_n3312_ | ~new_n2167_ | ~new_n2168_;
  assign po186 = ~new_n3302_ | ~new_n2165_ | ~new_n2166_;
  assign po185 = ~new_n3292_ | ~new_n2163_ | ~new_n2164_;
  assign po184 = ~new_n3282_ | ~new_n2161_ | ~new_n2162_;
  assign po183 = ~new_n3272_ | ~new_n2159_ | ~new_n2160_;
  assign po182 = ~new_n3262_ | ~new_n2157_ | ~new_n2158_;
  assign po181 = ~new_n3251_ | ~new_n2320_ | ~new_n3250_;
  assign po180 = ~new_n3249_ | ~new_n2319_ | ~new_n3248_;
  assign po178 = ~new_n2316_ | ~new_n3241_ | ~new_n2150_ | ~new_n2151_;
  assign po177 = ~new_n2315_ | ~new_n3236_ | ~new_n2148_ | ~new_n2149_;
  assign po176 = ~new_n2314_ | ~new_n3231_ | ~new_n2146_ | ~new_n2147_;
  assign po175 = ~new_n2313_ | ~new_n3226_ | ~new_n2144_ | ~new_n2145_;
  assign po174 = ~new_n2312_ | ~new_n3221_ | ~new_n2142_ | ~new_n2143_;
  assign po173 = ~new_n2311_ | ~new_n3216_ | ~new_n2140_ | ~new_n2141_;
  assign po172 = ~new_n2310_ | ~new_n3211_ | ~new_n2138_ | ~new_n2139_;
  assign po171 = ~new_n2309_ | ~new_n3206_ | ~new_n2136_ | ~new_n2137_;
  assign po170 = ~new_n2308_ | ~new_n3201_ | ~new_n2134_ | ~new_n2135_;
  assign po169 = ~new_n2307_ | ~new_n3196_ | ~new_n2132_ | ~new_n2133_;
  assign po168 = ~new_n2306_ | ~new_n2131_ | ~new_n2130_;
  assign po167 = ~new_n2305_ | ~new_n2129_ | ~new_n2128_;
  assign po166 = ~new_n2304_ | ~new_n3181_ | ~new_n2126_ | ~new_n2127_;
  assign po165 = ~new_n2303_ | ~new_n3176_ | ~new_n2124_ | ~new_n2125_;
  assign po164 = ~new_n2302_ | ~new_n2123_ | ~new_n2122_;
  assign po163 = ~new_n2301_ | ~new_n2121_ | ~new_n2120_;
  assign po162 = ~new_n2300_ | ~new_n2119_ | ~new_n2118_;
  assign po161 = ~new_n2299_ | ~new_n2117_ | ~new_n2116_;
  assign po160 = ~new_n2298_ | ~new_n3151_ | ~new_n2114_ | ~new_n2115_;
  assign po159 = ~new_n2297_ | ~new_n3146_ | ~new_n2112_ | ~new_n2113_;
  assign po158 = ~new_n2296_ | ~new_n2111_ | ~new_n2110_;
  assign po157 = ~new_n2295_ | ~new_n2109_ | ~new_n2108_;
  assign po156 = ~new_n2294_ | ~new_n2107_ | ~new_n2106_;
  assign po155 = ~new_n2293_ | ~new_n2105_ | ~new_n2104_;
  assign po154 = ~new_n2103_ | ~new_n2102_;
  assign po153 = ~new_n2101_ | ~new_n2100_;
  assign po152 = ~new_n2099_ | ~new_n2098_;
  assign po151 = ~new_n2097_ | ~new_n2096_;
  assign po150 = ~new_n2095_ | ~new_n2094_;
  assign po085 = pi096 & new_n2284_;
  assign po084 = pi095 & new_n2284_;
  assign po083 = pi094 & new_n2284_;
  assign po082 = pi093 & new_n2284_;
  assign po081 = pi092 & new_n2284_;
  assign po080 = pi091 & new_n2284_;
  assign po079 = pi090 & new_n2284_;
  assign po078 = pi089 & new_n2284_;
  assign po077 = pi088 & new_n2284_;
  assign po076 = pi087 & new_n2284_;
  assign po075 = pi086 & new_n2284_;
  assign po074 = pi085 & new_n2284_;
  assign po073 = pi084 & new_n2284_;
  assign po072 = pi083 & new_n2284_;
  assign po071 = pi082 & new_n2284_;
  assign po070 = pi081 & new_n2284_;
  assign po069 = pi080 & new_n2284_;
  assign po068 = pi079 & new_n2284_;
  assign po067 = pi078 & new_n2284_;
  assign po066 = pi077 & new_n2284_;
  assign po065 = pi076 & new_n2284_;
  assign po064 = pi075 & new_n2284_;
  assign po063 = pi074 & new_n2284_;
  assign po062 = pi073 & new_n2284_;
  assign po061 = pi072 & new_n2284_;
  assign po060 = pi071 & new_n2284_;
  assign po059 = pi070 & new_n2284_;
  assign po058 = pi069 & new_n2284_;
  assign po057 = pi068 & new_n2284_;
  assign po056 = pi067 & new_n2284_;
  assign po053 = ~new_n2470_ | ~new_n2471_ | ~new_n2472_;
  assign po052 = ~new_n2467_ | ~new_n2468_ | ~new_n2469_;
  assign po051 = ~new_n2464_ | ~new_n2465_ | ~new_n2466_;
  assign po050 = ~new_n2461_ | ~new_n2462_ | ~new_n2463_;
  assign po049 = ~new_n2458_ | ~new_n2459_ | ~new_n2460_;
  assign po048 = ~new_n2455_ | ~new_n2456_ | ~new_n2457_;
  assign po047 = ~new_n2452_ | ~new_n2453_ | ~new_n2454_;
  assign po046 = ~new_n2449_ | ~new_n2450_ | ~new_n2451_;
  assign po045 = ~new_n2446_ | ~new_n2447_ | ~new_n2448_;
  assign po044 = ~new_n2443_ | ~new_n2444_ | ~new_n2445_;
  assign po043 = ~new_n2440_ | ~new_n2441_ | ~new_n2442_;
  assign po042 = ~new_n2437_ | ~new_n2438_ | ~new_n2439_;
  assign po041 = ~new_n2434_ | ~new_n2435_ | ~new_n2436_;
  assign po040 = ~new_n2431_ | ~new_n2432_ | ~new_n2433_;
  assign po039 = ~new_n2428_ | ~new_n2429_ | ~new_n2430_;
  assign po038 = ~new_n2425_ | ~new_n2426_ | ~new_n2427_;
  assign po037 = ~new_n2422_ | ~new_n2423_ | ~new_n2424_;
  assign po036 = ~new_n2419_ | ~new_n2420_ | ~new_n2421_;
  assign po035 = ~new_n2416_ | ~new_n2417_ | ~new_n2418_;
  assign po034 = ~new_n2413_ | ~new_n2414_ | ~new_n2415_;
  assign po033 = ~new_n2410_ | ~new_n2411_ | ~new_n2412_;
  assign po032 = ~new_n2407_ | ~new_n2408_ | ~new_n2409_;
  assign po031 = ~new_n2404_ | ~new_n2405_ | ~new_n2406_;
  assign po030 = ~new_n2401_ | ~new_n2402_ | ~new_n2403_;
  assign po029 = ~new_n2398_ | ~new_n2399_ | ~new_n2400_;
  assign po028 = ~new_n2395_ | ~new_n2396_ | ~new_n2397_;
  assign po027 = ~new_n2392_ | ~new_n2393_ | ~new_n2394_;
  assign po026 = ~new_n2389_ | ~new_n2390_ | ~new_n2391_;
  assign po025 = ~new_n2386_ | ~new_n2387_ | ~new_n2388_;
  assign po024 = ~new_n2383_ | ~new_n2384_ | ~new_n2385_;
  assign po023 = ~new_n2380_ | ~new_n2381_ | ~new_n2382_;
  assign po022 = ~new_n2377_ | ~new_n2378_ | ~new_n2379_;
  assign new_n1693_ = new_n1782_ & new_n1778_;
  assign po179 = ~new_n2317_ | ~new_n3245_ | ~new_n3247_ | ~new_n3246_ | ~new_n3244_;
  assign new_n1695_ = ~pi275 | ~new_n2283_;
  assign new_n1696_ = ~new_n1777_ | ~new_n4034_;
  assign new_n1697_ = ~pi245;
  assign new_n1698_ = ~new_n1777_ | ~new_n4039_ | ~new_n4038_;
  assign new_n1699_ = ~new_n1387_ | ~new_n1783_;
  assign new_n1700_ = ~new_n1783_ | ~new_n1781_ | ~new_n1782_;
  assign new_n1701_ = ~new_n1781_ | ~new_n4052_;
  assign new_n1702_ = ~new_n2373_ | ~new_n1783_;
  assign new_n1703_ = ~new_n1787_ | ~new_n1781_ | ~new_n1782_;
  assign new_n1704_ = ~new_n2373_ | ~new_n1787_;
  assign new_n1705_ = ~new_n4055_ | ~new_n4052_;
  assign new_n1706_ = ~new_n2374_ | ~new_n1783_;
  assign new_n1707_ = ~new_n2332_ | ~new_n4058_;
  assign new_n1708_ = ~new_n2374_ | ~new_n1787_;
  assign new_n1709_ = ~new_n2328_ | ~new_n4049_;
  assign new_n1710_ = ~new_n4049_ | ~new_n1782_;
  assign new_n1711_ = ~new_n1783_ | ~new_n1787_;
  assign new_n1712_ = ~new_n1958_ | ~new_n1959_ | ~new_n2521_ | ~new_n2520_ | ~new_n2519_;
  assign new_n1713_ = ~pi161;
  assign new_n1714_ = ~new_n1976_ | ~new_n1974_ | ~new_n2539_ | ~new_n2538_;
  assign new_n1715_ = ~new_n1980_ | ~new_n1978_ | ~new_n2558_ | ~new_n2557_;
  assign new_n1716_ = ~new_n1984_ | ~new_n1982_ | ~new_n2577_ | ~new_n2576_;
  assign new_n1717_ = ~new_n1988_ | ~new_n1986_ | ~new_n2596_ | ~new_n2595_;
  assign new_n1718_ = ~new_n1992_ | ~new_n1990_ | ~new_n2615_ | ~new_n2614_;
  assign new_n1719_ = ~new_n1996_ | ~new_n1994_ | ~new_n2634_ | ~new_n2633_;
  assign new_n1720_ = ~new_n2000_ | ~new_n1998_ | ~new_n2653_ | ~new_n2652_;
  assign new_n1721_ = ~new_n2004_ | ~new_n2002_ | ~new_n2672_ | ~new_n2671_;
  assign new_n1722_ = ~new_n2008_ | ~new_n2006_ | ~new_n2691_ | ~new_n2690_;
  assign new_n1723_ = ~new_n2012_ | ~new_n2010_ | ~new_n2710_ | ~new_n2709_;
  assign new_n1724_ = ~new_n2016_ | ~new_n2014_ | ~new_n2729_ | ~new_n2728_;
  assign new_n1725_ = ~new_n2020_ | ~new_n2018_ | ~new_n2748_ | ~new_n2747_;
  assign new_n1726_ = ~new_n2024_ | ~new_n2022_ | ~new_n2767_ | ~new_n2766_;
  assign new_n1727_ = ~new_n2028_ | ~new_n2026_ | ~new_n2786_ | ~new_n2785_;
  assign new_n1728_ = ~new_n2032_ | ~new_n2030_ | ~new_n2805_ | ~new_n2804_;
  assign new_n1729_ = ~new_n2036_ | ~new_n2034_ | ~new_n2824_ | ~new_n2823_;
  assign new_n1730_ = ~new_n2040_ | ~new_n2038_ | ~new_n2843_ | ~new_n2842_;
  assign new_n1731_ = ~new_n2044_ | ~new_n2042_ | ~new_n2862_ | ~new_n2861_;
  assign new_n1732_ = ~new_n2048_ | ~new_n2046_ | ~new_n2881_ | ~new_n2880_;
  assign new_n1733_ = ~new_n1090_ | ~new_n2285_;
  assign new_n1734_ = ~new_n2052_ | ~new_n2050_ | ~new_n2900_ | ~new_n2899_;
  assign new_n1735_ = ~new_n1089_ | ~new_n2285_;
  assign new_n1736_ = ~new_n2056_ | ~new_n2054_ | ~new_n2919_ | ~new_n2918_;
  assign new_n1737_ = ~new_n1088_ | ~new_n2285_;
  assign new_n1738_ = ~new_n2060_ | ~new_n2058_ | ~new_n2938_ | ~new_n2937_;
  assign new_n1739_ = ~new_n1087_ | ~new_n2285_;
  assign new_n1740_ = ~new_n2064_ | ~new_n2062_ | ~new_n2957_ | ~new_n2956_;
  assign new_n1741_ = ~new_n1086_ | ~new_n2285_;
  assign new_n1742_ = ~new_n2068_ | ~new_n2066_ | ~new_n2976_ | ~new_n2975_;
  assign new_n1743_ = ~new_n1085_ | ~new_n2285_;
  assign new_n1744_ = ~new_n2072_ | ~new_n2070_ | ~new_n2995_ | ~new_n2994_;
  assign new_n1745_ = ~new_n1084_ | ~new_n2285_;
  assign new_n1746_ = ~new_n2076_ | ~new_n2074_ | ~new_n3014_ | ~new_n3013_;
  assign new_n1747_ = ~new_n1083_ | ~new_n2285_;
  assign new_n1748_ = ~new_n2080_ | ~new_n2078_ | ~new_n3033_ | ~new_n3032_;
  assign new_n1749_ = ~new_n1082_ | ~new_n2285_;
  assign new_n1750_ = ~new_n2084_ | ~new_n2082_ | ~new_n3052_ | ~new_n3051_;
  assign new_n1751_ = ~new_n1081_ | ~new_n2285_;
  assign new_n1752_ = ~new_n2089_ | ~new_n2087_;
  assign new_n1753_ = ~new_n1079_ | ~new_n2285_;
  assign new_n1754_ = ~new_n1078_ | ~new_n2285_;
  assign new_n1755_ = ~new_n2325_ | ~new_n4058_;
  assign new_n1756_ = ~new_n1361_ | ~new_n3096_;
  assign new_n1757_ = ~new_n2360_ | ~new_n4055_;
  assign new_n1758_ = ~new_n1387_ | ~new_n1787_;
  assign new_n1759_ = ~new_n1362_ | ~new_n4052_;
  assign new_n1760_ = ~new_n1389_ | ~new_n1776_;
  assign new_n1761_ = ~new_n2338_ | ~new_n3097_;
  assign new_n1762_ = ~new_n1763_ | ~new_n3260_;
  assign new_n1763_ = ~new_n2474_ | ~new_n4042_;
  assign new_n1764_ = ~new_n2371_ | ~pi275;
  assign new_n1765_ = ~new_n1783_ | ~new_n1778_;
  assign new_n1766_ = ~new_n1353_ | ~new_n1354_;
  assign new_n1767_ = ~new_n1778_ | ~new_n4052_;
  assign new_n1768_ = ~new_n10877_;
  assign new_n1769_ = ~new_n1361_ | ~new_n1761_;
  assign new_n1770_ = ~new_n2215_ | ~new_n1355_;
  assign new_n1771_ = ~new_n1353_ | ~new_n1361_;
  assign new_n1772_ = ~new_n2218_ | ~new_n3472_;
  assign new_n1773_ = ~new_n1782_ | ~new_n4058_;
  assign new_n1774_ = ~new_n3742_ | ~new_n3741_;
  assign new_n1775_ = ~new_n4030_ | ~new_n4029_;
  assign new_n1776_ = ~new_n4033_ | ~new_n4032_;
  assign new_n1777_ = ~new_n4036_ | ~new_n4035_;
  assign new_n1778_ = ~new_n4041_ | ~new_n4040_;
  assign po054 = ~new_n4044_ | ~new_n4043_;
  assign po055 = ~new_n4046_ | ~new_n4045_;
  assign new_n1781_ = ~new_n4054_ | ~new_n4053_;
  assign new_n1782_ = ~new_n4051_ | ~new_n4050_;
  assign new_n1783_ = ~new_n4048_ | ~new_n4047_;
  assign new_n1784_ = ~new_n4060_ | ~new_n4059_;
  assign new_n1785_ = ~new_n4063_ | ~new_n4062_;
  assign new_n1786_ = ~new_n4066_ | ~new_n4065_;
  assign new_n1787_ = ~new_n4057_ | ~new_n4056_;
  assign new_n1788_ = ~new_n4069_ | ~new_n4068_;
  assign new_n1789_ = ~new_n4072_ | ~new_n4071_;
  assign new_n1790_ = ~new_n4075_ | ~new_n4074_;
  assign new_n1791_ = ~new_n4083_ | ~new_n4082_;
  assign new_n1792_ = ~new_n4080_ | ~new_n4079_;
  assign po086 = ~new_n4086_ | ~new_n4085_;
  assign new_n1794_ = ~new_n4088_ | ~new_n4087_;
  assign new_n1795_ = ~new_n4090_ | ~new_n4089_;
  assign po087 = ~new_n4093_ | ~new_n4092_;
  assign new_n1797_ = ~new_n4095_ | ~new_n4094_;
  assign new_n1798_ = ~new_n4097_ | ~new_n4096_;
  assign po088 = ~new_n4100_ | ~new_n4099_;
  assign new_n1800_ = ~new_n4102_ | ~new_n4101_;
  assign new_n1801_ = ~new_n4104_ | ~new_n4103_;
  assign po089 = ~new_n4107_ | ~new_n4106_;
  assign new_n1803_ = ~new_n4109_ | ~new_n4108_;
  assign new_n1804_ = ~new_n4111_ | ~new_n4110_;
  assign po090 = ~new_n4114_ | ~new_n4113_;
  assign new_n1806_ = ~new_n4116_ | ~new_n4115_;
  assign new_n1807_ = ~new_n4118_ | ~new_n4117_;
  assign po091 = ~new_n4121_ | ~new_n4120_;
  assign new_n1809_ = ~new_n4123_ | ~new_n4122_;
  assign new_n1810_ = ~new_n4125_ | ~new_n4124_;
  assign po092 = ~new_n4128_ | ~new_n4127_;
  assign new_n1812_ = ~new_n4130_ | ~new_n4129_;
  assign new_n1813_ = ~new_n4132_ | ~new_n4131_;
  assign po093 = ~new_n4135_ | ~new_n4134_;
  assign new_n1815_ = ~new_n4137_ | ~new_n4136_;
  assign new_n1816_ = ~new_n4139_ | ~new_n4138_;
  assign po094 = ~new_n4142_ | ~new_n4141_;
  assign new_n1818_ = ~new_n4144_ | ~new_n4143_;
  assign new_n1819_ = ~new_n4146_ | ~new_n4145_;
  assign po095 = ~new_n4149_ | ~new_n4148_;
  assign new_n1821_ = ~new_n4151_ | ~new_n4150_;
  assign new_n1822_ = ~new_n4153_ | ~new_n4152_;
  assign po096 = ~new_n4156_ | ~new_n4155_;
  assign new_n1824_ = ~new_n4158_ | ~new_n4157_;
  assign new_n1825_ = ~new_n4160_ | ~new_n4159_;
  assign po097 = ~new_n4163_ | ~new_n4162_;
  assign new_n1827_ = ~new_n4165_ | ~new_n4164_;
  assign new_n1828_ = ~new_n4167_ | ~new_n4166_;
  assign po098 = ~new_n4170_ | ~new_n4169_;
  assign new_n1830_ = ~new_n4172_ | ~new_n4171_;
  assign new_n1831_ = ~new_n4174_ | ~new_n4173_;
  assign po099 = ~new_n4177_ | ~new_n4176_;
  assign new_n1833_ = ~new_n4179_ | ~new_n4178_;
  assign new_n1834_ = ~new_n4181_ | ~new_n4180_;
  assign po100 = ~new_n4184_ | ~new_n4183_;
  assign new_n1836_ = ~new_n4186_ | ~new_n4185_;
  assign new_n1837_ = ~new_n4188_ | ~new_n4187_;
  assign po101 = ~new_n4191_ | ~new_n4190_;
  assign new_n1839_ = ~new_n4193_ | ~new_n4192_;
  assign new_n1840_ = ~new_n4195_ | ~new_n4194_;
  assign po102 = ~new_n4198_ | ~new_n4197_;
  assign new_n1842_ = ~new_n4200_ | ~new_n4199_;
  assign new_n1843_ = ~new_n4202_ | ~new_n4201_;
  assign po103 = ~new_n4205_ | ~new_n4204_;
  assign new_n1845_ = ~new_n4207_ | ~new_n4206_;
  assign new_n1846_ = ~new_n4209_ | ~new_n4208_;
  assign po104 = ~new_n4212_ | ~new_n4211_;
  assign new_n1848_ = ~new_n4214_ | ~new_n4213_;
  assign po105 = ~new_n4217_ | ~new_n4216_;
  assign po106 = ~new_n4219_ | ~new_n4218_;
  assign po107 = ~new_n4221_ | ~new_n4220_;
  assign po108 = ~new_n4223_ | ~new_n4222_;
  assign po109 = ~new_n4225_ | ~new_n4224_;
  assign po110 = ~new_n4227_ | ~new_n4226_;
  assign po111 = ~new_n4229_ | ~new_n4228_;
  assign po112 = ~new_n4231_ | ~new_n4230_;
  assign po113 = ~new_n4233_ | ~new_n4232_;
  assign po114 = ~new_n4235_ | ~new_n4234_;
  assign po115 = ~new_n4237_ | ~new_n4236_;
  assign po116 = ~new_n4239_ | ~new_n4238_;
  assign po117 = ~new_n4241_ | ~new_n4240_;
  assign po118 = ~new_n4243_ | ~new_n4242_;
  assign po119 = ~new_n4245_ | ~new_n4244_;
  assign po120 = ~new_n4247_ | ~new_n4246_;
  assign po121 = ~new_n4249_ | ~new_n4248_;
  assign po122 = ~new_n4251_ | ~new_n4250_;
  assign po123 = ~new_n4253_ | ~new_n4252_;
  assign po124 = ~new_n4255_ | ~new_n4254_;
  assign po125 = ~new_n4257_ | ~new_n4256_;
  assign po126 = ~new_n4259_ | ~new_n4258_;
  assign po127 = ~new_n4261_ | ~new_n4260_;
  assign po128 = ~new_n4263_ | ~new_n4262_;
  assign po129 = ~new_n4265_ | ~new_n4264_;
  assign po130 = ~new_n4267_ | ~new_n4266_;
  assign po131 = ~new_n4269_ | ~new_n4268_;
  assign po132 = ~new_n4271_ | ~new_n4270_;
  assign po133 = ~new_n4273_ | ~new_n4272_;
  assign po134 = ~new_n4275_ | ~new_n4274_;
  assign po135 = ~new_n4277_ | ~new_n4276_;
  assign po136 = ~new_n4279_ | ~new_n4278_;
  assign po137 = ~new_n4281_ | ~new_n4280_;
  assign po138 = ~new_n4283_ | ~new_n4282_;
  assign po139 = ~new_n4285_ | ~new_n4284_;
  assign po140 = ~new_n4287_ | ~new_n4286_;
  assign po141 = ~new_n4289_ | ~new_n4288_;
  assign po142 = ~new_n4291_ | ~new_n4290_;
  assign po143 = ~new_n4293_ | ~new_n4292_;
  assign po144 = ~new_n4295_ | ~new_n4294_;
  assign po145 = ~new_n4297_ | ~new_n4296_;
  assign po146 = ~new_n4299_ | ~new_n4298_;
  assign po147 = ~new_n4301_ | ~new_n4300_;
  assign po148 = ~new_n4303_ | ~new_n4302_;
  assign po149 = ~new_n4305_ | ~new_n4304_;
  assign po202 = ~new_n4371_ | ~new_n4370_;
  assign po203 = ~new_n4373_ | ~new_n4372_;
  assign po204 = ~new_n4375_ | ~new_n4374_;
  assign po205 = ~new_n4377_ | ~new_n4376_;
  assign po206 = ~new_n4379_ | ~new_n4378_;
  assign po207 = ~new_n4381_ | ~new_n4380_;
  assign po208 = ~new_n4383_ | ~new_n4382_;
  assign po209 = ~new_n4385_ | ~new_n4384_;
  assign po210 = ~new_n4387_ | ~new_n4386_;
  assign po211 = ~new_n4389_ | ~new_n4388_;
  assign po212 = ~new_n4391_ | ~new_n4390_;
  assign po213 = ~new_n4393_ | ~new_n4392_;
  assign po214 = ~new_n4395_ | ~new_n4394_;
  assign po215 = ~new_n4397_ | ~new_n4396_;
  assign po216 = ~new_n4399_ | ~new_n4398_;
  assign po217 = ~new_n4401_ | ~new_n4400_;
  assign po218 = ~new_n4403_ | ~new_n4402_;
  assign po219 = ~new_n4405_ | ~new_n4404_;
  assign po220 = ~new_n4407_ | ~new_n4406_;
  assign po221 = ~new_n4409_ | ~new_n4408_;
  assign po222 = ~new_n4411_ | ~new_n4410_;
  assign po223 = ~new_n4413_ | ~new_n4412_;
  assign po224 = ~new_n4415_ | ~new_n4414_;
  assign po225 = ~new_n4417_ | ~new_n4416_;
  assign po226 = ~new_n4419_ | ~new_n4418_;
  assign po227 = ~new_n4421_ | ~new_n4420_;
  assign po228 = ~new_n4423_ | ~new_n4422_;
  assign po229 = ~new_n4425_ | ~new_n4424_;
  assign po230 = ~new_n4427_ | ~new_n4426_;
  assign po231 = ~new_n4429_ | ~new_n4428_;
  assign po232 = ~new_n4431_ | ~new_n4430_;
  assign po233 = ~new_n4433_ | ~new_n4432_;
  assign new_n1926_ = ~new_n4541_ | ~new_n4540_;
  assign new_n1927_ = ~new_n4543_ | ~new_n4542_;
  assign new_n1928_ = ~new_n4545_ | ~new_n4544_;
  assign new_n1929_ = ~new_n4547_ | ~new_n4546_;
  assign new_n1930_ = ~new_n4549_ | ~new_n4548_;
  assign new_n1931_ = ~new_n4551_ | ~new_n4550_;
  assign new_n1932_ = ~new_n4553_ | ~new_n4552_;
  assign new_n1933_ = ~new_n4555_ | ~new_n4554_;
  assign new_n1934_ = ~new_n4557_ | ~new_n4556_;
  assign new_n1935_ = ~new_n4559_ | ~new_n4558_;
  assign new_n1936_ = ~new_n4561_ | ~new_n4560_;
  assign new_n1937_ = ~new_n4563_ | ~new_n4562_;
  assign new_n1938_ = ~new_n4565_ | ~new_n4564_;
  assign new_n1939_ = ~new_n4567_ | ~new_n4566_;
  assign new_n1940_ = ~new_n4569_ | ~new_n4568_;
  assign new_n1941_ = ~new_n4571_ | ~new_n4570_;
  assign new_n1942_ = ~new_n4573_ | ~new_n4572_;
  assign new_n1943_ = ~new_n4575_ | ~new_n4574_;
  assign new_n1944_ = ~new_n4577_ | ~new_n4576_;
  assign new_n1945_ = ~new_n4579_ | ~new_n4578_;
  assign new_n1946_ = ~new_n4581_ | ~new_n4580_;
  assign new_n1947_ = ~new_n4583_ | ~new_n4582_;
  assign new_n1948_ = ~new_n4585_ | ~new_n4584_;
  assign new_n1949_ = ~new_n4587_ | ~new_n4586_;
  assign new_n1950_ = ~new_n4589_ | ~new_n4588_;
  assign new_n1951_ = ~new_n4591_ | ~new_n4590_;
  assign new_n1952_ = ~new_n4593_ | ~new_n4592_;
  assign new_n1953_ = ~new_n4595_ | ~new_n4594_;
  assign new_n1954_ = ~new_n4597_ | ~new_n4596_;
  assign new_n1955_ = ~new_n4599_ | ~new_n4598_;
  assign new_n1956_ = ~new_n4601_ | ~new_n4600_;
  assign new_n1957_ = ~new_n4603_ | ~new_n4602_;
  assign new_n1958_ = new_n2516_ & new_n2515_;
  assign new_n1959_ = new_n2518_ & new_n2517_;
  assign new_n1960_ = new_n2525_ & new_n2523_;
  assign new_n1961_ = new_n1960_ & new_n2526_ & new_n2524_;
  assign new_n1962_ = new_n2477_ & new_n2478_ & new_n2480_ & new_n2479_;
  assign new_n1963_ = new_n2481_ & new_n2482_ & new_n2484_ & new_n2483_;
  assign new_n1964_ = new_n2485_ & new_n2486_ & new_n2488_ & new_n2487_;
  assign new_n1965_ = new_n2491_ & new_n2490_ & new_n2489_;
  assign new_n1966_ = new_n1962_ & new_n1963_ & new_n1965_ & new_n1964_;
  assign new_n1967_ = new_n2492_ & new_n2493_ & new_n2495_ & new_n2494_;
  assign new_n1968_ = new_n2496_ & new_n2497_ & new_n2499_ & new_n2498_;
  assign new_n1969_ = new_n2500_ & new_n2501_ & new_n2503_ & new_n2502_;
  assign new_n1970_ = new_n2506_ & new_n2505_ & new_n2504_;
  assign new_n1971_ = new_n1967_ & new_n1968_ & new_n1970_ & new_n1969_;
  assign new_n1972_ = new_n4081_ & new_n2508_;
  assign new_n1973_ = new_n4084_ & new_n1361_;
  assign new_n1974_ = new_n2541_ & new_n2540_;
  assign new_n1975_ = new_n2543_ & new_n2542_;
  assign new_n1976_ = new_n1975_ & new_n2545_ & new_n2544_;
  assign new_n1977_ = new_n2547_ & new_n2550_ & new_n2548_ & new_n2549_;
  assign new_n1978_ = new_n2560_ & new_n2559_;
  assign new_n1979_ = new_n2562_ & new_n2561_;
  assign new_n1980_ = new_n1979_ & new_n2564_ & new_n2563_;
  assign new_n1981_ = new_n2566_ & new_n2569_ & new_n2567_ & new_n2568_;
  assign new_n1982_ = new_n2579_ & new_n2578_;
  assign new_n1983_ = new_n2581_ & new_n2580_;
  assign new_n1984_ = new_n1983_ & new_n2583_ & new_n2582_;
  assign new_n1985_ = new_n2585_ & new_n2588_ & new_n2586_ & new_n2587_;
  assign new_n1986_ = new_n2598_ & new_n2597_;
  assign new_n1987_ = new_n2600_ & new_n2599_;
  assign new_n1988_ = new_n1987_ & new_n2602_ & new_n2601_;
  assign new_n1989_ = new_n2604_ & new_n2607_ & new_n2605_ & new_n2606_;
  assign new_n1990_ = new_n2617_ & new_n2616_;
  assign new_n1991_ = new_n2619_ & new_n2618_;
  assign new_n1992_ = new_n1991_ & new_n2621_ & new_n2620_;
  assign new_n1993_ = new_n2623_ & new_n2626_ & new_n2624_ & new_n2625_;
  assign new_n1994_ = new_n2636_ & new_n2635_;
  assign new_n1995_ = new_n2638_ & new_n2637_;
  assign new_n1996_ = new_n1995_ & new_n2640_ & new_n2639_;
  assign new_n1997_ = new_n2642_ & new_n2645_ & new_n2643_ & new_n2644_;
  assign new_n1998_ = new_n2655_ & new_n2654_;
  assign new_n1999_ = new_n2657_ & new_n2656_;
  assign new_n2000_ = new_n1999_ & new_n2659_ & new_n2658_;
  assign new_n2001_ = new_n2661_ & new_n2664_ & new_n2662_ & new_n2663_;
  assign new_n2002_ = new_n2674_ & new_n2673_;
  assign new_n2003_ = new_n2676_ & new_n2675_;
  assign new_n2004_ = new_n2003_ & new_n2678_ & new_n2677_;
  assign new_n2005_ = new_n2680_ & new_n2683_ & new_n2681_ & new_n2682_;
  assign new_n2006_ = new_n2693_ & new_n2692_;
  assign new_n2007_ = new_n2695_ & new_n2694_;
  assign new_n2008_ = new_n2007_ & new_n2697_ & new_n2696_;
  assign new_n2009_ = new_n2699_ & new_n2702_ & new_n2700_ & new_n2701_;
  assign new_n2010_ = new_n2712_ & new_n2711_;
  assign new_n2011_ = new_n2714_ & new_n2713_;
  assign new_n2012_ = new_n2011_ & new_n2716_ & new_n2715_;
  assign new_n2013_ = new_n2718_ & new_n2721_ & new_n2719_ & new_n2720_;
  assign new_n2014_ = new_n2731_ & new_n2730_;
  assign new_n2015_ = new_n2733_ & new_n2732_;
  assign new_n2016_ = new_n2015_ & new_n2735_ & new_n2734_;
  assign new_n2017_ = new_n2737_ & new_n2738_ & new_n2740_ & new_n2739_;
  assign new_n2018_ = new_n2750_ & new_n2749_;
  assign new_n2019_ = new_n2752_ & new_n2751_;
  assign new_n2020_ = new_n2019_ & new_n2754_ & new_n2753_;
  assign new_n2021_ = new_n2756_ & new_n2757_ & new_n2759_ & new_n2758_;
  assign new_n2022_ = new_n2769_ & new_n2768_;
  assign new_n2023_ = new_n2771_ & new_n2770_;
  assign new_n2024_ = new_n2023_ & new_n2773_ & new_n2772_;
  assign new_n2025_ = new_n2775_ & new_n2776_ & new_n2778_ & new_n2777_;
  assign new_n2026_ = new_n2788_ & new_n2787_;
  assign new_n2027_ = new_n2790_ & new_n2789_;
  assign new_n2028_ = new_n2027_ & new_n2792_ & new_n2791_;
  assign new_n2029_ = new_n2796_ & new_n2795_ & new_n2797_ & new_n2794_;
  assign new_n2030_ = new_n2807_ & new_n2806_;
  assign new_n2031_ = new_n2809_ & new_n2808_;
  assign new_n2032_ = new_n2031_ & new_n2811_ & new_n2810_;
  assign new_n2033_ = new_n2813_ & new_n2816_ & new_n2814_ & new_n2815_;
  assign new_n2034_ = new_n2826_ & new_n2825_;
  assign new_n2035_ = new_n2828_ & new_n2827_;
  assign new_n2036_ = new_n2035_ & new_n2830_ & new_n2829_;
  assign new_n2037_ = new_n2832_ & new_n2835_ & new_n2833_ & new_n2834_;
  assign new_n2038_ = new_n2845_ & new_n2844_;
  assign new_n2039_ = new_n2847_ & new_n2846_;
  assign new_n2040_ = new_n2039_ & new_n2849_ & new_n2848_;
  assign new_n2041_ = new_n2853_ & new_n2852_ & new_n2854_ & new_n2851_;
  assign new_n2042_ = new_n2864_ & new_n2863_;
  assign new_n2043_ = new_n2866_ & new_n2865_;
  assign new_n2044_ = new_n2043_ & new_n2868_ & new_n2867_;
  assign new_n2045_ = new_n2872_ & new_n2871_ & new_n2873_ & new_n2870_;
  assign new_n2046_ = new_n2883_ & new_n2882_;
  assign new_n2047_ = new_n2885_ & new_n2884_;
  assign new_n2048_ = new_n2047_ & new_n2887_ & new_n2886_;
  assign new_n2049_ = new_n2889_ & new_n2892_ & new_n2890_ & new_n2891_;
  assign new_n2050_ = new_n2902_ & new_n2901_;
  assign new_n2051_ = new_n2904_ & new_n2903_;
  assign new_n2052_ = new_n2051_ & new_n2906_ & new_n2905_;
  assign new_n2053_ = new_n2908_ & new_n2911_ & new_n2909_ & new_n2910_;
  assign new_n2054_ = new_n2921_ & new_n2920_;
  assign new_n2055_ = new_n2923_ & new_n2922_;
  assign new_n2056_ = new_n2055_ & new_n2925_ & new_n2924_;
  assign new_n2057_ = new_n2927_ & new_n2930_ & new_n2928_ & new_n2929_;
  assign new_n2058_ = new_n2940_ & new_n2939_;
  assign new_n2059_ = new_n2942_ & new_n2941_;
  assign new_n2060_ = new_n2059_ & new_n2944_ & new_n2943_;
  assign new_n2061_ = new_n2946_ & new_n2949_ & new_n2947_ & new_n2948_;
  assign new_n2062_ = new_n2959_ & new_n2958_;
  assign new_n2063_ = new_n2961_ & new_n2960_;
  assign new_n2064_ = new_n2063_ & new_n2963_ & new_n2962_;
  assign new_n2065_ = new_n2965_ & new_n2968_ & new_n2966_ & new_n2967_;
  assign new_n2066_ = new_n2978_ & new_n2977_;
  assign new_n2067_ = new_n2980_ & new_n2979_;
  assign new_n2068_ = new_n2067_ & new_n2982_ & new_n2981_;
  assign new_n2069_ = new_n2984_ & new_n2987_ & new_n2985_ & new_n2986_;
  assign new_n2070_ = new_n2997_ & new_n2996_;
  assign new_n2071_ = new_n2999_ & new_n2998_;
  assign new_n2072_ = new_n2071_ & new_n3001_ & new_n3000_;
  assign new_n2073_ = new_n3003_ & new_n3006_ & new_n3004_ & new_n3005_;
  assign new_n2074_ = new_n3016_ & new_n3015_;
  assign new_n2075_ = new_n3018_ & new_n3017_;
  assign new_n2076_ = new_n2075_ & new_n3020_ & new_n3019_;
  assign new_n2077_ = new_n3022_ & new_n3025_ & new_n3023_ & new_n3024_;
  assign new_n2078_ = new_n3035_ & new_n3034_;
  assign new_n2079_ = new_n3037_ & new_n3036_;
  assign new_n2080_ = new_n2079_ & new_n3039_ & new_n3038_;
  assign new_n2081_ = new_n3041_ & new_n3044_ & new_n3042_ & new_n3043_;
  assign new_n2082_ = new_n3054_ & new_n3053_;
  assign new_n2083_ = new_n3056_ & new_n3055_;
  assign new_n2084_ = new_n2083_ & new_n3058_ & new_n3057_;
  assign new_n2085_ = new_n3060_ & new_n3063_ & new_n3061_ & new_n3062_;
  assign new_n2086_ = new_n3070_ & new_n2359_;
  assign new_n2087_ = new_n3075_ & new_n3074_ & new_n3073_ & new_n3072_ & new_n3071_;
  assign new_n2088_ = new_n3077_ & new_n3076_;
  assign new_n2089_ = new_n2088_ & new_n3079_ & new_n3078_;
  assign new_n2090_ = new_n3081_ & new_n3082_ & new_n3083_;
  assign new_n2091_ = new_n2359_ & new_n3070_;
  assign new_n2092_ = new_n1361_ & new_n1791_;
  assign new_n2093_ = new_n1792_ & new_n4084_ & new_n2341_;
  assign new_n2094_ = new_n3101_ & new_n3100_ & new_n3099_;
  assign new_n2095_ = new_n2288_ & new_n3103_ & new_n3102_;
  assign new_n2096_ = new_n3106_ & new_n3105_ & new_n3104_;
  assign new_n2097_ = new_n2289_ & new_n3108_ & new_n3107_;
  assign new_n2098_ = new_n3111_ & new_n3110_ & new_n3109_;
  assign new_n2099_ = new_n2290_ & new_n3113_ & new_n3112_;
  assign new_n2100_ = new_n3116_ & new_n3115_ & new_n3114_;
  assign new_n2101_ = new_n2291_ & new_n3118_ & new_n3117_;
  assign new_n2102_ = new_n3121_ & new_n3120_ & new_n3119_;
  assign new_n2103_ = new_n2292_ & new_n3123_ & new_n3122_;
  assign new_n2104_ = new_n3126_ & new_n3125_ & new_n3124_;
  assign new_n2105_ = new_n3128_ & new_n3127_;
  assign new_n2106_ = new_n3131_ & new_n3130_ & new_n3129_;
  assign new_n2107_ = new_n3133_ & new_n3132_;
  assign new_n2108_ = new_n3136_ & new_n3135_ & new_n3134_;
  assign new_n2109_ = new_n3138_ & new_n3137_;
  assign new_n2110_ = new_n3141_ & new_n3140_ & new_n3139_;
  assign new_n2111_ = new_n3143_ & new_n3142_;
  assign new_n2112_ = new_n3145_ & new_n3144_;
  assign new_n2113_ = new_n3148_ & new_n3147_;
  assign new_n2114_ = new_n3150_ & new_n3149_;
  assign new_n2115_ = new_n3153_ & new_n3152_;
  assign new_n2116_ = new_n3156_ & new_n3155_ & new_n3154_;
  assign new_n2117_ = new_n3158_ & new_n3157_;
  assign new_n2118_ = new_n3161_ & new_n3160_ & new_n3159_;
  assign new_n2119_ = new_n3163_ & new_n3162_;
  assign new_n2120_ = new_n3166_ & new_n3165_ & new_n3164_;
  assign new_n2121_ = new_n3168_ & new_n3167_;
  assign new_n2122_ = new_n3171_ & new_n3170_ & new_n3169_;
  assign new_n2123_ = new_n3173_ & new_n3172_;
  assign new_n2124_ = new_n3175_ & new_n3174_;
  assign new_n2125_ = new_n3178_ & new_n3177_;
  assign new_n2126_ = new_n3180_ & new_n3179_;
  assign new_n2127_ = new_n3183_ & new_n3182_;
  assign new_n2128_ = new_n3186_ & new_n3185_ & new_n3184_;
  assign new_n2129_ = new_n3188_ & new_n3187_;
  assign new_n2130_ = new_n3191_ & new_n3190_ & new_n3189_;
  assign new_n2131_ = new_n3193_ & new_n3192_;
  assign new_n2132_ = new_n3195_ & new_n3194_;
  assign new_n2133_ = new_n3198_ & new_n3197_;
  assign new_n2134_ = new_n3200_ & new_n3199_;
  assign new_n2135_ = new_n3203_ & new_n3202_;
  assign new_n2136_ = new_n3205_ & new_n3204_;
  assign new_n2137_ = new_n3208_ & new_n3207_;
  assign new_n2138_ = new_n3210_ & new_n3209_;
  assign new_n2139_ = new_n3213_ & new_n3212_;
  assign new_n2140_ = new_n3215_ & new_n3214_;
  assign new_n2141_ = new_n3218_ & new_n3217_;
  assign new_n2142_ = new_n3220_ & new_n3219_;
  assign new_n2143_ = new_n3223_ & new_n3222_;
  assign new_n2144_ = new_n3225_ & new_n3224_;
  assign new_n2145_ = new_n3228_ & new_n3227_;
  assign new_n2146_ = new_n3230_ & new_n3229_;
  assign new_n2147_ = new_n3233_ & new_n3232_;
  assign new_n2148_ = new_n3235_ & new_n3234_;
  assign new_n2149_ = new_n3238_ & new_n3237_;
  assign new_n2150_ = new_n3240_ & new_n3239_;
  assign new_n2151_ = new_n3243_ & new_n3242_;
  assign new_n2152_ = new_n1704_ & new_n1758_ & new_n1708_;
  assign new_n2153_ = new_n1699_ & new_n1706_ & new_n1703_;
  assign new_n2154_ = new_n1700_ & new_n1702_;
  assign new_n2155_ = new_n2154_ & new_n1759_;
  assign new_n2156_ = new_n1778_ & pi275;
  assign new_n2157_ = new_n3263_ & new_n3264_;
  assign new_n2158_ = new_n3266_ & new_n3267_ & new_n3265_;
  assign new_n2159_ = new_n3273_ & new_n3274_;
  assign new_n2160_ = new_n3276_ & new_n3277_ & new_n3275_;
  assign new_n2161_ = new_n3283_ & new_n3284_;
  assign new_n2162_ = new_n3286_ & new_n3287_ & new_n3285_;
  assign new_n2163_ = new_n3293_ & new_n3294_;
  assign new_n2164_ = new_n3296_ & new_n3297_ & new_n3295_;
  assign new_n2165_ = new_n3303_ & new_n3304_;
  assign new_n2166_ = new_n3306_ & new_n3307_ & new_n3305_;
  assign new_n2167_ = new_n3313_ & new_n3314_;
  assign new_n2168_ = new_n3316_ & new_n3317_ & new_n3315_;
  assign new_n2169_ = new_n3323_ & new_n3324_;
  assign new_n2170_ = new_n3326_ & new_n3327_ & new_n3325_;
  assign new_n2171_ = new_n3333_ & new_n3334_;
  assign new_n2172_ = new_n3336_ & new_n3337_ & new_n3335_;
  assign new_n2173_ = new_n3343_ & new_n3344_;
  assign new_n2174_ = new_n3346_ & new_n3347_ & new_n3345_;
  assign new_n2175_ = new_n3353_ & new_n3354_;
  assign new_n2176_ = new_n3356_ & new_n3357_ & new_n3355_;
  assign new_n2177_ = new_n3363_ & new_n3364_;
  assign new_n2178_ = new_n3366_ & new_n3367_ & new_n3365_;
  assign new_n2179_ = new_n3373_ & new_n3374_;
  assign new_n2180_ = new_n3376_ & new_n3377_ & new_n3375_;
  assign new_n2181_ = new_n3383_ & new_n3384_;
  assign new_n2182_ = new_n3387_ & new_n3386_ & new_n3385_;
  assign new_n2183_ = new_n3392_ & new_n3393_ & new_n3394_;
  assign new_n2184_ = new_n3397_ & new_n3396_ & new_n3395_;
  assign new_n2185_ = new_n3402_ & new_n3403_ & new_n3404_;
  assign new_n2186_ = new_n3407_ & new_n3406_ & new_n3405_;
  assign new_n2187_ = new_n3412_ & new_n2370_;
  assign new_n2188_ = new_n2187_ & new_n3414_ & new_n3413_;
  assign new_n2189_ = new_n3417_ & new_n3416_ & new_n3415_;
  assign new_n2190_ = new_n3422_ & new_n3423_ & new_n3424_;
  assign new_n2191_ = new_n3427_ & new_n3426_ & new_n3425_;
  assign new_n2192_ = new_n3432_ & new_n2370_;
  assign new_n2193_ = new_n2192_ & new_n3434_ & new_n3433_;
  assign new_n2194_ = new_n3437_ & new_n3436_ & new_n3435_;
  assign new_n2195_ = new_n3442_ & new_n3443_ & new_n3444_;
  assign new_n2196_ = new_n3447_ & new_n3446_ & new_n3445_;
  assign new_n2197_ = new_n3452_ & new_n3453_ & new_n3454_;
  assign new_n2198_ = new_n3457_ & new_n3456_ & new_n3455_;
  assign new_n2199_ = pi275 & new_n1765_;
  assign new_n2200_ = new_n2199_ & new_n1763_;
  assign new_n2201_ = new_n4469_ & new_n4466_ & new_n4463_;
  assign new_n2202_ = new_n4481_ & new_n2203_ & new_n2201_;
  assign new_n2203_ = new_n4472_ & new_n4478_ & new_n4475_;
  assign new_n2204_ = new_n4493_ & new_n4490_ & new_n4487_;
  assign new_n2205_ = new_n4502_ & new_n4499_ & new_n4496_;
  assign new_n2206_ = new_n4484_ & new_n2205_ & new_n2204_;
  assign new_n2207_ = new_n4505_ & new_n4460_ & new_n2206_ & new_n2202_;
  assign new_n2208_ = new_n4529_ & new_n4526_;
  assign new_n2209_ = new_n4523_ & new_n4511_ & new_n4514_ & new_n4520_ & new_n4517_;
  assign new_n2210_ = new_n2209_ & new_n4508_;
  assign new_n2211_ = new_n4442_ & new_n4445_ & new_n4451_ & new_n4448_;
  assign new_n2212_ = new_n4457_ & new_n4454_;
  assign new_n2213_ = new_n4436_ & new_n4439_ & new_n2212_ & new_n2211_;
  assign new_n2214_ = new_n4026_ & new_n2323_ & new_n4028_ & new_n3462_;
  assign new_n2215_ = new_n1791_ & new_n1792_;
  assign new_n2216_ = new_n1759_ & new_n1709_ & new_n1707_;
  assign new_n2217_ = new_n4042_ & new_n2341_;
  assign new_n2218_ = new_n1763_ & new_n2217_;
  assign new_n2219_ = new_n1361_ & new_n3471_;
  assign new_n2220_ = new_n2221_ & new_n3514_;
  assign new_n2221_ = new_n3518_ & new_n3517_;
  assign new_n2222_ = new_n2366_ & new_n1415_;
  assign new_n2223_ = new_n3559_ & new_n3558_;
  assign new_n2224_ = new_n3562_ & new_n3561_;
  assign new_n2225_ = new_n2226_ & new_n3576_;
  assign new_n2226_ = new_n3580_ & new_n3579_;
  assign new_n2227_ = new_n3607_ & new_n3606_;
  assign new_n2228_ = new_n2229_ & new_n3648_;
  assign new_n2229_ = new_n3652_ & new_n3651_;
  assign new_n2230_ = new_n2231_ & new_n3684_;
  assign new_n2231_ = new_n3688_ & new_n3687_;
  assign new_n2232_ = new_n1773_ & new_n3737_;
  assign new_n2233_ = new_n3802_ & new_n3803_;
  assign new_n2234_ = new_n3862_ & new_n3860_;
  assign new_n2235_ = new_n1778_ & new_n3874_;
  assign new_n2236_ = new_n1778_ & new_n3880_;
  assign new_n2237_ = new_n3883_ & new_n1778_;
  assign new_n2238_ = new_n3885_ & new_n1778_;
  assign new_n2239_ = new_n3887_ & new_n1778_;
  assign new_n2240_ = new_n3889_ & new_n1778_;
  assign new_n2241_ = new_n3891_ & new_n1778_;
  assign new_n2242_ = new_n3893_ & new_n1778_;
  assign new_n2243_ = new_n3895_ & new_n1778_;
  assign new_n2244_ = new_n3897_ & new_n1778_;
  assign new_n2245_ = new_n3899_ & new_n1778_;
  assign new_n2246_ = new_n3901_ & new_n1778_;
  assign new_n2247_ = new_n1778_ & new_n3902_;
  assign new_n2248_ = new_n1778_ & new_n3904_;
  assign new_n2249_ = new_n1778_ & new_n3906_;
  assign new_n2250_ = new_n1778_ & new_n3908_;
  assign new_n2251_ = new_n1778_ & new_n3910_;
  assign new_n2252_ = new_n1778_ & new_n3912_;
  assign new_n2253_ = new_n1778_ & new_n3914_;
  assign new_n2254_ = new_n1778_ & new_n3916_;
  assign new_n2255_ = new_n1778_ & new_n3918_;
  assign new_n2256_ = new_n1778_ & new_n3920_;
  assign new_n2257_ = new_n1778_ & new_n3922_;
  assign new_n2258_ = new_n1778_ & new_n3924_;
  assign new_n2259_ = new_n1778_ & new_n3926_;
  assign new_n2260_ = new_n3945_ & new_n3943_;
  assign new_n2261_ = new_n3952_ & new_n3950_;
  assign new_n2262_ = new_n3958_ & new_n3956_;
  assign new_n2263_ = new_n3961_ & new_n3959_;
  assign new_n2264_ = new_n3964_ & new_n3962_;
  assign new_n2265_ = new_n3967_ & new_n3965_;
  assign new_n2266_ = new_n3970_ & new_n3968_;
  assign new_n2267_ = new_n3973_ & new_n3971_;
  assign new_n2268_ = new_n3976_ & new_n3974_;
  assign new_n2269_ = new_n3979_ & new_n3977_;
  assign new_n2270_ = new_n3982_ & new_n3980_;
  assign new_n2271_ = new_n3985_ & new_n3983_;
  assign new_n2272_ = new_n3988_ & new_n3986_;
  assign new_n2273_ = new_n3991_ & new_n3989_;
  assign new_n2274_ = new_n3994_ & new_n3992_;
  assign new_n2275_ = new_n3997_ & new_n3995_;
  assign new_n2276_ = new_n4000_ & new_n3998_;
  assign new_n2277_ = new_n4003_ & new_n4001_;
  assign new_n2278_ = new_n4006_ & new_n4004_;
  assign new_n2279_ = new_n4009_ & new_n4007_;
  assign new_n2280_ = new_n4012_ & new_n4010_;
  assign new_n2281_ = new_n4015_ & new_n4013_;
  assign new_n2282_ = new_n4018_ & new_n4016_;
  assign new_n2283_ = ~pi064;
  assign new_n2284_ = ~new_n1361_ | ~new_n1698_;
  assign new_n2285_ = ~new_n4073_ | ~new_n4067_;
  assign new_n2286_ = ~new_n1973_ | ~new_n1386_;
  assign new_n2287_ = ~new_n2092_ | ~new_n1386_;
  assign new_n2288_ = new_n4307_ & new_n4306_;
  assign new_n2289_ = new_n4309_ & new_n4308_;
  assign new_n2290_ = new_n4311_ & new_n4310_;
  assign new_n2291_ = new_n4313_ & new_n4312_;
  assign new_n2292_ = new_n4315_ & new_n4314_;
  assign new_n2293_ = new_n4317_ & new_n4316_;
  assign new_n2294_ = new_n4319_ & new_n4318_;
  assign new_n2295_ = new_n4321_ & new_n4320_;
  assign new_n2296_ = new_n4323_ & new_n4322_;
  assign new_n2297_ = new_n4325_ & new_n4324_;
  assign new_n2298_ = new_n4327_ & new_n4326_;
  assign new_n2299_ = new_n4329_ & new_n4328_;
  assign new_n2300_ = new_n4331_ & new_n4330_;
  assign new_n2301_ = new_n4333_ & new_n4332_;
  assign new_n2302_ = new_n4335_ & new_n4334_;
  assign new_n2303_ = new_n4337_ & new_n4336_;
  assign new_n2304_ = new_n4339_ & new_n4338_;
  assign new_n2305_ = new_n4341_ & new_n4340_;
  assign new_n2306_ = new_n4343_ & new_n4342_;
  assign new_n2307_ = new_n4345_ & new_n4344_;
  assign new_n2308_ = new_n4347_ & new_n4346_;
  assign new_n2309_ = new_n4349_ & new_n4348_;
  assign new_n2310_ = new_n4351_ & new_n4350_;
  assign new_n2311_ = new_n4353_ & new_n4352_;
  assign new_n2312_ = new_n4355_ & new_n4354_;
  assign new_n2313_ = new_n4357_ & new_n4356_;
  assign new_n2314_ = new_n4359_ & new_n4358_;
  assign new_n2315_ = new_n4361_ & new_n4360_;
  assign new_n2316_ = new_n4363_ & new_n4362_;
  assign new_n2317_ = new_n4365_ & new_n4364_;
  assign new_n2318_ = ~new_n2091_ | ~new_n1393_;
  assign new_n2319_ = new_n4367_ & new_n4366_;
  assign new_n2320_ = new_n4369_ & new_n4368_;
  assign new_n2321_ = ~new_n2213_ | ~new_n2208_ | ~new_n2210_ | ~new_n2207_;
  assign new_n2322_ = ~new_n13286_;
  assign new_n2323_ = new_n4539_ & new_n4538_;
  assign new_n2324_ = ~new_n11071_;
  assign new_n2325_ = ~new_n1710_;
  assign new_n2326_ = ~new_n1767_;
  assign new_n2327_ = ~new_n1765_;
  assign new_n2328_ = ~new_n1708_;
  assign new_n2329_ = ~new_n1758_;
  assign new_n2330_ = ~new_n1704_;
  assign new_n2331_ = ~new_n1703_;
  assign new_n2332_ = ~new_n1706_;
  assign new_n2333_ = ~new_n1699_;
  assign new_n2334_ = ~new_n1702_;
  assign new_n2335_ = ~new_n1700_;
  assign new_n2336_ = ~new_n1759_;
  assign new_n2337_ = ~new_n1757_;
  assign new_n2338_ = ~new_n1388_ | ~new_n2373_;
  assign new_n2339_ = ~new_n1709_;
  assign new_n2340_ = ~new_n1707_;
  assign new_n2341_ = ~new_n2359_ | ~new_n1705_;
  assign new_n2342_ = ~new_n1388_ | ~new_n1760_;
  assign new_n2343_ = ~new_n2285_;
  assign new_n2344_ = ~new_n1770_;
  assign po266 = ~new_n1764_;
  assign new_n2346_ = ~new_n1749_;
  assign new_n2347_ = ~new_n1747_;
  assign new_n2348_ = ~new_n1745_;
  assign new_n2349_ = ~new_n1743_;
  assign new_n2350_ = ~new_n1741_;
  assign new_n2351_ = ~new_n1739_;
  assign new_n2352_ = ~new_n1737_;
  assign new_n2353_ = ~new_n1735_;
  assign new_n2354_ = ~new_n1733_;
  assign new_n2355_ = ~new_n1754_;
  assign new_n2356_ = ~new_n1753_;
  assign new_n2357_ = ~new_n1751_;
  assign new_n2358_ = ~new_n1766_;
  assign new_n2359_ = ~new_n1711_;
  assign new_n2360_ = ~new_n1755_;
  assign new_n2361_ = ~new_n1756_;
  assign new_n2362_ = ~new_n2287_;
  assign new_n2363_ = ~new_n2286_;
  assign new_n2364_ = ~new_n2284_;
  assign new_n2365_ = ~new_n2318_;
  assign new_n2366_ = ~new_n1771_;
  assign new_n2367_ = ~new_n1772_ | ~pi275;
  assign new_n2368_ = ~new_n2337_ | ~new_n1361_;
  assign new_n2369_ = ~new_n1769_;
  assign new_n2370_ = ~po266 | ~new_n1549_;
  assign new_n2371_ = ~new_n1763_;
  assign new_n2372_ = ~new_n1773_;
  assign new_n2373_ = ~new_n1701_;
  assign new_n2374_ = ~new_n1705_;
  assign new_n2375_ = ~new_n1696_;
  assign new_n2376_ = ~new_n1695_;
  assign new_n2377_ = ~new_n1102_ | ~po264;
  assign new_n2378_ = ~pi033 | ~new_n1367_;
  assign new_n2379_ = ~pi033 | ~new_n2376_;
  assign new_n2380_ = ~new_n1091_ | ~po264;
  assign new_n2381_ = ~new_n9224_ | ~new_n1367_;
  assign new_n2382_ = ~pi034 | ~new_n2376_;
  assign new_n2383_ = ~new_n1080_ | ~po264;
  assign new_n2384_ = ~new_n9205_ | ~new_n1367_;
  assign new_n2385_ = ~pi035 | ~new_n2376_;
  assign new_n2386_ = ~new_n1077_ | ~po264;
  assign new_n2387_ = ~new_n9206_ | ~new_n1367_;
  assign new_n2388_ = ~pi036 | ~new_n2376_;
  assign new_n2389_ = ~new_n1076_ | ~po264;
  assign new_n2390_ = ~new_n9207_ | ~new_n1367_;
  assign new_n2391_ = ~pi037 | ~new_n2376_;
  assign new_n2392_ = ~new_n1075_ | ~po264;
  assign new_n2393_ = ~new_n9346_ | ~new_n1367_;
  assign new_n2394_ = ~pi038 | ~new_n2376_;
  assign new_n2395_ = ~new_n1074_ | ~po264;
  assign new_n2396_ = ~new_n9208_ | ~new_n1367_;
  assign new_n2397_ = ~pi039 | ~new_n2376_;
  assign new_n2398_ = ~new_n1073_ | ~po264;
  assign new_n2399_ = ~new_n9209_ | ~new_n1367_;
  assign new_n2400_ = ~pi040 | ~new_n2376_;
  assign new_n2401_ = ~new_n1072_ | ~po264;
  assign new_n2402_ = ~new_n9210_ | ~new_n1367_;
  assign new_n2403_ = ~pi041 | ~new_n2376_;
  assign new_n2404_ = ~new_n1071_ | ~po264;
  assign new_n2405_ = ~new_n9344_ | ~new_n1367_;
  assign new_n2406_ = ~pi042 | ~new_n2376_;
  assign new_n2407_ = ~new_n1101_ | ~po264;
  assign new_n2408_ = ~new_n9190_ | ~new_n1367_;
  assign new_n2409_ = ~pi043 | ~new_n2376_;
  assign new_n2410_ = ~new_n1100_ | ~po264;
  assign new_n2411_ = ~new_n9191_ | ~new_n1367_;
  assign new_n2412_ = ~pi044 | ~new_n2376_;
  assign new_n2413_ = ~new_n1099_ | ~po264;
  assign new_n2414_ = ~new_n9192_ | ~new_n1367_;
  assign new_n2415_ = ~pi045 | ~new_n2376_;
  assign new_n2416_ = ~new_n1098_ | ~po264;
  assign new_n2417_ = ~new_n9363_ | ~new_n1367_;
  assign new_n2418_ = ~pi046 | ~new_n2376_;
  assign new_n2419_ = ~new_n1097_ | ~po264;
  assign new_n2420_ = ~new_n9193_ | ~new_n1367_;
  assign new_n2421_ = ~pi047 | ~new_n2376_;
  assign new_n2422_ = ~new_n1096_ | ~po264;
  assign new_n2423_ = ~new_n9194_ | ~new_n1367_;
  assign new_n2424_ = ~pi048 | ~new_n2376_;
  assign new_n2425_ = ~new_n1095_ | ~po264;
  assign new_n2426_ = ~new_n9195_ | ~new_n1367_;
  assign new_n2427_ = ~pi049 | ~new_n2376_;
  assign new_n2428_ = ~new_n1094_ | ~po264;
  assign new_n2429_ = ~new_n9361_ | ~new_n1367_;
  assign new_n2430_ = ~pi050 | ~new_n2376_;
  assign new_n2431_ = ~new_n1093_ | ~po264;
  assign new_n2432_ = ~new_n9196_ | ~new_n1367_;
  assign new_n2433_ = ~pi051 | ~new_n2376_;
  assign new_n2434_ = ~new_n1092_ | ~po264;
  assign new_n2435_ = ~new_n9197_ | ~new_n1367_;
  assign new_n2436_ = ~pi052 | ~new_n2376_;
  assign new_n2437_ = ~new_n1090_ | ~po264;
  assign new_n2438_ = ~new_n9198_ | ~new_n1367_;
  assign new_n2439_ = ~pi053 | ~new_n2376_;
  assign new_n2440_ = ~new_n1089_ | ~po264;
  assign new_n2441_ = ~new_n9357_ | ~new_n1367_;
  assign new_n2442_ = ~pi054 | ~new_n2376_;
  assign new_n2443_ = ~new_n1088_ | ~po264;
  assign new_n2444_ = ~new_n9199_ | ~new_n1367_;
  assign new_n2445_ = ~pi055 | ~new_n2376_;
  assign new_n2446_ = ~new_n1087_ | ~po264;
  assign new_n2447_ = ~new_n9200_ | ~new_n1367_;
  assign new_n2448_ = ~pi056 | ~new_n2376_;
  assign new_n2449_ = ~new_n1086_ | ~po264;
  assign new_n2450_ = ~new_n9201_ | ~new_n1367_;
  assign new_n2451_ = ~pi057 | ~new_n2376_;
  assign new_n2452_ = ~new_n1085_ | ~po264;
  assign new_n2453_ = ~new_n9354_ | ~new_n1367_;
  assign new_n2454_ = ~pi058 | ~new_n2376_;
  assign new_n2455_ = ~new_n1084_ | ~po264;
  assign new_n2456_ = ~new_n9202_ | ~new_n1367_;
  assign new_n2457_ = ~pi059 | ~new_n2376_;
  assign new_n2458_ = ~new_n1083_ | ~po264;
  assign new_n2459_ = ~new_n9226_ | ~new_n1367_;
  assign new_n2460_ = ~pi060 | ~new_n2376_;
  assign new_n2461_ = ~new_n1082_ | ~po264;
  assign new_n2462_ = ~new_n9203_ | ~new_n1367_;
  assign new_n2463_ = ~pi061 | ~new_n2376_;
  assign new_n2464_ = ~new_n1081_ | ~po264;
  assign new_n2465_ = ~new_n9204_ | ~new_n1367_;
  assign new_n2466_ = ~pi062 | ~new_n2376_;
  assign new_n2467_ = ~new_n1079_ | ~po264;
  assign new_n2468_ = ~new_n9349_ | ~new_n1367_;
  assign new_n2469_ = ~pi063 | ~new_n2376_;
  assign new_n2470_ = ~new_n1078_ | ~po264;
  assign new_n2471_ = ~new_n9225_ | ~new_n1367_;
  assign new_n2472_ = ~pi064 | ~new_n2376_;
  assign new_n2473_ = ~new_n1698_;
  assign new_n2474_ = ~new_n1760_;
  assign new_n2475_ = ~new_n1696_ | ~new_n4031_;
  assign new_n2476_ = ~new_n1696_ | ~new_n4034_;
  assign new_n2477_ = ~new_n2473_ | ~pi075;
  assign new_n2478_ = ~new_n2473_ | ~pi076;
  assign new_n2479_ = ~new_n2473_ | ~pi077;
  assign new_n2480_ = ~new_n2473_ | ~pi078;
  assign new_n2481_ = ~new_n2473_ | ~pi079;
  assign new_n2482_ = ~new_n2473_ | ~pi080;
  assign new_n2483_ = ~new_n2473_ | ~pi081;
  assign new_n2484_ = ~new_n2473_ | ~pi082;
  assign new_n2485_ = ~new_n2473_ | ~pi083;
  assign new_n2486_ = ~new_n2473_ | ~pi084;
  assign new_n2487_ = ~new_n2473_ | ~pi085;
  assign new_n2488_ = ~new_n2473_ | ~pi086;
  assign new_n2489_ = ~new_n2473_ | ~pi087;
  assign new_n2490_ = ~new_n2473_ | ~pi088;
  assign new_n2491_ = ~new_n2473_ | ~pi089;
  assign new_n2492_ = ~new_n2473_ | ~pi090;
  assign new_n2493_ = ~new_n2473_ | ~pi091;
  assign new_n2494_ = ~new_n2473_ | ~pi092;
  assign new_n2495_ = ~new_n2473_ | ~pi093;
  assign new_n2496_ = ~new_n2473_ | ~pi094;
  assign new_n2497_ = ~new_n2473_ | ~pi067;
  assign new_n2498_ = ~new_n2473_ | ~pi095;
  assign new_n2499_ = ~new_n2473_ | ~pi096;
  assign new_n2500_ = ~new_n2473_ | ~pi068;
  assign new_n2501_ = ~new_n2473_ | ~pi069;
  assign new_n2502_ = ~new_n2473_ | ~pi070;
  assign new_n2503_ = ~new_n2473_ | ~pi071;
  assign new_n2504_ = ~new_n2473_ | ~pi072;
  assign new_n2505_ = ~new_n2473_ | ~pi073;
  assign new_n2506_ = ~new_n2473_ | ~pi074;
  assign new_n2507_ = ~new_n4055_ | ~new_n4058_;
  assign new_n2508_ = ~new_n1705_ | ~new_n4078_ | ~new_n4077_;
  assign new_n2509_ = ~new_n1357_ | ~pi162;
  assign new_n2510_ = ~new_n1358_ | ~pi130;
  assign new_n2511_ = ~new_n1359_ | ~pi098;
  assign new_n2512_ = ~pi265 | ~new_n1356_;
  assign new_n2513_ = ~new_n1415_;
  assign new_n2514_ = ~new_n2338_ | ~new_n1755_;
  assign new_n2515_ = ~new_n2333_ | ~new_n12158_;
  assign new_n2516_ = ~new_n2335_ | ~new_n10413_;
  assign new_n2517_ = ~new_n2334_ | ~new_n14068_;
  assign new_n2518_ = ~new_n2331_ | ~new_n12629_;
  assign new_n2519_ = ~new_n2330_ | ~new_n11088_;
  assign new_n2520_ = ~new_n2340_ | ~new_n13570_;
  assign new_n2521_ = ~new_n2339_ | ~new_n9687_;
  assign new_n2522_ = ~new_n1712_;
  assign new_n2523_ = ~new_n14566_ | ~new_n1365_;
  assign new_n2524_ = ~new_n1364_ | ~new_n1415_;
  assign new_n2525_ = ~new_n1790_ | ~new_n1362_;
  assign new_n2526_ = ~new_n1790_ | ~new_n2514_;
  assign new_n2527_ = ~new_n1961_ | ~new_n2522_;
  assign new_n2528_ = ~pi163 | ~new_n1357_;
  assign new_n2529_ = ~pi131 | ~new_n1358_;
  assign new_n2530_ = ~pi099 | ~new_n1359_;
  assign new_n2531_ = ~pi250 | ~new_n1356_;
  assign new_n2532_ = ~new_n1405_;
  assign new_n2533_ = ~pi097 | ~new_n1359_;
  assign new_n2534_ = ~pi129 | ~new_n1358_;
  assign new_n2535_ = ~pi161 | ~new_n1357_;
  assign new_n2536_ = ~pi255 | ~new_n1356_;
  assign new_n2537_ = ~new_n1414_;
  assign new_n2538_ = ~new_n1372_ | ~new_n1414_;
  assign new_n2539_ = ~new_n12235_ | ~new_n2333_;
  assign new_n2540_ = ~new_n10490_ | ~new_n2335_;
  assign new_n2541_ = ~new_n14067_ | ~new_n2334_;
  assign new_n2542_ = ~new_n12706_ | ~new_n2331_;
  assign new_n2543_ = ~new_n11165_ | ~new_n2330_;
  assign new_n2544_ = ~new_n13569_ | ~new_n2340_;
  assign new_n2545_ = ~new_n9686_ | ~new_n2339_;
  assign new_n2546_ = ~new_n1714_;
  assign new_n2547_ = ~new_n14565_ | ~new_n1365_;
  assign new_n2548_ = ~new_n1364_ | ~new_n1405_;
  assign new_n2549_ = ~new_n9492_ | ~new_n1362_;
  assign new_n2550_ = ~new_n1795_ | ~new_n2514_;
  assign new_n2551_ = ~new_n1977_ | ~new_n2546_;
  assign new_n2552_ = ~pi164 | ~new_n1357_;
  assign new_n2553_ = ~pi132 | ~new_n1358_;
  assign new_n2554_ = ~pi100 | ~new_n1359_;
  assign new_n2555_ = ~new_n8735_ | ~new_n1356_;
  assign new_n2556_ = ~new_n1401_;
  assign new_n2557_ = ~new_n1372_ | ~new_n1415_;
  assign new_n2558_ = ~new_n12245_ | ~new_n2333_;
  assign new_n2559_ = ~new_n10500_ | ~new_n2335_;
  assign new_n2560_ = ~new_n13989_ | ~new_n2334_;
  assign new_n2561_ = ~new_n12716_ | ~new_n2331_;
  assign new_n2562_ = ~new_n11175_ | ~new_n2330_;
  assign new_n2563_ = ~new_n13491_ | ~new_n2340_;
  assign new_n2564_ = ~new_n9608_ | ~new_n2339_;
  assign new_n2565_ = ~new_n1715_;
  assign new_n2566_ = ~new_n14487_ | ~new_n1365_;
  assign new_n2567_ = ~new_n1364_ | ~new_n1401_;
  assign new_n2568_ = ~new_n9453_ | ~new_n1362_;
  assign new_n2569_ = ~new_n1798_ | ~new_n2514_;
  assign new_n2570_ = ~new_n1981_ | ~new_n2565_;
  assign new_n2571_ = ~pi165 | ~new_n1357_;
  assign new_n2572_ = ~pi133 | ~new_n1358_;
  assign new_n2573_ = ~pi101 | ~new_n1359_;
  assign new_n2574_ = ~new_n8790_ | ~new_n1356_;
  assign new_n2575_ = ~new_n1397_;
  assign new_n2576_ = ~new_n1372_ | ~new_n1405_;
  assign new_n2577_ = ~new_n12155_ | ~new_n2333_;
  assign new_n2578_ = ~new_n10410_ | ~new_n2335_;
  assign new_n2579_ = ~new_n14073_ | ~new_n2334_;
  assign new_n2580_ = ~new_n12626_ | ~new_n2331_;
  assign new_n2581_ = ~new_n11085_ | ~new_n2330_;
  assign new_n2582_ = ~new_n13575_ | ~new_n2340_;
  assign new_n2583_ = ~new_n9692_ | ~new_n2339_;
  assign new_n2584_ = ~new_n1716_;
  assign new_n2585_ = ~new_n14571_ | ~new_n1365_;
  assign new_n2586_ = ~new_n1364_ | ~new_n1397_;
  assign new_n2587_ = ~new_n9455_ | ~new_n1362_;
  assign new_n2588_ = ~new_n1801_ | ~new_n2514_;
  assign new_n2589_ = ~new_n1985_ | ~new_n2584_;
  assign new_n2590_ = ~pi166 | ~new_n1357_;
  assign new_n2591_ = ~pi134 | ~new_n1358_;
  assign new_n2592_ = ~pi102 | ~new_n1359_;
  assign new_n2593_ = ~new_n8789_ | ~new_n1356_;
  assign new_n2594_ = ~new_n1404_;
  assign new_n2595_ = ~new_n1372_ | ~new_n1401_;
  assign new_n2596_ = ~new_n12244_ | ~new_n2333_;
  assign new_n2597_ = ~new_n10499_ | ~new_n2335_;
  assign new_n2598_ = ~new_n14072_ | ~new_n2334_;
  assign new_n2599_ = ~new_n12715_ | ~new_n2331_;
  assign new_n2600_ = ~new_n11174_ | ~new_n2330_;
  assign new_n2601_ = ~new_n13574_ | ~new_n2340_;
  assign new_n2602_ = ~new_n9691_ | ~new_n2339_;
  assign new_n2603_ = ~new_n1717_;
  assign new_n2604_ = ~new_n14570_ | ~new_n1365_;
  assign new_n2605_ = ~new_n1364_ | ~new_n1404_;
  assign new_n2606_ = ~new_n9456_ | ~new_n1362_;
  assign new_n2607_ = ~new_n1804_ | ~new_n2514_;
  assign new_n2608_ = ~new_n1989_ | ~new_n2603_;
  assign new_n2609_ = ~pi167 | ~new_n1357_;
  assign new_n2610_ = ~pi135 | ~new_n1358_;
  assign new_n2611_ = ~pi103 | ~new_n1359_;
  assign new_n2612_ = ~new_n8788_ | ~new_n1356_;
  assign new_n2613_ = ~new_n1408_;
  assign new_n2614_ = ~new_n1372_ | ~new_n1397_;
  assign new_n2615_ = ~new_n12243_ | ~new_n2333_;
  assign new_n2616_ = ~new_n10498_ | ~new_n2335_;
  assign new_n2617_ = ~new_n13990_ | ~new_n2334_;
  assign new_n2618_ = ~new_n12714_ | ~new_n2331_;
  assign new_n2619_ = ~new_n11173_ | ~new_n2330_;
  assign new_n2620_ = ~new_n13492_ | ~new_n2340_;
  assign new_n2621_ = ~new_n9609_ | ~new_n2339_;
  assign new_n2622_ = ~new_n1718_;
  assign new_n2623_ = ~new_n14488_ | ~new_n1365_;
  assign new_n2624_ = ~new_n1364_ | ~new_n1408_;
  assign new_n2625_ = ~new_n9500_ | ~new_n1362_;
  assign new_n2626_ = ~new_n1807_ | ~new_n2514_;
  assign new_n2627_ = ~new_n1993_ | ~new_n2622_;
  assign new_n2628_ = ~pi168 | ~new_n1357_;
  assign new_n2629_ = ~pi136 | ~new_n1358_;
  assign new_n2630_ = ~pi104 | ~new_n1359_;
  assign new_n2631_ = ~new_n8787_ | ~new_n1356_;
  assign new_n2632_ = ~new_n1407_;
  assign new_n2633_ = ~new_n1372_ | ~new_n1404_;
  assign new_n2634_ = ~new_n12156_ | ~new_n2333_;
  assign new_n2635_ = ~new_n10411_ | ~new_n2335_;
  assign new_n2636_ = ~new_n14071_ | ~new_n2334_;
  assign new_n2637_ = ~new_n12627_ | ~new_n2331_;
  assign new_n2638_ = ~new_n11086_ | ~new_n2330_;
  assign new_n2639_ = ~new_n13573_ | ~new_n2340_;
  assign new_n2640_ = ~new_n9690_ | ~new_n2339_;
  assign new_n2641_ = ~new_n1719_;
  assign new_n2642_ = ~new_n14569_ | ~new_n1365_;
  assign new_n2643_ = ~new_n1364_ | ~new_n1407_;
  assign new_n2644_ = ~new_n9457_ | ~new_n1362_;
  assign new_n2645_ = ~new_n1810_ | ~new_n2514_;
  assign new_n2646_ = ~new_n1997_ | ~new_n2641_;
  assign new_n2647_ = ~pi169 | ~new_n1357_;
  assign new_n2648_ = ~pi137 | ~new_n1358_;
  assign new_n2649_ = ~pi105 | ~new_n1359_;
  assign new_n2650_ = ~new_n8786_ | ~new_n1356_;
  assign new_n2651_ = ~new_n1421_;
  assign new_n2652_ = ~new_n1372_ | ~new_n1408_;
  assign new_n2653_ = ~new_n12242_ | ~new_n2333_;
  assign new_n2654_ = ~new_n10497_ | ~new_n2335_;
  assign new_n2655_ = ~new_n13991_ | ~new_n2334_;
  assign new_n2656_ = ~new_n12713_ | ~new_n2331_;
  assign new_n2657_ = ~new_n11172_ | ~new_n2330_;
  assign new_n2658_ = ~new_n13493_ | ~new_n2340_;
  assign new_n2659_ = ~new_n9610_ | ~new_n2339_;
  assign new_n2660_ = ~new_n1720_;
  assign new_n2661_ = ~new_n14489_ | ~new_n1365_;
  assign new_n2662_ = ~new_n1364_ | ~new_n1421_;
  assign new_n2663_ = ~new_n9458_ | ~new_n1362_;
  assign new_n2664_ = ~new_n1813_ | ~new_n2514_;
  assign new_n2665_ = ~new_n2001_ | ~new_n2660_;
  assign new_n2666_ = ~pi170 | ~new_n1357_;
  assign new_n2667_ = ~pi138 | ~new_n1358_;
  assign new_n2668_ = ~pi106 | ~new_n1359_;
  assign new_n2669_ = ~new_n8785_ | ~new_n1356_;
  assign new_n2670_ = ~new_n1420_;
  assign new_n2671_ = ~new_n1372_ | ~new_n1407_;
  assign new_n2672_ = ~new_n12157_ | ~new_n2333_;
  assign new_n2673_ = ~new_n10412_ | ~new_n2335_;
  assign new_n2674_ = ~new_n14070_ | ~new_n2334_;
  assign new_n2675_ = ~new_n12628_ | ~new_n2331_;
  assign new_n2676_ = ~new_n11087_ | ~new_n2330_;
  assign new_n2677_ = ~new_n13572_ | ~new_n2340_;
  assign new_n2678_ = ~new_n9689_ | ~new_n2339_;
  assign new_n2679_ = ~new_n1721_;
  assign new_n2680_ = ~new_n14568_ | ~new_n1365_;
  assign new_n2681_ = ~new_n1364_ | ~new_n1420_;
  assign new_n2682_ = ~new_n9459_ | ~new_n1362_;
  assign new_n2683_ = ~new_n1816_ | ~new_n2514_;
  assign new_n2684_ = ~new_n2005_ | ~new_n2679_;
  assign new_n2685_ = ~pi171 | ~new_n1357_;
  assign new_n2686_ = ~pi139 | ~new_n1358_;
  assign new_n2687_ = ~pi107 | ~new_n1359_;
  assign new_n2688_ = ~new_n8809_ | ~new_n1356_;
  assign new_n2689_ = ~new_n1399_;
  assign new_n2690_ = ~new_n1372_ | ~new_n1421_;
  assign new_n2691_ = ~new_n12241_ | ~new_n2333_;
  assign new_n2692_ = ~new_n10496_ | ~new_n2335_;
  assign new_n2693_ = ~new_n14069_ | ~new_n2334_;
  assign new_n2694_ = ~new_n12712_ | ~new_n2331_;
  assign new_n2695_ = ~new_n11171_ | ~new_n2330_;
  assign new_n2696_ = ~new_n13571_ | ~new_n2340_;
  assign new_n2697_ = ~new_n9688_ | ~new_n2339_;
  assign new_n2698_ = ~new_n1722_;
  assign new_n2699_ = ~new_n14567_ | ~new_n1365_;
  assign new_n2700_ = ~new_n1364_ | ~new_n1399_;
  assign new_n2701_ = ~new_n9498_ | ~new_n1362_;
  assign new_n2702_ = ~new_n1819_ | ~new_n2514_;
  assign new_n2703_ = ~new_n2009_ | ~new_n2698_;
  assign new_n2704_ = ~pi172 | ~new_n1357_;
  assign new_n2705_ = ~pi140 | ~new_n1358_;
  assign new_n2706_ = ~pi108 | ~new_n1359_;
  assign new_n2707_ = ~new_n8808_ | ~new_n1356_;
  assign new_n2708_ = ~new_n1400_;
  assign new_n2709_ = ~new_n1372_ | ~new_n1420_;
  assign new_n2710_ = ~new_n12251_ | ~new_n2333_;
  assign new_n2711_ = ~new_n10506_ | ~new_n2335_;
  assign new_n2712_ = ~new_n13983_ | ~new_n2334_;
  assign new_n2713_ = ~new_n12722_ | ~new_n2331_;
  assign new_n2714_ = ~new_n11181_ | ~new_n2330_;
  assign new_n2715_ = ~new_n13485_ | ~new_n2340_;
  assign new_n2716_ = ~new_n9602_ | ~new_n2339_;
  assign new_n2717_ = ~new_n1723_;
  assign new_n2718_ = ~new_n14481_ | ~new_n1365_;
  assign new_n2719_ = ~new_n1364_ | ~new_n1400_;
  assign new_n2720_ = ~new_n9441_ | ~new_n1362_;
  assign new_n2721_ = ~new_n1822_ | ~new_n2514_;
  assign new_n2722_ = ~new_n2013_ | ~new_n2717_;
  assign new_n2723_ = ~pi173 | ~new_n1357_;
  assign new_n2724_ = ~pi141 | ~new_n1358_;
  assign new_n2725_ = ~pi109 | ~new_n1359_;
  assign new_n2726_ = ~new_n8807_ | ~new_n1356_;
  assign new_n2727_ = ~new_n1409_;
  assign new_n2728_ = ~new_n1372_ | ~new_n1399_;
  assign new_n2729_ = ~new_n12150_ | ~new_n2333_;
  assign new_n2730_ = ~new_n10405_ | ~new_n2335_;
  assign new_n2731_ = ~new_n14087_ | ~new_n2334_;
  assign new_n2732_ = ~new_n12621_ | ~new_n2331_;
  assign new_n2733_ = ~new_n11080_ | ~new_n2330_;
  assign new_n2734_ = ~new_n13589_ | ~new_n2340_;
  assign new_n2735_ = ~new_n9706_ | ~new_n2339_;
  assign new_n2736_ = ~new_n1724_;
  assign new_n2737_ = ~new_n14585_ | ~new_n1365_;
  assign new_n2738_ = ~new_n1364_ | ~new_n1409_;
  assign new_n2739_ = ~new_n9442_ | ~new_n1362_;
  assign new_n2740_ = ~new_n1825_ | ~new_n2514_;
  assign new_n2741_ = ~new_n2017_ | ~new_n2736_;
  assign new_n2742_ = ~pi174 | ~new_n1357_;
  assign new_n2743_ = ~pi142 | ~new_n1358_;
  assign new_n2744_ = ~pi110 | ~new_n1359_;
  assign new_n2745_ = ~new_n8806_ | ~new_n1356_;
  assign new_n2746_ = ~new_n1417_;
  assign new_n2747_ = ~new_n1372_ | ~new_n1400_;
  assign new_n2748_ = ~new_n12240_ | ~new_n2333_;
  assign new_n2749_ = ~new_n10495_ | ~new_n2335_;
  assign new_n2750_ = ~new_n14086_ | ~new_n2334_;
  assign new_n2751_ = ~new_n12711_ | ~new_n2331_;
  assign new_n2752_ = ~new_n11170_ | ~new_n2330_;
  assign new_n2753_ = ~new_n13588_ | ~new_n2340_;
  assign new_n2754_ = ~new_n9705_ | ~new_n2339_;
  assign new_n2755_ = ~new_n1725_;
  assign new_n2756_ = ~new_n14584_ | ~new_n1365_;
  assign new_n2757_ = ~new_n1364_ | ~new_n1417_;
  assign new_n2758_ = ~new_n9443_ | ~new_n1362_;
  assign new_n2759_ = ~new_n1828_ | ~new_n2514_;
  assign new_n2760_ = ~new_n2021_ | ~new_n2755_;
  assign new_n2761_ = ~pi175 | ~new_n1357_;
  assign new_n2762_ = ~pi143 | ~new_n1358_;
  assign new_n2763_ = ~pi111 | ~new_n1359_;
  assign new_n2764_ = ~new_n8805_ | ~new_n1356_;
  assign new_n2765_ = ~new_n1416_;
  assign new_n2766_ = ~new_n1372_ | ~new_n1409_;
  assign new_n2767_ = ~new_n12239_ | ~new_n2333_;
  assign new_n2768_ = ~new_n10494_ | ~new_n2335_;
  assign new_n2769_ = ~new_n13984_ | ~new_n2334_;
  assign new_n2770_ = ~new_n12710_ | ~new_n2331_;
  assign new_n2771_ = ~new_n11169_ | ~new_n2330_;
  assign new_n2772_ = ~new_n13486_ | ~new_n2340_;
  assign new_n2773_ = ~new_n9603_ | ~new_n2339_;
  assign new_n2774_ = ~new_n1726_;
  assign new_n2775_ = ~new_n14482_ | ~new_n1365_;
  assign new_n2776_ = ~new_n1364_ | ~new_n1416_;
  assign new_n2777_ = ~new_n9521_ | ~new_n1362_;
  assign new_n2778_ = ~new_n1831_ | ~new_n2514_;
  assign new_n2779_ = ~new_n2025_ | ~new_n2774_;
  assign new_n2780_ = ~pi176 | ~new_n1357_;
  assign new_n2781_ = ~pi144 | ~new_n1358_;
  assign new_n2782_ = ~pi112 | ~new_n1359_;
  assign new_n2783_ = ~new_n8804_ | ~new_n1356_;
  assign new_n2784_ = ~new_n1411_;
  assign new_n2785_ = ~new_n1372_ | ~new_n1417_;
  assign new_n2786_ = ~new_n12250_ | ~new_n2333_;
  assign new_n2787_ = ~new_n10505_ | ~new_n2335_;
  assign new_n2788_ = ~new_n14085_ | ~new_n2334_;
  assign new_n2789_ = ~new_n12721_ | ~new_n2331_;
  assign new_n2790_ = ~new_n11180_ | ~new_n2330_;
  assign new_n2791_ = ~new_n13587_ | ~new_n2340_;
  assign new_n2792_ = ~new_n9704_ | ~new_n2339_;
  assign new_n2793_ = ~new_n1727_;
  assign new_n2794_ = ~new_n14583_ | ~new_n1365_;
  assign new_n2795_ = ~new_n1364_ | ~new_n1411_;
  assign new_n2796_ = ~new_n9444_ | ~new_n1362_;
  assign new_n2797_ = ~new_n1834_ | ~new_n2514_;
  assign new_n2798_ = ~new_n2029_ | ~new_n2793_;
  assign new_n2799_ = ~pi177 | ~new_n1357_;
  assign new_n2800_ = ~pi145 | ~new_n1358_;
  assign new_n2801_ = ~pi113 | ~new_n1359_;
  assign new_n2802_ = ~new_n8803_ | ~new_n1356_;
  assign new_n2803_ = ~new_n1410_;
  assign new_n2804_ = ~new_n1372_ | ~new_n1416_;
  assign new_n2805_ = ~new_n12249_ | ~new_n2333_;
  assign new_n2806_ = ~new_n10504_ | ~new_n2335_;
  assign new_n2807_ = ~new_n14084_ | ~new_n2334_;
  assign new_n2808_ = ~new_n12720_ | ~new_n2331_;
  assign new_n2809_ = ~new_n11179_ | ~new_n2330_;
  assign new_n2810_ = ~new_n13586_ | ~new_n2340_;
  assign new_n2811_ = ~new_n9703_ | ~new_n2339_;
  assign new_n2812_ = ~new_n1728_;
  assign new_n2813_ = ~new_n14582_ | ~new_n1365_;
  assign new_n2814_ = ~new_n1364_ | ~new_n1410_;
  assign new_n2815_ = ~new_n9445_ | ~new_n1362_;
  assign new_n2816_ = ~new_n1837_ | ~new_n2514_;
  assign new_n2817_ = ~new_n2033_ | ~new_n2812_;
  assign new_n2818_ = ~pi178 | ~new_n1357_;
  assign new_n2819_ = ~pi146 | ~new_n1358_;
  assign new_n2820_ = ~pi114 | ~new_n1359_;
  assign new_n2821_ = ~new_n8802_ | ~new_n1356_;
  assign new_n2822_ = ~new_n1406_;
  assign new_n2823_ = ~new_n1372_ | ~new_n1411_;
  assign new_n2824_ = ~new_n12151_ | ~new_n2333_;
  assign new_n2825_ = ~new_n10406_ | ~new_n2335_;
  assign new_n2826_ = ~new_n14083_ | ~new_n2334_;
  assign new_n2827_ = ~new_n12622_ | ~new_n2331_;
  assign new_n2828_ = ~new_n11081_ | ~new_n2330_;
  assign new_n2829_ = ~new_n13585_ | ~new_n2340_;
  assign new_n2830_ = ~new_n9702_ | ~new_n2339_;
  assign new_n2831_ = ~new_n1729_;
  assign new_n2832_ = ~new_n14581_ | ~new_n1365_;
  assign new_n2833_ = ~new_n1364_ | ~new_n1406_;
  assign new_n2834_ = ~new_n9446_ | ~new_n1362_;
  assign new_n2835_ = ~new_n1840_ | ~new_n2514_;
  assign new_n2836_ = ~new_n2037_ | ~new_n2831_;
  assign new_n2837_ = ~pi179 | ~new_n1357_;
  assign new_n2838_ = ~pi147 | ~new_n1358_;
  assign new_n2839_ = ~pi115 | ~new_n1359_;
  assign new_n2840_ = ~new_n8801_ | ~new_n1356_;
  assign new_n2841_ = ~new_n1419_;
  assign new_n2842_ = ~new_n1372_ | ~new_n1410_;
  assign new_n2843_ = ~new_n12238_ | ~new_n2333_;
  assign new_n2844_ = ~new_n10493_ | ~new_n2335_;
  assign new_n2845_ = ~new_n13985_ | ~new_n2334_;
  assign new_n2846_ = ~new_n12709_ | ~new_n2331_;
  assign new_n2847_ = ~new_n11168_ | ~new_n2330_;
  assign new_n2848_ = ~new_n13487_ | ~new_n2340_;
  assign new_n2849_ = ~new_n9604_ | ~new_n2339_;
  assign new_n2850_ = ~new_n1730_;
  assign new_n2851_ = ~new_n14483_ | ~new_n1365_;
  assign new_n2852_ = ~new_n1364_ | ~new_n1419_;
  assign new_n2853_ = ~new_n9519_ | ~new_n1362_;
  assign new_n2854_ = ~new_n1843_ | ~new_n2514_;
  assign new_n2855_ = ~new_n2041_ | ~new_n2850_;
  assign new_n2856_ = ~pi180 | ~new_n1357_;
  assign new_n2857_ = ~pi148 | ~new_n1358_;
  assign new_n2858_ = ~pi116 | ~new_n1359_;
  assign new_n2859_ = ~new_n8800_ | ~new_n1356_;
  assign new_n2860_ = ~new_n1418_;
  assign new_n2861_ = ~new_n1372_ | ~new_n1406_;
  assign new_n2862_ = ~new_n12237_ | ~new_n2333_;
  assign new_n2863_ = ~new_n10492_ | ~new_n2335_;
  assign new_n2864_ = ~new_n14082_ | ~new_n2334_;
  assign new_n2865_ = ~new_n12708_ | ~new_n2331_;
  assign new_n2866_ = ~new_n11167_ | ~new_n2330_;
  assign new_n2867_ = ~new_n13584_ | ~new_n2340_;
  assign new_n2868_ = ~new_n9701_ | ~new_n2339_;
  assign new_n2869_ = ~new_n1731_;
  assign new_n2870_ = ~new_n14580_ | ~new_n1365_;
  assign new_n2871_ = ~new_n1364_ | ~new_n1418_;
  assign new_n2872_ = ~new_n9447_ | ~new_n1362_;
  assign new_n2873_ = ~new_n1846_ | ~new_n2514_;
  assign new_n2874_ = ~new_n2045_ | ~new_n2869_;
  assign new_n2875_ = ~pi181 | ~new_n1357_;
  assign new_n2876_ = ~pi149 | ~new_n1358_;
  assign new_n2877_ = ~pi117 | ~new_n1359_;
  assign new_n2878_ = ~new_n8799_ | ~new_n1356_;
  assign new_n2879_ = ~new_n1413_;
  assign new_n2880_ = ~new_n1372_ | ~new_n1419_;
  assign new_n2881_ = ~new_n12236_ | ~new_n2333_;
  assign new_n2882_ = ~new_n10491_ | ~new_n2335_;
  assign new_n2883_ = ~new_n14081_ | ~new_n2334_;
  assign new_n2884_ = ~new_n12707_ | ~new_n2331_;
  assign new_n2885_ = ~new_n11166_ | ~new_n2330_;
  assign new_n2886_ = ~new_n13583_ | ~new_n2340_;
  assign new_n2887_ = ~new_n9700_ | ~new_n2339_;
  assign new_n2888_ = ~new_n1732_;
  assign new_n2889_ = ~new_n14579_ | ~new_n1365_;
  assign new_n2890_ = ~new_n1364_ | ~new_n1413_;
  assign new_n2891_ = ~new_n9517_ | ~new_n1362_;
  assign new_n2892_ = ~new_n1848_ | ~new_n2514_;
  assign new_n2893_ = ~new_n2049_ | ~new_n2888_;
  assign new_n2894_ = ~pi182 | ~new_n1357_;
  assign new_n2895_ = ~pi150 | ~new_n1358_;
  assign new_n2896_ = ~pi118 | ~new_n1359_;
  assign new_n2897_ = ~new_n8798_ | ~new_n1356_;
  assign new_n2898_ = ~new_n1412_;
  assign new_n2899_ = ~new_n1372_ | ~new_n1418_;
  assign new_n2900_ = ~new_n12234_ | ~new_n2333_;
  assign new_n2901_ = ~new_n10489_ | ~new_n2335_;
  assign new_n2902_ = ~new_n13986_ | ~new_n2334_;
  assign new_n2903_ = ~new_n12705_ | ~new_n2331_;
  assign new_n2904_ = ~new_n11164_ | ~new_n2330_;
  assign new_n2905_ = ~new_n13488_ | ~new_n2340_;
  assign new_n2906_ = ~new_n9605_ | ~new_n2339_;
  assign new_n2907_ = ~new_n1734_;
  assign new_n2908_ = ~new_n14484_ | ~new_n1365_;
  assign new_n2909_ = ~new_n1364_ | ~new_n1412_;
  assign new_n2910_ = ~new_n9448_ | ~new_n1362_;
  assign new_n2911_ = ~new_n2354_ | ~new_n2514_;
  assign new_n2912_ = ~new_n2053_ | ~new_n2907_;
  assign new_n2913_ = ~pi183 | ~new_n1357_;
  assign new_n2914_ = ~pi151 | ~new_n1358_;
  assign new_n2915_ = ~pi119 | ~new_n1359_;
  assign new_n2916_ = ~new_n8797_ | ~new_n1356_;
  assign new_n2917_ = ~new_n1398_;
  assign new_n2918_ = ~new_n1372_ | ~new_n1413_;
  assign new_n2919_ = ~new_n12248_ | ~new_n2333_;
  assign new_n2920_ = ~new_n10503_ | ~new_n2335_;
  assign new_n2921_ = ~new_n13987_ | ~new_n2334_;
  assign new_n2922_ = ~new_n12719_ | ~new_n2331_;
  assign new_n2923_ = ~new_n11178_ | ~new_n2330_;
  assign new_n2924_ = ~new_n13489_ | ~new_n2340_;
  assign new_n2925_ = ~new_n9606_ | ~new_n2339_;
  assign new_n2926_ = ~new_n1736_;
  assign new_n2927_ = ~new_n14485_ | ~new_n1365_;
  assign new_n2928_ = ~new_n1364_ | ~new_n1398_;
  assign new_n2929_ = ~new_n9513_ | ~new_n1362_;
  assign new_n2930_ = ~new_n2353_ | ~new_n2514_;
  assign new_n2931_ = ~new_n2057_ | ~new_n2926_;
  assign new_n2932_ = ~pi184 | ~new_n1357_;
  assign new_n2933_ = ~pi152 | ~new_n1358_;
  assign new_n2934_ = ~pi120 | ~new_n1359_;
  assign new_n2935_ = ~new_n8796_ | ~new_n1356_;
  assign new_n2936_ = ~new_n1403_;
  assign new_n2937_ = ~new_n1372_ | ~new_n1412_;
  assign new_n2938_ = ~new_n12247_ | ~new_n2333_;
  assign new_n2939_ = ~new_n10502_ | ~new_n2335_;
  assign new_n2940_ = ~new_n14080_ | ~new_n2334_;
  assign new_n2941_ = ~new_n12718_ | ~new_n2331_;
  assign new_n2942_ = ~new_n11177_ | ~new_n2330_;
  assign new_n2943_ = ~new_n13582_ | ~new_n2340_;
  assign new_n2944_ = ~new_n9699_ | ~new_n2339_;
  assign new_n2945_ = ~new_n1738_;
  assign new_n2946_ = ~new_n14578_ | ~new_n1365_;
  assign new_n2947_ = ~new_n1364_ | ~new_n1403_;
  assign new_n2948_ = ~new_n9449_ | ~new_n1362_;
  assign new_n2949_ = ~new_n2352_ | ~new_n2514_;
  assign new_n2950_ = ~new_n2061_ | ~new_n2945_;
  assign new_n2951_ = ~pi185 | ~new_n1357_;
  assign new_n2952_ = ~pi153 | ~new_n1358_;
  assign new_n2953_ = ~pi121 | ~new_n1359_;
  assign new_n2954_ = ~new_n8795_ | ~new_n1356_;
  assign new_n2955_ = ~new_n1402_;
  assign new_n2956_ = ~new_n1372_ | ~new_n1398_;
  assign new_n2957_ = ~new_n12152_ | ~new_n2333_;
  assign new_n2958_ = ~new_n10407_ | ~new_n2335_;
  assign new_n2959_ = ~new_n14079_ | ~new_n2334_;
  assign new_n2960_ = ~new_n12623_ | ~new_n2331_;
  assign new_n2961_ = ~new_n11082_ | ~new_n2330_;
  assign new_n2962_ = ~new_n13581_ | ~new_n2340_;
  assign new_n2963_ = ~new_n9698_ | ~new_n2339_;
  assign new_n2964_ = ~new_n1740_;
  assign new_n2965_ = ~new_n14577_ | ~new_n1365_;
  assign new_n2966_ = ~new_n1364_ | ~new_n1402_;
  assign new_n2967_ = ~new_n9511_ | ~new_n1362_;
  assign new_n2968_ = ~new_n2351_ | ~new_n2514_;
  assign new_n2969_ = ~new_n2065_ | ~new_n2964_;
  assign new_n2970_ = ~pi186 | ~new_n1357_;
  assign new_n2971_ = ~pi154 | ~new_n1358_;
  assign new_n2972_ = ~pi122 | ~new_n1359_;
  assign new_n2973_ = ~new_n8794_ | ~new_n1356_;
  assign new_n2974_ = ~new_n1395_;
  assign new_n2975_ = ~new_n1372_ | ~new_n1403_;
  assign new_n2976_ = ~new_n12233_ | ~new_n2333_;
  assign new_n2977_ = ~new_n10488_ | ~new_n2335_;
  assign new_n2978_ = ~new_n14078_ | ~new_n2334_;
  assign new_n2979_ = ~new_n12704_ | ~new_n2331_;
  assign new_n2980_ = ~new_n11163_ | ~new_n2330_;
  assign new_n2981_ = ~new_n13580_ | ~new_n2340_;
  assign new_n2982_ = ~new_n9697_ | ~new_n2339_;
  assign new_n2983_ = ~new_n1742_;
  assign new_n2984_ = ~new_n14576_ | ~new_n1365_;
  assign new_n2985_ = ~new_n1364_ | ~new_n1395_;
  assign new_n2986_ = ~new_n9450_ | ~new_n1362_;
  assign new_n2987_ = ~new_n2350_ | ~new_n2514_;
  assign new_n2988_ = ~new_n2069_ | ~new_n2983_;
  assign new_n2989_ = ~pi187 | ~new_n1357_;
  assign new_n2990_ = ~pi155 | ~new_n1358_;
  assign new_n2991_ = ~pi123 | ~new_n1359_;
  assign new_n2992_ = ~new_n8793_ | ~new_n1356_;
  assign new_n2993_ = ~new_n1394_;
  assign new_n2994_ = ~new_n1372_ | ~new_n1402_;
  assign new_n2995_ = ~new_n12232_ | ~new_n2333_;
  assign new_n2996_ = ~new_n10487_ | ~new_n2335_;
  assign new_n2997_ = ~new_n14077_ | ~new_n2334_;
  assign new_n2998_ = ~new_n12703_ | ~new_n2331_;
  assign new_n2999_ = ~new_n11162_ | ~new_n2330_;
  assign new_n3000_ = ~new_n13579_ | ~new_n2340_;
  assign new_n3001_ = ~new_n9696_ | ~new_n2339_;
  assign new_n3002_ = ~new_n1744_;
  assign new_n3003_ = ~new_n14575_ | ~new_n1365_;
  assign new_n3004_ = ~new_n1364_ | ~new_n1394_;
  assign new_n3005_ = ~new_n9509_ | ~new_n1362_;
  assign new_n3006_ = ~new_n2349_ | ~new_n2514_;
  assign new_n3007_ = ~new_n2073_ | ~new_n3002_;
  assign new_n3008_ = ~pi188 | ~new_n1357_;
  assign new_n3009_ = ~pi156 | ~new_n1358_;
  assign new_n3010_ = ~pi124 | ~new_n1359_;
  assign new_n3011_ = ~new_n8792_ | ~new_n1356_;
  assign new_n3012_ = ~new_n1390_;
  assign new_n3013_ = ~new_n1372_ | ~new_n1395_;
  assign new_n3014_ = ~new_n12246_ | ~new_n2333_;
  assign new_n3015_ = ~new_n10501_ | ~new_n2335_;
  assign new_n3016_ = ~new_n13988_ | ~new_n2334_;
  assign new_n3017_ = ~new_n12717_ | ~new_n2331_;
  assign new_n3018_ = ~new_n11176_ | ~new_n2330_;
  assign new_n3019_ = ~new_n13490_ | ~new_n2340_;
  assign new_n3020_ = ~new_n9607_ | ~new_n2339_;
  assign new_n3021_ = ~new_n1746_;
  assign new_n3022_ = ~new_n14486_ | ~new_n1365_;
  assign new_n3023_ = ~new_n1364_ | ~new_n1390_;
  assign new_n3024_ = ~new_n9451_ | ~new_n1362_;
  assign new_n3025_ = ~new_n2348_ | ~new_n2514_;
  assign new_n3026_ = ~new_n2077_ | ~new_n3021_;
  assign new_n3027_ = ~pi189 | ~new_n1357_;
  assign new_n3028_ = ~pi157 | ~new_n1358_;
  assign new_n3029_ = ~pi125 | ~new_n1359_;
  assign new_n3030_ = ~new_n8791_ | ~new_n1356_;
  assign new_n3031_ = ~new_n1391_;
  assign new_n3032_ = ~new_n1372_ | ~new_n1394_;
  assign new_n3033_ = ~new_n12153_ | ~new_n2333_;
  assign new_n3034_ = ~new_n10408_ | ~new_n2335_;
  assign new_n3035_ = ~new_n14076_ | ~new_n2334_;
  assign new_n3036_ = ~new_n12624_ | ~new_n2331_;
  assign new_n3037_ = ~new_n11083_ | ~new_n2330_;
  assign new_n3038_ = ~new_n13578_ | ~new_n2340_;
  assign new_n3039_ = ~new_n9695_ | ~new_n2339_;
  assign new_n3040_ = ~new_n1748_;
  assign new_n3041_ = ~new_n14574_ | ~new_n1365_;
  assign new_n3042_ = ~new_n1364_ | ~new_n1391_;
  assign new_n3043_ = ~new_n9507_ | ~new_n1362_;
  assign new_n3044_ = ~new_n2347_ | ~new_n2514_;
  assign new_n3045_ = ~new_n2081_ | ~new_n3040_;
  assign new_n3046_ = ~new_n8736_ | ~new_n1356_;
  assign new_n3047_ = ~pi190 | ~new_n1357_;
  assign new_n3048_ = ~pi158 | ~new_n1358_;
  assign new_n3049_ = ~pi126 | ~new_n1359_;
  assign new_n3050_ = ~new_n1392_;
  assign new_n3051_ = ~new_n1372_ | ~new_n1390_;
  assign new_n3052_ = ~new_n12231_ | ~new_n2333_;
  assign new_n3053_ = ~new_n10486_ | ~new_n2335_;
  assign new_n3054_ = ~new_n14075_ | ~new_n2334_;
  assign new_n3055_ = ~new_n12702_ | ~new_n2331_;
  assign new_n3056_ = ~new_n11161_ | ~new_n2330_;
  assign new_n3057_ = ~new_n13577_ | ~new_n2340_;
  assign new_n3058_ = ~new_n9694_ | ~new_n2339_;
  assign new_n3059_ = ~new_n1750_;
  assign new_n3060_ = ~new_n14573_ | ~new_n1365_;
  assign new_n3061_ = ~new_n1364_ | ~new_n1392_;
  assign new_n3062_ = ~new_n9452_ | ~new_n1362_;
  assign new_n3063_ = ~new_n2346_ | ~new_n2514_;
  assign new_n3064_ = ~new_n2085_ | ~new_n3059_;
  assign new_n3065_ = ~pi191 | ~new_n1357_;
  assign new_n3066_ = ~pi159 | ~new_n1358_;
  assign new_n3067_ = ~pi127 | ~new_n1359_;
  assign new_n3068_ = ~new_n1396_;
  assign new_n3069_ = ~new_n4067_ | ~new_n1697_;
  assign new_n3070_ = ~new_n2285_ | ~new_n3069_;
  assign new_n3071_ = ~new_n2086_ | ~new_n1396_;
  assign new_n3072_ = ~new_n1372_ | ~new_n1391_;
  assign new_n3073_ = ~new_n12154_ | ~new_n2333_;
  assign new_n3074_ = ~new_n10409_ | ~new_n2335_;
  assign new_n3075_ = ~new_n14074_ | ~new_n2334_;
  assign new_n3076_ = ~new_n12625_ | ~new_n2331_;
  assign new_n3077_ = ~new_n11084_ | ~new_n2330_;
  assign new_n3078_ = ~new_n13576_ | ~new_n2340_;
  assign new_n3079_ = ~new_n9693_ | ~new_n2339_;
  assign new_n3080_ = ~new_n1752_;
  assign new_n3081_ = ~new_n14572_ | ~new_n1365_;
  assign new_n3082_ = ~new_n9505_ | ~new_n1362_;
  assign new_n3083_ = ~new_n2357_ | ~new_n2514_;
  assign new_n3084_ = ~new_n2090_ | ~new_n3080_;
  assign new_n3085_ = ~pi192 | ~new_n1357_;
  assign new_n3086_ = ~pi160 | ~new_n1358_;
  assign new_n3087_ = ~pi128 | ~new_n1359_;
  assign new_n3088_ = ~new_n1393_;
  assign new_n3089_ = ~new_n9454_ | ~new_n1362_;
  assign new_n3090_ = ~new_n2356_ | ~new_n2514_;
  assign new_n3091_ = ~new_n3089_ | ~new_n3090_ | ~new_n2318_;
  assign new_n3092_ = ~new_n9503_ | ~new_n1362_;
  assign new_n3093_ = ~new_n2355_ | ~new_n2514_;
  assign new_n3094_ = ~new_n3092_ | ~new_n3093_ | ~new_n2318_;
  assign new_n3095_ = ~new_n2093_ | ~new_n1355_;
  assign new_n3096_ = ~new_n1757_ | ~new_n3095_;
  assign new_n3097_ = ~new_n2360_ | ~new_n1781_;
  assign new_n3098_ = ~new_n1761_;
  assign new_n3099_ = ~new_n1374_ | ~new_n1415_;
  assign new_n3100_ = ~new_n1371_ | ~pi255;
  assign new_n3101_ = ~new_n1370_ | ~new_n14566_;
  assign new_n3102_ = ~new_n1369_ | ~new_n1790_;
  assign new_n3103_ = ~new_n1368_ | ~new_n1790_;
  assign new_n3104_ = ~new_n1374_ | ~new_n1405_;
  assign new_n3105_ = ~new_n1371_ | ~pi265;
  assign new_n3106_ = ~new_n1370_ | ~new_n14565_;
  assign new_n3107_ = ~new_n1369_ | ~new_n1795_;
  assign new_n3108_ = ~new_n1368_ | ~new_n9492_;
  assign new_n3109_ = ~new_n1374_ | ~new_n1401_;
  assign new_n3110_ = ~new_n1371_ | ~pi250;
  assign new_n3111_ = ~new_n1370_ | ~new_n14487_;
  assign new_n3112_ = ~new_n1369_ | ~new_n1798_;
  assign new_n3113_ = ~new_n1368_ | ~new_n9453_;
  assign new_n3114_ = ~new_n1374_ | ~new_n1397_;
  assign new_n3115_ = ~new_n1371_ | ~new_n8735_;
  assign new_n3116_ = ~new_n1370_ | ~new_n14571_;
  assign new_n3117_ = ~new_n1369_ | ~new_n1801_;
  assign new_n3118_ = ~new_n1368_ | ~new_n9455_;
  assign new_n3119_ = ~new_n1374_ | ~new_n1404_;
  assign new_n3120_ = ~new_n1371_ | ~new_n8790_;
  assign new_n3121_ = ~new_n1370_ | ~new_n14570_;
  assign new_n3122_ = ~new_n1369_ | ~new_n1804_;
  assign new_n3123_ = ~new_n1368_ | ~new_n9456_;
  assign new_n3124_ = ~new_n1374_ | ~new_n1408_;
  assign new_n3125_ = ~new_n1371_ | ~new_n8789_;
  assign new_n3126_ = ~new_n1370_ | ~new_n14488_;
  assign new_n3127_ = ~new_n1369_ | ~new_n1807_;
  assign new_n3128_ = ~new_n1368_ | ~new_n9500_;
  assign new_n3129_ = ~new_n1374_ | ~new_n1407_;
  assign new_n3130_ = ~new_n1371_ | ~new_n8788_;
  assign new_n3131_ = ~new_n1370_ | ~new_n14569_;
  assign new_n3132_ = ~new_n1369_ | ~new_n1810_;
  assign new_n3133_ = ~new_n1368_ | ~new_n9457_;
  assign new_n3134_ = ~new_n1374_ | ~new_n1421_;
  assign new_n3135_ = ~new_n1371_ | ~new_n8787_;
  assign new_n3136_ = ~new_n1370_ | ~new_n14489_;
  assign new_n3137_ = ~new_n1369_ | ~new_n1813_;
  assign new_n3138_ = ~new_n1368_ | ~new_n9458_;
  assign new_n3139_ = ~new_n1374_ | ~new_n1420_;
  assign new_n3140_ = ~new_n1371_ | ~new_n8786_;
  assign new_n3141_ = ~new_n1370_ | ~new_n14568_;
  assign new_n3142_ = ~new_n1369_ | ~new_n1816_;
  assign new_n3143_ = ~new_n1368_ | ~new_n9459_;
  assign new_n3144_ = ~new_n1374_ | ~new_n1399_;
  assign new_n3145_ = ~new_n1371_ | ~new_n8785_;
  assign new_n3146_ = ~new_n1370_ | ~new_n14567_;
  assign new_n3147_ = ~new_n1369_ | ~new_n1819_;
  assign new_n3148_ = ~new_n1368_ | ~new_n9498_;
  assign new_n3149_ = ~new_n1374_ | ~new_n1400_;
  assign new_n3150_ = ~new_n1371_ | ~new_n8809_;
  assign new_n3151_ = ~new_n1370_ | ~new_n14481_;
  assign new_n3152_ = ~new_n1369_ | ~new_n1822_;
  assign new_n3153_ = ~new_n1368_ | ~new_n9441_;
  assign new_n3154_ = ~new_n1374_ | ~new_n1409_;
  assign new_n3155_ = ~new_n1371_ | ~new_n8808_;
  assign new_n3156_ = ~new_n1370_ | ~new_n14585_;
  assign new_n3157_ = ~new_n1369_ | ~new_n1825_;
  assign new_n3158_ = ~new_n1368_ | ~new_n9442_;
  assign new_n3159_ = ~new_n1374_ | ~new_n1417_;
  assign new_n3160_ = ~new_n1371_ | ~new_n8807_;
  assign new_n3161_ = ~new_n1370_ | ~new_n14584_;
  assign new_n3162_ = ~new_n1369_ | ~new_n1828_;
  assign new_n3163_ = ~new_n1368_ | ~new_n9443_;
  assign new_n3164_ = ~new_n1374_ | ~new_n1416_;
  assign new_n3165_ = ~new_n1371_ | ~new_n8806_;
  assign new_n3166_ = ~new_n1370_ | ~new_n14482_;
  assign new_n3167_ = ~new_n1369_ | ~new_n1831_;
  assign new_n3168_ = ~new_n1368_ | ~new_n9521_;
  assign new_n3169_ = ~new_n1374_ | ~new_n1411_;
  assign new_n3170_ = ~new_n1371_ | ~new_n8805_;
  assign new_n3171_ = ~new_n1370_ | ~new_n14583_;
  assign new_n3172_ = ~new_n1369_ | ~new_n1834_;
  assign new_n3173_ = ~new_n1368_ | ~new_n9444_;
  assign new_n3174_ = ~new_n1374_ | ~new_n1410_;
  assign new_n3175_ = ~new_n1371_ | ~new_n8804_;
  assign new_n3176_ = ~new_n1370_ | ~new_n14582_;
  assign new_n3177_ = ~new_n1369_ | ~new_n1837_;
  assign new_n3178_ = ~new_n1368_ | ~new_n9445_;
  assign new_n3179_ = ~new_n1374_ | ~new_n1406_;
  assign new_n3180_ = ~new_n1371_ | ~new_n8803_;
  assign new_n3181_ = ~new_n1370_ | ~new_n14581_;
  assign new_n3182_ = ~new_n1369_ | ~new_n1840_;
  assign new_n3183_ = ~new_n1368_ | ~new_n9446_;
  assign new_n3184_ = ~new_n1374_ | ~new_n1419_;
  assign new_n3185_ = ~new_n1371_ | ~new_n8802_;
  assign new_n3186_ = ~new_n1370_ | ~new_n14483_;
  assign new_n3187_ = ~new_n1369_ | ~new_n1843_;
  assign new_n3188_ = ~new_n1368_ | ~new_n9519_;
  assign new_n3189_ = ~new_n1374_ | ~new_n1418_;
  assign new_n3190_ = ~new_n1371_ | ~new_n8801_;
  assign new_n3191_ = ~new_n1370_ | ~new_n14580_;
  assign new_n3192_ = ~new_n1369_ | ~new_n1846_;
  assign new_n3193_ = ~new_n1368_ | ~new_n9447_;
  assign new_n3194_ = ~new_n1374_ | ~new_n1413_;
  assign new_n3195_ = ~new_n1371_ | ~new_n8800_;
  assign new_n3196_ = ~new_n1370_ | ~new_n14579_;
  assign new_n3197_ = ~new_n1369_ | ~new_n1848_;
  assign new_n3198_ = ~new_n1368_ | ~new_n9517_;
  assign new_n3199_ = ~new_n1374_ | ~new_n1412_;
  assign new_n3200_ = ~new_n1371_ | ~new_n8799_;
  assign new_n3201_ = ~new_n1370_ | ~new_n14484_;
  assign new_n3202_ = ~new_n1369_ | ~new_n2354_;
  assign new_n3203_ = ~new_n1368_ | ~new_n9448_;
  assign new_n3204_ = ~new_n1374_ | ~new_n1398_;
  assign new_n3205_ = ~new_n1371_ | ~new_n8798_;
  assign new_n3206_ = ~new_n1370_ | ~new_n14485_;
  assign new_n3207_ = ~new_n1369_ | ~new_n2353_;
  assign new_n3208_ = ~new_n1368_ | ~new_n9513_;
  assign new_n3209_ = ~new_n1374_ | ~new_n1403_;
  assign new_n3210_ = ~new_n1371_ | ~new_n8797_;
  assign new_n3211_ = ~new_n1370_ | ~new_n14578_;
  assign new_n3212_ = ~new_n1369_ | ~new_n2352_;
  assign new_n3213_ = ~new_n1368_ | ~new_n9449_;
  assign new_n3214_ = ~new_n1374_ | ~new_n1402_;
  assign new_n3215_ = ~new_n1371_ | ~new_n8796_;
  assign new_n3216_ = ~new_n1370_ | ~new_n14577_;
  assign new_n3217_ = ~new_n1369_ | ~new_n2351_;
  assign new_n3218_ = ~new_n1368_ | ~new_n9511_;
  assign new_n3219_ = ~new_n1374_ | ~new_n1395_;
  assign new_n3220_ = ~new_n1371_ | ~new_n8795_;
  assign new_n3221_ = ~new_n1370_ | ~new_n14576_;
  assign new_n3222_ = ~new_n1369_ | ~new_n2350_;
  assign new_n3223_ = ~new_n1368_ | ~new_n9450_;
  assign new_n3224_ = ~new_n1374_ | ~new_n1394_;
  assign new_n3225_ = ~new_n1371_ | ~new_n8794_;
  assign new_n3226_ = ~new_n1370_ | ~new_n14575_;
  assign new_n3227_ = ~new_n1369_ | ~new_n2349_;
  assign new_n3228_ = ~new_n1368_ | ~new_n9509_;
  assign new_n3229_ = ~new_n1374_ | ~new_n1390_;
  assign new_n3230_ = ~new_n1371_ | ~new_n8793_;
  assign new_n3231_ = ~new_n1370_ | ~new_n14486_;
  assign new_n3232_ = ~new_n1369_ | ~new_n2348_;
  assign new_n3233_ = ~new_n1368_ | ~new_n9451_;
  assign new_n3234_ = ~new_n1374_ | ~new_n1391_;
  assign new_n3235_ = ~new_n1371_ | ~new_n8792_;
  assign new_n3236_ = ~new_n1370_ | ~new_n14574_;
  assign new_n3237_ = ~new_n1369_ | ~new_n2347_;
  assign new_n3238_ = ~new_n1368_ | ~new_n9507_;
  assign new_n3239_ = ~new_n1374_ | ~new_n1392_;
  assign new_n3240_ = ~new_n1371_ | ~new_n8791_;
  assign new_n3241_ = ~new_n1370_ | ~new_n14573_;
  assign new_n3242_ = ~new_n1369_ | ~new_n2346_;
  assign new_n3243_ = ~new_n1368_ | ~new_n9452_;
  assign new_n3244_ = ~new_n1371_ | ~new_n8736_;
  assign new_n3245_ = ~new_n1370_ | ~new_n14572_;
  assign new_n3246_ = ~new_n1369_ | ~new_n2357_;
  assign new_n3247_ = ~new_n1368_ | ~new_n9505_;
  assign new_n3248_ = ~new_n1369_ | ~new_n2356_;
  assign new_n3249_ = ~new_n1368_ | ~new_n9454_;
  assign new_n3250_ = ~new_n1369_ | ~new_n2355_;
  assign new_n3251_ = ~new_n1368_ | ~new_n9503_;
  assign new_n3252_ = ~new_n1757_ | ~new_n3098_ | ~new_n2155_ | ~new_n2153_ | ~new_n2152_;
  assign new_n3253_ = ~new_n8894_ | ~new_n1380_;
  assign new_n3254_ = ~new_n1378_ | ~new_n1782_;
  assign new_n3255_ = ~new_n10102_ | ~new_n1376_;
  assign new_n3256_ = ~new_n3255_ | ~new_n3254_ | ~new_n3253_;
  assign new_n3257_ = ~new_n1385_ | ~new_n1711_;
  assign new_n3258_ = ~new_n4042_ | ~new_n3257_;
  assign new_n3259_ = ~new_n3258_ | ~new_n2285_;
  assign new_n3260_ = ~po265;
  assign new_n3261_ = ~new_n1762_;
  assign new_n3262_ = ~new_n1382_ | ~new_n3256_;
  assign new_n3263_ = ~new_n1381_ | ~new_n8894_;
  assign new_n3264_ = ~pi268 | ~po264;
  assign new_n3265_ = ~new_n1379_ | ~new_n1782_;
  assign new_n3266_ = ~new_n1377_ | ~new_n10102_;
  assign new_n3267_ = ~pi193 | ~new_n3261_;
  assign new_n3268_ = ~new_n8956_ | ~new_n1380_;
  assign new_n3269_ = ~new_n1378_ | ~new_n1845_;
  assign new_n3270_ = ~new_n10164_ | ~new_n1376_;
  assign new_n3271_ = ~new_n3270_ | ~new_n3269_ | ~new_n3268_;
  assign new_n3272_ = ~new_n1382_ | ~new_n3271_;
  assign new_n3273_ = ~new_n8956_ | ~new_n1381_;
  assign new_n3274_ = ~pi249 | ~po264;
  assign new_n3275_ = ~new_n1379_ | ~new_n1845_;
  assign new_n3276_ = ~new_n10164_ | ~new_n1377_;
  assign new_n3277_ = ~pi194 | ~new_n3261_;
  assign new_n3278_ = ~new_n8893_ | ~new_n1380_;
  assign new_n3279_ = ~new_n1378_ | ~new_n1842_;
  assign new_n3280_ = ~new_n10101_ | ~new_n1376_;
  assign new_n3281_ = ~new_n3280_ | ~new_n3279_ | ~new_n3278_;
  assign new_n3282_ = ~new_n1382_ | ~new_n3281_;
  assign new_n3283_ = ~new_n8893_ | ~new_n1381_;
  assign new_n3284_ = ~pi259 | ~po264;
  assign new_n3285_ = ~new_n1379_ | ~new_n1842_;
  assign new_n3286_ = ~new_n10101_ | ~new_n1377_;
  assign new_n3287_ = ~pi195 | ~new_n3261_;
  assign new_n3288_ = ~new_n8957_ | ~new_n1380_;
  assign new_n3289_ = ~new_n1378_ | ~new_n1839_;
  assign new_n3290_ = ~new_n10165_ | ~new_n1376_;
  assign new_n3291_ = ~new_n3290_ | ~new_n3289_ | ~new_n3288_;
  assign new_n3292_ = ~new_n1382_ | ~new_n3291_;
  assign new_n3293_ = ~new_n8957_ | ~new_n1381_;
  assign new_n3294_ = ~pi261 | ~po264;
  assign new_n3295_ = ~new_n1379_ | ~new_n1839_;
  assign new_n3296_ = ~new_n10165_ | ~new_n1377_;
  assign new_n3297_ = ~pi196 | ~new_n3261_;
  assign new_n3298_ = ~new_n8958_ | ~new_n1380_;
  assign new_n3299_ = ~new_n1378_ | ~new_n1836_;
  assign new_n3300_ = ~new_n10166_ | ~new_n1376_;
  assign new_n3301_ = ~new_n3300_ | ~new_n3299_ | ~new_n3298_;
  assign new_n3302_ = ~new_n1382_ | ~new_n3301_;
  assign new_n3303_ = ~new_n8958_ | ~new_n1381_;
  assign new_n3304_ = ~pi246 | ~po264;
  assign new_n3305_ = ~new_n1379_ | ~new_n1836_;
  assign new_n3306_ = ~new_n10166_ | ~new_n1377_;
  assign new_n3307_ = ~pi197 | ~new_n3261_;
  assign new_n3308_ = ~new_n8959_ | ~new_n1380_;
  assign new_n3309_ = ~new_n1378_ | ~new_n1833_;
  assign new_n3310_ = ~new_n10167_ | ~new_n1376_;
  assign new_n3311_ = ~new_n3310_ | ~new_n3309_ | ~new_n3308_;
  assign new_n3312_ = ~new_n1382_ | ~new_n3311_;
  assign new_n3313_ = ~new_n8959_ | ~new_n1381_;
  assign new_n3314_ = ~pi272 | ~po264;
  assign new_n3315_ = ~new_n1379_ | ~new_n1833_;
  assign new_n3316_ = ~new_n10167_ | ~new_n1377_;
  assign new_n3317_ = ~pi198 | ~new_n3261_;
  assign new_n3318_ = ~new_n8892_ | ~new_n1380_;
  assign new_n3319_ = ~new_n1378_ | ~new_n1830_;
  assign new_n3320_ = ~new_n10100_ | ~new_n1376_;
  assign new_n3321_ = ~new_n3320_ | ~new_n3319_ | ~new_n3318_;
  assign new_n3322_ = ~new_n1382_ | ~new_n3321_;
  assign new_n3323_ = ~new_n8892_ | ~new_n1381_;
  assign new_n3324_ = ~pi253 | ~po264;
  assign new_n3325_ = ~new_n1379_ | ~new_n1830_;
  assign new_n3326_ = ~new_n10100_ | ~new_n1377_;
  assign new_n3327_ = ~pi199 | ~new_n3261_;
  assign new_n3328_ = ~new_n8960_ | ~new_n1380_;
  assign new_n3329_ = ~new_n1378_ | ~new_n1827_;
  assign new_n3330_ = ~new_n10168_ | ~new_n1376_;
  assign new_n3331_ = ~new_n3330_ | ~new_n3329_ | ~new_n3328_;
  assign new_n3332_ = ~new_n1382_ | ~new_n3331_;
  assign new_n3333_ = ~new_n8960_ | ~new_n1381_;
  assign new_n3334_ = ~pi263 | ~po264;
  assign new_n3335_ = ~new_n1379_ | ~new_n1827_;
  assign new_n3336_ = ~new_n10168_ | ~new_n1377_;
  assign new_n3337_ = ~pi200 | ~new_n3261_;
  assign new_n3338_ = ~new_n8961_ | ~new_n1380_;
  assign new_n3339_ = ~new_n1378_ | ~new_n1824_;
  assign new_n3340_ = ~new_n10169_ | ~new_n1376_;
  assign new_n3341_ = ~new_n3340_ | ~new_n3339_ | ~new_n3338_;
  assign new_n3342_ = ~new_n1382_ | ~new_n3341_;
  assign new_n3343_ = ~new_n8961_ | ~new_n1381_;
  assign new_n3344_ = ~pi251 | ~po264;
  assign new_n3345_ = ~new_n1379_ | ~new_n1824_;
  assign new_n3346_ = ~new_n10169_ | ~new_n1377_;
  assign new_n3347_ = ~pi201 | ~new_n3261_;
  assign new_n3348_ = ~new_n8891_ | ~new_n1380_;
  assign new_n3349_ = ~new_n1378_ | ~new_n1821_;
  assign new_n3350_ = ~new_n10099_ | ~new_n1376_;
  assign new_n3351_ = ~new_n3350_ | ~new_n3349_ | ~new_n3348_;
  assign new_n3352_ = ~new_n1382_ | ~new_n3351_;
  assign new_n3353_ = ~new_n8891_ | ~new_n1381_;
  assign new_n3354_ = ~pi270 | ~po264;
  assign new_n3355_ = ~new_n1379_ | ~new_n1821_;
  assign new_n3356_ = ~new_n10099_ | ~new_n1377_;
  assign new_n3357_ = ~pi202 | ~new_n3261_;
  assign new_n3358_ = ~new_n8951_ | ~new_n1380_;
  assign new_n3359_ = ~new_n1378_ | ~new_n1818_;
  assign new_n3360_ = ~new_n10159_ | ~new_n1376_;
  assign new_n3361_ = ~new_n3360_ | ~new_n3359_ | ~new_n3358_;
  assign new_n3362_ = ~new_n1382_ | ~new_n3361_;
  assign new_n3363_ = ~new_n8951_ | ~new_n1381_;
  assign new_n3364_ = ~pi256 | ~po264;
  assign new_n3365_ = ~new_n1379_ | ~new_n1818_;
  assign new_n3366_ = ~new_n10159_ | ~new_n1377_;
  assign new_n3367_ = ~pi203 | ~new_n3261_;
  assign new_n3368_ = ~new_n8952_ | ~new_n1380_;
  assign new_n3369_ = ~new_n1378_ | ~new_n1815_;
  assign new_n3370_ = ~new_n10160_ | ~new_n1376_;
  assign new_n3371_ = ~new_n3370_ | ~new_n3369_ | ~new_n3368_;
  assign new_n3372_ = ~new_n1382_ | ~new_n3371_;
  assign new_n3373_ = ~new_n8952_ | ~new_n1381_;
  assign new_n3374_ = ~pi266 | ~po264;
  assign new_n3375_ = ~new_n1379_ | ~new_n1815_;
  assign new_n3376_ = ~new_n10160_ | ~new_n1377_;
  assign new_n3377_ = ~pi204 | ~new_n3261_;
  assign new_n3378_ = ~new_n8897_ | ~new_n1380_;
  assign new_n3379_ = ~new_n1378_ | ~new_n1812_;
  assign new_n3380_ = ~new_n10105_ | ~new_n1376_;
  assign new_n3381_ = ~new_n3380_ | ~new_n3379_ | ~new_n3378_;
  assign new_n3382_ = ~new_n1382_ | ~new_n3381_;
  assign new_n3383_ = ~new_n8897_ | ~new_n1381_;
  assign new_n3384_ = ~pi274 | ~po264;
  assign new_n3385_ = ~new_n1379_ | ~new_n1812_;
  assign new_n3386_ = ~new_n10105_ | ~new_n1377_;
  assign new_n3387_ = ~pi205 | ~new_n3261_;
  assign new_n3388_ = ~new_n8953_ | ~new_n1380_;
  assign new_n3389_ = ~new_n1378_ | ~new_n1809_;
  assign new_n3390_ = ~new_n10161_ | ~new_n1376_;
  assign new_n3391_ = ~new_n3390_ | ~new_n3389_ | ~new_n3388_;
  assign new_n3392_ = ~new_n1382_ | ~new_n3391_;
  assign new_n3393_ = ~new_n8953_ | ~new_n1381_;
  assign new_n3394_ = ~pi248 | ~po264;
  assign new_n3395_ = ~new_n1379_ | ~new_n1809_;
  assign new_n3396_ = ~new_n10161_ | ~new_n1377_;
  assign new_n3397_ = ~pi206 | ~new_n3261_;
  assign new_n3398_ = ~new_n8896_ | ~new_n1380_;
  assign new_n3399_ = ~new_n1378_ | ~new_n1806_;
  assign new_n3400_ = ~new_n10104_ | ~new_n1376_;
  assign new_n3401_ = ~new_n3400_ | ~new_n3399_ | ~new_n3398_;
  assign new_n3402_ = ~new_n1382_ | ~new_n3401_;
  assign new_n3403_ = ~new_n8896_ | ~new_n1381_;
  assign new_n3404_ = ~pi260 | ~po264;
  assign new_n3405_ = ~new_n1379_ | ~new_n1806_;
  assign new_n3406_ = ~new_n10104_ | ~new_n1377_;
  assign new_n3407_ = ~pi207 | ~new_n3261_;
  assign new_n3408_ = ~new_n8954_ | ~new_n1380_;
  assign new_n3409_ = ~new_n1378_ | ~new_n1803_;
  assign new_n3410_ = ~new_n10162_ | ~new_n1376_;
  assign new_n3411_ = ~new_n3410_ | ~new_n3409_ | ~new_n3408_;
  assign new_n3412_ = ~new_n1382_ | ~new_n3411_;
  assign new_n3413_ = ~new_n8954_ | ~new_n1381_;
  assign new_n3414_ = ~pi257 | ~po264;
  assign new_n3415_ = ~new_n1379_ | ~new_n1803_;
  assign new_n3416_ = ~new_n10162_ | ~new_n1377_;
  assign new_n3417_ = ~pi208 | ~new_n3261_;
  assign new_n3418_ = ~new_n8955_ | ~new_n1380_;
  assign new_n3419_ = ~new_n1378_ | ~new_n1800_;
  assign new_n3420_ = ~new_n10163_ | ~new_n1376_;
  assign new_n3421_ = ~new_n3420_ | ~new_n3419_ | ~new_n3418_;
  assign new_n3422_ = ~new_n1382_ | ~new_n3421_;
  assign new_n3423_ = ~new_n8955_ | ~new_n1381_;
  assign new_n3424_ = ~pi269 | ~po264;
  assign new_n3425_ = ~new_n1379_ | ~new_n1800_;
  assign new_n3426_ = ~new_n10163_ | ~new_n1377_;
  assign new_n3427_ = ~pi209 | ~new_n3261_;
  assign new_n3428_ = ~new_n8895_ | ~new_n1380_;
  assign new_n3429_ = ~new_n1378_ | ~new_n1797_;
  assign new_n3430_ = ~new_n10103_ | ~new_n1376_;
  assign new_n3431_ = ~new_n3430_ | ~new_n3429_ | ~new_n3428_;
  assign new_n3432_ = ~new_n1382_ | ~new_n3431_;
  assign new_n3433_ = ~new_n8895_ | ~new_n1381_;
  assign new_n3434_ = ~pi250 | ~po264;
  assign new_n3435_ = ~new_n1379_ | ~new_n1797_;
  assign new_n3436_ = ~new_n10103_ | ~new_n1377_;
  assign new_n3437_ = ~pi210 | ~new_n3261_;
  assign new_n3438_ = ~new_n8949_ | ~new_n1380_;
  assign new_n3439_ = ~new_n1378_ | ~new_n1794_;
  assign new_n3440_ = ~new_n10157_ | ~new_n1376_;
  assign new_n3441_ = ~new_n3440_ | ~new_n3439_ | ~new_n3438_;
  assign new_n3442_ = ~new_n1382_ | ~new_n3441_;
  assign new_n3443_ = ~new_n8949_ | ~new_n1381_;
  assign new_n3444_ = ~pi265 | ~po264;
  assign new_n3445_ = ~new_n1379_ | ~new_n1794_;
  assign new_n3446_ = ~new_n10157_ | ~new_n1377_;
  assign new_n3447_ = ~pi211 | ~new_n3261_;
  assign new_n3448_ = ~new_n8950_ | ~new_n1380_;
  assign new_n3449_ = ~new_n1378_ | ~new_n1788_;
  assign new_n3450_ = ~new_n10158_ | ~new_n1376_;
  assign new_n3451_ = ~new_n3450_ | ~new_n3449_ | ~new_n3448_;
  assign new_n3452_ = ~new_n1382_ | ~new_n3451_;
  assign new_n3453_ = ~new_n8950_ | ~new_n1381_;
  assign new_n3454_ = ~pi255 | ~po264;
  assign new_n3455_ = ~new_n1379_ | ~new_n1788_;
  assign new_n3456_ = ~new_n10158_ | ~new_n1377_;
  assign new_n3457_ = ~pi212 | ~new_n3261_;
  assign new_n3458_ = ~new_n2321_;
  assign new_n3459_ = ~new_n2214_ | ~new_n4537_ | ~new_n4536_;
  assign new_n3460_ = ~new_n4042_ | ~new_n1766_;
  assign new_n3461_ = ~new_n2200_ | ~new_n3460_;
  assign new_n3462_ = ~pi245 | ~new_n3461_;
  assign new_n3463_ = ~new_n1375_ | ~new_n1416_;
  assign new_n3464_ = ~new_n1373_ | ~new_n1410_;
  assign new_n3465_ = ~new_n8804_ | ~new_n1770_;
  assign new_n3466_ = ~new_n3464_ | ~new_n3465_ | ~new_n3463_;
  assign new_n3467_ = ~new_n1700_ | ~new_n1702_ | ~new_n1699_;
  assign new_n3468_ = ~new_n1703_ | ~new_n1704_ | ~new_n1758_;
  assign new_n3469_ = ~new_n4049_ | ~new_n3468_;
  assign new_n3470_ = ~new_n4058_ | ~new_n3467_;
  assign new_n3471_ = ~new_n2216_ | ~new_n3470_ | ~new_n3469_;
  assign new_n3472_ = ~new_n3471_ | ~new_n1770_;
  assign new_n3473_ = ~new_n1772_;
  assign new_n3474_ = ~new_n1837_ | ~new_n4025_;
  assign new_n3475_ = ~new_n8804_ | ~new_n4024_;
  assign new_n3476_ = ~new_n2366_ | ~new_n3466_;
  assign new_n3477_ = ~new_n11644_ | ~new_n1366_;
  assign new_n3478_ = ~pi246 | ~po264;
  assign new_n3479_ = ~new_n1375_ | ~new_n1395_;
  assign new_n3480_ = ~new_n1373_ | ~new_n1390_;
  assign new_n3481_ = ~new_n8793_ | ~new_n1770_;
  assign new_n3482_ = ~new_n3480_ | ~new_n3481_ | ~new_n3479_;
  assign new_n3483_ = ~new_n1761_ | ~new_n1770_;
  assign new_n3484_ = ~new_n3473_ | ~new_n3483_;
  assign new_n3485_ = ~new_n2344_ | ~new_n1761_;
  assign new_n3486_ = ~new_n1757_ | ~new_n3485_;
  assign new_n3487_ = ~new_n1384_ | ~new_n2348_;
  assign new_n3488_ = ~new_n1383_ | ~new_n8793_;
  assign new_n3489_ = ~new_n2366_ | ~new_n3482_;
  assign new_n3490_ = ~new_n11553_ | ~new_n1366_;
  assign new_n3491_ = ~pi247 | ~po264;
  assign new_n3492_ = ~new_n1375_ | ~new_n1404_;
  assign new_n3493_ = ~new_n1373_ | ~new_n1407_;
  assign new_n3494_ = ~new_n8788_ | ~new_n1770_;
  assign new_n3495_ = ~new_n3494_ | ~new_n3493_ | ~new_n3492_;
  assign new_n3496_ = ~new_n1810_ | ~new_n4025_;
  assign new_n3497_ = ~new_n8788_ | ~new_n4024_;
  assign new_n3498_ = ~new_n2366_ | ~new_n3495_;
  assign new_n3499_ = ~new_n11629_ | ~new_n1366_;
  assign new_n3500_ = ~pi248 | ~po264;
  assign new_n3501_ = ~new_n1375_ | ~new_n1406_;
  assign new_n3502_ = ~new_n1373_ | ~new_n1418_;
  assign new_n3503_ = ~new_n8801_ | ~new_n1770_;
  assign new_n3504_ = ~new_n3502_ | ~new_n3503_ | ~new_n3501_;
  assign new_n3505_ = ~new_n1846_ | ~new_n4025_;
  assign new_n3506_ = ~new_n8801_ | ~new_n4024_;
  assign new_n3507_ = ~new_n2366_ | ~new_n3504_;
  assign new_n3508_ = ~new_n11642_ | ~new_n1366_;
  assign new_n3509_ = ~pi249 | ~po264;
  assign new_n3510_ = ~new_n1375_ | ~new_n1415_;
  assign new_n3511_ = ~new_n1373_ | ~new_n1401_;
  assign new_n3512_ = ~pi250 | ~new_n1770_;
  assign new_n3513_ = ~new_n3512_ | ~new_n3511_ | ~new_n3510_;
  assign new_n3514_ = ~new_n1798_ | ~new_n4025_;
  assign new_n3515_ = ~pi250 | ~new_n4024_;
  assign new_n3516_ = ~new_n2366_ | ~new_n3513_;
  assign new_n3517_ = ~new_n11632_ | ~new_n1366_;
  assign new_n3518_ = ~pi250 | ~po264;
  assign new_n3519_ = ~new_n1375_ | ~new_n1399_;
  assign new_n3520_ = ~new_n1373_ | ~new_n1409_;
  assign new_n3521_ = ~new_n8808_ | ~new_n1770_;
  assign new_n3522_ = ~new_n3521_ | ~new_n3520_ | ~new_n3519_;
  assign new_n3523_ = ~new_n1825_ | ~new_n4025_;
  assign new_n3524_ = ~new_n8808_ | ~new_n4024_;
  assign new_n3525_ = ~new_n2366_ | ~new_n3522_;
  assign new_n3526_ = ~new_n11647_ | ~new_n1366_;
  assign new_n3527_ = ~pi251 | ~po264;
  assign new_n3528_ = ~new_n1375_ | ~new_n1412_;
  assign new_n3529_ = ~new_n1373_ | ~new_n1403_;
  assign new_n3530_ = ~new_n8797_ | ~new_n1770_;
  assign new_n3531_ = ~new_n3529_ | ~new_n3530_ | ~new_n3528_;
  assign new_n3532_ = ~new_n1384_ | ~new_n2352_;
  assign new_n3533_ = ~new_n1383_ | ~new_n8797_;
  assign new_n3534_ = ~new_n2366_ | ~new_n3531_;
  assign new_n3535_ = ~new_n11638_ | ~new_n1366_;
  assign new_n3536_ = ~pi252 | ~po264;
  assign new_n3537_ = ~new_n1375_ | ~new_n1409_;
  assign new_n3538_ = ~new_n1373_ | ~new_n1416_;
  assign new_n3539_ = ~new_n8806_ | ~new_n1770_;
  assign new_n3540_ = ~new_n3538_ | ~new_n3539_ | ~new_n3537_;
  assign new_n3541_ = ~new_n1831_ | ~new_n4025_;
  assign new_n3542_ = ~new_n8806_ | ~new_n4024_;
  assign new_n3543_ = ~new_n2366_ | ~new_n3540_;
  assign new_n3544_ = ~new_n11550_ | ~new_n1366_;
  assign new_n3545_ = ~pi253 | ~po264;
  assign new_n3546_ = ~new_n1375_ | ~new_n1418_;
  assign new_n3547_ = ~new_n1373_ | ~new_n1412_;
  assign new_n3548_ = ~new_n8799_ | ~new_n1770_;
  assign new_n3549_ = ~new_n3547_ | ~new_n3548_ | ~new_n3546_;
  assign new_n3550_ = ~new_n1384_ | ~new_n2354_;
  assign new_n3551_ = ~new_n1383_ | ~new_n8799_;
  assign new_n3552_ = ~new_n2366_ | ~new_n3549_;
  assign new_n3553_ = ~new_n11639_ | ~new_n1366_;
  assign new_n3554_ = ~pi254 | ~po264;
  assign new_n3555_ = ~new_n1771_ | ~new_n1769_;
  assign new_n3556_ = ~new_n3555_ | ~new_n1770_;
  assign new_n3557_ = ~new_n2367_ | ~new_n3556_;
  assign new_n3558_ = ~new_n2222_ | ~new_n1373_;
  assign new_n3559_ = ~new_n1790_ | ~new_n4025_;
  assign new_n3560_ = ~pi255 | ~new_n3557_;
  assign new_n3561_ = ~new_n11626_ | ~new_n1366_;
  assign new_n3562_ = ~pi255 | ~po264;
  assign new_n3563_ = ~new_n1375_ | ~new_n1421_;
  assign new_n3564_ = ~new_n1373_ | ~new_n1399_;
  assign new_n3565_ = ~new_n8785_ | ~new_n1770_;
  assign new_n3566_ = ~new_n3565_ | ~new_n3564_ | ~new_n3563_;
  assign new_n3567_ = ~new_n1819_ | ~new_n4025_;
  assign new_n3568_ = ~new_n8785_ | ~new_n4024_;
  assign new_n3569_ = ~new_n2366_ | ~new_n3566_;
  assign new_n3570_ = ~new_n11627_ | ~new_n1366_;
  assign new_n3571_ = ~pi256 | ~po264;
  assign new_n3572_ = ~new_n1375_ | ~new_n1401_;
  assign new_n3573_ = ~new_n1373_ | ~new_n1404_;
  assign new_n3574_ = ~new_n8790_ | ~new_n1770_;
  assign new_n3575_ = ~new_n3574_ | ~new_n3573_ | ~new_n3572_;
  assign new_n3576_ = ~new_n1804_ | ~new_n4025_;
  assign new_n3577_ = ~new_n8790_ | ~new_n4024_;
  assign new_n3578_ = ~new_n2366_ | ~new_n3575_;
  assign new_n3579_ = ~new_n11631_ | ~new_n1366_;
  assign new_n3580_ = ~pi257 | ~po264;
  assign new_n3581_ = ~new_n1375_ | ~new_n1403_;
  assign new_n3582_ = ~new_n1373_ | ~new_n1395_;
  assign new_n3583_ = ~new_n8795_ | ~new_n1770_;
  assign new_n3584_ = ~new_n3582_ | ~new_n3583_ | ~new_n3581_;
  assign new_n3585_ = ~new_n1384_ | ~new_n2350_;
  assign new_n3586_ = ~new_n1383_ | ~new_n8795_;
  assign new_n3587_ = ~new_n2366_ | ~new_n3584_;
  assign new_n3588_ = ~new_n11636_ | ~new_n1366_;
  assign new_n3589_ = ~pi258 | ~po264;
  assign new_n3590_ = ~new_n1375_ | ~new_n1410_;
  assign new_n3591_ = ~new_n1373_ | ~new_n1419_;
  assign new_n3592_ = ~new_n8802_ | ~new_n1770_;
  assign new_n3593_ = ~new_n3591_ | ~new_n3592_ | ~new_n3590_;
  assign new_n3594_ = ~new_n1843_ | ~new_n4025_;
  assign new_n3595_ = ~new_n8802_ | ~new_n4024_;
  assign new_n3596_ = ~new_n2366_ | ~new_n3593_;
  assign new_n3597_ = ~new_n11551_ | ~new_n1366_;
  assign new_n3598_ = ~pi259 | ~po264;
  assign new_n3599_ = ~new_n1375_ | ~new_n1397_;
  assign new_n3600_ = ~new_n1373_ | ~new_n1408_;
  assign new_n3601_ = ~new_n8789_ | ~new_n1770_;
  assign new_n3602_ = ~new_n3601_ | ~new_n3600_ | ~new_n3599_;
  assign new_n3603_ = ~new_n1807_ | ~new_n4025_;
  assign new_n3604_ = ~new_n8789_ | ~new_n4024_;
  assign new_n3605_ = ~new_n2366_ | ~new_n3602_;
  assign new_n3606_ = ~new_n11630_ | ~new_n1366_;
  assign new_n3607_ = ~pi260 | ~po264;
  assign new_n3608_ = ~new_n1375_ | ~new_n1411_;
  assign new_n3609_ = ~new_n1373_ | ~new_n1406_;
  assign new_n3610_ = ~new_n8803_ | ~new_n1770_;
  assign new_n3611_ = ~new_n3609_ | ~new_n3610_ | ~new_n3608_;
  assign new_n3612_ = ~new_n1840_ | ~new_n4025_;
  assign new_n3613_ = ~new_n8803_ | ~new_n4024_;
  assign new_n3614_ = ~new_n2366_ | ~new_n3611_;
  assign new_n3615_ = ~new_n11643_ | ~new_n1366_;
  assign new_n3616_ = ~pi261 | ~po264;
  assign new_n3617_ = ~new_n1375_ | ~new_n1402_;
  assign new_n3618_ = ~new_n1373_ | ~new_n1394_;
  assign new_n3619_ = ~new_n8794_ | ~new_n1770_;
  assign new_n3620_ = ~new_n3618_ | ~new_n3619_ | ~new_n3617_;
  assign new_n3621_ = ~new_n1384_ | ~new_n2349_;
  assign new_n3622_ = ~new_n1383_ | ~new_n8794_;
  assign new_n3623_ = ~new_n2366_ | ~new_n3620_;
  assign new_n3624_ = ~new_n11635_ | ~new_n1366_;
  assign new_n3625_ = ~pi262 | ~po264;
  assign new_n3626_ = ~new_n1375_ | ~new_n1400_;
  assign new_n3627_ = ~new_n1373_ | ~new_n1417_;
  assign new_n3628_ = ~new_n8807_ | ~new_n1770_;
  assign new_n3629_ = ~new_n3627_ | ~new_n3628_ | ~new_n3626_;
  assign new_n3630_ = ~new_n1828_ | ~new_n4025_;
  assign new_n3631_ = ~new_n8807_ | ~new_n4024_;
  assign new_n3632_ = ~new_n2366_ | ~new_n3629_;
  assign new_n3633_ = ~new_n11646_ | ~new_n1366_;
  assign new_n3634_ = ~pi263 | ~po264;
  assign new_n3635_ = ~new_n1375_ | ~new_n1413_;
  assign new_n3636_ = ~new_n1373_ | ~new_n1398_;
  assign new_n3637_ = ~new_n8798_ | ~new_n1770_;
  assign new_n3638_ = ~new_n3636_ | ~new_n3637_ | ~new_n3635_;
  assign new_n3639_ = ~new_n1384_ | ~new_n2353_;
  assign new_n3640_ = ~new_n1383_ | ~new_n8798_;
  assign new_n3641_ = ~new_n2366_ | ~new_n3638_;
  assign new_n3642_ = ~new_n11552_ | ~new_n1366_;
  assign new_n3643_ = ~pi264 | ~po264;
  assign new_n3644_ = ~new_n1375_ | ~new_n1414_;
  assign new_n3645_ = ~new_n1373_ | ~new_n1405_;
  assign new_n3646_ = ~pi265 | ~new_n1770_;
  assign new_n3647_ = ~new_n3646_ | ~new_n3645_ | ~new_n3644_;
  assign new_n3648_ = ~new_n1795_ | ~new_n4025_;
  assign new_n3649_ = ~pi265 | ~new_n4024_;
  assign new_n3650_ = ~new_n2366_ | ~new_n3647_;
  assign new_n3651_ = ~new_n11640_ | ~new_n1366_;
  assign new_n3652_ = ~pi265 | ~po264;
  assign new_n3653_ = ~new_n1375_ | ~new_n1407_;
  assign new_n3654_ = ~new_n1373_ | ~new_n1420_;
  assign new_n3655_ = ~new_n8786_ | ~new_n1770_;
  assign new_n3656_ = ~new_n3655_ | ~new_n3654_ | ~new_n3653_;
  assign new_n3657_ = ~new_n1816_ | ~new_n4025_;
  assign new_n3658_ = ~new_n8786_ | ~new_n4024_;
  assign new_n3659_ = ~new_n2366_ | ~new_n3656_;
  assign new_n3660_ = ~new_n11628_ | ~new_n1366_;
  assign new_n3661_ = ~pi266 | ~po264;
  assign new_n3662_ = ~new_n1375_ | ~new_n1390_;
  assign new_n3663_ = ~new_n1373_ | ~new_n1392_;
  assign new_n3664_ = ~new_n8791_ | ~new_n1770_;
  assign new_n3665_ = ~new_n3664_ | ~new_n3663_ | ~new_n3662_;
  assign new_n3666_ = ~new_n1384_ | ~new_n2346_;
  assign new_n3667_ = ~new_n1383_ | ~new_n8791_;
  assign new_n3668_ = ~new_n2366_ | ~new_n3665_;
  assign new_n3669_ = ~new_n11633_ | ~new_n1366_;
  assign new_n3670_ = ~pi267 | ~po264;
  assign new_n3671_ = ~new_n1375_ | ~new_n1419_;
  assign new_n3672_ = ~new_n1373_ | ~new_n1413_;
  assign new_n3673_ = ~new_n8800_ | ~new_n1770_;
  assign new_n3674_ = ~new_n3672_ | ~new_n3673_ | ~new_n3671_;
  assign new_n3675_ = ~new_n1848_ | ~new_n4025_;
  assign new_n3676_ = ~new_n8800_ | ~new_n4024_;
  assign new_n3677_ = ~new_n2366_ | ~new_n3674_;
  assign new_n3678_ = ~new_n11641_ | ~new_n1366_;
  assign new_n3679_ = ~pi268 | ~po264;
  assign new_n3680_ = ~new_n1375_ | ~new_n1405_;
  assign new_n3681_ = ~new_n1373_ | ~new_n1397_;
  assign new_n3682_ = ~new_n8735_ | ~new_n1770_;
  assign new_n3683_ = ~new_n3682_ | ~new_n3681_ | ~new_n3680_;
  assign new_n3684_ = ~new_n1801_ | ~new_n4025_;
  assign new_n3685_ = ~new_n8735_ | ~new_n4024_;
  assign new_n3686_ = ~new_n2366_ | ~new_n3683_;
  assign new_n3687_ = ~new_n11554_ | ~new_n1366_;
  assign new_n3688_ = ~pi269 | ~po264;
  assign new_n3689_ = ~new_n1375_ | ~new_n1420_;
  assign new_n3690_ = ~new_n1373_ | ~new_n1400_;
  assign new_n3691_ = ~new_n8809_ | ~new_n1770_;
  assign new_n3692_ = ~new_n3691_ | ~new_n3690_ | ~new_n3689_;
  assign new_n3693_ = ~new_n1822_ | ~new_n4025_;
  assign new_n3694_ = ~new_n8809_ | ~new_n4024_;
  assign new_n3695_ = ~new_n2366_ | ~new_n3692_;
  assign new_n3696_ = ~new_n11648_ | ~new_n1366_;
  assign new_n3697_ = ~pi270 | ~po264;
  assign new_n3698_ = ~new_n1375_ | ~new_n1398_;
  assign new_n3699_ = ~new_n1373_ | ~new_n1402_;
  assign new_n3700_ = ~new_n8796_ | ~new_n1770_;
  assign new_n3701_ = ~new_n3699_ | ~new_n3700_ | ~new_n3698_;
  assign new_n3702_ = ~new_n1384_ | ~new_n2351_;
  assign new_n3703_ = ~new_n1383_ | ~new_n8796_;
  assign new_n3704_ = ~new_n2366_ | ~new_n3701_;
  assign new_n3705_ = ~new_n11637_ | ~new_n1366_;
  assign new_n3706_ = ~pi271 | ~po264;
  assign new_n3707_ = ~new_n1375_ | ~new_n1417_;
  assign new_n3708_ = ~new_n1373_ | ~new_n1411_;
  assign new_n3709_ = ~new_n8805_ | ~new_n1770_;
  assign new_n3710_ = ~new_n3708_ | ~new_n3709_ | ~new_n3707_;
  assign new_n3711_ = ~new_n1834_ | ~new_n4025_;
  assign new_n3712_ = ~new_n8805_ | ~new_n4024_;
  assign new_n3713_ = ~new_n2366_ | ~new_n3710_;
  assign new_n3714_ = ~new_n11645_ | ~new_n1366_;
  assign new_n3715_ = ~pi272 | ~po264;
  assign new_n3716_ = ~new_n1375_ | ~new_n1394_;
  assign new_n3717_ = ~new_n1373_ | ~new_n1391_;
  assign new_n3718_ = ~new_n8792_ | ~new_n1770_;
  assign new_n3719_ = ~new_n3717_ | ~new_n3718_ | ~new_n3716_;
  assign new_n3720_ = ~new_n1384_ | ~new_n2347_;
  assign new_n3721_ = ~new_n1383_ | ~new_n8792_;
  assign new_n3722_ = ~new_n2366_ | ~new_n3719_;
  assign new_n3723_ = ~new_n11634_ | ~new_n1366_;
  assign new_n3724_ = ~pi273 | ~po264;
  assign new_n3725_ = ~new_n1375_ | ~new_n1408_;
  assign new_n3726_ = ~new_n1373_ | ~new_n1421_;
  assign new_n3727_ = ~new_n8787_ | ~new_n1770_;
  assign new_n3728_ = ~new_n3727_ | ~new_n3726_ | ~new_n3725_;
  assign new_n3729_ = ~new_n1813_ | ~new_n4025_;
  assign new_n3730_ = ~new_n8787_ | ~new_n4024_;
  assign new_n3731_ = ~new_n2366_ | ~new_n3728_;
  assign new_n3732_ = ~new_n11555_ | ~new_n1366_;
  assign new_n3733_ = ~pi274 | ~po264;
  assign new_n3734_ = ~new_n1789_ | ~new_n1713_;
  assign new_n3735_ = ~new_n1786_ | ~new_n3734_;
  assign new_n3736_ = ~new_n11626_ | ~new_n4073_ | ~new_n1786_;
  assign new_n3737_ = ~new_n1787_ | ~new_n1781_;
  assign new_n3738_ = ~new_n2232_ | ~new_n2342_;
  assign new_n3739_ = ~new_n1708_ | ~new_n1758_;
  assign new_n3740_ = ~new_n1703_ | ~new_n1706_ | ~new_n1701_;
  assign new_n3741_ = ~new_n2372_ | ~new_n1760_;
  assign new_n3742_ = ~new_n3740_ | ~new_n1760_;
  assign new_n3743_ = ~new_n1774_;
  assign new_n3744_ = ~new_n3743_ | ~new_n2342_;
  assign new_n3745_ = ~new_n1819_ | ~new_n3744_;
  assign new_n3746_ = ~new_n1360_ | ~new_n1420_;
  assign new_n3747_ = ~new_n1816_ | ~new_n3744_;
  assign new_n3748_ = ~new_n1360_ | ~new_n1421_;
  assign new_n3749_ = ~new_n1813_ | ~new_n3744_;
  assign new_n3750_ = ~new_n1360_ | ~new_n1407_;
  assign new_n3751_ = ~new_n1810_ | ~new_n3744_;
  assign new_n3752_ = ~new_n1360_ | ~new_n1408_;
  assign new_n3753_ = ~new_n1807_ | ~new_n3744_;
  assign new_n3754_ = ~new_n1360_ | ~new_n1404_;
  assign new_n3755_ = ~new_n1804_ | ~new_n3744_;
  assign new_n3756_ = ~new_n1360_ | ~new_n1397_;
  assign new_n3757_ = ~new_n1801_ | ~new_n3744_;
  assign new_n3758_ = ~new_n1360_ | ~new_n1401_;
  assign new_n3759_ = ~new_n2346_ | ~new_n3744_;
  assign new_n3760_ = ~new_n1360_ | ~new_n1391_;
  assign new_n3761_ = ~new_n2347_ | ~new_n3744_;
  assign new_n3762_ = ~new_n1360_ | ~new_n1390_;
  assign new_n3763_ = ~new_n2348_ | ~new_n3744_;
  assign new_n3764_ = ~new_n1360_ | ~new_n1394_;
  assign new_n3765_ = ~new_n2349_ | ~new_n3744_;
  assign new_n3766_ = ~new_n1360_ | ~new_n1395_;
  assign new_n3767_ = ~new_n2350_ | ~new_n3744_;
  assign new_n3768_ = ~new_n1360_ | ~new_n1402_;
  assign new_n3769_ = ~new_n2351_ | ~new_n3744_;
  assign new_n3770_ = ~new_n1360_ | ~new_n1403_;
  assign new_n3771_ = ~new_n2352_ | ~new_n3744_;
  assign new_n3772_ = ~new_n1360_ | ~new_n1398_;
  assign new_n3773_ = ~new_n2353_ | ~new_n3744_;
  assign new_n3774_ = ~new_n1360_ | ~new_n1412_;
  assign new_n3775_ = ~new_n2354_ | ~new_n3744_;
  assign new_n3776_ = ~new_n1360_ | ~new_n1413_;
  assign new_n3777_ = ~new_n1798_ | ~new_n3744_;
  assign new_n3778_ = ~new_n1360_ | ~new_n1405_;
  assign new_n3779_ = ~new_n1848_ | ~new_n3744_;
  assign new_n3780_ = ~new_n1360_ | ~new_n1418_;
  assign new_n3781_ = ~new_n1846_ | ~new_n3744_;
  assign new_n3782_ = ~new_n1360_ | ~new_n1419_;
  assign new_n3783_ = ~new_n1843_ | ~new_n3744_;
  assign new_n3784_ = ~new_n1360_ | ~new_n1406_;
  assign new_n3785_ = ~new_n1840_ | ~new_n3744_;
  assign new_n3786_ = ~new_n1360_ | ~new_n1410_;
  assign new_n3787_ = ~new_n1837_ | ~new_n3744_;
  assign new_n3788_ = ~new_n1360_ | ~new_n1411_;
  assign new_n3789_ = ~new_n1834_ | ~new_n3744_;
  assign new_n3790_ = ~new_n1360_ | ~new_n1416_;
  assign new_n3791_ = ~new_n1831_ | ~new_n3744_;
  assign new_n3792_ = ~new_n1360_ | ~new_n1417_;
  assign new_n3793_ = ~new_n1828_ | ~new_n3744_;
  assign new_n3794_ = ~new_n1360_ | ~new_n1409_;
  assign new_n3795_ = ~new_n1825_ | ~new_n3744_;
  assign new_n3796_ = ~new_n1360_ | ~new_n1400_;
  assign new_n3797_ = ~new_n1822_ | ~new_n3744_;
  assign new_n3798_ = ~new_n1360_ | ~new_n1399_;
  assign new_n3799_ = ~new_n1795_ | ~new_n3744_;
  assign new_n3800_ = ~new_n1360_ | ~new_n1415_;
  assign new_n3801_ = ~new_n1790_ | ~new_n3744_;
  assign new_n3802_ = ~new_n1360_ | ~new_n1414_;
  assign new_n3803_ = ~new_n2474_ | ~pi129;
  assign new_n3804_ = ~new_n1360_ | ~new_n1819_;
  assign new_n3805_ = ~new_n1774_ | ~new_n1420_;
  assign new_n3806_ = ~new_n1360_ | ~new_n1816_;
  assign new_n3807_ = ~new_n1774_ | ~new_n1421_;
  assign new_n3808_ = ~new_n1360_ | ~new_n1813_;
  assign new_n3809_ = ~new_n1774_ | ~new_n1407_;
  assign new_n3810_ = ~new_n1360_ | ~new_n1810_;
  assign new_n3811_ = ~new_n1774_ | ~new_n1408_;
  assign new_n3812_ = ~new_n1360_ | ~new_n1807_;
  assign new_n3813_ = ~new_n1774_ | ~new_n1404_;
  assign new_n3814_ = ~new_n1360_ | ~new_n1804_;
  assign new_n3815_ = ~new_n1774_ | ~new_n1397_;
  assign new_n3816_ = ~new_n1360_ | ~new_n1801_;
  assign new_n3817_ = ~new_n1774_ | ~new_n1401_;
  assign new_n3818_ = ~new_n1360_ | ~new_n2346_;
  assign new_n3819_ = ~new_n1774_ | ~new_n1391_;
  assign new_n3820_ = ~new_n1360_ | ~new_n2347_;
  assign new_n3821_ = ~new_n1774_ | ~new_n1390_;
  assign new_n3822_ = ~new_n1360_ | ~new_n2348_;
  assign new_n3823_ = ~new_n1774_ | ~new_n1394_;
  assign new_n3824_ = ~new_n1360_ | ~new_n2349_;
  assign new_n3825_ = ~new_n1774_ | ~new_n1395_;
  assign new_n3826_ = ~new_n1360_ | ~new_n2350_;
  assign new_n3827_ = ~new_n1774_ | ~new_n1402_;
  assign new_n3828_ = ~new_n1360_ | ~new_n2351_;
  assign new_n3829_ = ~new_n1774_ | ~new_n1403_;
  assign new_n3830_ = ~new_n1360_ | ~new_n2352_;
  assign new_n3831_ = ~new_n1774_ | ~new_n1398_;
  assign new_n3832_ = ~new_n1360_ | ~new_n2353_;
  assign new_n3833_ = ~new_n1774_ | ~new_n1412_;
  assign new_n3834_ = ~new_n1360_ | ~new_n2354_;
  assign new_n3835_ = ~new_n1774_ | ~new_n1413_;
  assign new_n3836_ = ~new_n1360_ | ~new_n1798_;
  assign new_n3837_ = ~new_n1774_ | ~new_n1405_;
  assign new_n3838_ = ~new_n1360_ | ~new_n1848_;
  assign new_n3839_ = ~new_n1774_ | ~new_n1418_;
  assign new_n3840_ = ~new_n1360_ | ~new_n1846_;
  assign new_n3841_ = ~new_n1774_ | ~new_n1419_;
  assign new_n3842_ = ~new_n1360_ | ~new_n1843_;
  assign new_n3843_ = ~new_n1774_ | ~new_n1406_;
  assign new_n3844_ = ~new_n1360_ | ~new_n1840_;
  assign new_n3845_ = ~new_n1774_ | ~new_n1410_;
  assign new_n3846_ = ~new_n1360_ | ~new_n1837_;
  assign new_n3847_ = ~new_n1774_ | ~new_n1411_;
  assign new_n3848_ = ~new_n1360_ | ~new_n1834_;
  assign new_n3849_ = ~new_n1774_ | ~new_n1416_;
  assign new_n3850_ = ~new_n1360_ | ~new_n1831_;
  assign new_n3851_ = ~new_n1774_ | ~new_n1417_;
  assign new_n3852_ = ~new_n1360_ | ~new_n1828_;
  assign new_n3853_ = ~new_n1774_ | ~new_n1409_;
  assign new_n3854_ = ~new_n1360_ | ~new_n1825_;
  assign new_n3855_ = ~new_n1774_ | ~new_n1400_;
  assign new_n3856_ = ~new_n1360_ | ~new_n1822_;
  assign new_n3857_ = ~new_n1774_ | ~new_n1399_;
  assign new_n3858_ = ~new_n1360_ | ~new_n1795_;
  assign new_n3859_ = ~new_n1774_ | ~new_n1415_;
  assign new_n3860_ = ~new_n1360_ | ~new_n1790_;
  assign new_n3861_ = ~new_n1774_ | ~new_n1414_;
  assign new_n3862_ = ~new_n2474_ | ~new_n1788_;
  assign new_n3863_ = ~new_n1767_ | ~new_n1765_;
  assign new_n3864_ = ~new_n2325_ | ~new_n1819_;
  assign new_n3865_ = ~new_n1926_ | ~new_n3863_;
  assign new_n3866_ = ~new_n2325_ | ~new_n1816_;
  assign new_n3867_ = ~new_n1927_ | ~new_n3863_;
  assign new_n3868_ = ~new_n2325_ | ~new_n1813_;
  assign new_n3869_ = ~new_n1928_ | ~new_n3863_;
  assign new_n3870_ = ~new_n2325_ | ~new_n1810_;
  assign new_n3871_ = ~new_n1929_ | ~new_n3863_;
  assign new_n3872_ = ~new_n2325_ | ~new_n1807_;
  assign new_n3873_ = ~new_n1930_ | ~new_n3863_;
  assign new_n3874_ = ~new_n2325_ | ~new_n1804_;
  assign new_n3875_ = ~new_n1931_ | ~new_n3863_;
  assign new_n3876_ = ~new_n1933_ | ~new_n3863_;
  assign new_n3877_ = ~new_n2355_ | ~new_n2325_;
  assign new_n3878_ = ~new_n1934_ | ~new_n3863_;
  assign new_n3879_ = ~new_n2356_ | ~new_n2325_;
  assign new_n3880_ = ~new_n2325_ | ~new_n1801_;
  assign new_n3881_ = ~new_n1932_ | ~new_n3863_;
  assign new_n3882_ = ~new_n1936_ | ~new_n3863_;
  assign new_n3883_ = ~new_n2357_ | ~new_n2325_;
  assign new_n3884_ = ~new_n1937_ | ~new_n3863_;
  assign new_n3885_ = ~new_n2346_ | ~new_n2325_;
  assign new_n3886_ = ~new_n1938_ | ~new_n3863_;
  assign new_n3887_ = ~new_n2347_ | ~new_n2325_;
  assign new_n3888_ = ~new_n1939_ | ~new_n3863_;
  assign new_n3889_ = ~new_n2348_ | ~new_n2325_;
  assign new_n3890_ = ~new_n1940_ | ~new_n3863_;
  assign new_n3891_ = ~new_n2349_ | ~new_n2325_;
  assign new_n3892_ = ~new_n1941_ | ~new_n3863_;
  assign new_n3893_ = ~new_n2350_ | ~new_n2325_;
  assign new_n3894_ = ~new_n1942_ | ~new_n3863_;
  assign new_n3895_ = ~new_n2351_ | ~new_n2325_;
  assign new_n3896_ = ~new_n1943_ | ~new_n3863_;
  assign new_n3897_ = ~new_n2352_ | ~new_n2325_;
  assign new_n3898_ = ~new_n1944_ | ~new_n3863_;
  assign new_n3899_ = ~new_n2353_ | ~new_n2325_;
  assign new_n3900_ = ~new_n1945_ | ~new_n3863_;
  assign new_n3901_ = ~new_n2354_ | ~new_n2325_;
  assign new_n3902_ = ~new_n2325_ | ~new_n1798_;
  assign new_n3903_ = ~new_n1935_ | ~new_n3863_;
  assign new_n3904_ = ~new_n2325_ | ~new_n1848_;
  assign new_n3905_ = ~new_n1947_ | ~new_n3863_;
  assign new_n3906_ = ~new_n2325_ | ~new_n1846_;
  assign new_n3907_ = ~new_n1948_ | ~new_n3863_;
  assign new_n3908_ = ~new_n2325_ | ~new_n1843_;
  assign new_n3909_ = ~new_n1949_ | ~new_n3863_;
  assign new_n3910_ = ~new_n2325_ | ~new_n1840_;
  assign new_n3911_ = ~new_n1950_ | ~new_n3863_;
  assign new_n3912_ = ~new_n2325_ | ~new_n1837_;
  assign new_n3913_ = ~new_n1951_ | ~new_n3863_;
  assign new_n3914_ = ~new_n2325_ | ~new_n1834_;
  assign new_n3915_ = ~new_n1952_ | ~new_n3863_;
  assign new_n3916_ = ~new_n2325_ | ~new_n1831_;
  assign new_n3917_ = ~new_n1953_ | ~new_n3863_;
  assign new_n3918_ = ~new_n2325_ | ~new_n1828_;
  assign new_n3919_ = ~new_n1954_ | ~new_n3863_;
  assign new_n3920_ = ~new_n2325_ | ~new_n1825_;
  assign new_n3921_ = ~new_n1955_ | ~new_n3863_;
  assign new_n3922_ = ~new_n2325_ | ~new_n1822_;
  assign new_n3923_ = ~new_n1956_ | ~new_n3863_;
  assign new_n3924_ = ~new_n2325_ | ~new_n1795_;
  assign new_n3925_ = ~new_n1946_ | ~new_n3863_;
  assign new_n3926_ = ~new_n2325_ | ~new_n1790_;
  assign new_n3927_ = ~new_n1957_ | ~new_n3863_;
  assign new_n3928_ = ~new_n1819_ | ~new_n3863_;
  assign new_n3929_ = ~new_n2325_ | ~new_n1926_;
  assign new_n3930_ = ~new_n4042_ | ~new_n1421_;
  assign new_n3931_ = ~new_n1816_ | ~new_n3863_;
  assign new_n3932_ = ~new_n2325_ | ~new_n1927_;
  assign new_n3933_ = ~new_n4042_ | ~new_n1407_;
  assign new_n3934_ = ~new_n1813_ | ~new_n3863_;
  assign new_n3935_ = ~new_n2325_ | ~new_n1928_;
  assign new_n3936_ = ~new_n4042_ | ~new_n1408_;
  assign new_n3937_ = ~new_n1810_ | ~new_n3863_;
  assign new_n3938_ = ~new_n2325_ | ~new_n1929_;
  assign new_n3939_ = ~new_n4042_ | ~new_n1404_;
  assign new_n3940_ = ~new_n1807_ | ~new_n3863_;
  assign new_n3941_ = ~new_n2325_ | ~new_n1930_;
  assign new_n3942_ = ~new_n4042_ | ~new_n1397_;
  assign new_n3943_ = ~new_n1804_ | ~new_n3863_;
  assign new_n3944_ = ~new_n2325_ | ~new_n1931_;
  assign new_n3945_ = ~new_n4042_ | ~new_n1401_;
  assign new_n3946_ = ~new_n2355_ | ~new_n3863_;
  assign new_n3947_ = ~new_n2325_ | ~new_n1933_;
  assign new_n3948_ = ~new_n2356_ | ~new_n3863_;
  assign new_n3949_ = ~new_n2325_ | ~new_n1934_;
  assign new_n3950_ = ~new_n1801_ | ~new_n3863_;
  assign new_n3951_ = ~new_n2325_ | ~new_n1932_;
  assign new_n3952_ = ~new_n4042_ | ~new_n1405_;
  assign new_n3953_ = ~new_n2357_ | ~new_n3863_;
  assign new_n3954_ = ~new_n2325_ | ~new_n1936_;
  assign new_n3955_ = ~new_n4042_ | ~new_n1391_;
  assign new_n3956_ = ~new_n2346_ | ~new_n3863_;
  assign new_n3957_ = ~new_n2325_ | ~new_n1937_;
  assign new_n3958_ = ~new_n4042_ | ~new_n1390_;
  assign new_n3959_ = ~new_n2347_ | ~new_n3863_;
  assign new_n3960_ = ~new_n2325_ | ~new_n1938_;
  assign new_n3961_ = ~new_n4042_ | ~new_n1394_;
  assign new_n3962_ = ~new_n2348_ | ~new_n3863_;
  assign new_n3963_ = ~new_n2325_ | ~new_n1939_;
  assign new_n3964_ = ~new_n4042_ | ~new_n1395_;
  assign new_n3965_ = ~new_n2349_ | ~new_n3863_;
  assign new_n3966_ = ~new_n2325_ | ~new_n1940_;
  assign new_n3967_ = ~new_n4042_ | ~new_n1402_;
  assign new_n3968_ = ~new_n2350_ | ~new_n3863_;
  assign new_n3969_ = ~new_n2325_ | ~new_n1941_;
  assign new_n3970_ = ~new_n4042_ | ~new_n1403_;
  assign new_n3971_ = ~new_n2351_ | ~new_n3863_;
  assign new_n3972_ = ~new_n2325_ | ~new_n1942_;
  assign new_n3973_ = ~new_n4042_ | ~new_n1398_;
  assign new_n3974_ = ~new_n2352_ | ~new_n3863_;
  assign new_n3975_ = ~new_n2325_ | ~new_n1943_;
  assign new_n3976_ = ~new_n4042_ | ~new_n1412_;
  assign new_n3977_ = ~new_n2353_ | ~new_n3863_;
  assign new_n3978_ = ~new_n2325_ | ~new_n1944_;
  assign new_n3979_ = ~new_n4042_ | ~new_n1413_;
  assign new_n3980_ = ~new_n2354_ | ~new_n3863_;
  assign new_n3981_ = ~new_n2325_ | ~new_n1945_;
  assign new_n3982_ = ~new_n4042_ | ~new_n1418_;
  assign new_n3983_ = ~new_n1798_ | ~new_n3863_;
  assign new_n3984_ = ~new_n2325_ | ~new_n1935_;
  assign new_n3985_ = ~new_n4042_ | ~new_n1415_;
  assign new_n3986_ = ~new_n1848_ | ~new_n3863_;
  assign new_n3987_ = ~new_n2325_ | ~new_n1947_;
  assign new_n3988_ = ~new_n4042_ | ~new_n1419_;
  assign new_n3989_ = ~new_n1846_ | ~new_n3863_;
  assign new_n3990_ = ~new_n2325_ | ~new_n1948_;
  assign new_n3991_ = ~new_n4042_ | ~new_n1406_;
  assign new_n3992_ = ~new_n1843_ | ~new_n3863_;
  assign new_n3993_ = ~new_n2325_ | ~new_n1949_;
  assign new_n3994_ = ~new_n4042_ | ~new_n1410_;
  assign new_n3995_ = ~new_n1840_ | ~new_n3863_;
  assign new_n3996_ = ~new_n2325_ | ~new_n1950_;
  assign new_n3997_ = ~new_n4042_ | ~new_n1411_;
  assign new_n3998_ = ~new_n1837_ | ~new_n3863_;
  assign new_n3999_ = ~new_n2325_ | ~new_n1951_;
  assign new_n4000_ = ~new_n4042_ | ~new_n1416_;
  assign new_n4001_ = ~new_n1834_ | ~new_n3863_;
  assign new_n4002_ = ~new_n2325_ | ~new_n1952_;
  assign new_n4003_ = ~new_n4042_ | ~new_n1417_;
  assign new_n4004_ = ~new_n1831_ | ~new_n3863_;
  assign new_n4005_ = ~new_n2325_ | ~new_n1953_;
  assign new_n4006_ = ~new_n4042_ | ~new_n1409_;
  assign new_n4007_ = ~new_n1828_ | ~new_n3863_;
  assign new_n4008_ = ~new_n2325_ | ~new_n1954_;
  assign new_n4009_ = ~new_n4042_ | ~new_n1400_;
  assign new_n4010_ = ~new_n1825_ | ~new_n3863_;
  assign new_n4011_ = ~new_n2325_ | ~new_n1955_;
  assign new_n4012_ = ~new_n4042_ | ~new_n1399_;
  assign new_n4013_ = ~new_n1822_ | ~new_n3863_;
  assign new_n4014_ = ~new_n2325_ | ~new_n1956_;
  assign new_n4015_ = ~new_n4042_ | ~new_n1420_;
  assign new_n4016_ = ~new_n1795_ | ~new_n3863_;
  assign new_n4017_ = ~new_n2325_ | ~new_n1946_;
  assign new_n4018_ = ~new_n4042_ | ~new_n1414_;
  assign new_n4019_ = ~new_n1790_ | ~new_n3863_;
  assign new_n4020_ = ~new_n2325_ | ~new_n1957_;
  assign new_n4021_ = ~new_n3462_ | ~po264;
  assign new_n4022_ = ~new_n2369_ | ~new_n1770_;
  assign new_n4023_ = ~new_n2344_ | ~new_n2369_;
  assign new_n4024_ = ~new_n4022_ | ~new_n2367_;
  assign new_n4025_ = ~new_n4023_ | ~new_n2368_;
  assign new_n4026_ = ~new_n1768_ | ~new_n1778_ | ~new_n1387_;
  assign new_n4027_ = ~new_n4031_ | ~new_n4037_;
  assign new_n4028_ = ~new_n13093_ | ~new_n2326_ | ~new_n2359_ | ~new_n1781_;
  assign new_n4029_ = ~pi057 | ~new_n2283_;
  assign new_n4030_ = ~pi064 | ~new_n9201_;
  assign new_n4031_ = ~new_n1775_;
  assign new_n4032_ = ~pi058 | ~new_n2283_;
  assign new_n4033_ = ~pi064 | ~new_n9354_;
  assign new_n4034_ = ~new_n1776_;
  assign new_n4035_ = ~pi059 | ~new_n2283_;
  assign new_n4036_ = ~pi064 | ~new_n9202_;
  assign new_n4037_ = ~new_n1777_;
  assign new_n4038_ = ~new_n1389_ | ~new_n1697_;
  assign new_n4039_ = ~pi245 | ~new_n2375_ | ~new_n4031_;
  assign new_n4040_ = ~pi056 | ~new_n2283_;
  assign new_n4041_ = ~pi064 | ~new_n9200_;
  assign new_n4042_ = ~new_n1778_;
  assign new_n4043_ = ~pi065 | ~new_n2284_;
  assign new_n4044_ = ~new_n2364_ | ~new_n2475_;
  assign new_n4045_ = ~pi066 | ~new_n2284_;
  assign new_n4046_ = ~new_n2364_ | ~new_n2476_;
  assign new_n4047_ = ~pi055 | ~new_n2283_;
  assign new_n4048_ = ~pi064 | ~new_n9199_;
  assign new_n4049_ = ~new_n1783_;
  assign new_n4050_ = ~pi052 | ~new_n2283_;
  assign new_n4051_ = ~pi064 | ~new_n9197_;
  assign new_n4052_ = ~new_n1782_;
  assign new_n4053_ = ~pi053 | ~new_n2283_;
  assign new_n4054_ = ~pi064 | ~new_n9198_;
  assign new_n4055_ = ~new_n1781_;
  assign new_n4056_ = ~pi054 | ~new_n2283_;
  assign new_n4057_ = ~pi064 | ~new_n9357_;
  assign new_n4058_ = ~new_n1787_;
  assign new_n4059_ = ~pi063 | ~new_n2283_;
  assign new_n4060_ = ~pi064 | ~new_n9349_;
  assign new_n4061_ = ~new_n1784_;
  assign new_n4062_ = ~pi062 | ~new_n2283_;
  assign new_n4063_ = ~pi064 | ~new_n9204_;
  assign new_n4064_ = ~new_n1785_;
  assign new_n4065_ = ~pi061 | ~new_n2283_;
  assign new_n4066_ = ~pi064 | ~new_n9203_;
  assign new_n4067_ = ~new_n1786_;
  assign new_n4068_ = ~pi033 | ~new_n2283_;
  assign new_n4069_ = ~pi064 | ~pi033;
  assign new_n4070_ = ~new_n1788_;
  assign new_n4071_ = ~pi060 | ~new_n2283_;
  assign new_n4072_ = ~pi064 | ~new_n9226_;
  assign new_n4073_ = ~new_n1789_;
  assign new_n4074_ = ~new_n1102_ | ~new_n2285_;
  assign new_n4075_ = ~new_n2343_ | ~new_n1788_;
  assign new_n4076_ = ~new_n1790_;
  assign new_n4077_ = ~new_n1783_ | ~new_n4058_;
  assign new_n4078_ = ~new_n4049_ | ~new_n2507_;
  assign new_n4079_ = ~pi066 | ~new_n2473_;
  assign new_n4080_ = ~new_n2476_ | ~new_n1698_;
  assign new_n4081_ = ~new_n1792_;
  assign new_n4082_ = ~new_n4027_ | ~new_n1698_;
  assign new_n4083_ = ~pi065 | ~new_n2473_;
  assign new_n4084_ = ~new_n1791_;
  assign new_n4085_ = ~pi097 | ~new_n2286_;
  assign new_n4086_ = ~new_n2363_ | ~new_n2527_;
  assign new_n4087_ = ~pi034 | ~new_n2283_;
  assign new_n4088_ = ~pi064 | ~new_n9224_;
  assign new_n4089_ = ~new_n1091_ | ~new_n2285_;
  assign new_n4090_ = ~new_n1794_ | ~new_n2343_;
  assign new_n4091_ = ~new_n1795_;
  assign new_n4092_ = ~pi098 | ~new_n2286_;
  assign new_n4093_ = ~new_n2363_ | ~new_n2551_;
  assign new_n4094_ = ~pi035 | ~new_n2283_;
  assign new_n4095_ = ~pi064 | ~new_n9205_;
  assign new_n4096_ = ~new_n1080_ | ~new_n2285_;
  assign new_n4097_ = ~new_n1797_ | ~new_n2343_;
  assign new_n4098_ = ~new_n1798_;
  assign new_n4099_ = ~pi099 | ~new_n2286_;
  assign new_n4100_ = ~new_n2363_ | ~new_n2570_;
  assign new_n4101_ = ~pi036 | ~new_n2283_;
  assign new_n4102_ = ~pi064 | ~new_n9206_;
  assign new_n4103_ = ~new_n1077_ | ~new_n2285_;
  assign new_n4104_ = ~new_n1800_ | ~new_n2343_;
  assign new_n4105_ = ~new_n1801_;
  assign new_n4106_ = ~pi100 | ~new_n2286_;
  assign new_n4107_ = ~new_n2363_ | ~new_n2589_;
  assign new_n4108_ = ~pi037 | ~new_n2283_;
  assign new_n4109_ = ~pi064 | ~new_n9207_;
  assign new_n4110_ = ~new_n1076_ | ~new_n2285_;
  assign new_n4111_ = ~new_n1803_ | ~new_n2343_;
  assign new_n4112_ = ~new_n1804_;
  assign new_n4113_ = ~pi101 | ~new_n2286_;
  assign new_n4114_ = ~new_n2363_ | ~new_n2608_;
  assign new_n4115_ = ~pi038 | ~new_n2283_;
  assign new_n4116_ = ~pi064 | ~new_n9346_;
  assign new_n4117_ = ~new_n1075_ | ~new_n2285_;
  assign new_n4118_ = ~new_n1806_ | ~new_n2343_;
  assign new_n4119_ = ~new_n1807_;
  assign new_n4120_ = ~pi102 | ~new_n2286_;
  assign new_n4121_ = ~new_n2363_ | ~new_n2627_;
  assign new_n4122_ = ~pi039 | ~new_n2283_;
  assign new_n4123_ = ~pi064 | ~new_n9208_;
  assign new_n4124_ = ~new_n1074_ | ~new_n2285_;
  assign new_n4125_ = ~new_n1809_ | ~new_n2343_;
  assign new_n4126_ = ~new_n1810_;
  assign new_n4127_ = ~pi103 | ~new_n2286_;
  assign new_n4128_ = ~new_n2363_ | ~new_n2646_;
  assign new_n4129_ = ~pi040 | ~new_n2283_;
  assign new_n4130_ = ~pi064 | ~new_n9209_;
  assign new_n4131_ = ~new_n1073_ | ~new_n2285_;
  assign new_n4132_ = ~new_n1812_ | ~new_n2343_;
  assign new_n4133_ = ~new_n1813_;
  assign new_n4134_ = ~pi104 | ~new_n2286_;
  assign new_n4135_ = ~new_n2363_ | ~new_n2665_;
  assign new_n4136_ = ~pi041 | ~new_n2283_;
  assign new_n4137_ = ~pi064 | ~new_n9210_;
  assign new_n4138_ = ~new_n1072_ | ~new_n2285_;
  assign new_n4139_ = ~new_n1815_ | ~new_n2343_;
  assign new_n4140_ = ~new_n1816_;
  assign new_n4141_ = ~pi105 | ~new_n2286_;
  assign new_n4142_ = ~new_n2363_ | ~new_n2684_;
  assign new_n4143_ = ~pi042 | ~new_n2283_;
  assign new_n4144_ = ~pi064 | ~new_n9344_;
  assign new_n4145_ = ~new_n1071_ | ~new_n2285_;
  assign new_n4146_ = ~new_n1818_ | ~new_n2343_;
  assign new_n4147_ = ~new_n1819_;
  assign new_n4148_ = ~pi106 | ~new_n2286_;
  assign new_n4149_ = ~new_n2363_ | ~new_n2703_;
  assign new_n4150_ = ~pi043 | ~new_n2283_;
  assign new_n4151_ = ~pi064 | ~new_n9190_;
  assign new_n4152_ = ~new_n1101_ | ~new_n2285_;
  assign new_n4153_ = ~new_n1821_ | ~new_n2343_;
  assign new_n4154_ = ~new_n1822_;
  assign new_n4155_ = ~pi107 | ~new_n2286_;
  assign new_n4156_ = ~new_n2363_ | ~new_n2722_;
  assign new_n4157_ = ~pi044 | ~new_n2283_;
  assign new_n4158_ = ~pi064 | ~new_n9191_;
  assign new_n4159_ = ~new_n1100_ | ~new_n2285_;
  assign new_n4160_ = ~new_n1824_ | ~new_n2343_;
  assign new_n4161_ = ~new_n1825_;
  assign new_n4162_ = ~pi108 | ~new_n2286_;
  assign new_n4163_ = ~new_n2363_ | ~new_n2741_;
  assign new_n4164_ = ~pi045 | ~new_n2283_;
  assign new_n4165_ = ~pi064 | ~new_n9192_;
  assign new_n4166_ = ~new_n1099_ | ~new_n2285_;
  assign new_n4167_ = ~new_n1827_ | ~new_n2343_;
  assign new_n4168_ = ~new_n1828_;
  assign new_n4169_ = ~pi109 | ~new_n2286_;
  assign new_n4170_ = ~new_n2363_ | ~new_n2760_;
  assign new_n4171_ = ~pi046 | ~new_n2283_;
  assign new_n4172_ = ~pi064 | ~new_n9363_;
  assign new_n4173_ = ~new_n1098_ | ~new_n2285_;
  assign new_n4174_ = ~new_n1830_ | ~new_n2343_;
  assign new_n4175_ = ~new_n1831_;
  assign new_n4176_ = ~pi110 | ~new_n2286_;
  assign new_n4177_ = ~new_n2363_ | ~new_n2779_;
  assign new_n4178_ = ~pi047 | ~new_n2283_;
  assign new_n4179_ = ~pi064 | ~new_n9193_;
  assign new_n4180_ = ~new_n1097_ | ~new_n2285_;
  assign new_n4181_ = ~new_n1833_ | ~new_n2343_;
  assign new_n4182_ = ~new_n1834_;
  assign new_n4183_ = ~pi111 | ~new_n2286_;
  assign new_n4184_ = ~new_n2363_ | ~new_n2798_;
  assign new_n4185_ = ~pi048 | ~new_n2283_;
  assign new_n4186_ = ~pi064 | ~new_n9194_;
  assign new_n4187_ = ~new_n1096_ | ~new_n2285_;
  assign new_n4188_ = ~new_n1836_ | ~new_n2343_;
  assign new_n4189_ = ~new_n1837_;
  assign new_n4190_ = ~pi112 | ~new_n2286_;
  assign new_n4191_ = ~new_n2363_ | ~new_n2817_;
  assign new_n4192_ = ~pi049 | ~new_n2283_;
  assign new_n4193_ = ~pi064 | ~new_n9195_;
  assign new_n4194_ = ~new_n1095_ | ~new_n2285_;
  assign new_n4195_ = ~new_n1839_ | ~new_n2343_;
  assign new_n4196_ = ~new_n1840_;
  assign new_n4197_ = ~pi113 | ~new_n2286_;
  assign new_n4198_ = ~new_n2363_ | ~new_n2836_;
  assign new_n4199_ = ~pi050 | ~new_n2283_;
  assign new_n4200_ = ~pi064 | ~new_n9361_;
  assign new_n4201_ = ~new_n1094_ | ~new_n2285_;
  assign new_n4202_ = ~new_n1842_ | ~new_n2343_;
  assign new_n4203_ = ~new_n1843_;
  assign new_n4204_ = ~pi114 | ~new_n2286_;
  assign new_n4205_ = ~new_n2363_ | ~new_n2855_;
  assign new_n4206_ = ~pi051 | ~new_n2283_;
  assign new_n4207_ = ~pi064 | ~new_n9196_;
  assign new_n4208_ = ~new_n1093_ | ~new_n2285_;
  assign new_n4209_ = ~new_n1845_ | ~new_n2343_;
  assign new_n4210_ = ~new_n1846_;
  assign new_n4211_ = ~pi115 | ~new_n2286_;
  assign new_n4212_ = ~new_n2363_ | ~new_n2874_;
  assign new_n4213_ = ~new_n1092_ | ~new_n2285_;
  assign new_n4214_ = ~new_n2343_ | ~new_n1782_;
  assign new_n4215_ = ~new_n1848_;
  assign new_n4216_ = ~pi116 | ~new_n2286_;
  assign new_n4217_ = ~new_n2363_ | ~new_n2893_;
  assign new_n4218_ = ~pi117 | ~new_n2286_;
  assign new_n4219_ = ~new_n2363_ | ~new_n2912_;
  assign new_n4220_ = ~pi118 | ~new_n2286_;
  assign new_n4221_ = ~new_n2363_ | ~new_n2931_;
  assign new_n4222_ = ~pi119 | ~new_n2286_;
  assign new_n4223_ = ~new_n2363_ | ~new_n2950_;
  assign new_n4224_ = ~pi120 | ~new_n2286_;
  assign new_n4225_ = ~new_n2363_ | ~new_n2969_;
  assign new_n4226_ = ~pi121 | ~new_n2286_;
  assign new_n4227_ = ~new_n2363_ | ~new_n2988_;
  assign new_n4228_ = ~pi122 | ~new_n2286_;
  assign new_n4229_ = ~new_n2363_ | ~new_n3007_;
  assign new_n4230_ = ~pi123 | ~new_n2286_;
  assign new_n4231_ = ~new_n2363_ | ~new_n3026_;
  assign new_n4232_ = ~pi124 | ~new_n2286_;
  assign new_n4233_ = ~new_n2363_ | ~new_n3045_;
  assign new_n4234_ = ~pi125 | ~new_n2286_;
  assign new_n4235_ = ~new_n2363_ | ~new_n3064_;
  assign new_n4236_ = ~pi126 | ~new_n2286_;
  assign new_n4237_ = ~new_n2363_ | ~new_n3084_;
  assign new_n4238_ = ~pi127 | ~new_n2286_;
  assign new_n4239_ = ~new_n2363_ | ~new_n3091_;
  assign new_n4240_ = ~pi128 | ~new_n2286_;
  assign new_n4241_ = ~new_n2363_ | ~new_n3094_;
  assign new_n4242_ = ~pi129 | ~new_n2287_;
  assign new_n4243_ = ~new_n2362_ | ~new_n2527_;
  assign new_n4244_ = ~pi130 | ~new_n2287_;
  assign new_n4245_ = ~new_n2362_ | ~new_n2551_;
  assign new_n4246_ = ~pi131 | ~new_n2287_;
  assign new_n4247_ = ~new_n2362_ | ~new_n2570_;
  assign new_n4248_ = ~pi132 | ~new_n2287_;
  assign new_n4249_ = ~new_n2362_ | ~new_n2589_;
  assign new_n4250_ = ~pi133 | ~new_n2287_;
  assign new_n4251_ = ~new_n2362_ | ~new_n2608_;
  assign new_n4252_ = ~pi134 | ~new_n2287_;
  assign new_n4253_ = ~new_n2362_ | ~new_n2627_;
  assign new_n4254_ = ~pi135 | ~new_n2287_;
  assign new_n4255_ = ~new_n2362_ | ~new_n2646_;
  assign new_n4256_ = ~pi136 | ~new_n2287_;
  assign new_n4257_ = ~new_n2362_ | ~new_n2665_;
  assign new_n4258_ = ~pi137 | ~new_n2287_;
  assign new_n4259_ = ~new_n2362_ | ~new_n2684_;
  assign new_n4260_ = ~pi138 | ~new_n2287_;
  assign new_n4261_ = ~new_n2362_ | ~new_n2703_;
  assign new_n4262_ = ~pi139 | ~new_n2287_;
  assign new_n4263_ = ~new_n2362_ | ~new_n2722_;
  assign new_n4264_ = ~pi140 | ~new_n2287_;
  assign new_n4265_ = ~new_n2362_ | ~new_n2741_;
  assign new_n4266_ = ~pi141 | ~new_n2287_;
  assign new_n4267_ = ~new_n2362_ | ~new_n2760_;
  assign new_n4268_ = ~pi142 | ~new_n2287_;
  assign new_n4269_ = ~new_n2362_ | ~new_n2779_;
  assign new_n4270_ = ~pi143 | ~new_n2287_;
  assign new_n4271_ = ~new_n2362_ | ~new_n2798_;
  assign new_n4272_ = ~pi144 | ~new_n2287_;
  assign new_n4273_ = ~new_n2362_ | ~new_n2817_;
  assign new_n4274_ = ~pi145 | ~new_n2287_;
  assign new_n4275_ = ~new_n2362_ | ~new_n2836_;
  assign new_n4276_ = ~pi146 | ~new_n2287_;
  assign new_n4277_ = ~new_n2362_ | ~new_n2855_;
  assign new_n4278_ = ~pi147 | ~new_n2287_;
  assign new_n4279_ = ~new_n2362_ | ~new_n2874_;
  assign new_n4280_ = ~pi148 | ~new_n2287_;
  assign new_n4281_ = ~new_n2362_ | ~new_n2893_;
  assign new_n4282_ = ~pi149 | ~new_n2287_;
  assign new_n4283_ = ~new_n2362_ | ~new_n2912_;
  assign new_n4284_ = ~pi150 | ~new_n2287_;
  assign new_n4285_ = ~new_n2362_ | ~new_n2931_;
  assign new_n4286_ = ~pi151 | ~new_n2287_;
  assign new_n4287_ = ~new_n2362_ | ~new_n2950_;
  assign new_n4288_ = ~pi152 | ~new_n2287_;
  assign new_n4289_ = ~new_n2362_ | ~new_n2969_;
  assign new_n4290_ = ~pi153 | ~new_n2287_;
  assign new_n4291_ = ~new_n2362_ | ~new_n2988_;
  assign new_n4292_ = ~pi154 | ~new_n2287_;
  assign new_n4293_ = ~new_n2362_ | ~new_n3007_;
  assign new_n4294_ = ~pi155 | ~new_n2287_;
  assign new_n4295_ = ~new_n2362_ | ~new_n3026_;
  assign new_n4296_ = ~pi156 | ~new_n2287_;
  assign new_n4297_ = ~new_n2362_ | ~new_n3045_;
  assign new_n4298_ = ~pi157 | ~new_n2287_;
  assign new_n4299_ = ~new_n2362_ | ~new_n3064_;
  assign new_n4300_ = ~pi158 | ~new_n2287_;
  assign new_n4301_ = ~new_n2362_ | ~new_n3084_;
  assign new_n4302_ = ~pi159 | ~new_n2287_;
  assign new_n4303_ = ~new_n2362_ | ~new_n3091_;
  assign new_n4304_ = ~pi160 | ~new_n2287_;
  assign new_n4305_ = ~new_n2362_ | ~new_n3094_;
  assign new_n4306_ = ~pi161 | ~new_n1756_;
  assign new_n4307_ = ~new_n2361_ | ~new_n1712_;
  assign new_n4308_ = ~pi162 | ~new_n1756_;
  assign new_n4309_ = ~new_n2361_ | ~new_n1714_;
  assign new_n4310_ = ~pi163 | ~new_n1756_;
  assign new_n4311_ = ~new_n2361_ | ~new_n1715_;
  assign new_n4312_ = ~pi164 | ~new_n1756_;
  assign new_n4313_ = ~new_n2361_ | ~new_n1716_;
  assign new_n4314_ = ~pi165 | ~new_n1756_;
  assign new_n4315_ = ~new_n2361_ | ~new_n1717_;
  assign new_n4316_ = ~pi166 | ~new_n1756_;
  assign new_n4317_ = ~new_n2361_ | ~new_n1718_;
  assign new_n4318_ = ~pi167 | ~new_n1756_;
  assign new_n4319_ = ~new_n2361_ | ~new_n1719_;
  assign new_n4320_ = ~pi168 | ~new_n1756_;
  assign new_n4321_ = ~new_n2361_ | ~new_n1720_;
  assign new_n4322_ = ~pi169 | ~new_n1756_;
  assign new_n4323_ = ~new_n2361_ | ~new_n1721_;
  assign new_n4324_ = ~pi170 | ~new_n1756_;
  assign new_n4325_ = ~new_n2361_ | ~new_n1722_;
  assign new_n4326_ = ~pi171 | ~new_n1756_;
  assign new_n4327_ = ~new_n2361_ | ~new_n1723_;
  assign new_n4328_ = ~pi172 | ~new_n1756_;
  assign new_n4329_ = ~new_n2361_ | ~new_n1724_;
  assign new_n4330_ = ~pi173 | ~new_n1756_;
  assign new_n4331_ = ~new_n2361_ | ~new_n1725_;
  assign new_n4332_ = ~pi174 | ~new_n1756_;
  assign new_n4333_ = ~new_n2361_ | ~new_n1726_;
  assign new_n4334_ = ~pi175 | ~new_n1756_;
  assign new_n4335_ = ~new_n2361_ | ~new_n1727_;
  assign new_n4336_ = ~pi176 | ~new_n1756_;
  assign new_n4337_ = ~new_n2361_ | ~new_n1728_;
  assign new_n4338_ = ~pi177 | ~new_n1756_;
  assign new_n4339_ = ~new_n2361_ | ~new_n1729_;
  assign new_n4340_ = ~pi178 | ~new_n1756_;
  assign new_n4341_ = ~new_n2361_ | ~new_n1730_;
  assign new_n4342_ = ~pi179 | ~new_n1756_;
  assign new_n4343_ = ~new_n2361_ | ~new_n1731_;
  assign new_n4344_ = ~pi180 | ~new_n1756_;
  assign new_n4345_ = ~new_n2361_ | ~new_n1732_;
  assign new_n4346_ = ~pi181 | ~new_n1756_;
  assign new_n4347_ = ~new_n2361_ | ~new_n1734_;
  assign new_n4348_ = ~pi182 | ~new_n1756_;
  assign new_n4349_ = ~new_n2361_ | ~new_n1736_;
  assign new_n4350_ = ~pi183 | ~new_n1756_;
  assign new_n4351_ = ~new_n2361_ | ~new_n1738_;
  assign new_n4352_ = ~pi184 | ~new_n1756_;
  assign new_n4353_ = ~new_n2361_ | ~new_n1740_;
  assign new_n4354_ = ~pi185 | ~new_n1756_;
  assign new_n4355_ = ~new_n2361_ | ~new_n1742_;
  assign new_n4356_ = ~pi186 | ~new_n1756_;
  assign new_n4357_ = ~new_n2361_ | ~new_n1744_;
  assign new_n4358_ = ~pi187 | ~new_n1756_;
  assign new_n4359_ = ~new_n2361_ | ~new_n1746_;
  assign new_n4360_ = ~pi188 | ~new_n1756_;
  assign new_n4361_ = ~new_n2361_ | ~new_n1748_;
  assign new_n4362_ = ~pi189 | ~new_n1756_;
  assign new_n4363_ = ~new_n2361_ | ~new_n1750_;
  assign new_n4364_ = ~pi190 | ~new_n1756_;
  assign new_n4365_ = ~new_n2361_ | ~new_n1752_;
  assign new_n4366_ = ~pi191 | ~new_n1756_;
  assign new_n4367_ = ~new_n2365_ | ~new_n2361_;
  assign new_n4368_ = ~pi192 | ~new_n1756_;
  assign new_n4369_ = ~new_n2365_ | ~new_n2361_;
  assign new_n4370_ = ~pi213 | ~new_n1764_;
  assign new_n4371_ = ~po266 | ~new_n1414_;
  assign new_n4372_ = ~pi214 | ~new_n1764_;
  assign new_n4373_ = ~po266 | ~new_n1415_;
  assign new_n4374_ = ~pi215 | ~new_n1764_;
  assign new_n4375_ = ~po266 | ~new_n1405_;
  assign new_n4376_ = ~pi216 | ~new_n1764_;
  assign new_n4377_ = ~po266 | ~new_n1401_;
  assign new_n4378_ = ~pi217 | ~new_n1764_;
  assign new_n4379_ = ~po266 | ~new_n1397_;
  assign new_n4380_ = ~pi218 | ~new_n1764_;
  assign new_n4381_ = ~po266 | ~new_n1404_;
  assign new_n4382_ = ~pi219 | ~new_n1764_;
  assign new_n4383_ = ~po266 | ~new_n1408_;
  assign new_n4384_ = ~pi220 | ~new_n1764_;
  assign new_n4385_ = ~po266 | ~new_n1407_;
  assign new_n4386_ = ~pi221 | ~new_n1764_;
  assign new_n4387_ = ~po266 | ~new_n1421_;
  assign new_n4388_ = ~pi222 | ~new_n1764_;
  assign new_n4389_ = ~po266 | ~new_n1420_;
  assign new_n4390_ = ~pi223 | ~new_n1764_;
  assign new_n4391_ = ~po266 | ~new_n1399_;
  assign new_n4392_ = ~pi224 | ~new_n1764_;
  assign new_n4393_ = ~po266 | ~new_n1400_;
  assign new_n4394_ = ~pi225 | ~new_n1764_;
  assign new_n4395_ = ~po266 | ~new_n1409_;
  assign new_n4396_ = ~pi226 | ~new_n1764_;
  assign new_n4397_ = ~po266 | ~new_n1417_;
  assign new_n4398_ = ~pi227 | ~new_n1764_;
  assign new_n4399_ = ~po266 | ~new_n1416_;
  assign new_n4400_ = ~pi228 | ~new_n1764_;
  assign new_n4401_ = ~po266 | ~new_n1411_;
  assign new_n4402_ = ~pi229 | ~new_n1764_;
  assign new_n4403_ = ~po266 | ~new_n1410_;
  assign new_n4404_ = ~pi230 | ~new_n1764_;
  assign new_n4405_ = ~po266 | ~new_n1406_;
  assign new_n4406_ = ~pi231 | ~new_n1764_;
  assign new_n4407_ = ~po266 | ~new_n1419_;
  assign new_n4408_ = ~pi232 | ~new_n1764_;
  assign new_n4409_ = ~po266 | ~new_n1418_;
  assign new_n4410_ = ~pi233 | ~new_n1764_;
  assign new_n4411_ = ~po266 | ~new_n1413_;
  assign new_n4412_ = ~pi234 | ~new_n1764_;
  assign new_n4413_ = ~po266 | ~new_n1412_;
  assign new_n4414_ = ~pi235 | ~new_n1764_;
  assign new_n4415_ = ~po266 | ~new_n1398_;
  assign new_n4416_ = ~pi236 | ~new_n1764_;
  assign new_n4417_ = ~po266 | ~new_n1403_;
  assign new_n4418_ = ~pi237 | ~new_n1764_;
  assign new_n4419_ = ~po266 | ~new_n1402_;
  assign new_n4420_ = ~pi238 | ~new_n1764_;
  assign new_n4421_ = ~po266 | ~new_n1395_;
  assign new_n4422_ = ~pi239 | ~new_n1764_;
  assign new_n4423_ = ~po266 | ~new_n1394_;
  assign new_n4424_ = ~pi240 | ~new_n1764_;
  assign new_n4425_ = ~po266 | ~new_n1390_;
  assign new_n4426_ = ~pi241 | ~new_n1764_;
  assign new_n4427_ = ~po266 | ~new_n1391_;
  assign new_n4428_ = ~pi242 | ~new_n1764_;
  assign new_n4429_ = ~po266 | ~new_n1392_;
  assign new_n4430_ = ~pi243 | ~new_n1764_;
  assign new_n4431_ = ~po266 | ~new_n1396_;
  assign new_n4432_ = ~pi244 | ~new_n1764_;
  assign new_n4433_ = ~po266 | ~new_n1393_;
  assign new_n4434_ = ~new_n2346_ | ~new_n1391_;
  assign new_n4435_ = ~new_n1749_ | ~new_n3031_;
  assign new_n4436_ = ~new_n4435_ | ~new_n4434_;
  assign new_n4437_ = ~new_n2347_ | ~new_n1390_;
  assign new_n4438_ = ~new_n1747_ | ~new_n3012_;
  assign new_n4439_ = ~new_n4438_ | ~new_n4437_;
  assign new_n4440_ = ~new_n2350_ | ~new_n1402_;
  assign new_n4441_ = ~new_n1741_ | ~new_n2955_;
  assign new_n4442_ = ~new_n4441_ | ~new_n4440_;
  assign new_n4443_ = ~new_n2351_ | ~new_n1403_;
  assign new_n4444_ = ~new_n1739_ | ~new_n2936_;
  assign new_n4445_ = ~new_n4444_ | ~new_n4443_;
  assign new_n4446_ = ~new_n2353_ | ~new_n1412_;
  assign new_n4447_ = ~new_n1735_ | ~new_n2898_;
  assign new_n4448_ = ~new_n4447_ | ~new_n4446_;
  assign new_n4449_ = ~new_n2352_ | ~new_n1398_;
  assign new_n4450_ = ~new_n1737_ | ~new_n2917_;
  assign new_n4451_ = ~new_n4450_ | ~new_n4449_;
  assign new_n4452_ = ~new_n2349_ | ~new_n1395_;
  assign new_n4453_ = ~new_n1743_ | ~new_n2974_;
  assign new_n4454_ = ~new_n4453_ | ~new_n4452_;
  assign new_n4455_ = ~new_n2348_ | ~new_n1394_;
  assign new_n4456_ = ~new_n1745_ | ~new_n2993_;
  assign new_n4457_ = ~new_n4456_ | ~new_n4455_;
  assign new_n4458_ = ~new_n4203_ | ~new_n2822_;
  assign new_n4459_ = ~new_n1843_ | ~new_n1406_;
  assign new_n4460_ = ~new_n4459_ | ~new_n4458_;
  assign new_n4461_ = ~new_n4140_ | ~new_n2651_;
  assign new_n4462_ = ~new_n1816_ | ~new_n1421_;
  assign new_n4463_ = ~new_n4462_ | ~new_n4461_;
  assign new_n4464_ = ~new_n4147_ | ~new_n2670_;
  assign new_n4465_ = ~new_n1819_ | ~new_n1420_;
  assign new_n4466_ = ~new_n4465_ | ~new_n4464_;
  assign new_n4467_ = ~new_n4175_ | ~new_n2746_;
  assign new_n4468_ = ~new_n1831_ | ~new_n1417_;
  assign new_n4469_ = ~new_n4468_ | ~new_n4467_;
  assign new_n4470_ = ~new_n4182_ | ~new_n2765_;
  assign new_n4471_ = ~new_n1834_ | ~new_n1416_;
  assign new_n4472_ = ~new_n4471_ | ~new_n4470_;
  assign new_n4473_ = ~new_n4076_ | ~new_n2537_;
  assign new_n4474_ = ~new_n1790_ | ~new_n1414_;
  assign new_n4475_ = ~new_n4474_ | ~new_n4473_;
  assign new_n4476_ = ~new_n4091_ | ~new_n2513_;
  assign new_n4477_ = ~new_n1795_ | ~new_n1415_;
  assign new_n4478_ = ~new_n4477_ | ~new_n4476_;
  assign new_n4479_ = ~new_n4189_ | ~new_n2784_;
  assign new_n4480_ = ~new_n1837_ | ~new_n1411_;
  assign new_n4481_ = ~new_n4480_ | ~new_n4479_;
  assign new_n4482_ = ~new_n4196_ | ~new_n2803_;
  assign new_n4483_ = ~new_n1840_ | ~new_n1410_;
  assign new_n4484_ = ~new_n4483_ | ~new_n4482_;
  assign new_n4485_ = ~new_n4126_ | ~new_n2613_;
  assign new_n4486_ = ~new_n1810_ | ~new_n1408_;
  assign new_n4487_ = ~new_n4486_ | ~new_n4485_;
  assign new_n4488_ = ~new_n4133_ | ~new_n2632_;
  assign new_n4489_ = ~new_n1813_ | ~new_n1407_;
  assign new_n4490_ = ~new_n4489_ | ~new_n4488_;
  assign new_n4491_ = ~new_n4168_ | ~new_n2727_;
  assign new_n4492_ = ~new_n1828_ | ~new_n1409_;
  assign new_n4493_ = ~new_n4492_ | ~new_n4491_;
  assign new_n4494_ = ~new_n4098_ | ~new_n2532_;
  assign new_n4495_ = ~new_n1798_ | ~new_n1405_;
  assign new_n4496_ = ~new_n4495_ | ~new_n4494_;
  assign new_n4497_ = ~new_n4105_ | ~new_n2556_;
  assign new_n4498_ = ~new_n1801_ | ~new_n1401_;
  assign new_n4499_ = ~new_n4498_ | ~new_n4497_;
  assign new_n4500_ = ~new_n4119_ | ~new_n2594_;
  assign new_n4501_ = ~new_n1807_ | ~new_n1404_;
  assign new_n4502_ = ~new_n4501_ | ~new_n4500_;
  assign new_n4503_ = ~new_n4210_ | ~new_n2841_;
  assign new_n4504_ = ~new_n1846_ | ~new_n1419_;
  assign new_n4505_ = ~new_n4504_ | ~new_n4503_;
  assign new_n4506_ = ~new_n2355_ | ~new_n1393_;
  assign new_n4507_ = ~new_n1754_ | ~new_n3088_;
  assign new_n4508_ = ~new_n4507_ | ~new_n4506_;
  assign new_n4509_ = ~new_n4215_ | ~new_n2860_;
  assign new_n4510_ = ~new_n1848_ | ~new_n1418_;
  assign new_n4511_ = ~new_n4510_ | ~new_n4509_;
  assign new_n4512_ = ~new_n4161_ | ~new_n2708_;
  assign new_n4513_ = ~new_n1825_ | ~new_n1400_;
  assign new_n4514_ = ~new_n4513_ | ~new_n4512_;
  assign new_n4515_ = ~new_n4112_ | ~new_n2575_;
  assign new_n4516_ = ~new_n1804_ | ~new_n1397_;
  assign new_n4517_ = ~new_n4516_ | ~new_n4515_;
  assign new_n4518_ = ~new_n4154_ | ~new_n2689_;
  assign new_n4519_ = ~new_n1822_ | ~new_n1399_;
  assign new_n4520_ = ~new_n4519_ | ~new_n4518_;
  assign new_n4521_ = ~new_n2354_ | ~new_n1413_;
  assign new_n4522_ = ~new_n1733_ | ~new_n2879_;
  assign new_n4523_ = ~new_n4522_ | ~new_n4521_;
  assign new_n4524_ = ~new_n2357_ | ~new_n1392_;
  assign new_n4525_ = ~new_n1751_ | ~new_n3050_;
  assign new_n4526_ = ~new_n4525_ | ~new_n4524_;
  assign new_n4527_ = ~new_n2356_ | ~new_n1396_;
  assign new_n4528_ = ~new_n1753_ | ~new_n3068_;
  assign new_n4529_ = ~new_n4528_ | ~new_n4527_;
  assign new_n4530_ = ~new_n3458_ | ~new_n2326_;
  assign new_n4531_ = ~new_n1693_ | ~new_n2321_;
  assign new_n4532_ = ~new_n4531_ | ~new_n4530_;
  assign new_n4533_ = ~new_n1787_ | ~new_n2322_ | ~new_n1778_ | ~new_n4049_;
  assign new_n4534_ = ~new_n4532_ | ~new_n4058_;
  assign new_n4535_ = ~new_n4534_ | ~new_n4533_;
  assign new_n4536_ = ~new_n4055_ | ~new_n10877_ | ~new_n2326_;
  assign new_n4537_ = ~new_n4535_ | ~new_n1781_;
  assign new_n4538_ = ~new_n2322_ | ~new_n2358_ | ~new_n1361_;
  assign new_n4539_ = ~new_n13286_ | ~new_n2327_ | ~new_n2331_;
  assign new_n4540_ = ~new_n1420_ | ~new_n11071_;
  assign new_n4541_ = ~new_n1420_ | ~new_n2324_;
  assign new_n4542_ = ~new_n1421_ | ~new_n11071_;
  assign new_n4543_ = ~new_n1421_ | ~new_n2324_;
  assign new_n4544_ = ~new_n1407_ | ~new_n11071_;
  assign new_n4545_ = ~new_n1407_ | ~new_n2324_;
  assign new_n4546_ = ~new_n1408_ | ~new_n11071_;
  assign new_n4547_ = ~new_n1408_ | ~new_n2324_;
  assign new_n4548_ = ~new_n1404_ | ~new_n11071_;
  assign new_n4549_ = ~new_n1404_ | ~new_n2324_;
  assign new_n4550_ = ~new_n1397_ | ~new_n11071_;
  assign new_n4551_ = ~new_n1397_ | ~new_n2324_;
  assign new_n4552_ = ~new_n1401_ | ~new_n11071_;
  assign new_n4553_ = ~new_n1401_ | ~new_n2324_;
  assign new_n4554_ = ~new_n9438_ | ~new_n11071_;
  assign new_n4555_ = ~new_n1393_ | ~new_n2324_;
  assign new_n4556_ = ~new_n9436_ | ~new_n11071_;
  assign new_n4557_ = ~new_n1396_ | ~new_n2324_;
  assign new_n4558_ = ~new_n1405_ | ~new_n11071_;
  assign new_n4559_ = ~new_n1405_ | ~new_n2324_;
  assign new_n4560_ = ~new_n1392_ | ~new_n11071_;
  assign new_n4561_ = ~new_n1392_ | ~new_n2324_;
  assign new_n4562_ = ~new_n1391_ | ~new_n11071_;
  assign new_n4563_ = ~new_n1391_ | ~new_n2324_;
  assign new_n4564_ = ~new_n1390_ | ~new_n11071_;
  assign new_n4565_ = ~new_n1390_ | ~new_n2324_;
  assign new_n4566_ = ~new_n1394_ | ~new_n11071_;
  assign new_n4567_ = ~new_n1394_ | ~new_n2324_;
  assign new_n4568_ = ~new_n1395_ | ~new_n11071_;
  assign new_n4569_ = ~new_n1395_ | ~new_n2324_;
  assign new_n4570_ = ~new_n1402_ | ~new_n11071_;
  assign new_n4571_ = ~new_n1402_ | ~new_n2324_;
  assign new_n4572_ = ~new_n1403_ | ~new_n11071_;
  assign new_n4573_ = ~new_n1403_ | ~new_n2324_;
  assign new_n4574_ = ~new_n1398_ | ~new_n11071_;
  assign new_n4575_ = ~new_n1398_ | ~new_n2324_;
  assign new_n4576_ = ~new_n1412_ | ~new_n11071_;
  assign new_n4577_ = ~new_n1412_ | ~new_n2324_;
  assign new_n4578_ = ~new_n1413_ | ~new_n11071_;
  assign new_n4579_ = ~new_n1413_ | ~new_n2324_;
  assign new_n4580_ = ~new_n1415_ | ~new_n11071_;
  assign new_n4581_ = ~new_n1415_ | ~new_n2324_;
  assign new_n4582_ = ~new_n1418_ | ~new_n11071_;
  assign new_n4583_ = ~new_n1418_ | ~new_n2324_;
  assign new_n4584_ = ~new_n1419_ | ~new_n11071_;
  assign new_n4585_ = ~new_n1419_ | ~new_n2324_;
  assign new_n4586_ = ~new_n1406_ | ~new_n11071_;
  assign new_n4587_ = ~new_n1406_ | ~new_n2324_;
  assign new_n4588_ = ~new_n1410_ | ~new_n11071_;
  assign new_n4589_ = ~new_n1410_ | ~new_n2324_;
  assign new_n4590_ = ~new_n1411_ | ~new_n11071_;
  assign new_n4591_ = ~new_n1411_ | ~new_n2324_;
  assign new_n4592_ = ~new_n1416_ | ~new_n11071_;
  assign new_n4593_ = ~new_n1416_ | ~new_n2324_;
  assign new_n4594_ = ~new_n1417_ | ~new_n11071_;
  assign new_n4595_ = ~new_n1417_ | ~new_n2324_;
  assign new_n4596_ = ~new_n1409_ | ~new_n11071_;
  assign new_n4597_ = ~new_n1409_ | ~new_n2324_;
  assign new_n4598_ = ~new_n1400_ | ~new_n11071_;
  assign new_n4599_ = ~new_n1400_ | ~new_n2324_;
  assign new_n4600_ = ~new_n1399_ | ~new_n11071_;
  assign new_n4601_ = ~new_n1399_ | ~new_n2324_;
  assign new_n4602_ = ~new_n1414_ | ~new_n11071_;
  assign new_n4603_ = ~new_n1414_ | ~new_n2324_;
  assign new_n4604_ = ~new_n1788_ | ~new_n3735_;
  assign new_n4605_ = ~new_n4070_ | ~new_n1354_ | ~pi161;
  assign new_n4606_ = ~new_n4696_ | ~new_n20698_;
  assign new_n4607_ = ~new_n5105_ | ~new_n20699_;
  assign new_n4608_ = ~new_n20902_ | ~new_n20816_;
  assign new_n4609_ = ~new_n20979_ | ~new_n20817_;
  assign new_n4610_ = ~new_n4695_ | ~new_n20701_;
  assign new_n4611_ = ~new_n5108_ | ~new_n20704_;
  assign new_n4612_ = ~new_n20815_ | ~new_n20970_;
  assign new_n4613_ = ~new_n20978_ | ~new_n20731_;
  assign new_n4614_ = ~new_n4690_ | ~new_n20690_;
  assign new_n4615_ = ~new_n5111_ | ~new_n20703_;
  assign new_n4616_ = ~new_n4617_ | ~new_n4618_;
  assign new_n4617_ = ~new_n4689_ | ~new_n20700_;
  assign new_n4618_ = ~new_n5114_ | ~new_n20702_;
  assign new_n4619_ = ~new_n20784_ | ~new_n20814_;
  assign new_n4620_ = ~new_n20912_ | ~new_n4621_;
  assign new_n4621_ = ~new_n20784_;
  assign new_n4622_ = ~new_n4685_ | ~new_n20706_;
  assign new_n4623_ = ~new_n5117_ | ~new_n20707_;
  assign new_n4624_ = ~new_n20783_ | ~new_n20813_;
  assign new_n4625_ = ~new_n20916_ | ~new_n4626_;
  assign new_n4626_ = ~new_n20783_;
  assign new_n4627_ = ~new_n4698_ | ~new_n20812_;
  assign new_n4628_ = ~new_n5120_ | ~new_n20708_;
  assign new_n4629_ = ~new_n20782_ | ~new_n20811_;
  assign new_n4630_ = new_n5055_ & new_n7327_ & new_n5057_;
  assign new_n4631_ = new_n5061_ & new_n5055_ & new_n5057_;
  assign new_n4632_ = new_n5570_ & new_n7330_;
  assign new_n4633_ = new_n5577_ & new_n5056_;
  assign new_n4634_ = new_n5056_ & new_n5055_ & new_n5061_;
  assign new_n4635_ = new_n7290_ & new_n5055_;
  assign new_n4636_ = new_n5245_ & new_n5240_;
  assign new_n4637_ = new_n7349_ & new_n5060_;
  assign new_n4638_ = new_n5063_ & new_n5060_;
  assign new_n4639_ = new_n5058_ & new_n5059_;
  assign new_n4640_ = new_n7339_ & new_n5059_;
  assign new_n4641_ = new_n7336_ & new_n5058_;
  assign new_n4642_ = new_n7339_ & new_n7336_;
  assign new_n4643_ = new_n4664_ & pi520;
  assign new_n4644_ = new_n4666_ & new_n7324_;
  assign new_n4645_ = new_n5427_ & new_n5040_;
  assign new_n4646_ = new_n5598_ & new_n7344_;
  assign new_n4647_ = new_n5565_ & new_n7330_;
  assign new_n4648_ = new_n5506_ & new_n5581_;
  assign new_n4649_ = new_n4975_ & pi520;
  assign new_n4650_ = new_n5572_ & new_n5599_;
  assign new_n4651_ = new_n5599_ & new_n6329_;
  assign new_n4652_ = new_n5573_ & new_n5599_;
  assign new_n4653_ = new_n5367_ & new_n5599_;
  assign new_n4654_ = new_n5598_ & new_n5060_;
  assign new_n4655_ = new_n5581_ & new_n7344_;
  assign new_n4656_ = new_n5599_ & new_n4646_;
  assign new_n4657_ = new_n5581_ & new_n5060_;
  assign new_n4658_ = new_n4645_ & new_n7349_;
  assign new_n4659_ = new_n4645_ & new_n7344_;
  assign new_n4660_ = new_n4645_ & new_n4638_;
  assign new_n4661_ = new_n4643_ & new_n5040_;
  assign new_n4662_ = new_n6812_ & pi520;
  assign new_n4663_ = new_n4643_ & new_n6814_;
  assign new_n4664_ = new_n7317_ & new_n5036_;
  assign new_n4665_ = new_n5246_ & new_n4636_;
  assign new_n4666_ = new_n7330_ & new_n5061_;
  assign new_n4667_ = new_n5566_ & new_n6325_;
  assign new_n4668_ = new_n5038_ & pi520;
  assign new_n4669_ = ~new_n6241_ | ~new_n6238_ | ~new_n6239_ | ~new_n6240_;
  assign new_n4670_ = ~new_n6260_ | ~new_n6257_ | ~new_n6258_ | ~new_n6259_;
  assign new_n4671_ = ~new_n6276_ | ~new_n6277_ | ~new_n6279_ | ~new_n6278_;
  assign new_n4672_ = ~new_n6315_ | ~new_n6316_ | ~new_n6317_;
  assign new_n4673_ = ~new_n6222_ | ~new_n6219_ | ~new_n6220_ | ~new_n6221_;
  assign new_n4674_ = ~new_n6203_ | ~new_n6200_ | ~new_n6201_ | ~new_n6202_;
  assign new_n4675_ = ~new_n6295_ | ~new_n6296_ | ~new_n6297_;
  assign new_n4676_ = ~new_n5801_ | ~new_n5802_ | ~new_n5804_ | ~new_n5803_;
  assign new_n4677_ = ~new_n6146_ | ~new_n6143_ | ~new_n6144_ | ~new_n6145_;
  assign new_n4678_ = ~new_n5915_ | ~new_n5916_ | ~new_n5918_ | ~new_n5917_;
  assign new_n4679_ = ~new_n5934_ | ~new_n5935_ | ~new_n5937_ | ~new_n5936_;
  assign new_n4680_ = ~new_n5782_ | ~new_n5783_ | ~new_n5785_ | ~new_n5784_;
  assign new_n4681_ = ~new_n6184_ | ~new_n6181_ | ~new_n6182_ | ~new_n6183_;
  assign new_n4682_ = ~new_n6165_ | ~new_n6162_ | ~new_n6163_ | ~new_n6164_;
  assign new_n4683_ = ~new_n5820_ | ~new_n5821_ | ~new_n5823_ | ~new_n5822_;
  assign new_n4684_ = ~new_n7370_ | ~new_n7371_ | ~new_n5763_ | ~new_n5762_;
  assign new_n4685_ = ~new_n6051_ | ~new_n6048_ | ~new_n6049_ | ~new_n6050_;
  assign new_n4686_ = ~new_n5858_ | ~new_n5859_ | ~new_n5861_ | ~new_n5860_;
  assign new_n4687_ = ~new_n5839_ | ~new_n5840_ | ~new_n5842_ | ~new_n5841_;
  assign new_n4688_ = ~new_n5953_ | ~new_n5954_ | ~new_n5956_ | ~new_n5955_;
  assign new_n4689_ = ~new_n6029_ | ~new_n6030_ | ~new_n6032_ | ~new_n6031_;
  assign new_n4690_ = ~new_n6010_ | ~new_n6011_ | ~new_n6013_ | ~new_n6012_;
  assign new_n4691_ = ~new_n6127_ | ~new_n6124_ | ~new_n6125_ | ~new_n6126_;
  assign new_n4692_ = ~new_n6108_ | ~new_n6105_ | ~new_n6106_ | ~new_n6107_;
  assign new_n4693_ = ~new_n7363_ | ~new_n7364_ | ~new_n5766_ | ~new_n5765_;
  assign new_n4694_ = ~new_n7340_ | ~new_n7341_ | ~new_n5745_ | ~new_n5744_;
  assign new_n4695_ = ~new_n5991_ | ~new_n5992_ | ~new_n5994_ | ~new_n5993_;
  assign new_n4696_ = ~new_n5972_ | ~new_n5973_ | ~new_n5975_ | ~new_n5974_;
  assign new_n4697_ = ~new_n6089_ | ~new_n6086_ | ~new_n6087_ | ~new_n6088_;
  assign new_n4698_ = ~new_n6070_ | ~new_n6067_ | ~new_n6068_ | ~new_n6069_;
  assign new_n4699_ = ~new_n5896_ | ~new_n5897_ | ~new_n5899_ | ~new_n5898_;
  assign new_n4700_ = ~new_n5877_ | ~new_n5878_ | ~new_n5880_ | ~new_n5879_;
  assign new_n4701_ = ~new_n7212_ | ~new_n7211_;
  assign new_n4702_ = ~new_n7214_ | ~new_n7213_;
  assign new_n4703_ = ~new_n7218_ | ~new_n7219_ | ~new_n7220_;
  assign new_n4704_ = ~new_n7221_ | ~new_n7222_ | ~new_n7223_;
  assign new_n4705_ = ~new_n7224_ | ~new_n7225_ | ~new_n7226_;
  assign new_n4706_ = ~new_n7227_ | ~new_n7228_ | ~new_n7229_;
  assign new_n4707_ = ~new_n7230_ | ~new_n7231_ | ~new_n7232_;
  assign new_n4708_ = ~new_n7233_ | ~new_n7234_ | ~new_n7235_;
  assign new_n4709_ = ~new_n7236_ | ~new_n7237_ | ~new_n7238_;
  assign new_n4710_ = ~new_n7239_ | ~new_n7240_ | ~new_n7241_;
  assign new_n4711_ = ~new_n7242_ | ~new_n7243_ | ~new_n7244_;
  assign new_n4712_ = ~new_n7245_ | ~new_n7246_ | ~new_n7247_;
  assign new_n4713_ = ~new_n7251_ | ~new_n7252_ | ~new_n7253_;
  assign new_n4714_ = ~new_n7254_ | ~new_n7255_ | ~new_n7256_;
  assign new_n4715_ = ~new_n7257_ | ~new_n7258_ | ~new_n7259_;
  assign new_n4716_ = ~new_n7260_ | ~new_n7261_ | ~new_n7262_;
  assign new_n4717_ = ~new_n7263_ | ~new_n7264_ | ~new_n7265_;
  assign new_n4718_ = ~new_n7266_ | ~new_n7267_ | ~new_n7268_;
  assign new_n4719_ = ~new_n7269_ | ~new_n7270_ | ~new_n7271_;
  assign new_n4720_ = ~new_n7272_ | ~new_n7273_ | ~new_n7274_;
  assign new_n4721_ = ~new_n7277_ | ~new_n7276_ | ~new_n7275_;
  assign new_n4722_ = ~new_n7280_ | ~new_n7279_ | ~new_n7278_;
  assign new_n4723_ = ~new_n7195_ | ~new_n7194_ | ~new_n7193_;
  assign new_n4724_ = ~new_n7198_ | ~new_n7197_ | ~new_n7196_;
  assign new_n4725_ = ~new_n7201_ | ~new_n7200_ | ~new_n7199_;
  assign new_n4726_ = ~new_n7204_ | ~new_n7203_ | ~new_n7202_;
  assign new_n4727_ = ~new_n7207_ | ~new_n7206_ | ~new_n7205_;
  assign new_n4728_ = ~new_n7210_ | ~new_n7209_ | ~new_n7208_;
  assign new_n4729_ = ~new_n7216_ | ~new_n7217_ | ~new_n7215_;
  assign new_n4730_ = ~new_n7250_ | ~new_n7249_ | ~new_n7248_;
  assign new_n4731_ = ~new_n7283_ | ~new_n7282_ | ~new_n7281_;
  assign new_n4732_ = ~new_n7285_ | ~new_n7284_;
  assign new_n4733_ = ~new_n7143_ | ~new_n7142_;
  assign new_n4734_ = new_n7289_ & new_n7288_;
  assign new_n4735_ = ~new_n7148_ | ~new_n5052_ | ~new_n7147_;
  assign new_n4736_ = ~new_n7150_ | ~new_n5052_ | ~new_n7149_;
  assign new_n4737_ = ~new_n7152_ | ~new_n5052_ | ~new_n7151_;
  assign new_n4738_ = ~new_n7154_ | ~new_n5052_ | ~new_n7153_;
  assign new_n4739_ = ~new_n7156_ | ~new_n5052_ | ~new_n7155_;
  assign new_n4740_ = ~new_n7158_ | ~new_n5052_ | ~new_n7157_;
  assign new_n4741_ = ~new_n7160_ | ~new_n5052_ | ~new_n7159_;
  assign new_n4742_ = ~new_n7162_ | ~new_n5052_ | ~new_n7161_;
  assign new_n4743_ = ~new_n7164_ | ~new_n5052_ | ~new_n7163_;
  assign new_n4744_ = ~new_n7166_ | ~new_n5052_ | ~new_n7165_;
  assign new_n4745_ = ~new_n7169_ | ~new_n7170_ | ~new_n5052_;
  assign new_n4746_ = ~new_n7171_ | ~new_n7172_ | ~new_n5052_;
  assign new_n4747_ = ~new_n7173_ | ~new_n7174_ | ~new_n5052_;
  assign new_n4748_ = ~new_n7175_ | ~new_n7176_ | ~new_n5052_;
  assign new_n4749_ = ~new_n7177_ | ~new_n7178_ | ~new_n5052_;
  assign new_n4750_ = ~new_n7179_ | ~new_n7180_ | ~new_n5052_;
  assign new_n4751_ = ~new_n7181_ | ~new_n7182_ | ~new_n5052_;
  assign new_n4752_ = ~new_n7183_ | ~new_n7184_ | ~new_n5052_;
  assign new_n4753_ = ~new_n7186_ | ~new_n5052_ | ~new_n7185_;
  assign new_n4754_ = ~new_n7188_ | ~new_n5052_ | ~new_n7187_;
  assign new_n4755_ = ~new_n7131_ | ~new_n5052_ | ~new_n7130_;
  assign new_n4756_ = ~new_n7133_ | ~new_n5052_ | ~new_n7132_;
  assign new_n4757_ = ~new_n7135_ | ~new_n5052_ | ~new_n7134_;
  assign new_n4758_ = ~new_n7137_ | ~new_n5052_ | ~new_n7136_;
  assign new_n4759_ = ~new_n7139_ | ~new_n5052_ | ~new_n7138_;
  assign new_n4760_ = ~new_n7141_ | ~new_n5052_ | ~new_n7140_;
  assign new_n4761_ = ~new_n7146_ | ~new_n5052_ | ~new_n7145_;
  assign new_n4762_ = ~new_n7168_ | ~new_n5052_ | ~new_n7167_;
  assign new_n4763_ = ~new_n7190_ | ~new_n5052_ | ~new_n7189_;
  assign new_n4764_ = ~new_n7192_ | ~new_n5052_ | ~new_n7191_;
  assign new_n4765_ = ~new_n5056_ | ~new_n5052_ | ~new_n7127_;
  assign new_n4766_ = ~new_n5521_ | ~new_n5598_;
  assign po510 = ~new_n5519_ | ~new_n7062_;
  assign po509 = ~pi520;
  assign new_n4769_ = ~new_n7079_ | ~new_n7078_;
  assign new_n4770_ = ~new_n7081_ | ~new_n7080_;
  assign new_n4771_ = ~new_n7085_ | ~new_n7084_;
  assign new_n4772_ = ~new_n7087_ | ~new_n7086_;
  assign new_n4773_ = ~new_n7089_ | ~new_n7088_;
  assign new_n4774_ = ~new_n7091_ | ~new_n7090_;
  assign new_n4775_ = ~new_n7093_ | ~new_n7092_;
  assign new_n4776_ = ~new_n7095_ | ~new_n7094_;
  assign new_n4777_ = ~new_n7097_ | ~new_n7096_;
  assign new_n4778_ = ~new_n7099_ | ~new_n7098_;
  assign new_n4779_ = ~new_n7101_ | ~new_n7100_;
  assign new_n4780_ = ~new_n7103_ | ~new_n7102_;
  assign new_n4781_ = ~new_n7106_ | ~new_n7105_;
  assign new_n4782_ = ~new_n7108_ | ~new_n7107_;
  assign new_n4783_ = ~new_n7110_ | ~new_n7109_;
  assign new_n4784_ = ~new_n7112_ | ~new_n7111_;
  assign new_n4785_ = ~new_n7114_ | ~new_n7113_;
  assign new_n4786_ = ~new_n7116_ | ~new_n7115_;
  assign new_n4787_ = ~new_n7118_ | ~new_n7117_;
  assign new_n4788_ = ~new_n7120_ | ~new_n7119_;
  assign new_n4789_ = ~new_n7122_ | ~new_n7121_;
  assign new_n4790_ = ~new_n7124_ | ~new_n7123_;
  assign new_n4791_ = ~new_n7067_ | ~new_n7066_;
  assign new_n4792_ = ~new_n7069_ | ~new_n7068_;
  assign new_n4793_ = ~new_n7071_ | ~new_n7070_;
  assign new_n4794_ = ~new_n7073_ | ~new_n7072_;
  assign new_n4795_ = ~new_n7075_ | ~new_n7074_;
  assign new_n4796_ = ~new_n7077_ | ~new_n7076_;
  assign new_n4797_ = ~new_n7083_ | ~new_n7082_;
  assign new_n4798_ = new_n7299_ & new_n7295_;
  assign new_n4799_ = new_n7298_ & new_n7296_;
  assign new_n4800_ = new_n7300_ & new_n7297_;
  assign new_n4801_ = new_n7064_ & new_n4670_;
  assign new_n4802_ = new_n7064_ & new_n4669_;
  assign new_n4803_ = new_n7064_ & new_n4673_;
  assign new_n4804_ = new_n7064_ & new_n4674_;
  assign new_n4805_ = new_n7064_ & new_n4681_;
  assign new_n4806_ = new_n7064_ & new_n4682_;
  assign new_n4807_ = new_n7064_ & new_n4677_;
  assign new_n4808_ = new_n7064_ & new_n4691_;
  assign new_n4809_ = new_n7064_ & new_n4692_;
  assign new_n4810_ = new_n7064_ & new_n4697_;
  assign new_n4811_ = new_n7064_ & new_n4698_;
  assign new_n4812_ = new_n7064_ & new_n4685_;
  assign new_n4813_ = new_n7064_ & new_n4689_;
  assign new_n4814_ = new_n7064_ & new_n4690_;
  assign new_n4815_ = new_n7064_ & new_n4695_;
  assign new_n4816_ = new_n7064_ & new_n4696_;
  assign new_n4817_ = new_n7064_ & new_n4688_;
  assign new_n4818_ = new_n7064_ & new_n4679_;
  assign new_n4819_ = new_n7064_ & new_n4678_;
  assign new_n4820_ = new_n7064_ & new_n4699_;
  assign new_n4821_ = new_n7064_ & new_n4700_;
  assign new_n4822_ = new_n7064_ & new_n4686_;
  assign new_n4823_ = new_n7064_ & new_n4687_;
  assign new_n4824_ = new_n7064_ & new_n4683_;
  assign new_n4825_ = new_n7064_ & new_n4676_;
  assign new_n4826_ = new_n7064_ & new_n4680_;
  assign new_n4827_ = new_n7064_ & new_n4684_;
  assign new_n4828_ = new_n7064_ & new_n4694_;
  assign new_n4829_ = new_n7064_ & new_n4693_;
  assign new_n4830_ = ~new_n4986_ | ~new_n7886_ | ~new_n7885_;
  assign po508 = ~new_n7060_ | ~new_n7059_ | ~new_n7061_ | ~new_n7058_ | ~new_n7057_;
  assign po507 = ~new_n7051_ | ~new_n7048_ | ~new_n7052_ | ~new_n7049_ | ~new_n7050_;
  assign po506 = ~new_n7042_ | ~new_n7041_ | ~new_n7043_ | ~new_n7040_ | ~new_n7039_;
  assign po505 = ~new_n7033_ | ~new_n7030_ | ~new_n7034_ | ~new_n7031_ | ~new_n7032_;
  assign po504 = ~new_n7024_ | ~new_n7023_ | ~new_n7025_ | ~new_n7022_ | ~new_n7021_;
  assign po503 = ~new_n7014_ | ~new_n5517_ | ~new_n7013_;
  assign po502 = ~new_n7006_ | ~new_n5516_ | ~new_n7004_ | ~new_n7005_;
  assign po501 = ~new_n6997_ | ~new_n6994_ | ~new_n6998_ | ~new_n6995_ | ~new_n6996_;
  assign po500 = ~new_n6988_ | ~new_n6987_ | ~new_n6989_ | ~new_n6986_ | ~new_n6985_;
  assign po499 = ~new_n6978_ | ~new_n5514_ | ~new_n6977_;
  assign po498 = ~new_n6970_ | ~new_n6967_ | ~new_n6971_ | ~new_n6968_ | ~new_n6969_;
  assign po497 = ~new_n6961_ | ~new_n6960_ | ~new_n6962_ | ~new_n6959_ | ~new_n6958_;
  assign po496 = ~new_n6952_ | ~new_n6949_ | ~new_n6953_ | ~new_n6950_ | ~new_n6951_;
  assign po495 = ~new_n6943_ | ~new_n6942_ | ~new_n6944_ | ~new_n6941_ | ~new_n6940_;
  assign po494 = ~new_n5513_ | ~new_n6933_ | ~new_n6932_ | ~new_n6931_;
  assign po493 = ~new_n6925_ | ~new_n6924_ | ~new_n6926_ | ~new_n6923_ | ~new_n6922_;
  assign po492 = ~new_n6916_ | ~new_n6913_ | ~new_n6917_ | ~new_n6914_ | ~new_n6915_;
  assign po491 = ~new_n6906_ | ~new_n5512_ | ~new_n6905_ | ~new_n6904_;
  assign po490 = ~new_n6898_ | ~new_n6897_ | ~new_n6899_ | ~new_n6896_ | ~new_n6895_;
  assign po489 = ~new_n5510_ | ~new_n5511_ | ~new_n6888_;
  assign po488 = ~new_n6881_ | ~new_n6878_ | ~new_n6882_ | ~new_n6879_ | ~new_n6880_;
  assign po487 = ~new_n6872_ | ~new_n6871_ | ~new_n6873_ | ~new_n6870_ | ~new_n6869_;
  assign po486 = ~new_n6863_ | ~new_n6860_ | ~new_n6864_ | ~new_n6861_ | ~new_n6862_;
  assign po485 = ~new_n6854_ | ~new_n6853_ | ~new_n6855_ | ~new_n6852_ | ~new_n6851_;
  assign po484 = ~new_n6844_ | ~new_n5507_ | ~new_n6843_;
  assign po483 = ~new_n6836_ | ~new_n6835_ | ~new_n6837_ | ~new_n6834_ | ~new_n6833_;
  assign po482 = ~new_n6827_ | ~new_n6826_ | ~new_n6828_ | ~new_n6825_ | ~new_n6824_;
  assign po481 = ~new_n6818_ | ~new_n6815_ | ~new_n6819_ | ~new_n6816_ | ~new_n6817_;
  assign po480 = ~new_n6805_ | ~new_n6804_ | ~new_n6806_ | ~new_n6803_ | ~new_n6802_;
  assign po479 = new_n7287_ & new_n6790_;
  assign po446 = ~new_n5488_ | ~new_n5487_;
  assign po445 = ~new_n5484_ | ~new_n5483_;
  assign po444 = ~new_n5481_ | ~new_n5480_;
  assign po443 = ~new_n5478_ | ~new_n5477_;
  assign po442 = ~new_n5475_ | ~new_n5474_;
  assign po441 = ~new_n5472_ | ~new_n5471_;
  assign po440 = ~new_n5469_ | ~new_n5468_;
  assign po439 = ~new_n5466_ | ~new_n5465_;
  assign po438 = ~new_n5463_ | ~new_n5462_;
  assign po437 = ~new_n5458_ | ~new_n5459_ | ~new_n5460_;
  assign po436 = ~new_n5455_ | ~new_n5456_ | ~new_n5457_;
  assign po435 = ~new_n5452_ | ~new_n5453_ | ~new_n5454_;
  assign po434 = ~new_n5449_ | ~new_n5450_ | ~new_n5451_;
  assign po433 = ~new_n5446_ | ~new_n5447_ | ~new_n5448_;
  assign po432 = ~new_n5443_ | ~new_n5444_ | ~new_n5445_;
  assign po431 = ~new_n5440_ | ~new_n5441_ | ~new_n5442_;
  assign po430 = ~new_n5437_ | ~new_n5438_ | ~new_n5439_;
  assign po429 = ~new_n5434_ | ~new_n5435_ | ~new_n5436_;
  assign po428 = ~new_n5431_ | ~new_n5432_ | ~new_n5433_;
  assign po427 = ~new_n5428_ | ~new_n5429_ | ~new_n5430_;
  assign po426 = ~new_n6482_ | ~new_n5560_ | ~new_n6481_;
  assign po425 = ~new_n6480_ | ~new_n5559_ | ~new_n6479_;
  assign po424 = ~new_n5557_ | ~new_n6475_ | ~new_n6478_ | ~new_n6476_ | ~new_n6477_;
  assign po423 = ~new_n5556_ | ~new_n6471_ | ~new_n5424_ | ~new_n5425_;
  assign po422 = ~new_n5555_ | ~new_n6466_ | ~new_n5422_ | ~new_n5423_;
  assign po421 = ~new_n5554_ | ~new_n6461_ | ~new_n5420_ | ~new_n5421_;
  assign po420 = ~new_n5553_ | ~new_n6456_ | ~new_n5418_ | ~new_n5419_;
  assign po419 = ~new_n5552_ | ~new_n6451_ | ~new_n5416_ | ~new_n5417_;
  assign po418 = ~new_n5551_ | ~new_n6446_ | ~new_n5414_ | ~new_n5415_;
  assign po417 = ~new_n5550_ | ~new_n6441_ | ~new_n5412_ | ~new_n5413_;
  assign po416 = ~new_n5549_ | ~new_n6436_ | ~new_n5410_ | ~new_n5411_;
  assign po415 = ~new_n5548_ | ~new_n6431_ | ~new_n5408_ | ~new_n5409_;
  assign po414 = ~new_n5547_ | ~new_n6426_ | ~new_n5406_ | ~new_n5407_;
  assign po413 = ~new_n5546_ | ~new_n6421_ | ~new_n5404_ | ~new_n5405_;
  assign po412 = ~new_n5545_ | ~new_n6416_ | ~new_n5402_ | ~new_n5403_;
  assign po411 = ~new_n5544_ | ~new_n6411_ | ~new_n5400_ | ~new_n5401_;
  assign po410 = ~new_n5543_ | ~new_n6406_ | ~new_n5398_ | ~new_n5399_;
  assign po409 = ~new_n5542_ | ~new_n6401_ | ~new_n5396_ | ~new_n5397_;
  assign po408 = ~new_n5541_ | ~new_n6396_ | ~new_n5394_ | ~new_n5395_;
  assign po407 = ~new_n5540_ | ~new_n6391_ | ~new_n5392_ | ~new_n5393_;
  assign po406 = ~new_n5539_ | ~new_n5391_ | ~new_n5390_;
  assign po405 = ~new_n5538_ | ~new_n6381_ | ~new_n5388_ | ~new_n5389_;
  assign po404 = ~new_n5537_ | ~new_n5387_ | ~new_n5386_;
  assign po403 = ~new_n5536_ | ~new_n5385_ | ~new_n5384_;
  assign po402 = ~new_n5535_ | ~new_n5383_ | ~new_n5382_;
  assign po401 = ~new_n5534_ | ~new_n5381_ | ~new_n5380_;
  assign po400 = ~new_n5533_ | ~new_n5379_ | ~new_n5378_;
  assign po399 = ~new_n5377_ | ~new_n5376_;
  assign po398 = ~new_n5375_ | ~new_n5374_;
  assign po397 = ~new_n5373_ | ~new_n5372_;
  assign po396 = ~new_n5371_ | ~new_n5370_;
  assign po395 = ~new_n5369_ | ~new_n5368_;
  assign po330 = pi341 & new_n5524_;
  assign po329 = pi340 & new_n5524_;
  assign po328 = pi339 & new_n5524_;
  assign po327 = pi338 & new_n5524_;
  assign po326 = pi337 & new_n5524_;
  assign po325 = pi336 & new_n5524_;
  assign po324 = pi335 & new_n5524_;
  assign po323 = pi334 & new_n5524_;
  assign po322 = pi333 & new_n5524_;
  assign po321 = pi332 & new_n5524_;
  assign po320 = pi331 & new_n5524_;
  assign po319 = pi330 & new_n5524_;
  assign po318 = pi329 & new_n5524_;
  assign po317 = pi328 & new_n5524_;
  assign po316 = pi327 & new_n5524_;
  assign po315 = pi326 & new_n5524_;
  assign po314 = pi325 & new_n5524_;
  assign po313 = pi324 & new_n5524_;
  assign po312 = pi323 & new_n5524_;
  assign po311 = pi322 & new_n5524_;
  assign po310 = pi321 & new_n5524_;
  assign po309 = pi320 & new_n5524_;
  assign po308 = pi319 & new_n5524_;
  assign po307 = pi318 & new_n5524_;
  assign po306 = pi317 & new_n5524_;
  assign po305 = pi316 & new_n5524_;
  assign po304 = pi315 & new_n5524_;
  assign po303 = pi314 & new_n5524_;
  assign po302 = pi313 & new_n5524_;
  assign po301 = pi312 & new_n5524_;
  assign po298 = ~new_n5706_ | ~new_n5707_ | ~new_n5708_;
  assign po297 = ~new_n5703_ | ~new_n5704_ | ~new_n5705_;
  assign po296 = ~new_n5700_ | ~new_n5701_ | ~new_n5702_;
  assign po295 = ~new_n5697_ | ~new_n5698_ | ~new_n5699_;
  assign po294 = ~new_n5694_ | ~new_n5695_ | ~new_n5696_;
  assign po293 = ~new_n5691_ | ~new_n5692_ | ~new_n5693_;
  assign po292 = ~new_n5688_ | ~new_n5689_ | ~new_n5690_;
  assign po291 = ~new_n5685_ | ~new_n5686_ | ~new_n5687_;
  assign po290 = ~new_n5682_ | ~new_n5683_ | ~new_n5684_;
  assign po289 = ~new_n5679_ | ~new_n5680_ | ~new_n5681_;
  assign po288 = ~new_n5676_ | ~new_n5677_ | ~new_n5678_;
  assign po287 = ~new_n5673_ | ~new_n5674_ | ~new_n5675_;
  assign po286 = ~new_n5670_ | ~new_n5671_ | ~new_n5672_;
  assign po285 = ~new_n5667_ | ~new_n5668_ | ~new_n5669_;
  assign po284 = ~new_n5664_ | ~new_n5665_ | ~new_n5666_;
  assign po283 = ~new_n5661_ | ~new_n5662_ | ~new_n5663_;
  assign po282 = ~new_n5658_ | ~new_n5659_ | ~new_n5660_;
  assign po281 = ~new_n5655_ | ~new_n5656_ | ~new_n5657_;
  assign po280 = ~new_n5652_ | ~new_n5653_ | ~new_n5654_;
  assign po279 = ~new_n5649_ | ~new_n5650_ | ~new_n5651_;
  assign po278 = ~new_n5646_ | ~new_n5647_ | ~new_n5648_;
  assign po277 = ~new_n5643_ | ~new_n5644_ | ~new_n5645_;
  assign po276 = ~new_n5640_ | ~new_n5641_ | ~new_n5642_;
  assign po275 = ~new_n5637_ | ~new_n5638_ | ~new_n5639_;
  assign po274 = ~new_n5634_ | ~new_n5635_ | ~new_n5636_;
  assign po273 = ~new_n5631_ | ~new_n5632_ | ~new_n5633_;
  assign po272 = ~new_n5628_ | ~new_n5629_ | ~new_n5630_;
  assign po271 = ~new_n5625_ | ~new_n5626_ | ~new_n5627_;
  assign po270 = ~new_n5622_ | ~new_n5623_ | ~new_n5624_;
  assign po269 = ~new_n5619_ | ~new_n5620_ | ~new_n5621_;
  assign po268 = ~new_n5616_ | ~new_n5617_ | ~new_n5618_;
  assign po267 = ~new_n5613_ | ~new_n5614_ | ~new_n5615_;
  assign new_n4975_ = ~pi520 | ~new_n5523_;
  assign new_n4976_ = ~pi490;
  assign new_n4977_ = ~new_n5051_ | ~new_n7308_;
  assign new_n4978_ = ~new_n5051_ | ~new_n5709_;
  assign new_n4979_ = ~new_n4666_ | ~new_n5057_;
  assign new_n4980_ = ~new_n5056_ | ~new_n7327_ | ~new_n5055_;
  assign new_n4981_ = ~new_n7330_ | ~new_n7327_;
  assign new_n4982_ = ~new_n5610_ | ~new_n5057_;
  assign new_n4983_ = ~new_n5577_ | ~new_n7333_;
  assign new_n4984_ = ~new_n7324_ | ~new_n7327_;
  assign new_n4985_ = ~new_n5567_ | ~new_n5056_;
  assign new_n4986_ = ~new_n7324_ | ~new_n7333_;
  assign new_n4987_ = ~new_n5056_ | ~new_n5057_;
  assign new_n4988_ = ~new_n7333_ | ~new_n7327_ | ~new_n5055_;
  assign new_n4989_ = ~new_n5232_ | ~new_n5233_ | ~new_n5755_ | ~new_n5754_ | ~new_n5753_;
  assign new_n4990_ = ~new_n5250_ | ~new_n5248_ | ~new_n5769_ | ~new_n5768_;
  assign new_n4991_ = ~new_n5254_ | ~new_n5252_ | ~new_n5788_ | ~new_n5787_;
  assign new_n4992_ = ~new_n5258_ | ~new_n5256_ | ~new_n5807_ | ~new_n5806_;
  assign new_n4993_ = ~new_n5262_ | ~new_n5260_ | ~new_n5826_ | ~new_n5825_;
  assign new_n4994_ = ~new_n5266_ | ~new_n5264_ | ~new_n5845_ | ~new_n5844_;
  assign new_n4995_ = ~new_n5270_ | ~new_n5268_ | ~new_n5864_ | ~new_n5863_;
  assign new_n4996_ = ~new_n5274_ | ~new_n5272_ | ~new_n5883_ | ~new_n5882_;
  assign new_n4997_ = ~new_n5278_ | ~new_n5276_ | ~new_n5902_ | ~new_n5901_;
  assign new_n4998_ = ~new_n5282_ | ~new_n5280_ | ~new_n5921_ | ~new_n5920_;
  assign new_n4999_ = ~new_n5286_ | ~new_n5284_ | ~new_n5940_ | ~new_n5939_;
  assign new_n5000_ = ~new_n5290_ | ~new_n5288_ | ~new_n5959_ | ~new_n5958_;
  assign new_n5001_ = ~new_n5294_ | ~new_n5292_ | ~new_n5978_ | ~new_n5977_;
  assign new_n5002_ = ~new_n5298_ | ~new_n5296_ | ~new_n5997_ | ~new_n5996_;
  assign new_n5003_ = ~new_n5302_ | ~new_n5300_ | ~new_n6016_ | ~new_n6015_;
  assign new_n5004_ = ~new_n5306_ | ~new_n5304_ | ~new_n6035_ | ~new_n6034_;
  assign new_n5005_ = ~new_n5310_ | ~new_n5308_ | ~new_n6054_ | ~new_n6053_;
  assign new_n5006_ = ~new_n5314_ | ~new_n5312_ | ~new_n6073_ | ~new_n6072_;
  assign new_n5007_ = ~new_n5318_ | ~new_n5316_ | ~new_n6092_ | ~new_n6091_;
  assign new_n5008_ = ~new_n5322_ | ~new_n5320_ | ~new_n6111_ | ~new_n6110_;
  assign new_n5009_ = ~new_n1058_ | ~new_n5525_;
  assign new_n5010_ = ~new_n5326_ | ~new_n5324_ | ~new_n6130_ | ~new_n6129_;
  assign new_n5011_ = ~new_n1057_ | ~new_n5525_;
  assign new_n5012_ = ~new_n5330_ | ~new_n5328_ | ~new_n6149_ | ~new_n6148_;
  assign new_n5013_ = ~new_n1056_ | ~new_n5525_;
  assign new_n5014_ = ~new_n5334_ | ~new_n5332_ | ~new_n6168_ | ~new_n6167_;
  assign new_n5015_ = ~new_n1055_ | ~new_n5525_;
  assign new_n5016_ = ~new_n5338_ | ~new_n5336_ | ~new_n6187_ | ~new_n6186_;
  assign new_n5017_ = ~new_n1054_ | ~new_n5525_;
  assign new_n5018_ = ~new_n5342_ | ~new_n5340_ | ~new_n6206_ | ~new_n6205_;
  assign new_n5019_ = ~new_n1053_ | ~new_n5525_;
  assign new_n5020_ = ~new_n5346_ | ~new_n5344_ | ~new_n6225_ | ~new_n6224_;
  assign new_n5021_ = ~new_n1052_ | ~new_n5525_;
  assign new_n5022_ = ~new_n5350_ | ~new_n5348_ | ~new_n6244_ | ~new_n6243_;
  assign new_n5023_ = ~new_n1051_ | ~new_n5525_;
  assign new_n5024_ = ~new_n5354_ | ~new_n5352_ | ~new_n6263_ | ~new_n6262_;
  assign new_n5025_ = ~new_n1050_ | ~new_n5525_;
  assign new_n5026_ = ~new_n5357_ | ~new_n6284_ | ~new_n6283_ | ~new_n6282_ | ~new_n6281_;
  assign new_n5027_ = ~new_n1049_ | ~new_n5525_;
  assign new_n5028_ = ~new_n5362_ | ~new_n5360_ | ~new_n6303_ | ~new_n6302_ | ~new_n6301_;
  assign new_n5029_ = ~new_n1047_ | ~new_n5525_;
  assign new_n5030_ = ~new_n1046_ | ~new_n5525_;
  assign new_n5031_ = ~new_n5061_ | ~new_n7333_;
  assign new_n5032_ = ~new_n7290_ | ~new_n7330_;
  assign new_n5033_ = ~new_n4643_ | ~new_n6327_;
  assign new_n5034_ = ~new_n5576_ | ~new_n7324_;
  assign new_n5035_ = ~new_n4647_ | ~new_n7327_;
  assign new_n5036_ = ~new_n5049_ | ~new_n5050_ | ~new_n5051_;
  assign new_n5037_ = ~new_n4987_ | ~new_n5525_;
  assign new_n5038_ = ~new_n5597_ | ~new_n7317_;
  assign new_n5039_ = ~new_n5611_ | ~pi520;
  assign new_n5040_ = ~new_n5426_ | ~new_n4668_;
  assign new_n5041_ = ~new_n4633_ | ~new_n4638_;
  assign new_n5042_ = ~new_n4643_ | ~new_n6329_;
  assign new_n5043_ = ~new_n5503_ | ~new_n4636_;
  assign new_n5044_ = ~new_n7324_ | ~new_n5056_;
  assign new_n5045_ = ~new_n4633_ | ~new_n4643_;
  assign new_n5046_ = ~new_n6800_ | ~new_n5505_;
  assign new_n5047_ = ~new_n5567_ | ~new_n4985_;
  assign new_n5048_ = ~new_n5609_ | ~new_n5061_;
  assign new_n5049_ = ~new_n7304_ | ~new_n7303_;
  assign new_n5050_ = ~new_n7307_ | ~new_n7306_;
  assign new_n5051_ = ~new_n7310_ | ~new_n7309_;
  assign new_n5052_ = ~new_n7316_ | ~new_n7315_;
  assign po299 = ~new_n7319_ | ~new_n7318_;
  assign po300 = ~new_n7321_ | ~new_n7320_;
  assign new_n5055_ = ~new_n7329_ | ~new_n7328_;
  assign new_n5056_ = ~new_n7332_ | ~new_n7331_;
  assign new_n5057_ = ~new_n7323_ | ~new_n7322_;
  assign new_n5058_ = ~new_n7338_ | ~new_n7337_;
  assign new_n5059_ = ~new_n7335_ | ~new_n7334_;
  assign new_n5060_ = ~new_n7343_ | ~new_n7342_;
  assign new_n5061_ = ~new_n7326_ | ~new_n7325_;
  assign new_n5062_ = ~new_n7346_ | ~new_n7345_;
  assign new_n5063_ = ~new_n7348_ | ~new_n7347_;
  assign new_n5064_ = ~new_n7351_ | ~new_n7350_;
  assign new_n5065_ = ~new_n7359_ | ~new_n7358_;
  assign new_n5066_ = ~new_n7356_ | ~new_n7355_;
  assign po331 = ~new_n7362_ | ~new_n7361_;
  assign new_n5068_ = ~new_n7366_ | ~new_n7365_;
  assign new_n5069_ = ~new_n7368_ | ~new_n7367_;
  assign po332 = ~new_n7373_ | ~new_n7372_;
  assign new_n5071_ = ~new_n7375_ | ~new_n7374_;
  assign new_n5072_ = ~new_n7377_ | ~new_n7376_;
  assign po333 = ~new_n7380_ | ~new_n7379_;
  assign new_n5074_ = ~new_n7382_ | ~new_n7381_;
  assign new_n5075_ = ~new_n7384_ | ~new_n7383_;
  assign po334 = ~new_n7387_ | ~new_n7386_;
  assign new_n5077_ = ~new_n7389_ | ~new_n7388_;
  assign new_n5078_ = ~new_n7391_ | ~new_n7390_;
  assign po335 = ~new_n7394_ | ~new_n7393_;
  assign new_n5080_ = ~new_n7396_ | ~new_n7395_;
  assign new_n5081_ = ~new_n7398_ | ~new_n7397_;
  assign po336 = ~new_n7401_ | ~new_n7400_;
  assign new_n5083_ = ~new_n7403_ | ~new_n7402_;
  assign new_n5084_ = ~new_n7405_ | ~new_n7404_;
  assign po337 = ~new_n7408_ | ~new_n7407_;
  assign new_n5086_ = ~new_n7410_ | ~new_n7409_;
  assign new_n5087_ = ~new_n7412_ | ~new_n7411_;
  assign po338 = ~new_n7415_ | ~new_n7414_;
  assign new_n5089_ = ~new_n7417_ | ~new_n7416_;
  assign new_n5090_ = ~new_n7419_ | ~new_n7418_;
  assign po339 = ~new_n7422_ | ~new_n7421_;
  assign new_n5092_ = ~new_n7424_ | ~new_n7423_;
  assign new_n5093_ = ~new_n7426_ | ~new_n7425_;
  assign po340 = ~new_n7429_ | ~new_n7428_;
  assign new_n5095_ = ~new_n7431_ | ~new_n7430_;
  assign new_n5096_ = ~new_n7433_ | ~new_n7432_;
  assign po341 = ~new_n7436_ | ~new_n7435_;
  assign new_n5098_ = ~new_n7438_ | ~new_n7437_;
  assign new_n5099_ = ~new_n7440_ | ~new_n7439_;
  assign po342 = ~new_n7443_ | ~new_n7442_;
  assign new_n5101_ = ~new_n7445_ | ~new_n7444_;
  assign new_n5102_ = ~new_n7447_ | ~new_n7446_;
  assign po343 = ~new_n7450_ | ~new_n7449_;
  assign new_n5104_ = ~new_n7452_ | ~new_n7451_;
  assign new_n5105_ = ~new_n7454_ | ~new_n7453_;
  assign po344 = ~new_n7457_ | ~new_n7456_;
  assign new_n5107_ = ~new_n7459_ | ~new_n7458_;
  assign new_n5108_ = ~new_n7461_ | ~new_n7460_;
  assign po345 = ~new_n7464_ | ~new_n7463_;
  assign new_n5110_ = ~new_n7466_ | ~new_n7465_;
  assign new_n5111_ = ~new_n7468_ | ~new_n7467_;
  assign po346 = ~new_n7471_ | ~new_n7470_;
  assign new_n5113_ = ~new_n7473_ | ~new_n7472_;
  assign new_n5114_ = ~new_n7475_ | ~new_n7474_;
  assign po347 = ~new_n7478_ | ~new_n7477_;
  assign new_n5116_ = ~new_n7480_ | ~new_n7479_;
  assign new_n5117_ = ~new_n7482_ | ~new_n7481_;
  assign po348 = ~new_n7485_ | ~new_n7484_;
  assign new_n5119_ = ~new_n7487_ | ~new_n7486_;
  assign new_n5120_ = ~new_n7489_ | ~new_n7488_;
  assign po349 = ~new_n7492_ | ~new_n7491_;
  assign new_n5122_ = ~new_n7494_ | ~new_n7493_;
  assign po350 = ~new_n7497_ | ~new_n7496_;
  assign po351 = ~new_n7499_ | ~new_n7498_;
  assign po352 = ~new_n7501_ | ~new_n7500_;
  assign po353 = ~new_n7503_ | ~new_n7502_;
  assign po354 = ~new_n7505_ | ~new_n7504_;
  assign po355 = ~new_n7507_ | ~new_n7506_;
  assign po356 = ~new_n7509_ | ~new_n7508_;
  assign po357 = ~new_n7511_ | ~new_n7510_;
  assign po358 = ~new_n7513_ | ~new_n7512_;
  assign po359 = ~new_n7515_ | ~new_n7514_;
  assign po360 = ~new_n7517_ | ~new_n7516_;
  assign po361 = ~new_n7519_ | ~new_n7518_;
  assign po362 = ~new_n7521_ | ~new_n7520_;
  assign po363 = ~new_n7523_ | ~new_n7522_;
  assign po364 = ~new_n7525_ | ~new_n7524_;
  assign po365 = ~new_n7527_ | ~new_n7526_;
  assign po366 = ~new_n7529_ | ~new_n7528_;
  assign po367 = ~new_n7531_ | ~new_n7530_;
  assign po368 = ~new_n7533_ | ~new_n7532_;
  assign po369 = ~new_n7535_ | ~new_n7534_;
  assign po370 = ~new_n7537_ | ~new_n7536_;
  assign po371 = ~new_n7539_ | ~new_n7538_;
  assign po372 = ~new_n7541_ | ~new_n7540_;
  assign po373 = ~new_n7543_ | ~new_n7542_;
  assign po374 = ~new_n7545_ | ~new_n7544_;
  assign po375 = ~new_n7547_ | ~new_n7546_;
  assign po376 = ~new_n7549_ | ~new_n7548_;
  assign po377 = ~new_n7551_ | ~new_n7550_;
  assign po378 = ~new_n7553_ | ~new_n7552_;
  assign po379 = ~new_n7555_ | ~new_n7554_;
  assign po380 = ~new_n7557_ | ~new_n7556_;
  assign po381 = ~new_n7559_ | ~new_n7558_;
  assign po382 = ~new_n7561_ | ~new_n7560_;
  assign po383 = ~new_n7563_ | ~new_n7562_;
  assign po384 = ~new_n7565_ | ~new_n7564_;
  assign po385 = ~new_n7567_ | ~new_n7566_;
  assign po386 = ~new_n7569_ | ~new_n7568_;
  assign po387 = ~new_n7571_ | ~new_n7570_;
  assign po388 = ~new_n7573_ | ~new_n7572_;
  assign po389 = ~new_n7575_ | ~new_n7574_;
  assign po390 = ~new_n7577_ | ~new_n7576_;
  assign po391 = ~new_n7579_ | ~new_n7578_;
  assign po392 = ~new_n7581_ | ~new_n7580_;
  assign po393 = ~new_n7583_ | ~new_n7582_;
  assign po394 = ~new_n7585_ | ~new_n7584_;
  assign po447 = ~new_n7651_ | ~new_n7650_;
  assign po448 = ~new_n7653_ | ~new_n7652_;
  assign po449 = ~new_n7655_ | ~new_n7654_;
  assign po450 = ~new_n7657_ | ~new_n7656_;
  assign po451 = ~new_n7659_ | ~new_n7658_;
  assign po452 = ~new_n7661_ | ~new_n7660_;
  assign po453 = ~new_n7663_ | ~new_n7662_;
  assign po454 = ~new_n7665_ | ~new_n7664_;
  assign po455 = ~new_n7667_ | ~new_n7666_;
  assign po456 = ~new_n7669_ | ~new_n7668_;
  assign po457 = ~new_n7671_ | ~new_n7670_;
  assign po458 = ~new_n7673_ | ~new_n7672_;
  assign po459 = ~new_n7675_ | ~new_n7674_;
  assign po460 = ~new_n7677_ | ~new_n7676_;
  assign po461 = ~new_n7679_ | ~new_n7678_;
  assign po462 = ~new_n7681_ | ~new_n7680_;
  assign po463 = ~new_n7683_ | ~new_n7682_;
  assign po464 = ~new_n7685_ | ~new_n7684_;
  assign po465 = ~new_n7687_ | ~new_n7686_;
  assign po466 = ~new_n7689_ | ~new_n7688_;
  assign po467 = ~new_n7691_ | ~new_n7690_;
  assign po468 = ~new_n7693_ | ~new_n7692_;
  assign po469 = ~new_n7695_ | ~new_n7694_;
  assign po470 = ~new_n7697_ | ~new_n7696_;
  assign po471 = ~new_n7699_ | ~new_n7698_;
  assign po472 = ~new_n7701_ | ~new_n7700_;
  assign po473 = ~new_n7703_ | ~new_n7702_;
  assign po474 = ~new_n7705_ | ~new_n7704_;
  assign po475 = ~new_n7707_ | ~new_n7706_;
  assign po476 = ~new_n7709_ | ~new_n7708_;
  assign po477 = ~new_n7711_ | ~new_n7710_;
  assign po478 = ~new_n7713_ | ~new_n7712_;
  assign new_n5200_ = ~new_n7819_ | ~new_n7818_;
  assign new_n5201_ = ~new_n7821_ | ~new_n7820_;
  assign new_n5202_ = ~new_n7823_ | ~new_n7822_;
  assign new_n5203_ = ~new_n7825_ | ~new_n7824_;
  assign new_n5204_ = ~new_n7827_ | ~new_n7826_;
  assign new_n5205_ = ~new_n7829_ | ~new_n7828_;
  assign new_n5206_ = ~new_n7831_ | ~new_n7830_;
  assign new_n5207_ = ~new_n7833_ | ~new_n7832_;
  assign new_n5208_ = ~new_n7835_ | ~new_n7834_;
  assign new_n5209_ = ~new_n7837_ | ~new_n7836_;
  assign new_n5210_ = ~new_n7840_ | ~new_n7839_;
  assign new_n5211_ = ~new_n7842_ | ~new_n7841_;
  assign new_n5212_ = ~new_n7844_ | ~new_n7843_;
  assign new_n5213_ = ~new_n7846_ | ~new_n7845_;
  assign new_n5214_ = ~new_n7848_ | ~new_n7847_;
  assign new_n5215_ = ~new_n7850_ | ~new_n7849_;
  assign new_n5216_ = ~new_n7852_ | ~new_n7851_;
  assign new_n5217_ = ~new_n7854_ | ~new_n7853_;
  assign new_n5218_ = ~new_n7856_ | ~new_n7855_;
  assign new_n5219_ = ~new_n7858_ | ~new_n7857_;
  assign new_n5220_ = ~new_n7860_ | ~new_n7859_;
  assign new_n5221_ = ~new_n7863_ | ~new_n7862_;
  assign new_n5222_ = ~new_n7865_ | ~new_n7864_;
  assign new_n5223_ = ~new_n7867_ | ~new_n7866_;
  assign new_n5224_ = ~new_n7869_ | ~new_n7868_;
  assign new_n5225_ = ~new_n7871_ | ~new_n7870_;
  assign new_n5226_ = ~new_n7873_ | ~new_n7872_;
  assign new_n5227_ = ~new_n7875_ | ~new_n7874_;
  assign new_n5228_ = ~new_n7877_ | ~new_n7876_;
  assign new_n5229_ = ~new_n7879_ | ~new_n7878_;
  assign new_n5230_ = ~new_n7881_ | ~new_n7880_;
  assign new_n5231_ = ~new_n7883_ | ~new_n7882_;
  assign new_n5232_ = new_n5750_ & new_n5749_;
  assign new_n5233_ = new_n5752_ & new_n5751_;
  assign new_n5234_ = new_n5759_ & new_n5757_;
  assign new_n5235_ = new_n5234_ & new_n5760_ & new_n5758_;
  assign new_n5236_ = new_n5713_ & new_n5714_ & new_n5716_ & new_n5715_;
  assign new_n5237_ = new_n5717_ & new_n5718_ & new_n5720_ & new_n5719_;
  assign new_n5238_ = new_n5721_ & new_n5722_ & new_n5724_ & new_n5723_;
  assign new_n5239_ = new_n5727_ & new_n5726_ & new_n5725_;
  assign new_n5240_ = new_n5236_ & new_n5237_ & new_n5239_ & new_n5238_;
  assign new_n5241_ = new_n5728_ & new_n5729_ & new_n5731_ & new_n5730_;
  assign new_n5242_ = new_n5732_ & new_n5733_ & new_n5735_ & new_n5734_;
  assign new_n5243_ = new_n5736_ & new_n5737_ & new_n5739_ & new_n5738_;
  assign new_n5244_ = new_n5742_ & new_n5741_ & new_n5740_;
  assign new_n5245_ = new_n5241_ & new_n5242_ & new_n5244_ & new_n5243_;
  assign new_n5246_ = new_n7357_ & new_n5743_;
  assign new_n5247_ = new_n7360_ & new_n4643_;
  assign new_n5248_ = new_n5771_ & new_n5770_;
  assign new_n5249_ = new_n5773_ & new_n5772_;
  assign new_n5250_ = new_n5249_ & new_n5775_ & new_n5774_;
  assign new_n5251_ = new_n5779_ & new_n5780_ & new_n5778_ & new_n5777_;
  assign new_n5252_ = new_n5790_ & new_n5789_;
  assign new_n5253_ = new_n5792_ & new_n5791_;
  assign new_n5254_ = new_n5253_ & new_n5794_ & new_n5793_;
  assign new_n5255_ = new_n5798_ & new_n5799_ & new_n5797_ & new_n5796_;
  assign new_n5256_ = new_n5809_ & new_n5808_;
  assign new_n5257_ = new_n5811_ & new_n5810_;
  assign new_n5258_ = new_n5257_ & new_n5813_ & new_n5812_;
  assign new_n5259_ = new_n5817_ & new_n5818_ & new_n5816_ & new_n5815_;
  assign new_n5260_ = new_n5828_ & new_n5827_;
  assign new_n5261_ = new_n5830_ & new_n5829_;
  assign new_n5262_ = new_n5261_ & new_n5832_ & new_n5831_;
  assign new_n5263_ = new_n5836_ & new_n5837_ & new_n5835_ & new_n5834_;
  assign new_n5264_ = new_n5847_ & new_n5846_;
  assign new_n5265_ = new_n5849_ & new_n5848_;
  assign new_n5266_ = new_n5265_ & new_n5851_ & new_n5850_;
  assign new_n5267_ = new_n5855_ & new_n5856_ & new_n5854_ & new_n5853_;
  assign new_n5268_ = new_n5866_ & new_n5865_;
  assign new_n5269_ = new_n5868_ & new_n5867_;
  assign new_n5270_ = new_n5269_ & new_n5870_ & new_n5869_;
  assign new_n5271_ = new_n5874_ & new_n5875_ & new_n5873_ & new_n5872_;
  assign new_n5272_ = new_n5885_ & new_n5884_;
  assign new_n5273_ = new_n5887_ & new_n5886_;
  assign new_n5274_ = new_n5273_ & new_n5889_ & new_n5888_;
  assign new_n5275_ = new_n5893_ & new_n5894_ & new_n5892_ & new_n5891_;
  assign new_n5276_ = new_n5904_ & new_n5903_;
  assign new_n5277_ = new_n5906_ & new_n5905_;
  assign new_n5278_ = new_n5277_ & new_n5908_ & new_n5907_;
  assign new_n5279_ = new_n5912_ & new_n5913_ & new_n5911_ & new_n5910_;
  assign new_n5280_ = new_n5923_ & new_n5922_;
  assign new_n5281_ = new_n5925_ & new_n5924_;
  assign new_n5282_ = new_n5281_ & new_n5927_ & new_n5926_;
  assign new_n5283_ = new_n5931_ & new_n5932_ & new_n5930_ & new_n5929_;
  assign new_n5284_ = new_n5942_ & new_n5941_;
  assign new_n5285_ = new_n5944_ & new_n5943_;
  assign new_n5286_ = new_n5285_ & new_n5946_ & new_n5945_;
  assign new_n5287_ = new_n5950_ & new_n5951_ & new_n5949_ & new_n5948_;
  assign new_n5288_ = new_n5961_ & new_n5960_;
  assign new_n5289_ = new_n5963_ & new_n5962_;
  assign new_n5290_ = new_n5289_ & new_n5965_ & new_n5964_;
  assign new_n5291_ = new_n5969_ & new_n5970_ & new_n5968_ & new_n5967_;
  assign new_n5292_ = new_n5980_ & new_n5979_;
  assign new_n5293_ = new_n5982_ & new_n5981_;
  assign new_n5294_ = new_n5293_ & new_n5984_ & new_n5983_;
  assign new_n5295_ = new_n5988_ & new_n5989_ & new_n5987_ & new_n5986_;
  assign new_n5296_ = new_n5999_ & new_n5998_;
  assign new_n5297_ = new_n6001_ & new_n6000_;
  assign new_n5298_ = new_n5297_ & new_n6003_ & new_n6002_;
  assign new_n5299_ = new_n6007_ & new_n6008_ & new_n6006_ & new_n6005_;
  assign new_n5300_ = new_n6018_ & new_n6017_;
  assign new_n5301_ = new_n6020_ & new_n6019_;
  assign new_n5302_ = new_n5301_ & new_n6022_ & new_n6021_;
  assign new_n5303_ = new_n6026_ & new_n6027_ & new_n6025_ & new_n6024_;
  assign new_n5304_ = new_n6037_ & new_n6036_;
  assign new_n5305_ = new_n6039_ & new_n6038_;
  assign new_n5306_ = new_n5305_ & new_n6041_ & new_n6040_;
  assign new_n5307_ = new_n6045_ & new_n6046_ & new_n6044_ & new_n6043_;
  assign new_n5308_ = new_n6056_ & new_n6055_;
  assign new_n5309_ = new_n6058_ & new_n6057_;
  assign new_n5310_ = new_n5309_ & new_n6060_ & new_n6059_;
  assign new_n5311_ = new_n6064_ & new_n6065_ & new_n6063_ & new_n6062_;
  assign new_n5312_ = new_n6075_ & new_n6074_;
  assign new_n5313_ = new_n6077_ & new_n6076_;
  assign new_n5314_ = new_n5313_ & new_n6079_ & new_n6078_;
  assign new_n5315_ = new_n6083_ & new_n6084_ & new_n6082_ & new_n6081_;
  assign new_n5316_ = new_n6094_ & new_n6093_;
  assign new_n5317_ = new_n6096_ & new_n6095_;
  assign new_n5318_ = new_n5317_ & new_n6098_ & new_n6097_;
  assign new_n5319_ = new_n6102_ & new_n6103_ & new_n6101_ & new_n6100_;
  assign new_n5320_ = new_n6113_ & new_n6112_;
  assign new_n5321_ = new_n6115_ & new_n6114_;
  assign new_n5322_ = new_n5321_ & new_n6117_ & new_n6116_;
  assign new_n5323_ = new_n6121_ & new_n6122_ & new_n6120_ & new_n6119_;
  assign new_n5324_ = new_n6132_ & new_n6131_;
  assign new_n5325_ = new_n6134_ & new_n6133_;
  assign new_n5326_ = new_n5325_ & new_n6136_ & new_n6135_;
  assign new_n5327_ = new_n6140_ & new_n6141_ & new_n6139_ & new_n6138_;
  assign new_n5328_ = new_n6151_ & new_n6150_;
  assign new_n5329_ = new_n6153_ & new_n6152_;
  assign new_n5330_ = new_n5329_ & new_n6155_ & new_n6154_;
  assign new_n5331_ = new_n6159_ & new_n6160_ & new_n6158_ & new_n6157_;
  assign new_n5332_ = new_n6170_ & new_n6169_;
  assign new_n5333_ = new_n6172_ & new_n6171_;
  assign new_n5334_ = new_n5333_ & new_n6174_ & new_n6173_;
  assign new_n5335_ = new_n6178_ & new_n6179_ & new_n6177_ & new_n6176_;
  assign new_n5336_ = new_n6189_ & new_n6188_;
  assign new_n5337_ = new_n6191_ & new_n6190_;
  assign new_n5338_ = new_n5337_ & new_n6193_ & new_n6192_;
  assign new_n5339_ = new_n6197_ & new_n6198_ & new_n6196_ & new_n6195_;
  assign new_n5340_ = new_n6208_ & new_n6207_;
  assign new_n5341_ = new_n6210_ & new_n6209_;
  assign new_n5342_ = new_n5341_ & new_n6212_ & new_n6211_;
  assign new_n5343_ = new_n6216_ & new_n6217_ & new_n6215_ & new_n6214_;
  assign new_n5344_ = new_n6227_ & new_n6226_;
  assign new_n5345_ = new_n6229_ & new_n6228_;
  assign new_n5346_ = new_n5345_ & new_n6231_ & new_n6230_;
  assign new_n5347_ = new_n6235_ & new_n6236_ & new_n6234_ & new_n6233_;
  assign new_n5348_ = new_n6246_ & new_n6245_;
  assign new_n5349_ = new_n6248_ & new_n6247_;
  assign new_n5350_ = new_n5349_ & new_n6250_ & new_n6249_;
  assign new_n5351_ = new_n6254_ & new_n6255_ & new_n6253_ & new_n6252_;
  assign new_n5352_ = new_n6265_ & new_n6264_;
  assign new_n5353_ = new_n6267_ & new_n6266_;
  assign new_n5354_ = new_n5353_ & new_n6269_ & new_n6268_;
  assign new_n5355_ = new_n6273_ & new_n6274_ & new_n6272_ & new_n6271_;
  assign new_n5356_ = new_n6286_ & new_n6285_;
  assign new_n5357_ = new_n5356_ & new_n6288_ & new_n6287_;
  assign new_n5358_ = new_n6292_ & new_n6293_ & new_n6291_ & new_n6290_;
  assign new_n5359_ = new_n6300_ & new_n5598_;
  assign new_n5360_ = new_n6305_ & new_n6304_;
  assign new_n5361_ = new_n6307_ & new_n6306_;
  assign new_n5362_ = new_n5361_ & new_n6309_ & new_n6308_;
  assign new_n5363_ = new_n6312_ & new_n6313_ & new_n6311_;
  assign new_n5364_ = new_n5598_ & new_n6300_;
  assign new_n5365_ = new_n4643_ & new_n5065_;
  assign new_n5366_ = new_n5066_ & new_n7360_ & new_n4667_;
  assign new_n5367_ = new_n5056_ & new_n5061_ & new_n7330_;
  assign new_n5368_ = new_n6332_ & new_n6331_ & new_n6330_;
  assign new_n5369_ = new_n5528_ & new_n6334_ & new_n6333_;
  assign new_n5370_ = new_n6337_ & new_n6336_ & new_n6335_;
  assign new_n5371_ = new_n5529_ & new_n6339_ & new_n6338_;
  assign new_n5372_ = new_n6342_ & new_n6341_ & new_n6340_;
  assign new_n5373_ = new_n5530_ & new_n6344_ & new_n6343_;
  assign new_n5374_ = new_n6347_ & new_n6346_ & new_n6345_;
  assign new_n5375_ = new_n5531_ & new_n6349_ & new_n6348_;
  assign new_n5376_ = new_n6352_ & new_n6351_ & new_n6350_;
  assign new_n5377_ = new_n5532_ & new_n6354_ & new_n6353_;
  assign new_n5378_ = new_n6357_ & new_n6356_ & new_n6355_;
  assign new_n5379_ = new_n6359_ & new_n6358_;
  assign new_n5380_ = new_n6362_ & new_n6361_ & new_n6360_;
  assign new_n5381_ = new_n6364_ & new_n6363_;
  assign new_n5382_ = new_n6367_ & new_n6366_ & new_n6365_;
  assign new_n5383_ = new_n6369_ & new_n6368_;
  assign new_n5384_ = new_n6372_ & new_n6371_ & new_n6370_;
  assign new_n5385_ = new_n6374_ & new_n6373_;
  assign new_n5386_ = new_n6377_ & new_n6376_ & new_n6375_;
  assign new_n5387_ = new_n6379_ & new_n6378_;
  assign new_n5388_ = new_n6382_ & new_n6380_;
  assign new_n5389_ = new_n6384_ & new_n6383_;
  assign new_n5390_ = new_n6387_ & new_n6386_ & new_n6385_;
  assign new_n5391_ = new_n6389_ & new_n6388_;
  assign new_n5392_ = new_n6392_ & new_n6390_;
  assign new_n5393_ = new_n6394_ & new_n6393_;
  assign new_n5394_ = new_n6397_ & new_n6395_;
  assign new_n5395_ = new_n6399_ & new_n6398_;
  assign new_n5396_ = new_n6402_ & new_n6400_;
  assign new_n5397_ = new_n6404_ & new_n6403_;
  assign new_n5398_ = new_n6407_ & new_n6405_;
  assign new_n5399_ = new_n6409_ & new_n6408_;
  assign new_n5400_ = new_n6412_ & new_n6410_;
  assign new_n5401_ = new_n6414_ & new_n6413_;
  assign new_n5402_ = new_n6417_ & new_n6415_;
  assign new_n5403_ = new_n6419_ & new_n6418_;
  assign new_n5404_ = new_n6422_ & new_n6420_;
  assign new_n5405_ = new_n6424_ & new_n6423_;
  assign new_n5406_ = new_n6427_ & new_n6425_;
  assign new_n5407_ = new_n6429_ & new_n6428_;
  assign new_n5408_ = new_n6432_ & new_n6430_;
  assign new_n5409_ = new_n6434_ & new_n6433_;
  assign new_n5410_ = new_n6437_ & new_n6435_;
  assign new_n5411_ = new_n6439_ & new_n6438_;
  assign new_n5412_ = new_n6442_ & new_n6440_;
  assign new_n5413_ = new_n6444_ & new_n6443_;
  assign new_n5414_ = new_n6447_ & new_n6445_;
  assign new_n5415_ = new_n6449_ & new_n6448_;
  assign new_n5416_ = new_n6452_ & new_n6450_;
  assign new_n5417_ = new_n6454_ & new_n6453_;
  assign new_n5418_ = new_n6457_ & new_n6455_;
  assign new_n5419_ = new_n6459_ & new_n6458_;
  assign new_n5420_ = new_n6462_ & new_n6460_;
  assign new_n5421_ = new_n6464_ & new_n6463_;
  assign new_n5422_ = new_n6467_ & new_n6465_;
  assign new_n5423_ = new_n6469_ & new_n6468_;
  assign new_n5424_ = new_n6472_ & new_n6470_;
  assign new_n5425_ = new_n6474_ & new_n6473_;
  assign new_n5426_ = new_n7302_ & new_n5037_;
  assign new_n5427_ = new_n5052_ & pi520;
  assign new_n5428_ = new_n6493_ & new_n6492_;
  assign new_n5429_ = new_n6495_ & new_n6494_;
  assign new_n5430_ = new_n6497_ & new_n6498_ & new_n6496_;
  assign new_n5431_ = new_n6508_ & new_n6507_;
  assign new_n5432_ = new_n6510_ & new_n6509_;
  assign new_n5433_ = new_n6512_ & new_n6513_ & new_n6511_;
  assign new_n5434_ = new_n6523_ & new_n6522_;
  assign new_n5435_ = new_n6525_ & new_n6524_;
  assign new_n5436_ = new_n6527_ & new_n6528_ & new_n6526_;
  assign new_n5437_ = new_n6538_ & new_n6537_;
  assign new_n5438_ = new_n6540_ & new_n6539_;
  assign new_n5439_ = new_n6542_ & new_n6543_ & new_n6541_;
  assign new_n5440_ = new_n6553_ & new_n6552_;
  assign new_n5441_ = new_n6555_ & new_n6554_;
  assign new_n5442_ = new_n6557_ & new_n6558_ & new_n6556_;
  assign new_n5443_ = new_n6568_ & new_n6567_;
  assign new_n5444_ = new_n6570_ & new_n6569_;
  assign new_n5445_ = new_n6572_ & new_n6573_ & new_n6571_;
  assign new_n5446_ = new_n6583_ & new_n6582_;
  assign new_n5447_ = new_n6585_ & new_n6584_;
  assign new_n5448_ = new_n6587_ & new_n6588_ & new_n6586_;
  assign new_n5449_ = new_n6598_ & new_n6597_;
  assign new_n5450_ = new_n6600_ & new_n6599_;
  assign new_n5451_ = new_n6602_ & new_n6603_ & new_n6601_;
  assign new_n5452_ = new_n6613_ & new_n6612_;
  assign new_n5453_ = new_n6615_ & new_n6614_;
  assign new_n5454_ = new_n6617_ & new_n6618_ & new_n6616_;
  assign new_n5455_ = new_n6628_ & new_n6627_;
  assign new_n5456_ = new_n6630_ & new_n6629_;
  assign new_n5457_ = new_n6632_ & new_n6633_ & new_n6631_;
  assign new_n5458_ = new_n6643_ & new_n6642_;
  assign new_n5459_ = new_n6645_ & new_n6644_;
  assign new_n5460_ = new_n6647_ & new_n6648_ & new_n6646_;
  assign new_n5461_ = new_n6658_ & new_n6657_;
  assign new_n5462_ = new_n5461_ & new_n6660_ & new_n6659_;
  assign new_n5463_ = new_n6663_ & new_n6662_ & new_n6661_;
  assign new_n5464_ = new_n6673_ & new_n6672_;
  assign new_n5465_ = new_n5464_ & new_n6675_ & new_n6674_;
  assign new_n5466_ = new_n6678_ & new_n6677_ & new_n6676_;
  assign new_n5467_ = new_n6688_ & new_n6687_;
  assign new_n5468_ = new_n5467_ & new_n6690_ & new_n6689_;
  assign new_n5469_ = new_n6693_ & new_n6692_ & new_n6691_;
  assign new_n5470_ = new_n6703_ & new_n6702_;
  assign new_n5471_ = new_n5470_ & new_n6705_ & new_n6704_;
  assign new_n5472_ = new_n6708_ & new_n6707_ & new_n6706_;
  assign new_n5473_ = new_n6718_ & new_n6717_;
  assign new_n5474_ = new_n5473_ & new_n6720_ & new_n6719_;
  assign new_n5475_ = new_n6723_ & new_n6722_ & new_n6721_;
  assign new_n5476_ = new_n6733_ & new_n6732_;
  assign new_n5477_ = new_n5476_ & new_n6735_ & new_n6734_;
  assign new_n5478_ = new_n6738_ & new_n6737_ & new_n6736_;
  assign new_n5479_ = new_n6748_ & new_n6747_;
  assign new_n5480_ = new_n5479_ & new_n6750_ & new_n6749_;
  assign new_n5481_ = new_n6753_ & new_n6752_ & new_n6751_;
  assign new_n5482_ = new_n6763_ & new_n6762_;
  assign new_n5483_ = new_n5482_ & new_n6765_ & new_n6764_;
  assign new_n5484_ = new_n6768_ & new_n6767_ & new_n6766_;
  assign new_n5485_ = new_n6770_ & new_n6771_;
  assign new_n5486_ = new_n6778_ & new_n6777_;
  assign new_n5487_ = new_n5486_ & new_n6780_ & new_n6779_;
  assign new_n5488_ = new_n6783_ & new_n6782_ & new_n6781_;
  assign new_n5489_ = new_n7776_ & new_n7773_ & new_n7770_;
  assign new_n5490_ = new_n5489_ & new_n5491_;
  assign new_n5491_ = new_n7758_ & new_n7761_ & new_n7767_ & new_n7764_;
  assign new_n5492_ = new_n7788_ & new_n7785_ & new_n7782_;
  assign new_n5493_ = new_n7797_ & new_n7794_ & new_n7791_;
  assign new_n5494_ = new_n7779_ & new_n5493_ & new_n5492_;
  assign new_n5495_ = new_n7722_ & new_n7725_ & new_n7728_ & new_n5500_ & new_n5499_;
  assign new_n5496_ = new_n7815_ & new_n7803_ & new_n7806_ & new_n7812_ & new_n7809_;
  assign new_n5497_ = new_n5496_ & new_n7800_ & new_n7755_ & new_n5494_ & new_n5490_;
  assign new_n5498_ = new_n7749_ & new_n5495_;
  assign new_n5499_ = new_n7731_ & new_n7734_ & new_n7740_ & new_n7737_;
  assign new_n5500_ = new_n7746_ & new_n7743_;
  assign new_n5501_ = new_n6788_ & new_n6789_ & new_n6793_;
  assign new_n5502_ = new_n7286_ & new_n6792_;
  assign new_n5503_ = new_n5065_ & new_n5066_;
  assign new_n5504_ = new_n5048_ & new_n5568_;
  assign new_n5505_ = new_n5038_ & new_n7317_ & new_n4667_;
  assign new_n5506_ = new_n4643_ & new_n6799_;
  assign new_n5507_ = new_n5508_ & new_n6842_;
  assign new_n5508_ = new_n6846_ & new_n6845_;
  assign new_n5509_ = new_n5604_ & new_n4694_;
  assign new_n5510_ = new_n6887_ & new_n6886_;
  assign new_n5511_ = new_n6890_ & new_n6889_;
  assign new_n5512_ = new_n6908_ & new_n6907_;
  assign new_n5513_ = new_n6935_ & new_n6934_;
  assign new_n5514_ = new_n5515_ & new_n6976_;
  assign new_n5515_ = new_n6980_ & new_n6979_;
  assign new_n5516_ = new_n7007_ & new_n7003_;
  assign new_n5517_ = new_n5518_ & new_n7012_;
  assign new_n5518_ = new_n7016_ & new_n7015_;
  assign new_n5519_ = new_n7063_ & pi520;
  assign new_n5520_ = new_n7333_ & new_n5031_;
  assign new_n5521_ = new_n7327_ & new_n7317_;
  assign new_n5522_ = new_n5056_ & new_n7128_;
  assign new_n5523_ = ~pi309;
  assign new_n5524_ = ~new_n4643_ | ~new_n4978_;
  assign new_n5525_ = ~new_n7349_ | ~new_n7344_;
  assign new_n5526_ = ~new_n5247_ | ~new_n4665_;
  assign new_n5527_ = ~new_n5365_ | ~new_n4665_;
  assign new_n5528_ = new_n7587_ & new_n7586_;
  assign new_n5529_ = new_n7589_ & new_n7588_;
  assign new_n5530_ = new_n7591_ & new_n7590_;
  assign new_n5531_ = new_n7593_ & new_n7592_;
  assign new_n5532_ = new_n7595_ & new_n7594_;
  assign new_n5533_ = new_n7597_ & new_n7596_;
  assign new_n5534_ = new_n7599_ & new_n7598_;
  assign new_n5535_ = new_n7601_ & new_n7600_;
  assign new_n5536_ = new_n7603_ & new_n7602_;
  assign new_n5537_ = new_n7605_ & new_n7604_;
  assign new_n5538_ = new_n7607_ & new_n7606_;
  assign new_n5539_ = new_n7609_ & new_n7608_;
  assign new_n5540_ = new_n7611_ & new_n7610_;
  assign new_n5541_ = new_n7613_ & new_n7612_;
  assign new_n5542_ = new_n7615_ & new_n7614_;
  assign new_n5543_ = new_n7617_ & new_n7616_;
  assign new_n5544_ = new_n7619_ & new_n7618_;
  assign new_n5545_ = new_n7621_ & new_n7620_;
  assign new_n5546_ = new_n7623_ & new_n7622_;
  assign new_n5547_ = new_n7625_ & new_n7624_;
  assign new_n5548_ = new_n7627_ & new_n7626_;
  assign new_n5549_ = new_n7629_ & new_n7628_;
  assign new_n5550_ = new_n7631_ & new_n7630_;
  assign new_n5551_ = new_n7633_ & new_n7632_;
  assign new_n5552_ = new_n7635_ & new_n7634_;
  assign new_n5553_ = new_n7637_ & new_n7636_;
  assign new_n5554_ = new_n7639_ & new_n7638_;
  assign new_n5555_ = new_n7641_ & new_n7640_;
  assign new_n5556_ = new_n7643_ & new_n7642_;
  assign new_n5557_ = new_n7645_ & new_n7644_;
  assign new_n5558_ = ~new_n5364_ | ~new_n4672_;
  assign new_n5559_ = new_n7647_ & new_n7646_;
  assign new_n5560_ = new_n7649_ & new_n7648_;
  assign new_n5561_ = ~new_n15484_;
  assign new_n5562_ = new_n7719_ & new_n7718_;
  assign new_n5563_ = ~new_n5498_ | ~new_n5497_ | ~new_n7752_;
  assign new_n5564_ = ~new_n15467_;
  assign new_n5565_ = ~new_n4986_;
  assign new_n5566_ = ~new_n5598_ | ~new_n5061_;
  assign new_n5567_ = ~new_n4984_;
  assign new_n5568_ = ~new_n7290_ | ~new_n5057_;
  assign new_n5569_ = ~new_n5048_;
  assign new_n5570_ = ~new_n4985_;
  assign new_n5571_ = ~new_n4979_;
  assign new_n5572_ = ~new_n5035_;
  assign new_n5573_ = ~new_n5034_;
  assign new_n5574_ = ~new_n5578_ | ~new_n7324_;
  assign new_n5575_ = ~new_n4983_;
  assign new_n5576_ = ~new_n5032_;
  assign new_n5577_ = ~new_n4982_;
  assign new_n5578_ = ~new_n4988_;
  assign new_n5579_ = ~new_n4980_;
  assign new_n5580_ = ~new_n5525_;
  assign new_n5581_ = ~new_n5043_;
  assign po511 = ~new_n5039_;
  assign new_n5583_ = ~new_n5037_;
  assign new_n5584_ = ~new_n5025_;
  assign new_n5585_ = ~new_n5023_;
  assign new_n5586_ = ~new_n5021_;
  assign new_n5587_ = ~new_n5019_;
  assign new_n5588_ = ~new_n5017_;
  assign new_n5589_ = ~new_n5015_;
  assign new_n5590_ = ~new_n5013_;
  assign new_n5591_ = ~new_n5011_;
  assign new_n5592_ = ~new_n5009_;
  assign new_n5593_ = ~new_n5030_;
  assign new_n5594_ = ~new_n5029_;
  assign new_n5595_ = ~new_n5027_;
  assign new_n5596_ = ~new_n5041_;
  assign new_n5597_ = ~new_n5036_;
  assign new_n5598_ = ~new_n4987_;
  assign new_n5599_ = ~new_n5033_;
  assign new_n5600_ = ~new_n5527_;
  assign new_n5601_ = ~new_n5526_;
  assign new_n5602_ = ~new_n5524_;
  assign new_n5603_ = ~new_n5558_;
  assign new_n5604_ = ~new_n5045_;
  assign new_n5605_ = ~new_n5046_ | ~pi520;
  assign new_n5606_ = ~new_n5573_ | ~new_n4643_;
  assign new_n5607_ = ~new_n5042_;
  assign new_n5608_ = ~new_n4977_;
  assign new_n5609_ = ~new_n5044_;
  assign new_n5610_ = ~new_n4981_;
  assign new_n5611_ = ~new_n5038_;
  assign new_n5612_ = ~new_n4975_;
  assign new_n5613_ = ~new_n1070_ | ~po509;
  assign new_n5614_ = ~pi278 | ~new_n4649_;
  assign new_n5615_ = ~pi278 | ~new_n5612_;
  assign new_n5616_ = ~new_n1059_ | ~po509;
  assign new_n5617_ = ~new_n15342_ | ~new_n4649_;
  assign new_n5618_ = ~pi279 | ~new_n5612_;
  assign new_n5619_ = ~new_n1048_ | ~po509;
  assign new_n5620_ = ~new_n15317_ | ~new_n4649_;
  assign new_n5621_ = ~pi280 | ~new_n5612_;
  assign new_n5622_ = ~new_n1045_ | ~po509;
  assign new_n5623_ = ~new_n15318_ | ~new_n4649_;
  assign new_n5624_ = ~pi281 | ~new_n5612_;
  assign new_n5625_ = ~new_n1044_ | ~po509;
  assign new_n5626_ = ~new_n15319_ | ~new_n4649_;
  assign new_n5627_ = ~pi282 | ~new_n5612_;
  assign new_n5628_ = ~new_n1043_ | ~po509;
  assign new_n5629_ = ~new_n15367_ | ~new_n4649_;
  assign new_n5630_ = ~pi283 | ~new_n5612_;
  assign new_n5631_ = ~new_n1042_ | ~po509;
  assign new_n5632_ = ~new_n15320_ | ~new_n4649_;
  assign new_n5633_ = ~pi284 | ~new_n5612_;
  assign new_n5634_ = ~new_n1041_ | ~po509;
  assign new_n5635_ = ~new_n15321_ | ~new_n4649_;
  assign new_n5636_ = ~pi285 | ~new_n5612_;
  assign new_n5637_ = ~new_n1040_ | ~po509;
  assign new_n5638_ = ~new_n15322_ | ~new_n4649_;
  assign new_n5639_ = ~pi286 | ~new_n5612_;
  assign new_n5640_ = ~new_n1039_ | ~po509;
  assign new_n5641_ = ~new_n15365_ | ~new_n4649_;
  assign new_n5642_ = ~pi287 | ~new_n5612_;
  assign new_n5643_ = ~new_n1069_ | ~po509;
  assign new_n5644_ = ~new_n15304_ | ~new_n4649_;
  assign new_n5645_ = ~pi288 | ~new_n5612_;
  assign new_n5646_ = ~new_n1068_ | ~po509;
  assign new_n5647_ = ~new_n15305_ | ~new_n4649_;
  assign new_n5648_ = ~pi289 | ~new_n5612_;
  assign new_n5649_ = ~new_n1067_ | ~po509;
  assign new_n5650_ = ~new_n15306_ | ~new_n4649_;
  assign new_n5651_ = ~pi290 | ~new_n5612_;
  assign new_n5652_ = ~new_n1066_ | ~po509;
  assign new_n5653_ = ~new_n15392_ | ~new_n4649_;
  assign new_n5654_ = ~pi291 | ~new_n5612_;
  assign new_n5655_ = ~new_n1065_ | ~po509;
  assign new_n5656_ = ~new_n15307_ | ~new_n4649_;
  assign new_n5657_ = ~pi292 | ~new_n5612_;
  assign new_n5658_ = ~new_n1064_ | ~po509;
  assign new_n5659_ = ~new_n15308_ | ~new_n4649_;
  assign new_n5660_ = ~pi293 | ~new_n5612_;
  assign new_n5661_ = ~new_n1063_ | ~po509;
  assign new_n5662_ = ~new_n15309_ | ~new_n4649_;
  assign new_n5663_ = ~pi294 | ~new_n5612_;
  assign new_n5664_ = ~new_n1062_ | ~po509;
  assign new_n5665_ = ~new_n15390_ | ~new_n4649_;
  assign new_n5666_ = ~pi295 | ~new_n5612_;
  assign new_n5667_ = ~new_n1061_ | ~po509;
  assign new_n5668_ = ~new_n15310_ | ~new_n4649_;
  assign new_n5669_ = ~pi296 | ~new_n5612_;
  assign new_n5670_ = ~new_n1060_ | ~po509;
  assign new_n5671_ = ~new_n15311_ | ~new_n4649_;
  assign new_n5672_ = ~pi297 | ~new_n5612_;
  assign new_n5673_ = ~new_n1058_ | ~po509;
  assign new_n5674_ = ~new_n15312_ | ~new_n4649_;
  assign new_n5675_ = ~pi298 | ~new_n5612_;
  assign new_n5676_ = ~new_n1057_ | ~po509;
  assign new_n5677_ = ~new_n15385_ | ~new_n4649_;
  assign new_n5678_ = ~pi299 | ~new_n5612_;
  assign new_n5679_ = ~new_n1056_ | ~po509;
  assign new_n5680_ = ~new_n15313_ | ~new_n4649_;
  assign new_n5681_ = ~pi300 | ~new_n5612_;
  assign new_n5682_ = ~new_n1055_ | ~po509;
  assign new_n5683_ = ~new_n15314_ | ~new_n4649_;
  assign new_n5684_ = ~pi301 | ~new_n5612_;
  assign new_n5685_ = ~new_n1054_ | ~po509;
  assign new_n5686_ = ~new_n15383_ | ~new_n4649_;
  assign new_n5687_ = ~pi302 | ~new_n5612_;
  assign new_n5688_ = ~new_n1053_ | ~po509;
  assign new_n5689_ = ~new_n15315_ | ~new_n4649_;
  assign new_n5690_ = ~pi303 | ~new_n5612_;
  assign new_n5691_ = ~new_n1052_ | ~po509;
  assign new_n5692_ = ~new_n15316_ | ~new_n4649_;
  assign new_n5693_ = ~pi304 | ~new_n5612_;
  assign new_n5694_ = ~new_n1051_ | ~po509;
  assign new_n5695_ = ~new_n15380_ | ~new_n4649_;
  assign new_n5696_ = ~pi305 | ~new_n5612_;
  assign new_n5697_ = ~new_n1050_ | ~po509;
  assign new_n5698_ = ~new_n15377_ | ~new_n4649_;
  assign new_n5699_ = ~pi306 | ~new_n5612_;
  assign new_n5700_ = ~new_n1049_ | ~po509;
  assign new_n5701_ = ~new_n15374_ | ~new_n4649_;
  assign new_n5702_ = ~pi307 | ~new_n5612_;
  assign new_n5703_ = ~new_n1047_ | ~po509;
  assign new_n5704_ = ~new_n15372_ | ~new_n4649_;
  assign new_n5705_ = ~pi308 | ~new_n5612_;
  assign new_n5706_ = ~new_n1046_ | ~po509;
  assign new_n5707_ = ~new_n15370_ | ~new_n4649_;
  assign new_n5708_ = ~pi309 | ~new_n5612_;
  assign new_n5709_ = ~new_n5608_ | ~new_n7314_;
  assign new_n5710_ = ~new_n4978_;
  assign new_n5711_ = ~new_n4977_ | ~new_n7305_;
  assign new_n5712_ = ~new_n4977_ | ~new_n7308_;
  assign new_n5713_ = ~new_n5710_ | ~pi320;
  assign new_n5714_ = ~new_n5710_ | ~pi321;
  assign new_n5715_ = ~new_n5710_ | ~pi322;
  assign new_n5716_ = ~new_n5710_ | ~pi323;
  assign new_n5717_ = ~new_n5710_ | ~pi324;
  assign new_n5718_ = ~new_n5710_ | ~pi325;
  assign new_n5719_ = ~new_n5710_ | ~pi326;
  assign new_n5720_ = ~new_n5710_ | ~pi327;
  assign new_n5721_ = ~new_n5710_ | ~pi328;
  assign new_n5722_ = ~new_n5710_ | ~pi329;
  assign new_n5723_ = ~new_n5710_ | ~pi330;
  assign new_n5724_ = ~new_n5710_ | ~pi331;
  assign new_n5725_ = ~new_n5710_ | ~pi332;
  assign new_n5726_ = ~new_n5710_ | ~pi333;
  assign new_n5727_ = ~new_n5710_ | ~pi334;
  assign new_n5728_ = ~new_n5710_ | ~pi335;
  assign new_n5729_ = ~new_n5710_ | ~pi336;
  assign new_n5730_ = ~new_n5710_ | ~pi337;
  assign new_n5731_ = ~new_n5710_ | ~pi338;
  assign new_n5732_ = ~new_n5710_ | ~pi339;
  assign new_n5733_ = ~new_n5710_ | ~pi312;
  assign new_n5734_ = ~new_n5710_ | ~pi340;
  assign new_n5735_ = ~new_n5710_ | ~pi341;
  assign new_n5736_ = ~new_n5710_ | ~pi313;
  assign new_n5737_ = ~new_n5710_ | ~pi314;
  assign new_n5738_ = ~new_n5710_ | ~pi315;
  assign new_n5739_ = ~new_n5710_ | ~pi316;
  assign new_n5740_ = ~new_n5710_ | ~pi317;
  assign new_n5741_ = ~new_n5710_ | ~pi318;
  assign new_n5742_ = ~new_n5710_ | ~pi319;
  assign new_n5743_ = ~new_n7353_ | ~new_n7354_ | ~new_n4981_ | ~new_n5044_;
  assign new_n5744_ = ~new_n4641_ | ~pi375;
  assign new_n5745_ = ~new_n4642_ | ~pi343;
  assign new_n5746_ = ~new_n4694_;
  assign new_n5747_ = ~new_n5565_ | ~new_n5061_;
  assign new_n5748_ = ~new_n5574_ | ~new_n5747_;
  assign new_n5749_ = ~new_n5571_ | ~new_n19719_;
  assign new_n5750_ = ~new_n4631_ | ~new_n20663_;
  assign new_n5751_ = ~new_n4630_ | ~new_n19296_;
  assign new_n5752_ = ~new_n4634_ | ~new_n16644_;
  assign new_n5753_ = ~new_n5579_ | ~new_n20191_;
  assign new_n5754_ = ~new_n5575_ | ~new_n17695_;
  assign new_n5755_ = ~new_n4632_ | ~new_n18196_;
  assign new_n5756_ = ~new_n4989_;
  assign new_n5757_ = ~new_n5064_ | ~new_n4647_;
  assign new_n5758_ = ~new_n4646_ | ~new_n4694_;
  assign new_n5759_ = ~new_n17194_ | ~new_n4644_;
  assign new_n5760_ = ~new_n5064_ | ~new_n5748_;
  assign new_n5761_ = ~new_n5235_ | ~new_n5756_;
  assign new_n5762_ = ~pi376 | ~new_n4641_;
  assign new_n5763_ = ~pi344 | ~new_n4642_;
  assign new_n5764_ = ~new_n4684_;
  assign new_n5765_ = ~pi374 | ~new_n4641_;
  assign new_n5766_ = ~pi342 | ~new_n4642_;
  assign new_n5767_ = ~new_n4693_;
  assign new_n5768_ = ~new_n4654_ | ~new_n4693_;
  assign new_n5769_ = ~new_n19794_ | ~new_n5571_;
  assign new_n5770_ = ~new_n20738_ | ~new_n4631_;
  assign new_n5771_ = ~new_n19295_ | ~new_n4630_;
  assign new_n5772_ = ~new_n16719_ | ~new_n4634_;
  assign new_n5773_ = ~new_n20266_ | ~new_n5579_;
  assign new_n5774_ = ~new_n17694_ | ~new_n5575_;
  assign new_n5775_ = ~new_n18195_ | ~new_n4632_;
  assign new_n5776_ = ~new_n4990_;
  assign new_n5777_ = ~new_n16337_ | ~new_n4647_;
  assign new_n5778_ = ~new_n4646_ | ~new_n4684_;
  assign new_n5779_ = ~new_n17193_ | ~new_n4644_;
  assign new_n5780_ = ~new_n5069_ | ~new_n5748_;
  assign new_n5781_ = ~new_n5251_ | ~new_n5776_;
  assign new_n5782_ = ~new_n4640_ | ~pi409;
  assign new_n5783_ = ~pi377 | ~new_n4641_;
  assign new_n5784_ = ~pi345 | ~new_n4642_;
  assign new_n5785_ = ~new_n14972_ | ~new_n4639_;
  assign new_n5786_ = ~new_n4680_;
  assign new_n5787_ = ~new_n4654_ | ~new_n4694_;
  assign new_n5788_ = ~new_n19804_ | ~new_n5571_;
  assign new_n5789_ = ~new_n20748_ | ~new_n4631_;
  assign new_n5790_ = ~new_n19217_ | ~new_n4630_;
  assign new_n5791_ = ~new_n16729_ | ~new_n4634_;
  assign new_n5792_ = ~new_n20276_ | ~new_n5579_;
  assign new_n5793_ = ~new_n17616_ | ~new_n5575_;
  assign new_n5794_ = ~new_n18117_ | ~new_n4632_;
  assign new_n5795_ = ~new_n4991_;
  assign new_n5796_ = ~new_n16300_ | ~new_n4647_;
  assign new_n5797_ = ~new_n4646_ | ~new_n4680_;
  assign new_n5798_ = ~new_n17115_ | ~new_n4644_;
  assign new_n5799_ = ~new_n5072_ | ~new_n5748_;
  assign new_n5800_ = ~new_n5255_ | ~new_n5795_;
  assign new_n5801_ = ~pi410 | ~new_n4640_;
  assign new_n5802_ = ~pi378 | ~new_n4641_;
  assign new_n5803_ = ~pi346 | ~new_n4642_;
  assign new_n5804_ = ~new_n15022_ | ~new_n4639_;
  assign new_n5805_ = ~new_n4676_;
  assign new_n5806_ = ~new_n4654_ | ~new_n4684_;
  assign new_n5807_ = ~new_n19716_ | ~new_n5571_;
  assign new_n5808_ = ~new_n20660_ | ~new_n4631_;
  assign new_n5809_ = ~new_n19301_ | ~new_n4630_;
  assign new_n5810_ = ~new_n16641_ | ~new_n4634_;
  assign new_n5811_ = ~new_n20188_ | ~new_n5579_;
  assign new_n5812_ = ~new_n17700_ | ~new_n5575_;
  assign new_n5813_ = ~new_n18201_ | ~new_n4632_;
  assign new_n5814_ = ~new_n4992_;
  assign new_n5815_ = ~new_n16302_ | ~new_n4647_;
  assign new_n5816_ = ~new_n4646_ | ~new_n4676_;
  assign new_n5817_ = ~new_n17199_ | ~new_n4644_;
  assign new_n5818_ = ~new_n5075_ | ~new_n5748_;
  assign new_n5819_ = ~new_n5259_ | ~new_n5814_;
  assign new_n5820_ = ~pi411 | ~new_n4640_;
  assign new_n5821_ = ~pi379 | ~new_n4641_;
  assign new_n5822_ = ~pi347 | ~new_n4642_;
  assign new_n5823_ = ~new_n15021_ | ~new_n4639_;
  assign new_n5824_ = ~new_n4683_;
  assign new_n5825_ = ~new_n4654_ | ~new_n4680_;
  assign new_n5826_ = ~new_n19803_ | ~new_n5571_;
  assign new_n5827_ = ~new_n20747_ | ~new_n4631_;
  assign new_n5828_ = ~new_n19300_ | ~new_n4630_;
  assign new_n5829_ = ~new_n16728_ | ~new_n4634_;
  assign new_n5830_ = ~new_n20275_ | ~new_n5579_;
  assign new_n5831_ = ~new_n17699_ | ~new_n5575_;
  assign new_n5832_ = ~new_n18200_ | ~new_n4632_;
  assign new_n5833_ = ~new_n4993_;
  assign new_n5834_ = ~new_n16303_ | ~new_n4647_;
  assign new_n5835_ = ~new_n4646_ | ~new_n4683_;
  assign new_n5836_ = ~new_n17198_ | ~new_n4644_;
  assign new_n5837_ = ~new_n5078_ | ~new_n5748_;
  assign new_n5838_ = ~new_n5263_ | ~new_n5833_;
  assign new_n5839_ = ~pi412 | ~new_n4640_;
  assign new_n5840_ = ~pi380 | ~new_n4641_;
  assign new_n5841_ = ~pi348 | ~new_n4642_;
  assign new_n5842_ = ~new_n15020_ | ~new_n4639_;
  assign new_n5843_ = ~new_n4687_;
  assign new_n5844_ = ~new_n4654_ | ~new_n4676_;
  assign new_n5845_ = ~new_n19802_ | ~new_n5571_;
  assign new_n5846_ = ~new_n20746_ | ~new_n4631_;
  assign new_n5847_ = ~new_n19218_ | ~new_n4630_;
  assign new_n5848_ = ~new_n16727_ | ~new_n4634_;
  assign new_n5849_ = ~new_n20274_ | ~new_n5579_;
  assign new_n5850_ = ~new_n17617_ | ~new_n5575_;
  assign new_n5851_ = ~new_n18118_ | ~new_n4632_;
  assign new_n5852_ = ~new_n4994_;
  assign new_n5853_ = ~new_n16347_ | ~new_n4647_;
  assign new_n5854_ = ~new_n4646_ | ~new_n4687_;
  assign new_n5855_ = ~new_n17116_ | ~new_n4644_;
  assign new_n5856_ = ~new_n5081_ | ~new_n5748_;
  assign new_n5857_ = ~new_n5267_ | ~new_n5852_;
  assign new_n5858_ = ~pi413 | ~new_n4640_;
  assign new_n5859_ = ~pi381 | ~new_n4641_;
  assign new_n5860_ = ~pi349 | ~new_n4642_;
  assign new_n5861_ = ~new_n15019_ | ~new_n4639_;
  assign new_n5862_ = ~new_n4686_;
  assign new_n5863_ = ~new_n4654_ | ~new_n4683_;
  assign new_n5864_ = ~new_n19717_ | ~new_n5571_;
  assign new_n5865_ = ~new_n20661_ | ~new_n4631_;
  assign new_n5866_ = ~new_n19299_ | ~new_n4630_;
  assign new_n5867_ = ~new_n16642_ | ~new_n4634_;
  assign new_n5868_ = ~new_n20189_ | ~new_n5579_;
  assign new_n5869_ = ~new_n17698_ | ~new_n5575_;
  assign new_n5870_ = ~new_n18199_ | ~new_n4632_;
  assign new_n5871_ = ~new_n4995_;
  assign new_n5872_ = ~new_n16304_ | ~new_n4647_;
  assign new_n5873_ = ~new_n4646_ | ~new_n4686_;
  assign new_n5874_ = ~new_n17197_ | ~new_n4644_;
  assign new_n5875_ = ~new_n5084_ | ~new_n5748_;
  assign new_n5876_ = ~new_n5271_ | ~new_n5871_;
  assign new_n5877_ = ~pi414 | ~new_n4640_;
  assign new_n5878_ = ~pi382 | ~new_n4641_;
  assign new_n5879_ = ~pi350 | ~new_n4642_;
  assign new_n5880_ = ~new_n15018_ | ~new_n4639_;
  assign new_n5881_ = ~new_n4700_;
  assign new_n5882_ = ~new_n4654_ | ~new_n4687_;
  assign new_n5883_ = ~new_n19801_ | ~new_n5571_;
  assign new_n5884_ = ~new_n20745_ | ~new_n4631_;
  assign new_n5885_ = ~new_n19219_ | ~new_n4630_;
  assign new_n5886_ = ~new_n16726_ | ~new_n4634_;
  assign new_n5887_ = ~new_n20273_ | ~new_n5579_;
  assign new_n5888_ = ~new_n17618_ | ~new_n5575_;
  assign new_n5889_ = ~new_n18119_ | ~new_n4632_;
  assign new_n5890_ = ~new_n4996_;
  assign new_n5891_ = ~new_n16305_ | ~new_n4647_;
  assign new_n5892_ = ~new_n4646_ | ~new_n4700_;
  assign new_n5893_ = ~new_n17117_ | ~new_n4644_;
  assign new_n5894_ = ~new_n5087_ | ~new_n5748_;
  assign new_n5895_ = ~new_n5275_ | ~new_n5890_;
  assign new_n5896_ = ~pi415 | ~new_n4640_;
  assign new_n5897_ = ~pi383 | ~new_n4641_;
  assign new_n5898_ = ~pi351 | ~new_n4642_;
  assign new_n5899_ = ~new_n15017_ | ~new_n4639_;
  assign new_n5900_ = ~new_n4699_;
  assign new_n5901_ = ~new_n4654_ | ~new_n4686_;
  assign new_n5902_ = ~new_n19718_ | ~new_n5571_;
  assign new_n5903_ = ~new_n20662_ | ~new_n4631_;
  assign new_n5904_ = ~new_n19298_ | ~new_n4630_;
  assign new_n5905_ = ~new_n16643_ | ~new_n4634_;
  assign new_n5906_ = ~new_n20190_ | ~new_n5579_;
  assign new_n5907_ = ~new_n17697_ | ~new_n5575_;
  assign new_n5908_ = ~new_n18198_ | ~new_n4632_;
  assign new_n5909_ = ~new_n4997_;
  assign new_n5910_ = ~new_n16306_ | ~new_n4647_;
  assign new_n5911_ = ~new_n4646_ | ~new_n4699_;
  assign new_n5912_ = ~new_n17196_ | ~new_n4644_;
  assign new_n5913_ = ~new_n5090_ | ~new_n5748_;
  assign new_n5914_ = ~new_n5279_ | ~new_n5909_;
  assign new_n5915_ = ~pi416 | ~new_n4640_;
  assign new_n5916_ = ~pi384 | ~new_n4641_;
  assign new_n5917_ = ~pi352 | ~new_n4642_;
  assign new_n5918_ = ~new_n15041_ | ~new_n4639_;
  assign new_n5919_ = ~new_n4678_;
  assign new_n5920_ = ~new_n4654_ | ~new_n4700_;
  assign new_n5921_ = ~new_n19800_ | ~new_n5571_;
  assign new_n5922_ = ~new_n20744_ | ~new_n4631_;
  assign new_n5923_ = ~new_n19297_ | ~new_n4630_;
  assign new_n5924_ = ~new_n16725_ | ~new_n4634_;
  assign new_n5925_ = ~new_n20272_ | ~new_n5579_;
  assign new_n5926_ = ~new_n17696_ | ~new_n5575_;
  assign new_n5927_ = ~new_n18197_ | ~new_n4632_;
  assign new_n5928_ = ~new_n4998_;
  assign new_n5929_ = ~new_n16345_ | ~new_n4647_;
  assign new_n5930_ = ~new_n4646_ | ~new_n4678_;
  assign new_n5931_ = ~new_n17195_ | ~new_n4644_;
  assign new_n5932_ = ~new_n5093_ | ~new_n5748_;
  assign new_n5933_ = ~new_n5283_ | ~new_n5928_;
  assign new_n5934_ = ~pi417 | ~new_n4640_;
  assign new_n5935_ = ~pi385 | ~new_n4641_;
  assign new_n5936_ = ~pi353 | ~new_n4642_;
  assign new_n5937_ = ~new_n15040_ | ~new_n4639_;
  assign new_n5938_ = ~new_n4679_;
  assign new_n5939_ = ~new_n4654_ | ~new_n4699_;
  assign new_n5940_ = ~new_n19810_ | ~new_n5571_;
  assign new_n5941_ = ~new_n20754_ | ~new_n4631_;
  assign new_n5942_ = ~new_n19211_ | ~new_n4630_;
  assign new_n5943_ = ~new_n16735_ | ~new_n4634_;
  assign new_n5944_ = ~new_n20282_ | ~new_n5579_;
  assign new_n5945_ = ~new_n17610_ | ~new_n5575_;
  assign new_n5946_ = ~new_n18111_ | ~new_n4632_;
  assign new_n5947_ = ~new_n4999_;
  assign new_n5948_ = ~new_n16288_ | ~new_n4647_;
  assign new_n5949_ = ~new_n4646_ | ~new_n4679_;
  assign new_n5950_ = ~new_n17109_ | ~new_n4644_;
  assign new_n5951_ = ~new_n5096_ | ~new_n5748_;
  assign new_n5952_ = ~new_n5287_ | ~new_n5947_;
  assign new_n5953_ = ~pi418 | ~new_n4640_;
  assign new_n5954_ = ~pi386 | ~new_n4641_;
  assign new_n5955_ = ~pi354 | ~new_n4642_;
  assign new_n5956_ = ~new_n15039_ | ~new_n4639_;
  assign new_n5957_ = ~new_n4688_;
  assign new_n5958_ = ~new_n4654_ | ~new_n4678_;
  assign new_n5959_ = ~new_n19711_ | ~new_n5571_;
  assign new_n5960_ = ~new_n20655_ | ~new_n4631_;
  assign new_n5961_ = ~new_n19315_ | ~new_n4630_;
  assign new_n5962_ = ~new_n16636_ | ~new_n4634_;
  assign new_n5963_ = ~new_n20183_ | ~new_n5579_;
  assign new_n5964_ = ~new_n17714_ | ~new_n5575_;
  assign new_n5965_ = ~new_n18215_ | ~new_n4632_;
  assign new_n5966_ = ~new_n5000_;
  assign new_n5967_ = ~new_n16289_ | ~new_n4647_;
  assign new_n5968_ = ~new_n4646_ | ~new_n4688_;
  assign new_n5969_ = ~new_n17213_ | ~new_n4644_;
  assign new_n5970_ = ~new_n5099_ | ~new_n5748_;
  assign new_n5971_ = ~new_n5291_ | ~new_n5966_;
  assign new_n5972_ = ~pi419 | ~new_n4640_;
  assign new_n5973_ = ~pi387 | ~new_n4641_;
  assign new_n5974_ = ~pi355 | ~new_n4642_;
  assign new_n5975_ = ~new_n15038_ | ~new_n4639_;
  assign new_n5976_ = ~new_n4696_;
  assign new_n5977_ = ~new_n4654_ | ~new_n4679_;
  assign new_n5978_ = ~new_n19799_ | ~new_n5571_;
  assign new_n5979_ = ~new_n20743_ | ~new_n4631_;
  assign new_n5980_ = ~new_n19314_ | ~new_n4630_;
  assign new_n5981_ = ~new_n16724_ | ~new_n4634_;
  assign new_n5982_ = ~new_n20271_ | ~new_n5579_;
  assign new_n5983_ = ~new_n17713_ | ~new_n5575_;
  assign new_n5984_ = ~new_n18214_ | ~new_n4632_;
  assign new_n5985_ = ~new_n5001_;
  assign new_n5986_ = ~new_n16290_ | ~new_n4647_;
  assign new_n5987_ = ~new_n4646_ | ~new_n4696_;
  assign new_n5988_ = ~new_n17212_ | ~new_n4644_;
  assign new_n5989_ = ~new_n5102_ | ~new_n5748_;
  assign new_n5990_ = ~new_n5295_ | ~new_n5985_;
  assign new_n5991_ = ~pi420 | ~new_n4640_;
  assign new_n5992_ = ~pi388 | ~new_n4641_;
  assign new_n5993_ = ~pi356 | ~new_n4642_;
  assign new_n5994_ = ~new_n15037_ | ~new_n4639_;
  assign new_n5995_ = ~new_n4695_;
  assign new_n5996_ = ~new_n4654_ | ~new_n4688_;
  assign new_n5997_ = ~new_n19798_ | ~new_n5571_;
  assign new_n5998_ = ~new_n20742_ | ~new_n4631_;
  assign new_n5999_ = ~new_n19212_ | ~new_n4630_;
  assign new_n6000_ = ~new_n16723_ | ~new_n4634_;
  assign new_n6001_ = ~new_n20270_ | ~new_n5579_;
  assign new_n6002_ = ~new_n17611_ | ~new_n5575_;
  assign new_n6003_ = ~new_n18112_ | ~new_n4632_;
  assign new_n6004_ = ~new_n5002_;
  assign new_n6005_ = ~new_n16368_ | ~new_n4647_;
  assign new_n6006_ = ~new_n4646_ | ~new_n4695_;
  assign new_n6007_ = ~new_n17110_ | ~new_n4644_;
  assign new_n6008_ = ~new_n5105_ | ~new_n5748_;
  assign new_n6009_ = ~new_n5299_ | ~new_n6004_;
  assign new_n6010_ = ~pi421 | ~new_n4640_;
  assign new_n6011_ = ~pi389 | ~new_n4641_;
  assign new_n6012_ = ~pi357 | ~new_n4642_;
  assign new_n6013_ = ~new_n15036_ | ~new_n4639_;
  assign new_n6014_ = ~new_n4690_;
  assign new_n6015_ = ~new_n4654_ | ~new_n4696_;
  assign new_n6016_ = ~new_n19809_ | ~new_n5571_;
  assign new_n6017_ = ~new_n20753_ | ~new_n4631_;
  assign new_n6018_ = ~new_n19313_ | ~new_n4630_;
  assign new_n6019_ = ~new_n16734_ | ~new_n4634_;
  assign new_n6020_ = ~new_n20281_ | ~new_n5579_;
  assign new_n6021_ = ~new_n17712_ | ~new_n5575_;
  assign new_n6022_ = ~new_n18213_ | ~new_n4632_;
  assign new_n6023_ = ~new_n5003_;
  assign new_n6024_ = ~new_n16291_ | ~new_n4647_;
  assign new_n6025_ = ~new_n4646_ | ~new_n4690_;
  assign new_n6026_ = ~new_n17211_ | ~new_n4644_;
  assign new_n6027_ = ~new_n5108_ | ~new_n5748_;
  assign new_n6028_ = ~new_n5303_ | ~new_n6023_;
  assign new_n6029_ = ~pi422 | ~new_n4640_;
  assign new_n6030_ = ~pi390 | ~new_n4641_;
  assign new_n6031_ = ~pi358 | ~new_n4642_;
  assign new_n6032_ = ~new_n15035_ | ~new_n4639_;
  assign new_n6033_ = ~new_n4689_;
  assign new_n6034_ = ~new_n4654_ | ~new_n4695_;
  assign new_n6035_ = ~new_n19808_ | ~new_n5571_;
  assign new_n6036_ = ~new_n20752_ | ~new_n4631_;
  assign new_n6037_ = ~new_n19312_ | ~new_n4630_;
  assign new_n6038_ = ~new_n16733_ | ~new_n4634_;
  assign new_n6039_ = ~new_n20280_ | ~new_n5579_;
  assign new_n6040_ = ~new_n17711_ | ~new_n5575_;
  assign new_n6041_ = ~new_n18212_ | ~new_n4632_;
  assign new_n6042_ = ~new_n5004_;
  assign new_n6043_ = ~new_n16292_ | ~new_n4647_;
  assign new_n6044_ = ~new_n4646_ | ~new_n4689_;
  assign new_n6045_ = ~new_n17210_ | ~new_n4644_;
  assign new_n6046_ = ~new_n5111_ | ~new_n5748_;
  assign new_n6047_ = ~new_n5307_ | ~new_n6042_;
  assign new_n6048_ = ~pi423 | ~new_n4640_;
  assign new_n6049_ = ~pi391 | ~new_n4641_;
  assign new_n6050_ = ~pi359 | ~new_n4642_;
  assign new_n6051_ = ~new_n15034_ | ~new_n4639_;
  assign new_n6052_ = ~new_n4685_;
  assign new_n6053_ = ~new_n4654_ | ~new_n4690_;
  assign new_n6054_ = ~new_n19712_ | ~new_n5571_;
  assign new_n6055_ = ~new_n20656_ | ~new_n4631_;
  assign new_n6056_ = ~new_n19311_ | ~new_n4630_;
  assign new_n6057_ = ~new_n16637_ | ~new_n4634_;
  assign new_n6058_ = ~new_n20184_ | ~new_n5579_;
  assign new_n6059_ = ~new_n17710_ | ~new_n5575_;
  assign new_n6060_ = ~new_n18211_ | ~new_n4632_;
  assign new_n6061_ = ~new_n5005_;
  assign new_n6062_ = ~new_n16293_ | ~new_n4647_;
  assign new_n6063_ = ~new_n4646_ | ~new_n4685_;
  assign new_n6064_ = ~new_n17209_ | ~new_n4644_;
  assign new_n6065_ = ~new_n5114_ | ~new_n5748_;
  assign new_n6066_ = ~new_n5311_ | ~new_n6061_;
  assign new_n6067_ = ~pi424 | ~new_n4640_;
  assign new_n6068_ = ~pi392 | ~new_n4641_;
  assign new_n6069_ = ~pi360 | ~new_n4642_;
  assign new_n6070_ = ~new_n15033_ | ~new_n4639_;
  assign new_n6071_ = ~new_n4698_;
  assign new_n6072_ = ~new_n4654_ | ~new_n4689_;
  assign new_n6073_ = ~new_n19797_ | ~new_n5571_;
  assign new_n6074_ = ~new_n20741_ | ~new_n4631_;
  assign new_n6075_ = ~new_n19213_ | ~new_n4630_;
  assign new_n6076_ = ~new_n16722_ | ~new_n4634_;
  assign new_n6077_ = ~new_n20269_ | ~new_n5579_;
  assign new_n6078_ = ~new_n17612_ | ~new_n5575_;
  assign new_n6079_ = ~new_n18113_ | ~new_n4632_;
  assign new_n6080_ = ~new_n5006_;
  assign new_n6081_ = ~new_n16366_ | ~new_n4647_;
  assign new_n6082_ = ~new_n4646_ | ~new_n4698_;
  assign new_n6083_ = ~new_n17111_ | ~new_n4644_;
  assign new_n6084_ = ~new_n5117_ | ~new_n5748_;
  assign new_n6085_ = ~new_n5315_ | ~new_n6080_;
  assign new_n6086_ = ~pi425 | ~new_n4640_;
  assign new_n6087_ = ~pi393 | ~new_n4641_;
  assign new_n6088_ = ~pi361 | ~new_n4642_;
  assign new_n6089_ = ~new_n15032_ | ~new_n4639_;
  assign new_n6090_ = ~new_n4697_;
  assign new_n6091_ = ~new_n4654_ | ~new_n4685_;
  assign new_n6092_ = ~new_n19796_ | ~new_n5571_;
  assign new_n6093_ = ~new_n20740_ | ~new_n4631_;
  assign new_n6094_ = ~new_n19310_ | ~new_n4630_;
  assign new_n6095_ = ~new_n16721_ | ~new_n4634_;
  assign new_n6096_ = ~new_n20268_ | ~new_n5579_;
  assign new_n6097_ = ~new_n17709_ | ~new_n5575_;
  assign new_n6098_ = ~new_n18210_ | ~new_n4632_;
  assign new_n6099_ = ~new_n5007_;
  assign new_n6100_ = ~new_n16294_ | ~new_n4647_;
  assign new_n6101_ = ~new_n4646_ | ~new_n4697_;
  assign new_n6102_ = ~new_n17208_ | ~new_n4644_;
  assign new_n6103_ = ~new_n5120_ | ~new_n5748_;
  assign new_n6104_ = ~new_n5319_ | ~new_n6099_;
  assign new_n6105_ = ~pi426 | ~new_n4640_;
  assign new_n6106_ = ~pi394 | ~new_n4641_;
  assign new_n6107_ = ~pi362 | ~new_n4642_;
  assign new_n6108_ = ~new_n15031_ | ~new_n4639_;
  assign new_n6109_ = ~new_n4692_;
  assign new_n6110_ = ~new_n4654_ | ~new_n4698_;
  assign new_n6111_ = ~new_n19795_ | ~new_n5571_;
  assign new_n6112_ = ~new_n20739_ | ~new_n4631_;
  assign new_n6113_ = ~new_n19309_ | ~new_n4630_;
  assign new_n6114_ = ~new_n16720_ | ~new_n4634_;
  assign new_n6115_ = ~new_n20267_ | ~new_n5579_;
  assign new_n6116_ = ~new_n17708_ | ~new_n5575_;
  assign new_n6117_ = ~new_n18209_ | ~new_n4632_;
  assign new_n6118_ = ~new_n5008_;
  assign new_n6119_ = ~new_n16364_ | ~new_n4647_;
  assign new_n6120_ = ~new_n4646_ | ~new_n4692_;
  assign new_n6121_ = ~new_n17207_ | ~new_n4644_;
  assign new_n6122_ = ~new_n5122_ | ~new_n5748_;
  assign new_n6123_ = ~new_n5323_ | ~new_n6118_;
  assign new_n6124_ = ~pi427 | ~new_n4640_;
  assign new_n6125_ = ~pi395 | ~new_n4641_;
  assign new_n6126_ = ~pi363 | ~new_n4642_;
  assign new_n6127_ = ~new_n15030_ | ~new_n4639_;
  assign new_n6128_ = ~new_n4691_;
  assign new_n6129_ = ~new_n4654_ | ~new_n4697_;
  assign new_n6130_ = ~new_n19793_ | ~new_n5571_;
  assign new_n6131_ = ~new_n20737_ | ~new_n4631_;
  assign new_n6132_ = ~new_n19214_ | ~new_n4630_;
  assign new_n6133_ = ~new_n16718_ | ~new_n4634_;
  assign new_n6134_ = ~new_n20265_ | ~new_n5579_;
  assign new_n6135_ = ~new_n17613_ | ~new_n5575_;
  assign new_n6136_ = ~new_n18114_ | ~new_n4632_;
  assign new_n6137_ = ~new_n5010_;
  assign new_n6138_ = ~new_n16295_ | ~new_n4647_;
  assign new_n6139_ = ~new_n4646_ | ~new_n4691_;
  assign new_n6140_ = ~new_n17112_ | ~new_n4644_;
  assign new_n6141_ = ~new_n5592_ | ~new_n5748_;
  assign new_n6142_ = ~new_n5327_ | ~new_n6137_;
  assign new_n6143_ = ~pi428 | ~new_n4640_;
  assign new_n6144_ = ~pi396 | ~new_n4641_;
  assign new_n6145_ = ~pi364 | ~new_n4642_;
  assign new_n6146_ = ~new_n15029_ | ~new_n4639_;
  assign new_n6147_ = ~new_n4677_;
  assign new_n6148_ = ~new_n4654_ | ~new_n4692_;
  assign new_n6149_ = ~new_n19807_ | ~new_n5571_;
  assign new_n6150_ = ~new_n20751_ | ~new_n4631_;
  assign new_n6151_ = ~new_n19215_ | ~new_n4630_;
  assign new_n6152_ = ~new_n16732_ | ~new_n4634_;
  assign new_n6153_ = ~new_n20279_ | ~new_n5579_;
  assign new_n6154_ = ~new_n17614_ | ~new_n5575_;
  assign new_n6155_ = ~new_n18115_ | ~new_n4632_;
  assign new_n6156_ = ~new_n5012_;
  assign new_n6157_ = ~new_n16360_ | ~new_n4647_;
  assign new_n6158_ = ~new_n4646_ | ~new_n4677_;
  assign new_n6159_ = ~new_n17113_ | ~new_n4644_;
  assign new_n6160_ = ~new_n5591_ | ~new_n5748_;
  assign new_n6161_ = ~new_n5331_ | ~new_n6156_;
  assign new_n6162_ = ~pi429 | ~new_n4640_;
  assign new_n6163_ = ~pi397 | ~new_n4641_;
  assign new_n6164_ = ~pi365 | ~new_n4642_;
  assign new_n6165_ = ~new_n15028_ | ~new_n4639_;
  assign new_n6166_ = ~new_n4682_;
  assign new_n6167_ = ~new_n4654_ | ~new_n4691_;
  assign new_n6168_ = ~new_n19806_ | ~new_n5571_;
  assign new_n6169_ = ~new_n20750_ | ~new_n4631_;
  assign new_n6170_ = ~new_n19308_ | ~new_n4630_;
  assign new_n6171_ = ~new_n16731_ | ~new_n4634_;
  assign new_n6172_ = ~new_n20278_ | ~new_n5579_;
  assign new_n6173_ = ~new_n17707_ | ~new_n5575_;
  assign new_n6174_ = ~new_n18208_ | ~new_n4632_;
  assign new_n6175_ = ~new_n5014_;
  assign new_n6176_ = ~new_n16296_ | ~new_n4647_;
  assign new_n6177_ = ~new_n4646_ | ~new_n4682_;
  assign new_n6178_ = ~new_n17206_ | ~new_n4644_;
  assign new_n6179_ = ~new_n5590_ | ~new_n5748_;
  assign new_n6180_ = ~new_n5335_ | ~new_n6175_;
  assign new_n6181_ = ~pi430 | ~new_n4640_;
  assign new_n6182_ = ~pi398 | ~new_n4641_;
  assign new_n6183_ = ~pi366 | ~new_n4642_;
  assign new_n6184_ = ~new_n15027_ | ~new_n4639_;
  assign new_n6185_ = ~new_n4681_;
  assign new_n6186_ = ~new_n4654_ | ~new_n4677_;
  assign new_n6187_ = ~new_n19713_ | ~new_n5571_;
  assign new_n6188_ = ~new_n20657_ | ~new_n4631_;
  assign new_n6189_ = ~new_n19307_ | ~new_n4630_;
  assign new_n6190_ = ~new_n16638_ | ~new_n4634_;
  assign new_n6191_ = ~new_n20185_ | ~new_n5579_;
  assign new_n6192_ = ~new_n17706_ | ~new_n5575_;
  assign new_n6193_ = ~new_n18207_ | ~new_n4632_;
  assign new_n6194_ = ~new_n5016_;
  assign new_n6195_ = ~new_n16358_ | ~new_n4647_;
  assign new_n6196_ = ~new_n4646_ | ~new_n4681_;
  assign new_n6197_ = ~new_n17205_ | ~new_n4644_;
  assign new_n6198_ = ~new_n5589_ | ~new_n5748_;
  assign new_n6199_ = ~new_n5339_ | ~new_n6194_;
  assign new_n6200_ = ~pi431 | ~new_n4640_;
  assign new_n6201_ = ~pi399 | ~new_n4641_;
  assign new_n6202_ = ~pi367 | ~new_n4642_;
  assign new_n6203_ = ~new_n15026_ | ~new_n4639_;
  assign new_n6204_ = ~new_n4674_;
  assign new_n6205_ = ~new_n4654_ | ~new_n4682_;
  assign new_n6206_ = ~new_n19792_ | ~new_n5571_;
  assign new_n6207_ = ~new_n20736_ | ~new_n4631_;
  assign new_n6208_ = ~new_n19306_ | ~new_n4630_;
  assign new_n6209_ = ~new_n16717_ | ~new_n4634_;
  assign new_n6210_ = ~new_n20264_ | ~new_n5579_;
  assign new_n6211_ = ~new_n17705_ | ~new_n5575_;
  assign new_n6212_ = ~new_n18206_ | ~new_n4632_;
  assign new_n6213_ = ~new_n5018_;
  assign new_n6214_ = ~new_n16297_ | ~new_n4647_;
  assign new_n6215_ = ~new_n4646_ | ~new_n4674_;
  assign new_n6216_ = ~new_n17204_ | ~new_n4644_;
  assign new_n6217_ = ~new_n5588_ | ~new_n5748_;
  assign new_n6218_ = ~new_n5343_ | ~new_n6213_;
  assign new_n6219_ = ~pi432 | ~new_n4640_;
  assign new_n6220_ = ~pi400 | ~new_n4641_;
  assign new_n6221_ = ~pi368 | ~new_n4642_;
  assign new_n6222_ = ~new_n15025_ | ~new_n4639_;
  assign new_n6223_ = ~new_n4673_;
  assign new_n6224_ = ~new_n4654_ | ~new_n4681_;
  assign new_n6225_ = ~new_n19791_ | ~new_n5571_;
  assign new_n6226_ = ~new_n20735_ | ~new_n4631_;
  assign new_n6227_ = ~new_n19305_ | ~new_n4630_;
  assign new_n6228_ = ~new_n16716_ | ~new_n4634_;
  assign new_n6229_ = ~new_n20263_ | ~new_n5579_;
  assign new_n6230_ = ~new_n17704_ | ~new_n5575_;
  assign new_n6231_ = ~new_n18205_ | ~new_n4632_;
  assign new_n6232_ = ~new_n5020_;
  assign new_n6233_ = ~new_n16356_ | ~new_n4647_;
  assign new_n6234_ = ~new_n4646_ | ~new_n4673_;
  assign new_n6235_ = ~new_n17203_ | ~new_n4644_;
  assign new_n6236_ = ~new_n5587_ | ~new_n5748_;
  assign new_n6237_ = ~new_n5347_ | ~new_n6232_;
  assign new_n6238_ = ~pi433 | ~new_n4640_;
  assign new_n6239_ = ~pi401 | ~new_n4641_;
  assign new_n6240_ = ~pi369 | ~new_n4642_;
  assign new_n6241_ = ~new_n15024_ | ~new_n4639_;
  assign new_n6242_ = ~new_n4669_;
  assign new_n6243_ = ~new_n4654_ | ~new_n4674_;
  assign new_n6244_ = ~new_n19805_ | ~new_n5571_;
  assign new_n6245_ = ~new_n20749_ | ~new_n4631_;
  assign new_n6246_ = ~new_n19216_ | ~new_n4630_;
  assign new_n6247_ = ~new_n16730_ | ~new_n4634_;
  assign new_n6248_ = ~new_n20277_ | ~new_n5579_;
  assign new_n6249_ = ~new_n17615_ | ~new_n5575_;
  assign new_n6250_ = ~new_n18116_ | ~new_n4632_;
  assign new_n6251_ = ~new_n5022_;
  assign new_n6252_ = ~new_n16298_ | ~new_n4647_;
  assign new_n6253_ = ~new_n4646_ | ~new_n4669_;
  assign new_n6254_ = ~new_n17114_ | ~new_n4644_;
  assign new_n6255_ = ~new_n5586_ | ~new_n5748_;
  assign new_n6256_ = ~new_n5351_ | ~new_n6251_;
  assign new_n6257_ = ~pi434 | ~new_n4640_;
  assign new_n6258_ = ~pi402 | ~new_n4641_;
  assign new_n6259_ = ~pi370 | ~new_n4642_;
  assign new_n6260_ = ~new_n15023_ | ~new_n4639_;
  assign new_n6261_ = ~new_n4670_;
  assign new_n6262_ = ~new_n4654_ | ~new_n4673_;
  assign new_n6263_ = ~new_n19714_ | ~new_n5571_;
  assign new_n6264_ = ~new_n20658_ | ~new_n4631_;
  assign new_n6265_ = ~new_n19304_ | ~new_n4630_;
  assign new_n6266_ = ~new_n16639_ | ~new_n4634_;
  assign new_n6267_ = ~new_n20186_ | ~new_n5579_;
  assign new_n6268_ = ~new_n17703_ | ~new_n5575_;
  assign new_n6269_ = ~new_n18204_ | ~new_n4632_;
  assign new_n6270_ = ~new_n5024_;
  assign new_n6271_ = ~new_n16354_ | ~new_n4647_;
  assign new_n6272_ = ~new_n4646_ | ~new_n4670_;
  assign new_n6273_ = ~new_n17202_ | ~new_n4644_;
  assign new_n6274_ = ~new_n5585_ | ~new_n5748_;
  assign new_n6275_ = ~new_n5355_ | ~new_n6270_;
  assign new_n6276_ = ~new_n14973_ | ~new_n4639_;
  assign new_n6277_ = ~pi435 | ~new_n4640_;
  assign new_n6278_ = ~pi403 | ~new_n4641_;
  assign new_n6279_ = ~pi371 | ~new_n4642_;
  assign new_n6280_ = ~new_n4671_;
  assign new_n6281_ = ~new_n4654_ | ~new_n4669_;
  assign new_n6282_ = ~new_n19790_ | ~new_n5571_;
  assign new_n6283_ = ~new_n20734_ | ~new_n4631_;
  assign new_n6284_ = ~new_n19303_ | ~new_n4630_;
  assign new_n6285_ = ~new_n16715_ | ~new_n4634_;
  assign new_n6286_ = ~new_n20262_ | ~new_n5579_;
  assign new_n6287_ = ~new_n17702_ | ~new_n5575_;
  assign new_n6288_ = ~new_n18203_ | ~new_n4632_;
  assign new_n6289_ = ~new_n5026_;
  assign new_n6290_ = ~new_n16299_ | ~new_n4647_;
  assign new_n6291_ = ~new_n4646_ | ~new_n4671_;
  assign new_n6292_ = ~new_n17201_ | ~new_n4644_;
  assign new_n6293_ = ~new_n5584_ | ~new_n5748_;
  assign new_n6294_ = ~new_n5358_ | ~new_n6289_;
  assign new_n6295_ = ~pi436 | ~new_n4640_;
  assign new_n6296_ = ~pi404 | ~new_n4641_;
  assign new_n6297_ = ~pi372 | ~new_n4642_;
  assign new_n6298_ = ~new_n4675_;
  assign new_n6299_ = ~new_n7344_ | ~new_n4976_;
  assign new_n6300_ = ~new_n5525_ | ~new_n6299_;
  assign new_n6301_ = ~new_n5359_ | ~new_n4675_;
  assign new_n6302_ = ~new_n4654_ | ~new_n4670_;
  assign new_n6303_ = ~new_n19715_ | ~new_n5571_;
  assign new_n6304_ = ~new_n20659_ | ~new_n4631_;
  assign new_n6305_ = ~new_n19302_ | ~new_n4630_;
  assign new_n6306_ = ~new_n16640_ | ~new_n4634_;
  assign new_n6307_ = ~new_n20187_ | ~new_n5579_;
  assign new_n6308_ = ~new_n17701_ | ~new_n5575_;
  assign new_n6309_ = ~new_n18202_ | ~new_n4632_;
  assign new_n6310_ = ~new_n5028_;
  assign new_n6311_ = ~new_n16352_ | ~new_n4647_;
  assign new_n6312_ = ~new_n17200_ | ~new_n4644_;
  assign new_n6313_ = ~new_n5595_ | ~new_n5748_;
  assign new_n6314_ = ~new_n5363_ | ~new_n6310_;
  assign new_n6315_ = ~pi437 | ~new_n4640_;
  assign new_n6316_ = ~pi405 | ~new_n4641_;
  assign new_n6317_ = ~pi373 | ~new_n4642_;
  assign new_n6318_ = ~new_n4672_;
  assign new_n6319_ = ~new_n16301_ | ~new_n4647_;
  assign new_n6320_ = ~new_n5594_ | ~new_n5748_;
  assign new_n6321_ = ~new_n6319_ | ~new_n6320_ | ~new_n5558_;
  assign new_n6322_ = ~new_n16350_ | ~new_n4647_;
  assign new_n6323_ = ~new_n5593_ | ~new_n5748_;
  assign new_n6324_ = ~new_n6322_ | ~new_n6323_ | ~new_n5558_;
  assign new_n6325_ = ~new_n5598_ | ~new_n5055_;
  assign new_n6326_ = ~new_n4636_ | ~new_n5366_;
  assign new_n6327_ = ~new_n5034_ | ~new_n6326_;
  assign new_n6328_ = ~new_n4635_ | ~new_n7324_;
  assign new_n6329_ = ~new_n5574_ | ~new_n6328_;
  assign new_n6330_ = ~new_n4656_ | ~new_n4694_;
  assign new_n6331_ = ~new_n4653_ | ~new_n17194_;
  assign new_n6332_ = ~new_n4652_ | ~pi500;
  assign new_n6333_ = ~new_n4651_ | ~new_n5064_;
  assign new_n6334_ = ~new_n4650_ | ~new_n5064_;
  assign new_n6335_ = ~new_n4656_ | ~new_n4684_;
  assign new_n6336_ = ~new_n4653_ | ~new_n17193_;
  assign new_n6337_ = ~new_n4652_ | ~pi510;
  assign new_n6338_ = ~new_n4651_ | ~new_n5069_;
  assign new_n6339_ = ~new_n4650_ | ~new_n16337_;
  assign new_n6340_ = ~new_n4656_ | ~new_n4680_;
  assign new_n6341_ = ~new_n4653_ | ~new_n17115_;
  assign new_n6342_ = ~new_n4652_ | ~pi495;
  assign new_n6343_ = ~new_n4651_ | ~new_n5072_;
  assign new_n6344_ = ~new_n4650_ | ~new_n16300_;
  assign new_n6345_ = ~new_n4656_ | ~new_n4676_;
  assign new_n6346_ = ~new_n4653_ | ~new_n17199_;
  assign new_n6347_ = ~new_n4652_ | ~new_n14972_;
  assign new_n6348_ = ~new_n4651_ | ~new_n5075_;
  assign new_n6349_ = ~new_n4650_ | ~new_n16302_;
  assign new_n6350_ = ~new_n4656_ | ~new_n4683_;
  assign new_n6351_ = ~new_n4653_ | ~new_n17198_;
  assign new_n6352_ = ~new_n4652_ | ~new_n15022_;
  assign new_n6353_ = ~new_n4651_ | ~new_n5078_;
  assign new_n6354_ = ~new_n4650_ | ~new_n16303_;
  assign new_n6355_ = ~new_n4656_ | ~new_n4687_;
  assign new_n6356_ = ~new_n4653_ | ~new_n17116_;
  assign new_n6357_ = ~new_n4652_ | ~new_n15021_;
  assign new_n6358_ = ~new_n4651_ | ~new_n5081_;
  assign new_n6359_ = ~new_n4650_ | ~new_n16347_;
  assign new_n6360_ = ~new_n4656_ | ~new_n4686_;
  assign new_n6361_ = ~new_n4653_ | ~new_n17197_;
  assign new_n6362_ = ~new_n4652_ | ~new_n15020_;
  assign new_n6363_ = ~new_n4651_ | ~new_n5084_;
  assign new_n6364_ = ~new_n4650_ | ~new_n16304_;
  assign new_n6365_ = ~new_n4656_ | ~new_n4700_;
  assign new_n6366_ = ~new_n4653_ | ~new_n17117_;
  assign new_n6367_ = ~new_n4652_ | ~new_n15019_;
  assign new_n6368_ = ~new_n4651_ | ~new_n5087_;
  assign new_n6369_ = ~new_n4650_ | ~new_n16305_;
  assign new_n6370_ = ~new_n4656_ | ~new_n4699_;
  assign new_n6371_ = ~new_n4653_ | ~new_n17196_;
  assign new_n6372_ = ~new_n4652_ | ~new_n15018_;
  assign new_n6373_ = ~new_n4651_ | ~new_n5090_;
  assign new_n6374_ = ~new_n4650_ | ~new_n16306_;
  assign new_n6375_ = ~new_n4656_ | ~new_n4678_;
  assign new_n6376_ = ~new_n4653_ | ~new_n17195_;
  assign new_n6377_ = ~new_n4652_ | ~new_n15017_;
  assign new_n6378_ = ~new_n4651_ | ~new_n5093_;
  assign new_n6379_ = ~new_n4650_ | ~new_n16345_;
  assign new_n6380_ = ~new_n4656_ | ~new_n4679_;
  assign new_n6381_ = ~new_n4653_ | ~new_n17109_;
  assign new_n6382_ = ~new_n4652_ | ~new_n15041_;
  assign new_n6383_ = ~new_n4651_ | ~new_n5096_;
  assign new_n6384_ = ~new_n4650_ | ~new_n16288_;
  assign new_n6385_ = ~new_n4656_ | ~new_n4688_;
  assign new_n6386_ = ~new_n4653_ | ~new_n17213_;
  assign new_n6387_ = ~new_n4652_ | ~new_n15040_;
  assign new_n6388_ = ~new_n4651_ | ~new_n5099_;
  assign new_n6389_ = ~new_n4650_ | ~new_n16289_;
  assign new_n6390_ = ~new_n4656_ | ~new_n4696_;
  assign new_n6391_ = ~new_n4653_ | ~new_n17212_;
  assign new_n6392_ = ~new_n4652_ | ~new_n15039_;
  assign new_n6393_ = ~new_n4651_ | ~new_n5102_;
  assign new_n6394_ = ~new_n4650_ | ~new_n16290_;
  assign new_n6395_ = ~new_n4656_ | ~new_n4695_;
  assign new_n6396_ = ~new_n4653_ | ~new_n17110_;
  assign new_n6397_ = ~new_n4652_ | ~new_n15038_;
  assign new_n6398_ = ~new_n4651_ | ~new_n5105_;
  assign new_n6399_ = ~new_n4650_ | ~new_n16368_;
  assign new_n6400_ = ~new_n4656_ | ~new_n4690_;
  assign new_n6401_ = ~new_n4653_ | ~new_n17211_;
  assign new_n6402_ = ~new_n4652_ | ~new_n15037_;
  assign new_n6403_ = ~new_n4651_ | ~new_n5108_;
  assign new_n6404_ = ~new_n4650_ | ~new_n16291_;
  assign new_n6405_ = ~new_n4656_ | ~new_n4689_;
  assign new_n6406_ = ~new_n4653_ | ~new_n17210_;
  assign new_n6407_ = ~new_n4652_ | ~new_n15036_;
  assign new_n6408_ = ~new_n4651_ | ~new_n5111_;
  assign new_n6409_ = ~new_n4650_ | ~new_n16292_;
  assign new_n6410_ = ~new_n4656_ | ~new_n4685_;
  assign new_n6411_ = ~new_n4653_ | ~new_n17209_;
  assign new_n6412_ = ~new_n4652_ | ~new_n15035_;
  assign new_n6413_ = ~new_n4651_ | ~new_n5114_;
  assign new_n6414_ = ~new_n4650_ | ~new_n16293_;
  assign new_n6415_ = ~new_n4656_ | ~new_n4698_;
  assign new_n6416_ = ~new_n4653_ | ~new_n17111_;
  assign new_n6417_ = ~new_n4652_ | ~new_n15034_;
  assign new_n6418_ = ~new_n4651_ | ~new_n5117_;
  assign new_n6419_ = ~new_n4650_ | ~new_n16366_;
  assign new_n6420_ = ~new_n4656_ | ~new_n4697_;
  assign new_n6421_ = ~new_n4653_ | ~new_n17208_;
  assign new_n6422_ = ~new_n4652_ | ~new_n15033_;
  assign new_n6423_ = ~new_n4651_ | ~new_n5120_;
  assign new_n6424_ = ~new_n4650_ | ~new_n16294_;
  assign new_n6425_ = ~new_n4656_ | ~new_n4692_;
  assign new_n6426_ = ~new_n4653_ | ~new_n17207_;
  assign new_n6427_ = ~new_n4652_ | ~new_n15032_;
  assign new_n6428_ = ~new_n4651_ | ~new_n5122_;
  assign new_n6429_ = ~new_n4650_ | ~new_n16364_;
  assign new_n6430_ = ~new_n4656_ | ~new_n4691_;
  assign new_n6431_ = ~new_n4653_ | ~new_n17112_;
  assign new_n6432_ = ~new_n4652_ | ~new_n15031_;
  assign new_n6433_ = ~new_n4651_ | ~new_n5592_;
  assign new_n6434_ = ~new_n4650_ | ~new_n16295_;
  assign new_n6435_ = ~new_n4656_ | ~new_n4677_;
  assign new_n6436_ = ~new_n4653_ | ~new_n17113_;
  assign new_n6437_ = ~new_n4652_ | ~new_n15030_;
  assign new_n6438_ = ~new_n4651_ | ~new_n5591_;
  assign new_n6439_ = ~new_n4650_ | ~new_n16360_;
  assign new_n6440_ = ~new_n4656_ | ~new_n4682_;
  assign new_n6441_ = ~new_n4653_ | ~new_n17206_;
  assign new_n6442_ = ~new_n4652_ | ~new_n15029_;
  assign new_n6443_ = ~new_n4651_ | ~new_n5590_;
  assign new_n6444_ = ~new_n4650_ | ~new_n16296_;
  assign new_n6445_ = ~new_n4656_ | ~new_n4681_;
  assign new_n6446_ = ~new_n4653_ | ~new_n17205_;
  assign new_n6447_ = ~new_n4652_ | ~new_n15028_;
  assign new_n6448_ = ~new_n4651_ | ~new_n5589_;
  assign new_n6449_ = ~new_n4650_ | ~new_n16358_;
  assign new_n6450_ = ~new_n4656_ | ~new_n4674_;
  assign new_n6451_ = ~new_n4653_ | ~new_n17204_;
  assign new_n6452_ = ~new_n4652_ | ~new_n15027_;
  assign new_n6453_ = ~new_n4651_ | ~new_n5588_;
  assign new_n6454_ = ~new_n4650_ | ~new_n16297_;
  assign new_n6455_ = ~new_n4656_ | ~new_n4673_;
  assign new_n6456_ = ~new_n4653_ | ~new_n17203_;
  assign new_n6457_ = ~new_n4652_ | ~new_n15026_;
  assign new_n6458_ = ~new_n4651_ | ~new_n5587_;
  assign new_n6459_ = ~new_n4650_ | ~new_n16356_;
  assign new_n6460_ = ~new_n4656_ | ~new_n4669_;
  assign new_n6461_ = ~new_n4653_ | ~new_n17114_;
  assign new_n6462_ = ~new_n4652_ | ~new_n15025_;
  assign new_n6463_ = ~new_n4651_ | ~new_n5586_;
  assign new_n6464_ = ~new_n4650_ | ~new_n16298_;
  assign new_n6465_ = ~new_n4656_ | ~new_n4670_;
  assign new_n6466_ = ~new_n4653_ | ~new_n17202_;
  assign new_n6467_ = ~new_n4652_ | ~new_n15024_;
  assign new_n6468_ = ~new_n4651_ | ~new_n5585_;
  assign new_n6469_ = ~new_n4650_ | ~new_n16354_;
  assign new_n6470_ = ~new_n4656_ | ~new_n4671_;
  assign new_n6471_ = ~new_n4653_ | ~new_n17201_;
  assign new_n6472_ = ~new_n4652_ | ~new_n15023_;
  assign new_n6473_ = ~new_n4651_ | ~new_n5584_;
  assign new_n6474_ = ~new_n4650_ | ~new_n16299_;
  assign new_n6475_ = ~new_n4653_ | ~new_n17200_;
  assign new_n6476_ = ~new_n4652_ | ~new_n14973_;
  assign new_n6477_ = ~new_n4651_ | ~new_n5595_;
  assign new_n6478_ = ~new_n4650_ | ~new_n16352_;
  assign new_n6479_ = ~new_n4651_ | ~new_n5594_;
  assign new_n6480_ = ~new_n4650_ | ~new_n16301_;
  assign new_n6481_ = ~new_n4651_ | ~new_n5593_;
  assign new_n6482_ = ~new_n4650_ | ~new_n16350_;
  assign new_n6483_ = ~new_n15992_ | ~new_n4638_;
  assign new_n6484_ = ~new_n7344_ | ~new_n5061_;
  assign new_n6485_ = ~new_n15687_ | ~new_n7349_;
  assign new_n6486_ = ~new_n6485_ | ~new_n6484_ | ~new_n6483_;
  assign new_n6487_ = ~new_n15992_ | ~new_n4638_;
  assign new_n6488_ = ~new_n4637_ | ~new_n15687_;
  assign new_n6489_ = ~new_n7344_ | ~new_n5061_;
  assign new_n6490_ = ~new_n6489_ | ~new_n6488_ | ~new_n6487_;
  assign new_n6491_ = ~new_n5040_;
  assign new_n6492_ = ~new_n4661_ | ~new_n6486_;
  assign new_n6493_ = ~po511 | ~new_n6490_;
  assign new_n6494_ = ~new_n4660_ | ~new_n15992_;
  assign new_n6495_ = ~pi513 | ~po509;
  assign new_n6496_ = ~new_n4659_ | ~new_n5061_;
  assign new_n6497_ = ~new_n4658_ | ~new_n15687_;
  assign new_n6498_ = ~pi438 | ~new_n6491_;
  assign new_n6499_ = ~new_n16054_ | ~new_n4638_;
  assign new_n6500_ = ~new_n7344_ | ~new_n5119_;
  assign new_n6501_ = ~new_n15749_ | ~new_n7349_;
  assign new_n6502_ = ~new_n6501_ | ~new_n6500_ | ~new_n6499_;
  assign new_n6503_ = ~new_n16054_ | ~new_n4638_;
  assign new_n6504_ = ~new_n15749_ | ~new_n4637_;
  assign new_n6505_ = ~new_n7344_ | ~new_n5119_;
  assign new_n6506_ = ~new_n6505_ | ~new_n6504_ | ~new_n6503_;
  assign new_n6507_ = ~new_n4661_ | ~new_n6502_;
  assign new_n6508_ = ~po511 | ~new_n6506_;
  assign new_n6509_ = ~new_n16054_ | ~new_n4660_;
  assign new_n6510_ = ~pi494 | ~po509;
  assign new_n6511_ = ~new_n4659_ | ~new_n5119_;
  assign new_n6512_ = ~new_n15749_ | ~new_n4658_;
  assign new_n6513_ = ~pi439 | ~new_n6491_;
  assign new_n6514_ = ~new_n15991_ | ~new_n4638_;
  assign new_n6515_ = ~new_n7344_ | ~new_n5116_;
  assign new_n6516_ = ~new_n15686_ | ~new_n7349_;
  assign new_n6517_ = ~new_n6516_ | ~new_n6515_ | ~new_n6514_;
  assign new_n6518_ = ~new_n15991_ | ~new_n4638_;
  assign new_n6519_ = ~new_n15686_ | ~new_n4637_;
  assign new_n6520_ = ~new_n7344_ | ~new_n5116_;
  assign new_n6521_ = ~new_n6520_ | ~new_n6519_ | ~new_n6518_;
  assign new_n6522_ = ~new_n4661_ | ~new_n6517_;
  assign new_n6523_ = ~po511 | ~new_n6521_;
  assign new_n6524_ = ~new_n15991_ | ~new_n4660_;
  assign new_n6525_ = ~pi504 | ~po509;
  assign new_n6526_ = ~new_n4659_ | ~new_n5116_;
  assign new_n6527_ = ~new_n15686_ | ~new_n4658_;
  assign new_n6528_ = ~pi440 | ~new_n6491_;
  assign new_n6529_ = ~new_n16055_ | ~new_n4638_;
  assign new_n6530_ = ~new_n7344_ | ~new_n5113_;
  assign new_n6531_ = ~new_n15750_ | ~new_n7349_;
  assign new_n6532_ = ~new_n6531_ | ~new_n6530_ | ~new_n6529_;
  assign new_n6533_ = ~new_n16055_ | ~new_n4638_;
  assign new_n6534_ = ~new_n15750_ | ~new_n4637_;
  assign new_n6535_ = ~new_n7344_ | ~new_n5113_;
  assign new_n6536_ = ~new_n6535_ | ~new_n6534_ | ~new_n6533_;
  assign new_n6537_ = ~new_n4661_ | ~new_n6532_;
  assign new_n6538_ = ~po511 | ~new_n6536_;
  assign new_n6539_ = ~new_n16055_ | ~new_n4660_;
  assign new_n6540_ = ~pi506 | ~po509;
  assign new_n6541_ = ~new_n4659_ | ~new_n5113_;
  assign new_n6542_ = ~new_n15750_ | ~new_n4658_;
  assign new_n6543_ = ~pi441 | ~new_n6491_;
  assign new_n6544_ = ~new_n16056_ | ~new_n4638_;
  assign new_n6545_ = ~new_n7344_ | ~new_n5110_;
  assign new_n6546_ = ~new_n15751_ | ~new_n7349_;
  assign new_n6547_ = ~new_n6546_ | ~new_n6545_ | ~new_n6544_;
  assign new_n6548_ = ~new_n16056_ | ~new_n4638_;
  assign new_n6549_ = ~new_n15751_ | ~new_n4637_;
  assign new_n6550_ = ~new_n7344_ | ~new_n5110_;
  assign new_n6551_ = ~new_n6550_ | ~new_n6549_ | ~new_n6548_;
  assign new_n6552_ = ~new_n4661_ | ~new_n6547_;
  assign new_n6553_ = ~po511 | ~new_n6551_;
  assign new_n6554_ = ~new_n16056_ | ~new_n4660_;
  assign new_n6555_ = ~pi491 | ~po509;
  assign new_n6556_ = ~new_n4659_ | ~new_n5110_;
  assign new_n6557_ = ~new_n15751_ | ~new_n4658_;
  assign new_n6558_ = ~pi442 | ~new_n6491_;
  assign new_n6559_ = ~new_n16057_ | ~new_n4638_;
  assign new_n6560_ = ~new_n7344_ | ~new_n5107_;
  assign new_n6561_ = ~new_n15752_ | ~new_n7349_;
  assign new_n6562_ = ~new_n6561_ | ~new_n6560_ | ~new_n6559_;
  assign new_n6563_ = ~new_n16057_ | ~new_n4638_;
  assign new_n6564_ = ~new_n15752_ | ~new_n4637_;
  assign new_n6565_ = ~new_n7344_ | ~new_n5107_;
  assign new_n6566_ = ~new_n6565_ | ~new_n6564_ | ~new_n6563_;
  assign new_n6567_ = ~new_n4661_ | ~new_n6562_;
  assign new_n6568_ = ~po511 | ~new_n6566_;
  assign new_n6569_ = ~new_n16057_ | ~new_n4660_;
  assign new_n6570_ = ~pi517 | ~po509;
  assign new_n6571_ = ~new_n4659_ | ~new_n5107_;
  assign new_n6572_ = ~new_n15752_ | ~new_n4658_;
  assign new_n6573_ = ~pi443 | ~new_n6491_;
  assign new_n6574_ = ~new_n15990_ | ~new_n4638_;
  assign new_n6575_ = ~new_n7344_ | ~new_n5104_;
  assign new_n6576_ = ~new_n15685_ | ~new_n7349_;
  assign new_n6577_ = ~new_n6576_ | ~new_n6575_ | ~new_n6574_;
  assign new_n6578_ = ~new_n15990_ | ~new_n4638_;
  assign new_n6579_ = ~new_n15685_ | ~new_n4637_;
  assign new_n6580_ = ~new_n7344_ | ~new_n5104_;
  assign new_n6581_ = ~new_n6580_ | ~new_n6579_ | ~new_n6578_;
  assign new_n6582_ = ~new_n4661_ | ~new_n6577_;
  assign new_n6583_ = ~po511 | ~new_n6581_;
  assign new_n6584_ = ~new_n15990_ | ~new_n4660_;
  assign new_n6585_ = ~pi498 | ~po509;
  assign new_n6586_ = ~new_n4659_ | ~new_n5104_;
  assign new_n6587_ = ~new_n15685_ | ~new_n4658_;
  assign new_n6588_ = ~pi444 | ~new_n6491_;
  assign new_n6589_ = ~new_n16058_ | ~new_n4638_;
  assign new_n6590_ = ~new_n7344_ | ~new_n5101_;
  assign new_n6591_ = ~new_n15753_ | ~new_n7349_;
  assign new_n6592_ = ~new_n6591_ | ~new_n6590_ | ~new_n6589_;
  assign new_n6593_ = ~new_n16058_ | ~new_n4638_;
  assign new_n6594_ = ~new_n15753_ | ~new_n4637_;
  assign new_n6595_ = ~new_n7344_ | ~new_n5101_;
  assign new_n6596_ = ~new_n6595_ | ~new_n6594_ | ~new_n6593_;
  assign new_n6597_ = ~new_n4661_ | ~new_n6592_;
  assign new_n6598_ = ~po511 | ~new_n6596_;
  assign new_n6599_ = ~new_n16058_ | ~new_n4660_;
  assign new_n6600_ = ~pi508 | ~po509;
  assign new_n6601_ = ~new_n4659_ | ~new_n5101_;
  assign new_n6602_ = ~new_n15753_ | ~new_n4658_;
  assign new_n6603_ = ~pi445 | ~new_n6491_;
  assign new_n6604_ = ~new_n16059_ | ~new_n4638_;
  assign new_n6605_ = ~new_n7344_ | ~new_n5098_;
  assign new_n6606_ = ~new_n15754_ | ~new_n7349_;
  assign new_n6607_ = ~new_n6606_ | ~new_n6605_ | ~new_n6604_;
  assign new_n6608_ = ~new_n16059_ | ~new_n4638_;
  assign new_n6609_ = ~new_n15754_ | ~new_n4637_;
  assign new_n6610_ = ~new_n7344_ | ~new_n5098_;
  assign new_n6611_ = ~new_n6610_ | ~new_n6609_ | ~new_n6608_;
  assign new_n6612_ = ~new_n4661_ | ~new_n6607_;
  assign new_n6613_ = ~po511 | ~new_n6611_;
  assign new_n6614_ = ~new_n16059_ | ~new_n4660_;
  assign new_n6615_ = ~pi496 | ~po509;
  assign new_n6616_ = ~new_n4659_ | ~new_n5098_;
  assign new_n6617_ = ~new_n15754_ | ~new_n4658_;
  assign new_n6618_ = ~pi446 | ~new_n6491_;
  assign new_n6619_ = ~new_n15989_ | ~new_n4638_;
  assign new_n6620_ = ~new_n7344_ | ~new_n5095_;
  assign new_n6621_ = ~new_n15684_ | ~new_n7349_;
  assign new_n6622_ = ~new_n6621_ | ~new_n6620_ | ~new_n6619_;
  assign new_n6623_ = ~new_n15989_ | ~new_n4638_;
  assign new_n6624_ = ~new_n15684_ | ~new_n4637_;
  assign new_n6625_ = ~new_n7344_ | ~new_n5095_;
  assign new_n6626_ = ~new_n6625_ | ~new_n6624_ | ~new_n6623_;
  assign new_n6627_ = ~new_n4661_ | ~new_n6622_;
  assign new_n6628_ = ~po511 | ~new_n6626_;
  assign new_n6629_ = ~new_n15989_ | ~new_n4660_;
  assign new_n6630_ = ~pi515 | ~po509;
  assign new_n6631_ = ~new_n4659_ | ~new_n5095_;
  assign new_n6632_ = ~new_n15684_ | ~new_n4658_;
  assign new_n6633_ = ~pi447 | ~new_n6491_;
  assign new_n6634_ = ~new_n16049_ | ~new_n4638_;
  assign new_n6635_ = ~new_n7344_ | ~new_n5092_;
  assign new_n6636_ = ~new_n15744_ | ~new_n7349_;
  assign new_n6637_ = ~new_n6636_ | ~new_n6635_ | ~new_n6634_;
  assign new_n6638_ = ~new_n16049_ | ~new_n4638_;
  assign new_n6639_ = ~new_n15744_ | ~new_n4637_;
  assign new_n6640_ = ~new_n7344_ | ~new_n5092_;
  assign new_n6641_ = ~new_n6640_ | ~new_n6639_ | ~new_n6638_;
  assign new_n6642_ = ~new_n4661_ | ~new_n6637_;
  assign new_n6643_ = ~po511 | ~new_n6641_;
  assign new_n6644_ = ~new_n16049_ | ~new_n4660_;
  assign new_n6645_ = ~pi501 | ~po509;
  assign new_n6646_ = ~new_n4659_ | ~new_n5092_;
  assign new_n6647_ = ~new_n15744_ | ~new_n4658_;
  assign new_n6648_ = ~pi448 | ~new_n6491_;
  assign new_n6649_ = ~new_n16050_ | ~new_n4638_;
  assign new_n6650_ = ~new_n7344_ | ~new_n5089_;
  assign new_n6651_ = ~new_n15745_ | ~new_n7349_;
  assign new_n6652_ = ~new_n6651_ | ~new_n6650_ | ~new_n6649_;
  assign new_n6653_ = ~new_n16050_ | ~new_n4638_;
  assign new_n6654_ = ~new_n15745_ | ~new_n4637_;
  assign new_n6655_ = ~new_n7344_ | ~new_n5089_;
  assign new_n6656_ = ~new_n6655_ | ~new_n6654_ | ~new_n6653_;
  assign new_n6657_ = ~new_n4661_ | ~new_n6652_;
  assign new_n6658_ = ~po511 | ~new_n6656_;
  assign new_n6659_ = ~new_n16050_ | ~new_n4660_;
  assign new_n6660_ = ~pi511 | ~po509;
  assign new_n6661_ = ~new_n4659_ | ~new_n5089_;
  assign new_n6662_ = ~new_n15745_ | ~new_n4658_;
  assign new_n6663_ = ~pi449 | ~new_n6491_;
  assign new_n6664_ = ~new_n15995_ | ~new_n4638_;
  assign new_n6665_ = ~new_n7344_ | ~new_n5086_;
  assign new_n6666_ = ~new_n15690_ | ~new_n7349_;
  assign new_n6667_ = ~new_n6666_ | ~new_n6665_ | ~new_n6664_;
  assign new_n6668_ = ~new_n15995_ | ~new_n4638_;
  assign new_n6669_ = ~new_n15690_ | ~new_n4637_;
  assign new_n6670_ = ~new_n7344_ | ~new_n5086_;
  assign new_n6671_ = ~new_n6670_ | ~new_n6669_ | ~new_n6668_;
  assign new_n6672_ = ~new_n4661_ | ~new_n6667_;
  assign new_n6673_ = ~po511 | ~new_n6671_;
  assign new_n6674_ = ~new_n15995_ | ~new_n4660_;
  assign new_n6675_ = ~pi519 | ~po509;
  assign new_n6676_ = ~new_n4659_ | ~new_n5086_;
  assign new_n6677_ = ~new_n15690_ | ~new_n4658_;
  assign new_n6678_ = ~pi450 | ~new_n6491_;
  assign new_n6679_ = ~new_n16051_ | ~new_n4638_;
  assign new_n6680_ = ~new_n7344_ | ~new_n5083_;
  assign new_n6681_ = ~new_n15746_ | ~new_n7349_;
  assign new_n6682_ = ~new_n6681_ | ~new_n6680_ | ~new_n6679_;
  assign new_n6683_ = ~new_n16051_ | ~new_n4638_;
  assign new_n6684_ = ~new_n15746_ | ~new_n4637_;
  assign new_n6685_ = ~new_n7344_ | ~new_n5083_;
  assign new_n6686_ = ~new_n6685_ | ~new_n6684_ | ~new_n6683_;
  assign new_n6687_ = ~new_n4661_ | ~new_n6682_;
  assign new_n6688_ = ~po511 | ~new_n6686_;
  assign new_n6689_ = ~new_n16051_ | ~new_n4660_;
  assign new_n6690_ = ~pi493 | ~po509;
  assign new_n6691_ = ~new_n4659_ | ~new_n5083_;
  assign new_n6692_ = ~new_n15746_ | ~new_n4658_;
  assign new_n6693_ = ~pi451 | ~new_n6491_;
  assign new_n6694_ = ~new_n15994_ | ~new_n4638_;
  assign new_n6695_ = ~new_n7344_ | ~new_n5080_;
  assign new_n6696_ = ~new_n15689_ | ~new_n7349_;
  assign new_n6697_ = ~new_n6696_ | ~new_n6695_ | ~new_n6694_;
  assign new_n6698_ = ~new_n15994_ | ~new_n4638_;
  assign new_n6699_ = ~new_n15689_ | ~new_n4637_;
  assign new_n6700_ = ~new_n7344_ | ~new_n5080_;
  assign new_n6701_ = ~new_n6700_ | ~new_n6699_ | ~new_n6698_;
  assign new_n6702_ = ~new_n4661_ | ~new_n6697_;
  assign new_n6703_ = ~po511 | ~new_n6701_;
  assign new_n6704_ = ~new_n15994_ | ~new_n4660_;
  assign new_n6705_ = ~pi505 | ~po509;
  assign new_n6706_ = ~new_n4659_ | ~new_n5080_;
  assign new_n6707_ = ~new_n15689_ | ~new_n4658_;
  assign new_n6708_ = ~pi452 | ~new_n6491_;
  assign new_n6709_ = ~new_n16052_ | ~new_n4638_;
  assign new_n6710_ = ~new_n7344_ | ~new_n5077_;
  assign new_n6711_ = ~new_n15747_ | ~new_n7349_;
  assign new_n6712_ = ~new_n6711_ | ~new_n6710_ | ~new_n6709_;
  assign new_n6713_ = ~new_n16052_ | ~new_n4638_;
  assign new_n6714_ = ~new_n15747_ | ~new_n4637_;
  assign new_n6715_ = ~new_n7344_ | ~new_n5077_;
  assign new_n6716_ = ~new_n6715_ | ~new_n6714_ | ~new_n6713_;
  assign new_n6717_ = ~new_n4661_ | ~new_n6712_;
  assign new_n6718_ = ~po511 | ~new_n6716_;
  assign new_n6719_ = ~new_n16052_ | ~new_n4660_;
  assign new_n6720_ = ~pi502 | ~po509;
  assign new_n6721_ = ~new_n4659_ | ~new_n5077_;
  assign new_n6722_ = ~new_n15747_ | ~new_n4658_;
  assign new_n6723_ = ~pi453 | ~new_n6491_;
  assign new_n6724_ = ~new_n16053_ | ~new_n4638_;
  assign new_n6725_ = ~new_n7344_ | ~new_n5074_;
  assign new_n6726_ = ~new_n15748_ | ~new_n7349_;
  assign new_n6727_ = ~new_n6726_ | ~new_n6725_ | ~new_n6724_;
  assign new_n6728_ = ~new_n16053_ | ~new_n4638_;
  assign new_n6729_ = ~new_n15748_ | ~new_n4637_;
  assign new_n6730_ = ~new_n7344_ | ~new_n5074_;
  assign new_n6731_ = ~new_n6730_ | ~new_n6729_ | ~new_n6728_;
  assign new_n6732_ = ~new_n4661_ | ~new_n6727_;
  assign new_n6733_ = ~po511 | ~new_n6731_;
  assign new_n6734_ = ~new_n16053_ | ~new_n4660_;
  assign new_n6735_ = ~pi514 | ~po509;
  assign new_n6736_ = ~new_n4659_ | ~new_n5074_;
  assign new_n6737_ = ~new_n15748_ | ~new_n4658_;
  assign new_n6738_ = ~pi454 | ~new_n6491_;
  assign new_n6739_ = ~new_n15993_ | ~new_n4638_;
  assign new_n6740_ = ~new_n7344_ | ~new_n5071_;
  assign new_n6741_ = ~new_n15688_ | ~new_n7349_;
  assign new_n6742_ = ~new_n6741_ | ~new_n6740_ | ~new_n6739_;
  assign new_n6743_ = ~new_n15993_ | ~new_n4638_;
  assign new_n6744_ = ~new_n15688_ | ~new_n4637_;
  assign new_n6745_ = ~new_n7344_ | ~new_n5071_;
  assign new_n6746_ = ~new_n6745_ | ~new_n6744_ | ~new_n6743_;
  assign new_n6747_ = ~new_n4661_ | ~new_n6742_;
  assign new_n6748_ = ~po511 | ~new_n6746_;
  assign new_n6749_ = ~new_n15993_ | ~new_n4660_;
  assign new_n6750_ = ~pi495 | ~po509;
  assign new_n6751_ = ~new_n4659_ | ~new_n5071_;
  assign new_n6752_ = ~new_n15688_ | ~new_n4658_;
  assign new_n6753_ = ~pi455 | ~new_n6491_;
  assign new_n6754_ = ~new_n16047_ | ~new_n4638_;
  assign new_n6755_ = ~new_n7344_ | ~new_n5068_;
  assign new_n6756_ = ~new_n15742_ | ~new_n7349_;
  assign new_n6757_ = ~new_n6756_ | ~new_n6755_ | ~new_n6754_;
  assign new_n6758_ = ~new_n16047_ | ~new_n4638_;
  assign new_n6759_ = ~new_n15742_ | ~new_n4637_;
  assign new_n6760_ = ~new_n7344_ | ~new_n5068_;
  assign new_n6761_ = ~new_n6760_ | ~new_n6759_ | ~new_n6758_;
  assign new_n6762_ = ~new_n4661_ | ~new_n6757_;
  assign new_n6763_ = ~po511 | ~new_n6761_;
  assign new_n6764_ = ~new_n16047_ | ~new_n4660_;
  assign new_n6765_ = ~pi510 | ~po509;
  assign new_n6766_ = ~new_n4659_ | ~new_n5068_;
  assign new_n6767_ = ~new_n15742_ | ~new_n4658_;
  assign new_n6768_ = ~pi456 | ~new_n6491_;
  assign new_n6769_ = ~new_n16048_ | ~new_n4638_;
  assign new_n6770_ = ~new_n7344_ | ~new_n5062_;
  assign new_n6771_ = ~new_n15743_ | ~new_n7349_;
  assign new_n6772_ = ~new_n5485_ | ~new_n6769_;
  assign new_n6773_ = ~new_n16048_ | ~new_n4638_;
  assign new_n6774_ = ~new_n15743_ | ~new_n4637_;
  assign new_n6775_ = ~new_n7344_ | ~new_n5062_;
  assign new_n6776_ = ~new_n6775_ | ~new_n6774_ | ~new_n6773_;
  assign new_n6777_ = ~new_n4661_ | ~new_n6772_;
  assign new_n6778_ = ~po511 | ~new_n6776_;
  assign new_n6779_ = ~new_n16048_ | ~new_n4660_;
  assign new_n6780_ = ~pi500 | ~po509;
  assign new_n6781_ = ~new_n4659_ | ~new_n5062_;
  assign new_n6782_ = ~new_n15743_ | ~new_n4658_;
  assign new_n6783_ = ~pi457 | ~new_n6491_;
  assign new_n6784_ = ~new_n5563_;
  assign new_n6785_ = ~new_n4979_ | ~new_n5032_;
  assign new_n6786_ = ~new_n4982_ | ~new_n5044_;
  assign new_n6787_ = ~new_n5035_ | ~new_n4980_;
  assign new_n6788_ = ~new_n4634_ | ~new_n7715_ | ~new_n7714_;
  assign new_n6789_ = ~new_n15125_ | ~new_n6787_;
  assign new_n6790_ = ~new_n5501_ | ~new_n5562_ | ~new_n7817_ | ~new_n7816_;
  assign new_n6791_ = ~new_n4668_ | ~new_n7717_ | ~new_n7716_;
  assign new_n6792_ = ~new_n5596_ | ~new_n4643_;
  assign new_n6793_ = ~pi490 | ~new_n6791_;
  assign new_n6794_ = ~new_n4657_ | ~new_n4695_;
  assign new_n6795_ = ~new_n4655_ | ~new_n4689_;
  assign new_n6796_ = ~new_n15036_ | ~new_n5043_;
  assign new_n6797_ = ~new_n6796_ | ~new_n6795_ | ~new_n6794_;
  assign new_n6798_ = ~new_n4630_ | ~new_n7333_;
  assign new_n6799_ = ~new_n5035_ | ~new_n5504_ | ~new_n6798_ | ~new_n4985_ | ~new_n4983_;
  assign new_n6800_ = ~new_n6799_ | ~new_n5043_;
  assign new_n6801_ = ~new_n5046_;
  assign new_n6802_ = ~new_n5111_ | ~new_n7294_;
  assign new_n6803_ = ~new_n15036_ | ~new_n7293_;
  assign new_n6804_ = ~new_n5604_ | ~new_n6797_;
  assign new_n6805_ = ~new_n18704_ | ~new_n4648_;
  assign new_n6806_ = ~pi491 | ~po509;
  assign new_n6807_ = ~new_n4657_ | ~new_n4674_;
  assign new_n6808_ = ~new_n4655_ | ~new_n4669_;
  assign new_n6809_ = ~new_n15025_ | ~new_n5043_;
  assign new_n6810_ = ~new_n6808_ | ~new_n6809_ | ~new_n6807_;
  assign new_n6811_ = ~new_n6329_ | ~new_n5043_;
  assign new_n6812_ = ~new_n6801_ | ~new_n6811_;
  assign new_n6813_ = ~new_n5581_ | ~new_n6329_;
  assign new_n6814_ = ~new_n5034_ | ~new_n6813_;
  assign new_n6815_ = ~new_n4663_ | ~new_n5586_;
  assign new_n6816_ = ~new_n4662_ | ~new_n15025_;
  assign new_n6817_ = ~new_n5604_ | ~new_n6810_;
  assign new_n6818_ = ~new_n18614_ | ~new_n4648_;
  assign new_n6819_ = ~pi492 | ~po509;
  assign new_n6820_ = ~new_n4657_ | ~new_n4683_;
  assign new_n6821_ = ~new_n4655_ | ~new_n4686_;
  assign new_n6822_ = ~new_n15020_ | ~new_n5043_;
  assign new_n6823_ = ~new_n6822_ | ~new_n6821_ | ~new_n6820_;
  assign new_n6824_ = ~new_n5084_ | ~new_n7294_;
  assign new_n6825_ = ~new_n15020_ | ~new_n7293_;
  assign new_n6826_ = ~new_n5604_ | ~new_n6823_;
  assign new_n6827_ = ~new_n18689_ | ~new_n4648_;
  assign new_n6828_ = ~pi493 | ~po509;
  assign new_n6829_ = ~new_n4657_ | ~new_n4685_;
  assign new_n6830_ = ~new_n4655_ | ~new_n4697_;
  assign new_n6831_ = ~new_n15033_ | ~new_n5043_;
  assign new_n6832_ = ~new_n6831_ | ~new_n6830_ | ~new_n6829_;
  assign new_n6833_ = ~new_n5120_ | ~new_n7294_;
  assign new_n6834_ = ~new_n15033_ | ~new_n7293_;
  assign new_n6835_ = ~new_n5604_ | ~new_n6832_;
  assign new_n6836_ = ~new_n18702_ | ~new_n4648_;
  assign new_n6837_ = ~pi494 | ~po509;
  assign new_n6838_ = ~new_n4657_ | ~new_n4694_;
  assign new_n6839_ = ~new_n4655_ | ~new_n4680_;
  assign new_n6840_ = ~pi495 | ~new_n5043_;
  assign new_n6841_ = ~new_n6840_ | ~new_n6839_ | ~new_n6838_;
  assign new_n6842_ = ~new_n5072_ | ~new_n7294_;
  assign new_n6843_ = ~pi495 | ~new_n7293_;
  assign new_n6844_ = ~new_n5604_ | ~new_n6841_;
  assign new_n6845_ = ~new_n18692_ | ~new_n4648_;
  assign new_n6846_ = ~pi495 | ~po509;
  assign new_n6847_ = ~new_n4657_ | ~new_n4678_;
  assign new_n6848_ = ~new_n4655_ | ~new_n4688_;
  assign new_n6849_ = ~new_n15040_ | ~new_n5043_;
  assign new_n6850_ = ~new_n6849_ | ~new_n6848_ | ~new_n6847_;
  assign new_n6851_ = ~new_n5099_ | ~new_n7294_;
  assign new_n6852_ = ~new_n15040_ | ~new_n7293_;
  assign new_n6853_ = ~new_n5604_ | ~new_n6850_;
  assign new_n6854_ = ~new_n18707_ | ~new_n4648_;
  assign new_n6855_ = ~pi496 | ~po509;
  assign new_n6856_ = ~new_n4657_ | ~new_n4691_;
  assign new_n6857_ = ~new_n4655_ | ~new_n4682_;
  assign new_n6858_ = ~new_n15029_ | ~new_n5043_;
  assign new_n6859_ = ~new_n6857_ | ~new_n6858_ | ~new_n6856_;
  assign new_n6860_ = ~new_n4663_ | ~new_n5590_;
  assign new_n6861_ = ~new_n4662_ | ~new_n15029_;
  assign new_n6862_ = ~new_n5604_ | ~new_n6859_;
  assign new_n6863_ = ~new_n18698_ | ~new_n4648_;
  assign new_n6864_ = ~pi497 | ~po509;
  assign new_n6865_ = ~new_n4657_ | ~new_n4688_;
  assign new_n6866_ = ~new_n4655_ | ~new_n4695_;
  assign new_n6867_ = ~new_n15038_ | ~new_n5043_;
  assign new_n6868_ = ~new_n6867_ | ~new_n6866_ | ~new_n6865_;
  assign new_n6869_ = ~new_n5105_ | ~new_n7294_;
  assign new_n6870_ = ~new_n15038_ | ~new_n7293_;
  assign new_n6871_ = ~new_n5604_ | ~new_n6868_;
  assign new_n6872_ = ~new_n18611_ | ~new_n4648_;
  assign new_n6873_ = ~pi498 | ~po509;
  assign new_n6874_ = ~new_n4657_ | ~new_n4697_;
  assign new_n6875_ = ~new_n4655_ | ~new_n4691_;
  assign new_n6876_ = ~new_n15031_ | ~new_n5043_;
  assign new_n6877_ = ~new_n6876_ | ~new_n6875_ | ~new_n6874_;
  assign new_n6878_ = ~new_n4663_ | ~new_n5592_;
  assign new_n6879_ = ~new_n4662_ | ~new_n15031_;
  assign new_n6880_ = ~new_n5604_ | ~new_n6877_;
  assign new_n6881_ = ~new_n18699_ | ~new_n4648_;
  assign new_n6882_ = ~pi499 | ~po509;
  assign new_n6883_ = ~new_n5045_ | ~new_n5042_;
  assign new_n6884_ = ~new_n6883_ | ~new_n5043_;
  assign new_n6885_ = ~new_n5605_ | ~new_n6884_;
  assign new_n6886_ = ~new_n5509_ | ~new_n4655_;
  assign new_n6887_ = ~new_n5064_ | ~new_n7294_;
  assign new_n6888_ = ~pi500 | ~new_n6885_;
  assign new_n6889_ = ~new_n18686_ | ~new_n4648_;
  assign new_n6890_ = ~pi500 | ~po509;
  assign new_n6891_ = ~new_n4657_ | ~new_n4700_;
  assign new_n6892_ = ~new_n4655_ | ~new_n4678_;
  assign new_n6893_ = ~new_n15017_ | ~new_n5043_;
  assign new_n6894_ = ~new_n6893_ | ~new_n6892_ | ~new_n6891_;
  assign new_n6895_ = ~new_n5093_ | ~new_n7294_;
  assign new_n6896_ = ~new_n15017_ | ~new_n7293_;
  assign new_n6897_ = ~new_n5604_ | ~new_n6894_;
  assign new_n6898_ = ~new_n18687_ | ~new_n4648_;
  assign new_n6899_ = ~pi501 | ~po509;
  assign new_n6900_ = ~new_n4657_ | ~new_n4680_;
  assign new_n6901_ = ~new_n4655_ | ~new_n4683_;
  assign new_n6902_ = ~new_n15022_ | ~new_n5043_;
  assign new_n6903_ = ~new_n6902_ | ~new_n6901_ | ~new_n6900_;
  assign new_n6904_ = ~new_n5078_ | ~new_n7294_;
  assign new_n6905_ = ~new_n15022_ | ~new_n7293_;
  assign new_n6906_ = ~new_n5604_ | ~new_n6903_;
  assign new_n6907_ = ~new_n18691_ | ~new_n4648_;
  assign new_n6908_ = ~pi502 | ~po509;
  assign new_n6909_ = ~new_n4657_ | ~new_n4682_;
  assign new_n6910_ = ~new_n4655_ | ~new_n4674_;
  assign new_n6911_ = ~new_n15027_ | ~new_n5043_;
  assign new_n6912_ = ~new_n6910_ | ~new_n6911_ | ~new_n6909_;
  assign new_n6913_ = ~new_n4663_ | ~new_n5588_;
  assign new_n6914_ = ~new_n4662_ | ~new_n15027_;
  assign new_n6915_ = ~new_n5604_ | ~new_n6912_;
  assign new_n6916_ = ~new_n18696_ | ~new_n4648_;
  assign new_n6917_ = ~pi503 | ~po509;
  assign new_n6918_ = ~new_n4657_ | ~new_n4689_;
  assign new_n6919_ = ~new_n4655_ | ~new_n4698_;
  assign new_n6920_ = ~new_n15034_ | ~new_n5043_;
  assign new_n6921_ = ~new_n6920_ | ~new_n6919_ | ~new_n6918_;
  assign new_n6922_ = ~new_n5117_ | ~new_n7294_;
  assign new_n6923_ = ~new_n15034_ | ~new_n7293_;
  assign new_n6924_ = ~new_n5604_ | ~new_n6921_;
  assign new_n6925_ = ~new_n18612_ | ~new_n4648_;
  assign new_n6926_ = ~pi504 | ~po509;
  assign new_n6927_ = ~new_n4657_ | ~new_n4676_;
  assign new_n6928_ = ~new_n4655_ | ~new_n4687_;
  assign new_n6929_ = ~new_n15021_ | ~new_n5043_;
  assign new_n6930_ = ~new_n6929_ | ~new_n6928_ | ~new_n6927_;
  assign new_n6931_ = ~new_n5081_ | ~new_n7294_;
  assign new_n6932_ = ~new_n15021_ | ~new_n7293_;
  assign new_n6933_ = ~new_n5604_ | ~new_n6930_;
  assign new_n6934_ = ~new_n18690_ | ~new_n4648_;
  assign new_n6935_ = ~pi505 | ~po509;
  assign new_n6936_ = ~new_n4657_ | ~new_n4690_;
  assign new_n6937_ = ~new_n4655_ | ~new_n4685_;
  assign new_n6938_ = ~new_n15035_ | ~new_n5043_;
  assign new_n6939_ = ~new_n6938_ | ~new_n6937_ | ~new_n6936_;
  assign new_n6940_ = ~new_n5114_ | ~new_n7294_;
  assign new_n6941_ = ~new_n15035_ | ~new_n7293_;
  assign new_n6942_ = ~new_n5604_ | ~new_n6939_;
  assign new_n6943_ = ~new_n18703_ | ~new_n4648_;
  assign new_n6944_ = ~pi506 | ~po509;
  assign new_n6945_ = ~new_n4657_ | ~new_n4681_;
  assign new_n6946_ = ~new_n4655_ | ~new_n4673_;
  assign new_n6947_ = ~new_n15026_ | ~new_n5043_;
  assign new_n6948_ = ~new_n6946_ | ~new_n6947_ | ~new_n6945_;
  assign new_n6949_ = ~new_n4663_ | ~new_n5587_;
  assign new_n6950_ = ~new_n4662_ | ~new_n15026_;
  assign new_n6951_ = ~new_n5604_ | ~new_n6948_;
  assign new_n6952_ = ~new_n18695_ | ~new_n4648_;
  assign new_n6953_ = ~pi507 | ~po509;
  assign new_n6954_ = ~new_n4657_ | ~new_n4679_;
  assign new_n6955_ = ~new_n4655_ | ~new_n4696_;
  assign new_n6956_ = ~new_n15039_ | ~new_n5043_;
  assign new_n6957_ = ~new_n6956_ | ~new_n6955_ | ~new_n6954_;
  assign new_n6958_ = ~new_n5102_ | ~new_n7294_;
  assign new_n6959_ = ~new_n15039_ | ~new_n7293_;
  assign new_n6960_ = ~new_n5604_ | ~new_n6957_;
  assign new_n6961_ = ~new_n18706_ | ~new_n4648_;
  assign new_n6962_ = ~pi508 | ~po509;
  assign new_n6963_ = ~new_n4657_ | ~new_n4692_;
  assign new_n6964_ = ~new_n4655_ | ~new_n4677_;
  assign new_n6965_ = ~new_n15030_ | ~new_n5043_;
  assign new_n6966_ = ~new_n6965_ | ~new_n6964_ | ~new_n6963_;
  assign new_n6967_ = ~new_n4663_ | ~new_n5591_;
  assign new_n6968_ = ~new_n4662_ | ~new_n15030_;
  assign new_n6969_ = ~new_n5604_ | ~new_n6966_;
  assign new_n6970_ = ~new_n18613_ | ~new_n4648_;
  assign new_n6971_ = ~pi509 | ~po509;
  assign new_n6972_ = ~new_n4657_ | ~new_n4693_;
  assign new_n6973_ = ~new_n4655_ | ~new_n4684_;
  assign new_n6974_ = ~pi510 | ~new_n5043_;
  assign new_n6975_ = ~new_n6974_ | ~new_n6973_ | ~new_n6972_;
  assign new_n6976_ = ~new_n5069_ | ~new_n7294_;
  assign new_n6977_ = ~pi510 | ~new_n7293_;
  assign new_n6978_ = ~new_n5604_ | ~new_n6975_;
  assign new_n6979_ = ~new_n18700_ | ~new_n4648_;
  assign new_n6980_ = ~pi510 | ~po509;
  assign new_n6981_ = ~new_n4657_ | ~new_n4686_;
  assign new_n6982_ = ~new_n4655_ | ~new_n4699_;
  assign new_n6983_ = ~new_n15018_ | ~new_n5043_;
  assign new_n6984_ = ~new_n6983_ | ~new_n6982_ | ~new_n6981_;
  assign new_n6985_ = ~new_n5090_ | ~new_n7294_;
  assign new_n6986_ = ~new_n15018_ | ~new_n7293_;
  assign new_n6987_ = ~new_n5604_ | ~new_n6984_;
  assign new_n6988_ = ~new_n18688_ | ~new_n4648_;
  assign new_n6989_ = ~pi511 | ~po509;
  assign new_n6990_ = ~new_n4657_ | ~new_n4669_;
  assign new_n6991_ = ~new_n4655_ | ~new_n4671_;
  assign new_n6992_ = ~new_n15023_ | ~new_n5043_;
  assign new_n6993_ = ~new_n6990_ | ~new_n6991_ | ~new_n6992_;
  assign new_n6994_ = ~new_n4663_ | ~new_n5584_;
  assign new_n6995_ = ~new_n4662_ | ~new_n15023_;
  assign new_n6996_ = ~new_n5604_ | ~new_n6993_;
  assign new_n6997_ = ~new_n18693_ | ~new_n4648_;
  assign new_n6998_ = ~pi512 | ~po509;
  assign new_n6999_ = ~new_n4657_ | ~new_n4698_;
  assign new_n7000_ = ~new_n4655_ | ~new_n4692_;
  assign new_n7001_ = ~new_n15032_ | ~new_n5043_;
  assign new_n7002_ = ~new_n7001_ | ~new_n7000_ | ~new_n6999_;
  assign new_n7003_ = ~new_n5122_ | ~new_n7294_;
  assign new_n7004_ = ~new_n15032_ | ~new_n7293_;
  assign new_n7005_ = ~new_n5604_ | ~new_n7002_;
  assign new_n7006_ = ~new_n18701_ | ~new_n4648_;
  assign new_n7007_ = ~pi513 | ~po509;
  assign new_n7008_ = ~new_n4657_ | ~new_n4684_;
  assign new_n7009_ = ~new_n4655_ | ~new_n4676_;
  assign new_n7010_ = ~new_n14972_ | ~new_n5043_;
  assign new_n7011_ = ~new_n7010_ | ~new_n7009_ | ~new_n7008_;
  assign new_n7012_ = ~new_n5075_ | ~new_n7294_;
  assign new_n7013_ = ~new_n14972_ | ~new_n7293_;
  assign new_n7014_ = ~new_n5604_ | ~new_n7011_;
  assign new_n7015_ = ~new_n18615_ | ~new_n4648_;
  assign new_n7016_ = ~pi514 | ~po509;
  assign new_n7017_ = ~new_n4657_ | ~new_n4699_;
  assign new_n7018_ = ~new_n4655_ | ~new_n4679_;
  assign new_n7019_ = ~new_n15041_ | ~new_n5043_;
  assign new_n7020_ = ~new_n7019_ | ~new_n7018_ | ~new_n7017_;
  assign new_n7021_ = ~new_n5096_ | ~new_n7294_;
  assign new_n7022_ = ~new_n15041_ | ~new_n7293_;
  assign new_n7023_ = ~new_n5604_ | ~new_n7020_;
  assign new_n7024_ = ~new_n18708_ | ~new_n4648_;
  assign new_n7025_ = ~pi515 | ~po509;
  assign new_n7026_ = ~new_n4657_ | ~new_n4677_;
  assign new_n7027_ = ~new_n4655_ | ~new_n4681_;
  assign new_n7028_ = ~new_n15028_ | ~new_n5043_;
  assign new_n7029_ = ~new_n7027_ | ~new_n7028_ | ~new_n7026_;
  assign new_n7030_ = ~new_n4663_ | ~new_n5589_;
  assign new_n7031_ = ~new_n4662_ | ~new_n15028_;
  assign new_n7032_ = ~new_n5604_ | ~new_n7029_;
  assign new_n7033_ = ~new_n18697_ | ~new_n4648_;
  assign new_n7034_ = ~pi516 | ~po509;
  assign new_n7035_ = ~new_n4657_ | ~new_n4696_;
  assign new_n7036_ = ~new_n4655_ | ~new_n4690_;
  assign new_n7037_ = ~new_n15037_ | ~new_n5043_;
  assign new_n7038_ = ~new_n7037_ | ~new_n7036_ | ~new_n7035_;
  assign new_n7039_ = ~new_n5108_ | ~new_n7294_;
  assign new_n7040_ = ~new_n15037_ | ~new_n7293_;
  assign new_n7041_ = ~new_n5604_ | ~new_n7038_;
  assign new_n7042_ = ~new_n18705_ | ~new_n4648_;
  assign new_n7043_ = ~pi517 | ~po509;
  assign new_n7044_ = ~new_n4657_ | ~new_n4673_;
  assign new_n7045_ = ~new_n4655_ | ~new_n4670_;
  assign new_n7046_ = ~new_n15024_ | ~new_n5043_;
  assign new_n7047_ = ~new_n7045_ | ~new_n7046_ | ~new_n7044_;
  assign new_n7048_ = ~new_n4663_ | ~new_n5585_;
  assign new_n7049_ = ~new_n4662_ | ~new_n15024_;
  assign new_n7050_ = ~new_n5604_ | ~new_n7047_;
  assign new_n7051_ = ~new_n18694_ | ~new_n4648_;
  assign new_n7052_ = ~pi518 | ~po509;
  assign new_n7053_ = ~new_n4657_ | ~new_n4687_;
  assign new_n7054_ = ~new_n4655_ | ~new_n4700_;
  assign new_n7055_ = ~new_n15019_ | ~new_n5043_;
  assign new_n7056_ = ~new_n7055_ | ~new_n7054_ | ~new_n7053_;
  assign new_n7057_ = ~new_n5087_ | ~new_n7294_;
  assign new_n7058_ = ~new_n15019_ | ~new_n7293_;
  assign new_n7059_ = ~new_n5604_ | ~new_n7056_;
  assign new_n7060_ = ~new_n18616_ | ~new_n4648_;
  assign new_n7061_ = ~pi519 | ~po509;
  assign new_n7062_ = ~new_n5583_ | ~new_n4664_;
  assign new_n7063_ = ~new_n5052_ | ~new_n5525_;
  assign new_n7064_ = ~new_n5520_ | ~new_n4988_ | ~new_n4982_;
  assign new_n7065_ = ~new_n5047_;
  assign new_n7066_ = ~new_n5200_ | ~new_n5047_;
  assign new_n7067_ = ~new_n7333_ | ~new_n4699_;
  assign new_n7068_ = ~new_n5201_ | ~new_n5047_;
  assign new_n7069_ = ~new_n7333_ | ~new_n4700_;
  assign new_n7070_ = ~new_n5202_ | ~new_n5047_;
  assign new_n7071_ = ~new_n7333_ | ~new_n4686_;
  assign new_n7072_ = ~new_n5203_ | ~new_n5047_;
  assign new_n7073_ = ~new_n7333_ | ~new_n4687_;
  assign new_n7074_ = ~new_n5204_ | ~new_n5047_;
  assign new_n7075_ = ~new_n7333_ | ~new_n4683_;
  assign new_n7076_ = ~new_n5205_ | ~new_n5047_;
  assign new_n7077_ = ~new_n7333_ | ~new_n4676_;
  assign new_n7078_ = ~new_n5207_ | ~new_n5047_;
  assign new_n7079_ = ~new_n7333_ | ~new_n4672_;
  assign new_n7080_ = ~new_n5208_ | ~new_n5047_;
  assign new_n7081_ = ~new_n7333_ | ~new_n4675_;
  assign new_n7082_ = ~new_n5206_ | ~new_n5047_;
  assign new_n7083_ = ~new_n7333_ | ~new_n4680_;
  assign new_n7084_ = ~new_n5210_ | ~new_n5047_;
  assign new_n7085_ = ~new_n7333_ | ~new_n4671_;
  assign new_n7086_ = ~new_n5211_ | ~new_n5047_;
  assign new_n7087_ = ~new_n7333_ | ~new_n4670_;
  assign new_n7088_ = ~new_n5212_ | ~new_n5047_;
  assign new_n7089_ = ~new_n7333_ | ~new_n4669_;
  assign new_n7090_ = ~new_n5213_ | ~new_n5047_;
  assign new_n7091_ = ~new_n7333_ | ~new_n4673_;
  assign new_n7092_ = ~new_n5214_ | ~new_n5047_;
  assign new_n7093_ = ~new_n7333_ | ~new_n4674_;
  assign new_n7094_ = ~new_n5215_ | ~new_n5047_;
  assign new_n7095_ = ~new_n7333_ | ~new_n4681_;
  assign new_n7096_ = ~new_n5216_ | ~new_n5047_;
  assign new_n7097_ = ~new_n7333_ | ~new_n4682_;
  assign new_n7098_ = ~new_n5217_ | ~new_n5047_;
  assign new_n7099_ = ~new_n7333_ | ~new_n4677_;
  assign new_n7100_ = ~new_n5218_ | ~new_n5047_;
  assign new_n7101_ = ~new_n7333_ | ~new_n4691_;
  assign new_n7102_ = ~new_n5219_ | ~new_n5047_;
  assign new_n7103_ = ~new_n7333_ | ~new_n4692_;
  assign new_n7104_ = ~new_n7333_ | ~new_n4684_;
  assign new_n7105_ = ~new_n5221_ | ~new_n5047_;
  assign new_n7106_ = ~new_n7333_ | ~new_n4697_;
  assign new_n7107_ = ~new_n5222_ | ~new_n5047_;
  assign new_n7108_ = ~new_n7333_ | ~new_n4698_;
  assign new_n7109_ = ~new_n5223_ | ~new_n5047_;
  assign new_n7110_ = ~new_n7333_ | ~new_n4685_;
  assign new_n7111_ = ~new_n5224_ | ~new_n5047_;
  assign new_n7112_ = ~new_n7333_ | ~new_n4689_;
  assign new_n7113_ = ~new_n5225_ | ~new_n5047_;
  assign new_n7114_ = ~new_n7333_ | ~new_n4690_;
  assign new_n7115_ = ~new_n5226_ | ~new_n5047_;
  assign new_n7116_ = ~new_n7333_ | ~new_n4695_;
  assign new_n7117_ = ~new_n5227_ | ~new_n5047_;
  assign new_n7118_ = ~new_n7333_ | ~new_n4696_;
  assign new_n7119_ = ~new_n5228_ | ~new_n5047_;
  assign new_n7120_ = ~new_n7333_ | ~new_n4688_;
  assign new_n7121_ = ~new_n5229_ | ~new_n5047_;
  assign new_n7122_ = ~new_n7333_ | ~new_n4679_;
  assign new_n7123_ = ~new_n5230_ | ~new_n5047_;
  assign new_n7124_ = ~new_n7333_ | ~new_n4678_;
  assign new_n7125_ = ~new_n7333_ | ~new_n4694_;
  assign new_n7126_ = ~new_n7333_ | ~new_n4693_;
  assign new_n7127_ = ~new_n7324_ | ~new_n5061_;
  assign new_n7128_ = ~new_n5052_ | ~new_n7327_;
  assign new_n7129_ = ~new_n5522_ | ~new_n4984_ | ~new_n5566_;
  assign new_n7130_ = ~new_n5569_ | ~new_n5093_;
  assign new_n7131_ = ~new_n7129_ | ~new_n4699_;
  assign new_n7132_ = ~new_n5569_ | ~new_n5090_;
  assign new_n7133_ = ~new_n7129_ | ~new_n4700_;
  assign new_n7134_ = ~new_n5569_ | ~new_n5087_;
  assign new_n7135_ = ~new_n7129_ | ~new_n4686_;
  assign new_n7136_ = ~new_n5569_ | ~new_n5084_;
  assign new_n7137_ = ~new_n7129_ | ~new_n4687_;
  assign new_n7138_ = ~new_n5569_ | ~new_n5081_;
  assign new_n7139_ = ~new_n7129_ | ~new_n4683_;
  assign new_n7140_ = ~new_n5569_ | ~new_n5078_;
  assign new_n7141_ = ~new_n7129_ | ~new_n4676_;
  assign new_n7142_ = ~new_n7129_ | ~new_n4672_;
  assign new_n7143_ = ~new_n5569_ | ~new_n5593_;
  assign new_n7144_ = ~new_n7129_ | ~new_n4675_;
  assign new_n7145_ = ~new_n5569_ | ~new_n5075_;
  assign new_n7146_ = ~new_n7129_ | ~new_n4680_;
  assign new_n7147_ = ~new_n7129_ | ~new_n4671_;
  assign new_n7148_ = ~new_n5569_ | ~new_n5595_;
  assign new_n7149_ = ~new_n7129_ | ~new_n4670_;
  assign new_n7150_ = ~new_n5569_ | ~new_n5584_;
  assign new_n7151_ = ~new_n7129_ | ~new_n4669_;
  assign new_n7152_ = ~new_n5569_ | ~new_n5585_;
  assign new_n7153_ = ~new_n7129_ | ~new_n4673_;
  assign new_n7154_ = ~new_n5569_ | ~new_n5586_;
  assign new_n7155_ = ~new_n7129_ | ~new_n4674_;
  assign new_n7156_ = ~new_n5569_ | ~new_n5587_;
  assign new_n7157_ = ~new_n7129_ | ~new_n4681_;
  assign new_n7158_ = ~new_n5569_ | ~new_n5588_;
  assign new_n7159_ = ~new_n7129_ | ~new_n4682_;
  assign new_n7160_ = ~new_n5569_ | ~new_n5589_;
  assign new_n7161_ = ~new_n7129_ | ~new_n4677_;
  assign new_n7162_ = ~new_n5569_ | ~new_n5590_;
  assign new_n7163_ = ~new_n7129_ | ~new_n4691_;
  assign new_n7164_ = ~new_n5569_ | ~new_n5591_;
  assign new_n7165_ = ~new_n7129_ | ~new_n4692_;
  assign new_n7166_ = ~new_n5569_ | ~new_n5592_;
  assign new_n7167_ = ~new_n5569_ | ~new_n5072_;
  assign new_n7168_ = ~new_n7129_ | ~new_n4684_;
  assign new_n7169_ = ~new_n5569_ | ~new_n5122_;
  assign new_n7170_ = ~new_n7129_ | ~new_n4697_;
  assign new_n7171_ = ~new_n5569_ | ~new_n5120_;
  assign new_n7172_ = ~new_n7129_ | ~new_n4698_;
  assign new_n7173_ = ~new_n5569_ | ~new_n5117_;
  assign new_n7174_ = ~new_n7129_ | ~new_n4685_;
  assign new_n7175_ = ~new_n5569_ | ~new_n5114_;
  assign new_n7176_ = ~new_n7129_ | ~new_n4689_;
  assign new_n7177_ = ~new_n5569_ | ~new_n5111_;
  assign new_n7178_ = ~new_n7129_ | ~new_n4690_;
  assign new_n7179_ = ~new_n5569_ | ~new_n5108_;
  assign new_n7180_ = ~new_n7129_ | ~new_n4695_;
  assign new_n7181_ = ~new_n5569_ | ~new_n5105_;
  assign new_n7182_ = ~new_n7129_ | ~new_n4696_;
  assign new_n7183_ = ~new_n5569_ | ~new_n5102_;
  assign new_n7184_ = ~new_n7129_ | ~new_n4688_;
  assign new_n7185_ = ~new_n5569_ | ~new_n5099_;
  assign new_n7186_ = ~new_n7129_ | ~new_n4679_;
  assign new_n7187_ = ~new_n5569_ | ~new_n5096_;
  assign new_n7188_ = ~new_n7129_ | ~new_n4678_;
  assign new_n7189_ = ~new_n5569_ | ~new_n5069_;
  assign new_n7190_ = ~new_n7129_ | ~new_n4694_;
  assign new_n7191_ = ~new_n5569_ | ~new_n5064_;
  assign new_n7192_ = ~new_n7129_ | ~new_n4693_;
  assign new_n7193_ = ~new_n5093_ | ~new_n7129_;
  assign new_n7194_ = ~new_n5569_ | ~new_n4699_;
  assign new_n7195_ = ~new_n7317_ | ~new_n4700_;
  assign new_n7196_ = ~new_n5090_ | ~new_n7129_;
  assign new_n7197_ = ~new_n5569_ | ~new_n4700_;
  assign new_n7198_ = ~new_n7317_ | ~new_n4686_;
  assign new_n7199_ = ~new_n5087_ | ~new_n7129_;
  assign new_n7200_ = ~new_n5569_ | ~new_n4686_;
  assign new_n7201_ = ~new_n7317_ | ~new_n4687_;
  assign new_n7202_ = ~new_n5084_ | ~new_n7129_;
  assign new_n7203_ = ~new_n5569_ | ~new_n4687_;
  assign new_n7204_ = ~new_n7317_ | ~new_n4683_;
  assign new_n7205_ = ~new_n5081_ | ~new_n7129_;
  assign new_n7206_ = ~new_n5569_ | ~new_n4683_;
  assign new_n7207_ = ~new_n7317_ | ~new_n4676_;
  assign new_n7208_ = ~new_n5078_ | ~new_n7129_;
  assign new_n7209_ = ~new_n5569_ | ~new_n4676_;
  assign new_n7210_ = ~new_n7317_ | ~new_n4680_;
  assign new_n7211_ = ~new_n5593_ | ~new_n7129_;
  assign new_n7212_ = ~new_n5569_ | ~new_n4672_;
  assign new_n7213_ = ~new_n5594_ | ~new_n7129_;
  assign new_n7214_ = ~new_n5569_ | ~new_n4675_;
  assign new_n7215_ = ~new_n5075_ | ~new_n7129_;
  assign new_n7216_ = ~new_n5569_ | ~new_n4680_;
  assign new_n7217_ = ~new_n7317_ | ~new_n4684_;
  assign new_n7218_ = ~new_n5595_ | ~new_n7129_;
  assign new_n7219_ = ~new_n5569_ | ~new_n4671_;
  assign new_n7220_ = ~new_n7317_ | ~new_n4670_;
  assign new_n7221_ = ~new_n5584_ | ~new_n7129_;
  assign new_n7222_ = ~new_n5569_ | ~new_n4670_;
  assign new_n7223_ = ~new_n7317_ | ~new_n4669_;
  assign new_n7224_ = ~new_n5585_ | ~new_n7129_;
  assign new_n7225_ = ~new_n5569_ | ~new_n4669_;
  assign new_n7226_ = ~new_n7317_ | ~new_n4673_;
  assign new_n7227_ = ~new_n5586_ | ~new_n7129_;
  assign new_n7228_ = ~new_n5569_ | ~new_n4673_;
  assign new_n7229_ = ~new_n7317_ | ~new_n4674_;
  assign new_n7230_ = ~new_n5587_ | ~new_n7129_;
  assign new_n7231_ = ~new_n5569_ | ~new_n4674_;
  assign new_n7232_ = ~new_n7317_ | ~new_n4681_;
  assign new_n7233_ = ~new_n5588_ | ~new_n7129_;
  assign new_n7234_ = ~new_n5569_ | ~new_n4681_;
  assign new_n7235_ = ~new_n7317_ | ~new_n4682_;
  assign new_n7236_ = ~new_n5589_ | ~new_n7129_;
  assign new_n7237_ = ~new_n5569_ | ~new_n4682_;
  assign new_n7238_ = ~new_n7317_ | ~new_n4677_;
  assign new_n7239_ = ~new_n5590_ | ~new_n7129_;
  assign new_n7240_ = ~new_n5569_ | ~new_n4677_;
  assign new_n7241_ = ~new_n7317_ | ~new_n4691_;
  assign new_n7242_ = ~new_n5591_ | ~new_n7129_;
  assign new_n7243_ = ~new_n5569_ | ~new_n4691_;
  assign new_n7244_ = ~new_n7317_ | ~new_n4692_;
  assign new_n7245_ = ~new_n5592_ | ~new_n7129_;
  assign new_n7246_ = ~new_n5569_ | ~new_n4692_;
  assign new_n7247_ = ~new_n7317_ | ~new_n4697_;
  assign new_n7248_ = ~new_n5072_ | ~new_n7129_;
  assign new_n7249_ = ~new_n5569_ | ~new_n4684_;
  assign new_n7250_ = ~new_n7317_ | ~new_n4694_;
  assign new_n7251_ = ~new_n5122_ | ~new_n7129_;
  assign new_n7252_ = ~new_n5569_ | ~new_n4697_;
  assign new_n7253_ = ~new_n7317_ | ~new_n4698_;
  assign new_n7254_ = ~new_n5120_ | ~new_n7129_;
  assign new_n7255_ = ~new_n5569_ | ~new_n4698_;
  assign new_n7256_ = ~new_n7317_ | ~new_n4685_;
  assign new_n7257_ = ~new_n5117_ | ~new_n7129_;
  assign new_n7258_ = ~new_n5569_ | ~new_n4685_;
  assign new_n7259_ = ~new_n7317_ | ~new_n4689_;
  assign new_n7260_ = ~new_n5114_ | ~new_n7129_;
  assign new_n7261_ = ~new_n5569_ | ~new_n4689_;
  assign new_n7262_ = ~new_n7317_ | ~new_n4690_;
  assign new_n7263_ = ~new_n5111_ | ~new_n7129_;
  assign new_n7264_ = ~new_n5569_ | ~new_n4690_;
  assign new_n7265_ = ~new_n7317_ | ~new_n4695_;
  assign new_n7266_ = ~new_n5108_ | ~new_n7129_;
  assign new_n7267_ = ~new_n5569_ | ~new_n4695_;
  assign new_n7268_ = ~new_n7317_ | ~new_n4696_;
  assign new_n7269_ = ~new_n5105_ | ~new_n7129_;
  assign new_n7270_ = ~new_n5569_ | ~new_n4696_;
  assign new_n7271_ = ~new_n7317_ | ~new_n4688_;
  assign new_n7272_ = ~new_n5102_ | ~new_n7129_;
  assign new_n7273_ = ~new_n5569_ | ~new_n4688_;
  assign new_n7274_ = ~new_n7317_ | ~new_n4679_;
  assign new_n7275_ = ~new_n5099_ | ~new_n7129_;
  assign new_n7276_ = ~new_n5569_ | ~new_n4679_;
  assign new_n7277_ = ~new_n7317_ | ~new_n4678_;
  assign new_n7278_ = ~new_n5096_ | ~new_n7129_;
  assign new_n7279_ = ~new_n5569_ | ~new_n4678_;
  assign new_n7280_ = ~new_n7317_ | ~new_n4699_;
  assign new_n7281_ = ~new_n5069_ | ~new_n7129_;
  assign new_n7282_ = ~new_n5569_ | ~new_n4694_;
  assign new_n7283_ = ~new_n7317_ | ~new_n4693_;
  assign new_n7284_ = ~new_n5064_ | ~new_n7129_;
  assign new_n7285_ = ~new_n5569_ | ~new_n4693_;
  assign new_n7286_ = ~new_n5052_ | ~pi520;
  assign new_n7287_ = ~new_n5502_ | ~new_n6793_;
  assign new_n7288_ = ~new_n7144_ | ~new_n5029_;
  assign new_n7289_ = ~new_n5048_ | ~new_n7144_;
  assign new_n7290_ = ~new_n5031_;
  assign new_n7291_ = ~new_n5607_ | ~new_n5043_;
  assign new_n7292_ = ~new_n5581_ | ~new_n5607_;
  assign new_n7293_ = ~new_n7291_ | ~new_n5605_;
  assign new_n7294_ = ~new_n7292_ | ~new_n5606_;
  assign new_n7295_ = ~new_n7838_ | ~new_n7104_;
  assign new_n7296_ = ~new_n7861_ | ~new_n7125_;
  assign new_n7297_ = ~new_n7884_ | ~new_n7126_;
  assign new_n7298_ = ~new_n7065_ | ~new_n7125_;
  assign new_n7299_ = ~new_n7065_ | ~new_n7104_;
  assign new_n7300_ = ~new_n7065_ | ~new_n7126_;
  assign new_n7301_ = ~new_n7311_ | ~new_n7305_;
  assign new_n7302_ = ~new_n5052_ | ~new_n5525_;
  assign new_n7303_ = ~pi302 | ~new_n5523_;
  assign new_n7304_ = ~pi309 | ~new_n15383_;
  assign new_n7305_ = ~new_n5049_;
  assign new_n7306_ = ~pi303 | ~new_n5523_;
  assign new_n7307_ = ~pi309 | ~new_n15315_;
  assign new_n7308_ = ~new_n5050_;
  assign new_n7309_ = ~pi304 | ~new_n5523_;
  assign new_n7310_ = ~pi309 | ~new_n15316_;
  assign new_n7311_ = ~new_n5051_;
  assign new_n7312_ = ~new_n7305_ | ~pi490;
  assign new_n7313_ = ~new_n5049_ | ~new_n4976_;
  assign new_n7314_ = ~new_n7313_ | ~new_n7312_;
  assign new_n7315_ = ~pi301 | ~new_n5523_;
  assign new_n7316_ = ~pi309 | ~new_n15314_;
  assign new_n7317_ = ~new_n5052_;
  assign new_n7318_ = ~pi310 | ~new_n5524_;
  assign new_n7319_ = ~new_n5602_ | ~new_n5711_;
  assign new_n7320_ = ~pi311 | ~new_n5524_;
  assign new_n7321_ = ~new_n5602_ | ~new_n5712_;
  assign new_n7322_ = ~pi300 | ~new_n5523_;
  assign new_n7323_ = ~pi309 | ~new_n15313_;
  assign new_n7324_ = ~new_n5057_;
  assign new_n7325_ = ~pi297 | ~new_n5523_;
  assign new_n7326_ = ~pi309 | ~new_n15311_;
  assign new_n7327_ = ~new_n5061_;
  assign new_n7328_ = ~pi298 | ~new_n5523_;
  assign new_n7329_ = ~pi309 | ~new_n15312_;
  assign new_n7330_ = ~new_n5055_;
  assign new_n7331_ = ~pi299 | ~new_n5523_;
  assign new_n7332_ = ~pi309 | ~new_n15385_;
  assign new_n7333_ = ~new_n5056_;
  assign new_n7334_ = ~pi308 | ~new_n5523_;
  assign new_n7335_ = ~pi309 | ~new_n15372_;
  assign new_n7336_ = ~new_n5059_;
  assign new_n7337_ = ~pi307 | ~new_n5523_;
  assign new_n7338_ = ~pi309 | ~new_n15374_;
  assign new_n7339_ = ~new_n5058_;
  assign new_n7340_ = ~new_n7339_ | ~pi407 | ~new_n5059_;
  assign new_n7341_ = ~new_n5058_ | ~pi510 | ~new_n5059_;
  assign new_n7342_ = ~pi306 | ~new_n5523_;
  assign new_n7343_ = ~pi309 | ~new_n15377_;
  assign new_n7344_ = ~new_n5060_;
  assign new_n7345_ = ~pi278 | ~new_n5523_;
  assign new_n7346_ = ~pi309 | ~pi278;
  assign new_n7347_ = ~pi305 | ~new_n5523_;
  assign new_n7348_ = ~pi309 | ~new_n15380_;
  assign new_n7349_ = ~new_n5063_;
  assign new_n7350_ = ~new_n1070_ | ~new_n5525_;
  assign new_n7351_ = ~new_n5580_ | ~new_n5062_;
  assign new_n7352_ = ~new_n5064_;
  assign new_n7353_ = ~new_n5057_ | ~new_n7333_;
  assign new_n7354_ = ~new_n5055_ | ~new_n7324_;
  assign new_n7355_ = ~pi311 | ~new_n5710_;
  assign new_n7356_ = ~new_n5712_ | ~new_n4978_;
  assign new_n7357_ = ~new_n5066_;
  assign new_n7358_ = ~new_n7301_ | ~new_n4978_;
  assign new_n7359_ = ~pi310 | ~new_n5710_;
  assign new_n7360_ = ~new_n5065_;
  assign new_n7361_ = ~pi342 | ~new_n5526_;
  assign new_n7362_ = ~new_n5601_ | ~new_n5761_;
  assign new_n7363_ = ~new_n7339_ | ~pi406 | ~new_n5059_;
  assign new_n7364_ = ~new_n5058_ | ~pi500 | ~new_n5059_;
  assign new_n7365_ = ~pi279 | ~new_n5523_;
  assign new_n7366_ = ~pi309 | ~new_n15342_;
  assign new_n7367_ = ~new_n1059_ | ~new_n5525_;
  assign new_n7368_ = ~new_n5068_ | ~new_n5580_;
  assign new_n7369_ = ~new_n5069_;
  assign new_n7370_ = ~new_n7339_ | ~pi408 | ~new_n5059_;
  assign new_n7371_ = ~new_n5058_ | ~pi495 | ~new_n5059_;
  assign new_n7372_ = ~pi343 | ~new_n5526_;
  assign new_n7373_ = ~new_n5601_ | ~new_n5781_;
  assign new_n7374_ = ~pi280 | ~new_n5523_;
  assign new_n7375_ = ~pi309 | ~new_n15317_;
  assign new_n7376_ = ~new_n1048_ | ~new_n5525_;
  assign new_n7377_ = ~new_n5071_ | ~new_n5580_;
  assign new_n7378_ = ~new_n5072_;
  assign new_n7379_ = ~pi344 | ~new_n5526_;
  assign new_n7380_ = ~new_n5601_ | ~new_n5800_;
  assign new_n7381_ = ~pi281 | ~new_n5523_;
  assign new_n7382_ = ~pi309 | ~new_n15318_;
  assign new_n7383_ = ~new_n1045_ | ~new_n5525_;
  assign new_n7384_ = ~new_n5074_ | ~new_n5580_;
  assign new_n7385_ = ~new_n5075_;
  assign new_n7386_ = ~pi345 | ~new_n5526_;
  assign new_n7387_ = ~new_n5601_ | ~new_n5819_;
  assign new_n7388_ = ~pi282 | ~new_n5523_;
  assign new_n7389_ = ~pi309 | ~new_n15319_;
  assign new_n7390_ = ~new_n1044_ | ~new_n5525_;
  assign new_n7391_ = ~new_n5077_ | ~new_n5580_;
  assign new_n7392_ = ~new_n5078_;
  assign new_n7393_ = ~pi346 | ~new_n5526_;
  assign new_n7394_ = ~new_n5601_ | ~new_n5838_;
  assign new_n7395_ = ~pi283 | ~new_n5523_;
  assign new_n7396_ = ~pi309 | ~new_n15367_;
  assign new_n7397_ = ~new_n1043_ | ~new_n5525_;
  assign new_n7398_ = ~new_n5080_ | ~new_n5580_;
  assign new_n7399_ = ~new_n5081_;
  assign new_n7400_ = ~pi347 | ~new_n5526_;
  assign new_n7401_ = ~new_n5601_ | ~new_n5857_;
  assign new_n7402_ = ~pi284 | ~new_n5523_;
  assign new_n7403_ = ~pi309 | ~new_n15320_;
  assign new_n7404_ = ~new_n1042_ | ~new_n5525_;
  assign new_n7405_ = ~new_n5083_ | ~new_n5580_;
  assign new_n7406_ = ~new_n5084_;
  assign new_n7407_ = ~pi348 | ~new_n5526_;
  assign new_n7408_ = ~new_n5601_ | ~new_n5876_;
  assign new_n7409_ = ~pi285 | ~new_n5523_;
  assign new_n7410_ = ~pi309 | ~new_n15321_;
  assign new_n7411_ = ~new_n1041_ | ~new_n5525_;
  assign new_n7412_ = ~new_n5086_ | ~new_n5580_;
  assign new_n7413_ = ~new_n5087_;
  assign new_n7414_ = ~pi349 | ~new_n5526_;
  assign new_n7415_ = ~new_n5601_ | ~new_n5895_;
  assign new_n7416_ = ~pi286 | ~new_n5523_;
  assign new_n7417_ = ~pi309 | ~new_n15322_;
  assign new_n7418_ = ~new_n1040_ | ~new_n5525_;
  assign new_n7419_ = ~new_n5089_ | ~new_n5580_;
  assign new_n7420_ = ~new_n5090_;
  assign new_n7421_ = ~pi350 | ~new_n5526_;
  assign new_n7422_ = ~new_n5601_ | ~new_n5914_;
  assign new_n7423_ = ~pi287 | ~new_n5523_;
  assign new_n7424_ = ~pi309 | ~new_n15365_;
  assign new_n7425_ = ~new_n1039_ | ~new_n5525_;
  assign new_n7426_ = ~new_n5092_ | ~new_n5580_;
  assign new_n7427_ = ~new_n5093_;
  assign new_n7428_ = ~pi351 | ~new_n5526_;
  assign new_n7429_ = ~new_n5601_ | ~new_n5933_;
  assign new_n7430_ = ~pi288 | ~new_n5523_;
  assign new_n7431_ = ~pi309 | ~new_n15304_;
  assign new_n7432_ = ~new_n1069_ | ~new_n5525_;
  assign new_n7433_ = ~new_n5095_ | ~new_n5580_;
  assign new_n7434_ = ~new_n5096_;
  assign new_n7435_ = ~pi352 | ~new_n5526_;
  assign new_n7436_ = ~new_n5601_ | ~new_n5952_;
  assign new_n7437_ = ~pi289 | ~new_n5523_;
  assign new_n7438_ = ~pi309 | ~new_n15305_;
  assign new_n7439_ = ~new_n1068_ | ~new_n5525_;
  assign new_n7440_ = ~new_n5098_ | ~new_n5580_;
  assign new_n7441_ = ~new_n5099_;
  assign new_n7442_ = ~pi353 | ~new_n5526_;
  assign new_n7443_ = ~new_n5601_ | ~new_n5971_;
  assign new_n7444_ = ~pi290 | ~new_n5523_;
  assign new_n7445_ = ~pi309 | ~new_n15306_;
  assign new_n7446_ = ~new_n1067_ | ~new_n5525_;
  assign new_n7447_ = ~new_n5101_ | ~new_n5580_;
  assign new_n7448_ = ~new_n5102_;
  assign new_n7449_ = ~pi354 | ~new_n5526_;
  assign new_n7450_ = ~new_n5601_ | ~new_n5990_;
  assign new_n7451_ = ~pi291 | ~new_n5523_;
  assign new_n7452_ = ~pi309 | ~new_n15392_;
  assign new_n7453_ = ~new_n1066_ | ~new_n5525_;
  assign new_n7454_ = ~new_n5104_ | ~new_n5580_;
  assign new_n7455_ = ~new_n5105_;
  assign new_n7456_ = ~pi355 | ~new_n5526_;
  assign new_n7457_ = ~new_n5601_ | ~new_n6009_;
  assign new_n7458_ = ~pi292 | ~new_n5523_;
  assign new_n7459_ = ~pi309 | ~new_n15307_;
  assign new_n7460_ = ~new_n1065_ | ~new_n5525_;
  assign new_n7461_ = ~new_n5107_ | ~new_n5580_;
  assign new_n7462_ = ~new_n5108_;
  assign new_n7463_ = ~pi356 | ~new_n5526_;
  assign new_n7464_ = ~new_n5601_ | ~new_n6028_;
  assign new_n7465_ = ~pi293 | ~new_n5523_;
  assign new_n7466_ = ~pi309 | ~new_n15308_;
  assign new_n7467_ = ~new_n1064_ | ~new_n5525_;
  assign new_n7468_ = ~new_n5110_ | ~new_n5580_;
  assign new_n7469_ = ~new_n5111_;
  assign new_n7470_ = ~pi357 | ~new_n5526_;
  assign new_n7471_ = ~new_n5601_ | ~new_n6047_;
  assign new_n7472_ = ~pi294 | ~new_n5523_;
  assign new_n7473_ = ~pi309 | ~new_n15309_;
  assign new_n7474_ = ~new_n1063_ | ~new_n5525_;
  assign new_n7475_ = ~new_n5113_ | ~new_n5580_;
  assign new_n7476_ = ~new_n5114_;
  assign new_n7477_ = ~pi358 | ~new_n5526_;
  assign new_n7478_ = ~new_n5601_ | ~new_n6066_;
  assign new_n7479_ = ~pi295 | ~new_n5523_;
  assign new_n7480_ = ~pi309 | ~new_n15390_;
  assign new_n7481_ = ~new_n1062_ | ~new_n5525_;
  assign new_n7482_ = ~new_n5116_ | ~new_n5580_;
  assign new_n7483_ = ~new_n5117_;
  assign new_n7484_ = ~pi359 | ~new_n5526_;
  assign new_n7485_ = ~new_n5601_ | ~new_n6085_;
  assign new_n7486_ = ~pi296 | ~new_n5523_;
  assign new_n7487_ = ~pi309 | ~new_n15310_;
  assign new_n7488_ = ~new_n1061_ | ~new_n5525_;
  assign new_n7489_ = ~new_n5119_ | ~new_n5580_;
  assign new_n7490_ = ~new_n5120_;
  assign new_n7491_ = ~pi360 | ~new_n5526_;
  assign new_n7492_ = ~new_n5601_ | ~new_n6104_;
  assign new_n7493_ = ~new_n1060_ | ~new_n5525_;
  assign new_n7494_ = ~new_n5580_ | ~new_n5061_;
  assign new_n7495_ = ~new_n5122_;
  assign new_n7496_ = ~pi361 | ~new_n5526_;
  assign new_n7497_ = ~new_n5601_ | ~new_n6123_;
  assign new_n7498_ = ~pi362 | ~new_n5526_;
  assign new_n7499_ = ~new_n5601_ | ~new_n6142_;
  assign new_n7500_ = ~pi363 | ~new_n5526_;
  assign new_n7501_ = ~new_n5601_ | ~new_n6161_;
  assign new_n7502_ = ~pi364 | ~new_n5526_;
  assign new_n7503_ = ~new_n5601_ | ~new_n6180_;
  assign new_n7504_ = ~pi365 | ~new_n5526_;
  assign new_n7505_ = ~new_n5601_ | ~new_n6199_;
  assign new_n7506_ = ~pi366 | ~new_n5526_;
  assign new_n7507_ = ~new_n5601_ | ~new_n6218_;
  assign new_n7508_ = ~pi367 | ~new_n5526_;
  assign new_n7509_ = ~new_n5601_ | ~new_n6237_;
  assign new_n7510_ = ~pi368 | ~new_n5526_;
  assign new_n7511_ = ~new_n5601_ | ~new_n6256_;
  assign new_n7512_ = ~pi369 | ~new_n5526_;
  assign new_n7513_ = ~new_n5601_ | ~new_n6275_;
  assign new_n7514_ = ~pi370 | ~new_n5526_;
  assign new_n7515_ = ~new_n5601_ | ~new_n6294_;
  assign new_n7516_ = ~pi371 | ~new_n5526_;
  assign new_n7517_ = ~new_n5601_ | ~new_n6314_;
  assign new_n7518_ = ~pi372 | ~new_n5526_;
  assign new_n7519_ = ~new_n5601_ | ~new_n6321_;
  assign new_n7520_ = ~pi373 | ~new_n5526_;
  assign new_n7521_ = ~new_n5601_ | ~new_n6324_;
  assign new_n7522_ = ~pi374 | ~new_n5527_;
  assign new_n7523_ = ~new_n5600_ | ~new_n5761_;
  assign new_n7524_ = ~pi375 | ~new_n5527_;
  assign new_n7525_ = ~new_n5600_ | ~new_n5781_;
  assign new_n7526_ = ~pi376 | ~new_n5527_;
  assign new_n7527_ = ~new_n5600_ | ~new_n5800_;
  assign new_n7528_ = ~pi377 | ~new_n5527_;
  assign new_n7529_ = ~new_n5600_ | ~new_n5819_;
  assign new_n7530_ = ~pi378 | ~new_n5527_;
  assign new_n7531_ = ~new_n5600_ | ~new_n5838_;
  assign new_n7532_ = ~pi379 | ~new_n5527_;
  assign new_n7533_ = ~new_n5600_ | ~new_n5857_;
  assign new_n7534_ = ~pi380 | ~new_n5527_;
  assign new_n7535_ = ~new_n5600_ | ~new_n5876_;
  assign new_n7536_ = ~pi381 | ~new_n5527_;
  assign new_n7537_ = ~new_n5600_ | ~new_n5895_;
  assign new_n7538_ = ~pi382 | ~new_n5527_;
  assign new_n7539_ = ~new_n5600_ | ~new_n5914_;
  assign new_n7540_ = ~pi383 | ~new_n5527_;
  assign new_n7541_ = ~new_n5600_ | ~new_n5933_;
  assign new_n7542_ = ~pi384 | ~new_n5527_;
  assign new_n7543_ = ~new_n5600_ | ~new_n5952_;
  assign new_n7544_ = ~pi385 | ~new_n5527_;
  assign new_n7545_ = ~new_n5600_ | ~new_n5971_;
  assign new_n7546_ = ~pi386 | ~new_n5527_;
  assign new_n7547_ = ~new_n5600_ | ~new_n5990_;
  assign new_n7548_ = ~pi387 | ~new_n5527_;
  assign new_n7549_ = ~new_n5600_ | ~new_n6009_;
  assign new_n7550_ = ~pi388 | ~new_n5527_;
  assign new_n7551_ = ~new_n5600_ | ~new_n6028_;
  assign new_n7552_ = ~pi389 | ~new_n5527_;
  assign new_n7553_ = ~new_n5600_ | ~new_n6047_;
  assign new_n7554_ = ~pi390 | ~new_n5527_;
  assign new_n7555_ = ~new_n5600_ | ~new_n6066_;
  assign new_n7556_ = ~pi391 | ~new_n5527_;
  assign new_n7557_ = ~new_n5600_ | ~new_n6085_;
  assign new_n7558_ = ~pi392 | ~new_n5527_;
  assign new_n7559_ = ~new_n5600_ | ~new_n6104_;
  assign new_n7560_ = ~pi393 | ~new_n5527_;
  assign new_n7561_ = ~new_n5600_ | ~new_n6123_;
  assign new_n7562_ = ~pi394 | ~new_n5527_;
  assign new_n7563_ = ~new_n5600_ | ~new_n6142_;
  assign new_n7564_ = ~pi395 | ~new_n5527_;
  assign new_n7565_ = ~new_n5600_ | ~new_n6161_;
  assign new_n7566_ = ~pi396 | ~new_n5527_;
  assign new_n7567_ = ~new_n5600_ | ~new_n6180_;
  assign new_n7568_ = ~pi397 | ~new_n5527_;
  assign new_n7569_ = ~new_n5600_ | ~new_n6199_;
  assign new_n7570_ = ~pi398 | ~new_n5527_;
  assign new_n7571_ = ~new_n5600_ | ~new_n6218_;
  assign new_n7572_ = ~pi399 | ~new_n5527_;
  assign new_n7573_ = ~new_n5600_ | ~new_n6237_;
  assign new_n7574_ = ~pi400 | ~new_n5527_;
  assign new_n7575_ = ~new_n5600_ | ~new_n6256_;
  assign new_n7576_ = ~pi401 | ~new_n5527_;
  assign new_n7577_ = ~new_n5600_ | ~new_n6275_;
  assign new_n7578_ = ~pi402 | ~new_n5527_;
  assign new_n7579_ = ~new_n5600_ | ~new_n6294_;
  assign new_n7580_ = ~pi403 | ~new_n5527_;
  assign new_n7581_ = ~new_n5600_ | ~new_n6314_;
  assign new_n7582_ = ~pi404 | ~new_n5527_;
  assign new_n7583_ = ~new_n5600_ | ~new_n6321_;
  assign new_n7584_ = ~pi405 | ~new_n5527_;
  assign new_n7585_ = ~new_n5600_ | ~new_n6324_;
  assign new_n7586_ = ~pi406 | ~new_n5033_;
  assign new_n7587_ = ~new_n5599_ | ~new_n4989_;
  assign new_n7588_ = ~pi407 | ~new_n5033_;
  assign new_n7589_ = ~new_n5599_ | ~new_n4990_;
  assign new_n7590_ = ~pi408 | ~new_n5033_;
  assign new_n7591_ = ~new_n5599_ | ~new_n4991_;
  assign new_n7592_ = ~pi409 | ~new_n5033_;
  assign new_n7593_ = ~new_n5599_ | ~new_n4992_;
  assign new_n7594_ = ~pi410 | ~new_n5033_;
  assign new_n7595_ = ~new_n5599_ | ~new_n4993_;
  assign new_n7596_ = ~pi411 | ~new_n5033_;
  assign new_n7597_ = ~new_n5599_ | ~new_n4994_;
  assign new_n7598_ = ~pi412 | ~new_n5033_;
  assign new_n7599_ = ~new_n5599_ | ~new_n4995_;
  assign new_n7600_ = ~pi413 | ~new_n5033_;
  assign new_n7601_ = ~new_n5599_ | ~new_n4996_;
  assign new_n7602_ = ~pi414 | ~new_n5033_;
  assign new_n7603_ = ~new_n5599_ | ~new_n4997_;
  assign new_n7604_ = ~pi415 | ~new_n5033_;
  assign new_n7605_ = ~new_n5599_ | ~new_n4998_;
  assign new_n7606_ = ~pi416 | ~new_n5033_;
  assign new_n7607_ = ~new_n5599_ | ~new_n4999_;
  assign new_n7608_ = ~pi417 | ~new_n5033_;
  assign new_n7609_ = ~new_n5599_ | ~new_n5000_;
  assign new_n7610_ = ~pi418 | ~new_n5033_;
  assign new_n7611_ = ~new_n5599_ | ~new_n5001_;
  assign new_n7612_ = ~pi419 | ~new_n5033_;
  assign new_n7613_ = ~new_n5599_ | ~new_n5002_;
  assign new_n7614_ = ~pi420 | ~new_n5033_;
  assign new_n7615_ = ~new_n5599_ | ~new_n5003_;
  assign new_n7616_ = ~pi421 | ~new_n5033_;
  assign new_n7617_ = ~new_n5599_ | ~new_n5004_;
  assign new_n7618_ = ~pi422 | ~new_n5033_;
  assign new_n7619_ = ~new_n5599_ | ~new_n5005_;
  assign new_n7620_ = ~pi423 | ~new_n5033_;
  assign new_n7621_ = ~new_n5599_ | ~new_n5006_;
  assign new_n7622_ = ~pi424 | ~new_n5033_;
  assign new_n7623_ = ~new_n5599_ | ~new_n5007_;
  assign new_n7624_ = ~pi425 | ~new_n5033_;
  assign new_n7625_ = ~new_n5599_ | ~new_n5008_;
  assign new_n7626_ = ~pi426 | ~new_n5033_;
  assign new_n7627_ = ~new_n5599_ | ~new_n5010_;
  assign new_n7628_ = ~pi427 | ~new_n5033_;
  assign new_n7629_ = ~new_n5599_ | ~new_n5012_;
  assign new_n7630_ = ~pi428 | ~new_n5033_;
  assign new_n7631_ = ~new_n5599_ | ~new_n5014_;
  assign new_n7632_ = ~pi429 | ~new_n5033_;
  assign new_n7633_ = ~new_n5599_ | ~new_n5016_;
  assign new_n7634_ = ~pi430 | ~new_n5033_;
  assign new_n7635_ = ~new_n5599_ | ~new_n5018_;
  assign new_n7636_ = ~pi431 | ~new_n5033_;
  assign new_n7637_ = ~new_n5599_ | ~new_n5020_;
  assign new_n7638_ = ~pi432 | ~new_n5033_;
  assign new_n7639_ = ~new_n5599_ | ~new_n5022_;
  assign new_n7640_ = ~pi433 | ~new_n5033_;
  assign new_n7641_ = ~new_n5599_ | ~new_n5024_;
  assign new_n7642_ = ~pi434 | ~new_n5033_;
  assign new_n7643_ = ~new_n5599_ | ~new_n5026_;
  assign new_n7644_ = ~pi435 | ~new_n5033_;
  assign new_n7645_ = ~new_n5599_ | ~new_n5028_;
  assign new_n7646_ = ~pi436 | ~new_n5033_;
  assign new_n7647_ = ~new_n5603_ | ~new_n5599_;
  assign new_n7648_ = ~pi437 | ~new_n5033_;
  assign new_n7649_ = ~new_n5603_ | ~new_n5599_;
  assign new_n7650_ = ~pi458 | ~new_n5039_;
  assign new_n7651_ = ~po511 | ~new_n4693_;
  assign new_n7652_ = ~pi459 | ~new_n5039_;
  assign new_n7653_ = ~po511 | ~new_n4694_;
  assign new_n7654_ = ~pi460 | ~new_n5039_;
  assign new_n7655_ = ~po511 | ~new_n4684_;
  assign new_n7656_ = ~pi461 | ~new_n5039_;
  assign new_n7657_ = ~po511 | ~new_n4680_;
  assign new_n7658_ = ~pi462 | ~new_n5039_;
  assign new_n7659_ = ~po511 | ~new_n4676_;
  assign new_n7660_ = ~pi463 | ~new_n5039_;
  assign new_n7661_ = ~po511 | ~new_n4683_;
  assign new_n7662_ = ~pi464 | ~new_n5039_;
  assign new_n7663_ = ~po511 | ~new_n4687_;
  assign new_n7664_ = ~pi465 | ~new_n5039_;
  assign new_n7665_ = ~po511 | ~new_n4686_;
  assign new_n7666_ = ~pi466 | ~new_n5039_;
  assign new_n7667_ = ~po511 | ~new_n4700_;
  assign new_n7668_ = ~pi467 | ~new_n5039_;
  assign new_n7669_ = ~po511 | ~new_n4699_;
  assign new_n7670_ = ~pi468 | ~new_n5039_;
  assign new_n7671_ = ~po511 | ~new_n4678_;
  assign new_n7672_ = ~pi469 | ~new_n5039_;
  assign new_n7673_ = ~po511 | ~new_n4679_;
  assign new_n7674_ = ~pi470 | ~new_n5039_;
  assign new_n7675_ = ~po511 | ~new_n4688_;
  assign new_n7676_ = ~pi471 | ~new_n5039_;
  assign new_n7677_ = ~po511 | ~new_n4696_;
  assign new_n7678_ = ~pi472 | ~new_n5039_;
  assign new_n7679_ = ~po511 | ~new_n4695_;
  assign new_n7680_ = ~pi473 | ~new_n5039_;
  assign new_n7681_ = ~po511 | ~new_n4690_;
  assign new_n7682_ = ~pi474 | ~new_n5039_;
  assign new_n7683_ = ~po511 | ~new_n4689_;
  assign new_n7684_ = ~pi475 | ~new_n5039_;
  assign new_n7685_ = ~po511 | ~new_n4685_;
  assign new_n7686_ = ~pi476 | ~new_n5039_;
  assign new_n7687_ = ~po511 | ~new_n4698_;
  assign new_n7688_ = ~pi477 | ~new_n5039_;
  assign new_n7689_ = ~po511 | ~new_n4697_;
  assign new_n7690_ = ~pi478 | ~new_n5039_;
  assign new_n7691_ = ~po511 | ~new_n4692_;
  assign new_n7692_ = ~pi479 | ~new_n5039_;
  assign new_n7693_ = ~po511 | ~new_n4691_;
  assign new_n7694_ = ~pi480 | ~new_n5039_;
  assign new_n7695_ = ~po511 | ~new_n4677_;
  assign new_n7696_ = ~pi481 | ~new_n5039_;
  assign new_n7697_ = ~po511 | ~new_n4682_;
  assign new_n7698_ = ~pi482 | ~new_n5039_;
  assign new_n7699_ = ~po511 | ~new_n4681_;
  assign new_n7700_ = ~pi483 | ~new_n5039_;
  assign new_n7701_ = ~po511 | ~new_n4674_;
  assign new_n7702_ = ~pi484 | ~new_n5039_;
  assign new_n7703_ = ~po511 | ~new_n4673_;
  assign new_n7704_ = ~pi485 | ~new_n5039_;
  assign new_n7705_ = ~po511 | ~new_n4669_;
  assign new_n7706_ = ~pi486 | ~new_n5039_;
  assign new_n7707_ = ~po511 | ~new_n4670_;
  assign new_n7708_ = ~pi487 | ~new_n5039_;
  assign new_n7709_ = ~po511 | ~new_n4671_;
  assign new_n7710_ = ~pi488 | ~new_n5039_;
  assign new_n7711_ = ~po511 | ~new_n4675_;
  assign new_n7712_ = ~pi489 | ~new_n5039_;
  assign new_n7713_ = ~po511 | ~new_n4672_;
  assign new_n7714_ = ~new_n7324_ | ~new_n15125_;
  assign new_n7715_ = ~new_n16447_ | ~new_n5057_;
  assign new_n7716_ = ~new_n7317_ | ~new_n5041_;
  assign new_n7717_ = ~new_n5057_ | ~new_n5052_;
  assign new_n7718_ = ~new_n15484_ | ~new_n6785_;
  assign new_n7719_ = ~new_n5561_ | ~new_n7330_ | ~new_n6786_;
  assign new_n7720_ = ~new_n5595_ | ~new_n4671_;
  assign new_n7721_ = ~new_n5027_ | ~new_n6280_;
  assign new_n7722_ = ~new_n7721_ | ~new_n7720_;
  assign new_n7723_ = ~new_n5584_ | ~new_n4670_;
  assign new_n7724_ = ~new_n5025_ | ~new_n6261_;
  assign new_n7725_ = ~new_n7724_ | ~new_n7723_;
  assign new_n7726_ = ~new_n5585_ | ~new_n4669_;
  assign new_n7727_ = ~new_n5023_ | ~new_n6242_;
  assign new_n7728_ = ~new_n7727_ | ~new_n7726_;
  assign new_n7729_ = ~new_n5588_ | ~new_n4681_;
  assign new_n7730_ = ~new_n5017_ | ~new_n6185_;
  assign new_n7731_ = ~new_n7730_ | ~new_n7729_;
  assign new_n7732_ = ~new_n5589_ | ~new_n4682_;
  assign new_n7733_ = ~new_n5015_ | ~new_n6166_;
  assign new_n7734_ = ~new_n7733_ | ~new_n7732_;
  assign new_n7735_ = ~new_n5591_ | ~new_n4691_;
  assign new_n7736_ = ~new_n5011_ | ~new_n6128_;
  assign new_n7737_ = ~new_n7736_ | ~new_n7735_;
  assign new_n7738_ = ~new_n5590_ | ~new_n4677_;
  assign new_n7739_ = ~new_n5013_ | ~new_n6147_;
  assign new_n7740_ = ~new_n7739_ | ~new_n7738_;
  assign new_n7741_ = ~new_n5587_ | ~new_n4674_;
  assign new_n7742_ = ~new_n5019_ | ~new_n6204_;
  assign new_n7743_ = ~new_n7742_ | ~new_n7741_;
  assign new_n7744_ = ~new_n5586_ | ~new_n4673_;
  assign new_n7745_ = ~new_n5021_ | ~new_n6223_;
  assign new_n7746_ = ~new_n7745_ | ~new_n7744_;
  assign new_n7747_ = ~new_n5594_ | ~new_n4675_;
  assign new_n7748_ = ~new_n5029_ | ~new_n6298_;
  assign new_n7749_ = ~new_n7748_ | ~new_n7747_;
  assign new_n7750_ = ~new_n5593_ | ~new_n4672_;
  assign new_n7751_ = ~new_n5030_ | ~new_n6318_;
  assign new_n7752_ = ~new_n7751_ | ~new_n7750_;
  assign new_n7753_ = ~new_n7483_ | ~new_n6052_;
  assign new_n7754_ = ~new_n5117_ | ~new_n4685_;
  assign new_n7755_ = ~new_n7754_ | ~new_n7753_;
  assign new_n7756_ = ~new_n7462_ | ~new_n5995_;
  assign new_n7757_ = ~new_n5108_ | ~new_n4695_;
  assign new_n7758_ = ~new_n7757_ | ~new_n7756_;
  assign new_n7759_ = ~new_n7369_ | ~new_n5746_;
  assign new_n7760_ = ~new_n5069_ | ~new_n4694_;
  assign new_n7761_ = ~new_n7760_ | ~new_n7759_;
  assign new_n7762_ = ~new_n7352_ | ~new_n5767_;
  assign new_n7763_ = ~new_n5064_ | ~new_n4693_;
  assign new_n7764_ = ~new_n7763_ | ~new_n7762_;
  assign new_n7765_ = ~new_n7469_ | ~new_n6014_;
  assign new_n7766_ = ~new_n5111_ | ~new_n4690_;
  assign new_n7767_ = ~new_n7766_ | ~new_n7765_;
  assign new_n7768_ = ~new_n7420_ | ~new_n5881_;
  assign new_n7769_ = ~new_n5090_ | ~new_n4700_;
  assign new_n7770_ = ~new_n7769_ | ~new_n7768_;
  assign new_n7771_ = ~new_n7427_ | ~new_n5900_;
  assign new_n7772_ = ~new_n5093_ | ~new_n4699_;
  assign new_n7773_ = ~new_n7772_ | ~new_n7771_;
  assign new_n7774_ = ~new_n7455_ | ~new_n5976_;
  assign new_n7775_ = ~new_n5105_ | ~new_n4696_;
  assign new_n7776_ = ~new_n7775_ | ~new_n7774_;
  assign new_n7777_ = ~new_n7476_ | ~new_n6033_;
  assign new_n7778_ = ~new_n5114_ | ~new_n4689_;
  assign new_n7779_ = ~new_n7778_ | ~new_n7777_;
  assign new_n7780_ = ~new_n7406_ | ~new_n5843_;
  assign new_n7781_ = ~new_n5084_ | ~new_n4687_;
  assign new_n7782_ = ~new_n7781_ | ~new_n7780_;
  assign new_n7783_ = ~new_n7413_ | ~new_n5862_;
  assign new_n7784_ = ~new_n5087_ | ~new_n4686_;
  assign new_n7785_ = ~new_n7784_ | ~new_n7783_;
  assign new_n7786_ = ~new_n7448_ | ~new_n5957_;
  assign new_n7787_ = ~new_n5102_ | ~new_n4688_;
  assign new_n7788_ = ~new_n7787_ | ~new_n7786_;
  assign new_n7789_ = ~new_n7399_ | ~new_n5824_;
  assign new_n7790_ = ~new_n5081_ | ~new_n4683_;
  assign new_n7791_ = ~new_n7790_ | ~new_n7789_;
  assign new_n7792_ = ~new_n7385_ | ~new_n5786_;
  assign new_n7793_ = ~new_n5075_ | ~new_n4680_;
  assign new_n7794_ = ~new_n7793_ | ~new_n7792_;
  assign new_n7795_ = ~new_n7378_ | ~new_n5764_;
  assign new_n7796_ = ~new_n5072_ | ~new_n4684_;
  assign new_n7797_ = ~new_n7796_ | ~new_n7795_;
  assign new_n7798_ = ~new_n7490_ | ~new_n6071_;
  assign new_n7799_ = ~new_n5120_ | ~new_n4698_;
  assign new_n7800_ = ~new_n7799_ | ~new_n7798_;
  assign new_n7801_ = ~new_n7495_ | ~new_n6090_;
  assign new_n7802_ = ~new_n5122_ | ~new_n4697_;
  assign new_n7803_ = ~new_n7802_ | ~new_n7801_;
  assign new_n7804_ = ~new_n7392_ | ~new_n5805_;
  assign new_n7805_ = ~new_n5078_ | ~new_n4676_;
  assign new_n7806_ = ~new_n7805_ | ~new_n7804_;
  assign new_n7807_ = ~new_n7441_ | ~new_n5938_;
  assign new_n7808_ = ~new_n5099_ | ~new_n4679_;
  assign new_n7809_ = ~new_n7808_ | ~new_n7807_;
  assign new_n7810_ = ~new_n7434_ | ~new_n5919_;
  assign new_n7811_ = ~new_n5096_ | ~new_n4678_;
  assign new_n7812_ = ~new_n7811_ | ~new_n7810_;
  assign new_n7813_ = ~new_n5592_ | ~new_n4692_;
  assign new_n7814_ = ~new_n5009_ | ~new_n6109_;
  assign new_n7815_ = ~new_n7814_ | ~new_n7813_;
  assign new_n7816_ = ~new_n4635_ | ~new_n5563_;
  assign new_n7817_ = ~new_n6784_ | ~new_n5578_;
  assign new_n7818_ = ~new_n4699_ | ~new_n15467_;
  assign new_n7819_ = ~new_n4699_ | ~new_n5564_;
  assign new_n7820_ = ~new_n4700_ | ~new_n15467_;
  assign new_n7821_ = ~new_n4700_ | ~new_n5564_;
  assign new_n7822_ = ~new_n4686_ | ~new_n15467_;
  assign new_n7823_ = ~new_n4686_ | ~new_n5564_;
  assign new_n7824_ = ~new_n4687_ | ~new_n15467_;
  assign new_n7825_ = ~new_n4687_ | ~new_n5564_;
  assign new_n7826_ = ~new_n4683_ | ~new_n15467_;
  assign new_n7827_ = ~new_n4683_ | ~new_n5564_;
  assign new_n7828_ = ~new_n4676_ | ~new_n15467_;
  assign new_n7829_ = ~new_n4676_ | ~new_n5564_;
  assign new_n7830_ = ~new_n4680_ | ~new_n15467_;
  assign new_n7831_ = ~new_n4680_ | ~new_n5564_;
  assign new_n7832_ = ~new_n15675_ | ~new_n15467_;
  assign new_n7833_ = ~new_n4672_ | ~new_n5564_;
  assign new_n7834_ = ~new_n15673_ | ~new_n15467_;
  assign new_n7835_ = ~new_n4675_ | ~new_n5564_;
  assign new_n7836_ = ~new_n4684_ | ~new_n15467_;
  assign new_n7837_ = ~new_n4684_ | ~new_n5564_;
  assign new_n7838_ = ~new_n5209_;
  assign new_n7839_ = ~new_n4671_ | ~new_n15467_;
  assign new_n7840_ = ~new_n4671_ | ~new_n5564_;
  assign new_n7841_ = ~new_n4670_ | ~new_n15467_;
  assign new_n7842_ = ~new_n4670_ | ~new_n5564_;
  assign new_n7843_ = ~new_n4669_ | ~new_n15467_;
  assign new_n7844_ = ~new_n4669_ | ~new_n5564_;
  assign new_n7845_ = ~new_n4673_ | ~new_n15467_;
  assign new_n7846_ = ~new_n4673_ | ~new_n5564_;
  assign new_n7847_ = ~new_n4674_ | ~new_n15467_;
  assign new_n7848_ = ~new_n4674_ | ~new_n5564_;
  assign new_n7849_ = ~new_n4681_ | ~new_n15467_;
  assign new_n7850_ = ~new_n4681_ | ~new_n5564_;
  assign new_n7851_ = ~new_n4682_ | ~new_n15467_;
  assign new_n7852_ = ~new_n4682_ | ~new_n5564_;
  assign new_n7853_ = ~new_n4677_ | ~new_n15467_;
  assign new_n7854_ = ~new_n4677_ | ~new_n5564_;
  assign new_n7855_ = ~new_n4691_ | ~new_n15467_;
  assign new_n7856_ = ~new_n4691_ | ~new_n5564_;
  assign new_n7857_ = ~new_n4692_ | ~new_n15467_;
  assign new_n7858_ = ~new_n4692_ | ~new_n5564_;
  assign new_n7859_ = ~new_n4694_ | ~new_n15467_;
  assign new_n7860_ = ~new_n4694_ | ~new_n5564_;
  assign new_n7861_ = ~new_n5220_;
  assign new_n7862_ = ~new_n4697_ | ~new_n15467_;
  assign new_n7863_ = ~new_n4697_ | ~new_n5564_;
  assign new_n7864_ = ~new_n4698_ | ~new_n15467_;
  assign new_n7865_ = ~new_n4698_ | ~new_n5564_;
  assign new_n7866_ = ~new_n4685_ | ~new_n15467_;
  assign new_n7867_ = ~new_n4685_ | ~new_n5564_;
  assign new_n7868_ = ~new_n4689_ | ~new_n15467_;
  assign new_n7869_ = ~new_n4689_ | ~new_n5564_;
  assign new_n7870_ = ~new_n4690_ | ~new_n15467_;
  assign new_n7871_ = ~new_n4690_ | ~new_n5564_;
  assign new_n7872_ = ~new_n4695_ | ~new_n15467_;
  assign new_n7873_ = ~new_n4695_ | ~new_n5564_;
  assign new_n7874_ = ~new_n4696_ | ~new_n15467_;
  assign new_n7875_ = ~new_n4696_ | ~new_n5564_;
  assign new_n7876_ = ~new_n4688_ | ~new_n15467_;
  assign new_n7877_ = ~new_n4688_ | ~new_n5564_;
  assign new_n7878_ = ~new_n4679_ | ~new_n15467_;
  assign new_n7879_ = ~new_n4679_ | ~new_n5564_;
  assign new_n7880_ = ~new_n4678_ | ~new_n15467_;
  assign new_n7881_ = ~new_n4678_ | ~new_n5564_;
  assign new_n7882_ = ~new_n4693_ | ~new_n15467_;
  assign new_n7883_ = ~new_n4693_ | ~new_n5564_;
  assign new_n7884_ = ~new_n5231_;
  assign new_n7885_ = ~new_n5061_ | ~new_n7333_;
  assign new_n7886_ = ~new_n5056_ | ~new_n5055_;
  assign new_n7887_ = ~new_n20918_ | ~new_n7888_;
  assign new_n7888_ = ~new_n20782_;
  assign new_n7889_ = ~new_n4697_ | ~new_n20709_;
  assign new_n7890_ = ~new_n5122_ | ~new_n20710_;
  assign new_n7891_ = ~new_n20781_ | ~new_n20810_;
  assign new_n7892_ = ~new_n20838_ | ~new_n7893_;
  assign new_n7893_ = ~new_n20781_;
  assign new_n7894_ = ~new_n4694_ | ~new_n20809_;
  assign new_n7895_ = ~new_n5069_ | ~new_n20668_;
  assign new_n7896_ = ~new_n20780_ | ~new_n20808_;
  assign new_n7897_ = ~new_n20922_ | ~new_n7898_;
  assign new_n7898_ = ~new_n20780_;
  assign new_n7899_ = ~new_n4692_ | ~new_n20711_;
  assign new_n7900_ = ~new_n5592_ | ~new_n20712_;
  assign new_n7901_ = ~new_n20926_ | ~new_n20806_;
  assign new_n7902_ = ~new_n20968_ | ~new_n20807_;
  assign new_n7903_ = ~new_n4691_ | ~new_n20714_;
  assign new_n7904_ = ~new_n5591_ | ~new_n20717_;
  assign new_n7905_ = ~new_n20805_ | ~new_n20959_;
  assign new_n7906_ = ~new_n20967_ | ~new_n20730_;
  assign new_n7907_ = ~pi193;
  assign po000 = new_n8063_ & new_n8059_;
  assign po018 = ~new_n8064_ | ~new_n8125_ | ~new_n8124_;
  assign new_n7910_ = ~pi212;
  assign new_n7911_ = ~pi457;
  assign new_n7912_ = ~pi456;
  assign new_n7913_ = ~pi457 | ~pi212;
  assign new_n7914_ = ~pi211;
  assign new_n7915_ = ~pi210;
  assign new_n7916_ = ~pi455;
  assign new_n7917_ = ~pi209;
  assign new_n7918_ = ~pi454;
  assign new_n7919_ = ~pi208;
  assign new_n7920_ = ~pi453;
  assign new_n7921_ = ~pi207;
  assign new_n7922_ = ~pi452;
  assign new_n7923_ = ~pi206;
  assign new_n7924_ = ~pi451;
  assign new_n7925_ = ~pi205;
  assign new_n7926_ = ~pi450;
  assign new_n7927_ = ~pi204;
  assign new_n7928_ = ~pi449;
  assign new_n7929_ = ~pi448;
  assign new_n7930_ = ~pi203;
  assign new_n7931_ = ~pi202;
  assign new_n7932_ = ~pi447;
  assign new_n7933_ = ~pi201;
  assign new_n7934_ = ~pi446;
  assign new_n7935_ = ~pi200;
  assign new_n7936_ = ~pi445;
  assign new_n7937_ = ~pi199;
  assign new_n7938_ = ~pi444;
  assign new_n7939_ = ~pi198;
  assign new_n7940_ = ~pi443;
  assign new_n7941_ = ~pi197;
  assign new_n7942_ = ~pi442;
  assign new_n7943_ = ~pi196;
  assign new_n7944_ = ~pi441;
  assign new_n7945_ = ~pi195;
  assign new_n7946_ = ~pi440;
  assign new_n7947_ = ~pi194;
  assign new_n7948_ = ~pi439;
  assign new_n7949_ = ~new_n8054_ | ~new_n8053_;
  assign po019 = ~new_n8195_ | ~new_n8194_;
  assign po010 = ~new_n8071_ | ~new_n8070_;
  assign po011 = ~new_n8078_ | ~new_n8077_;
  assign po012 = ~new_n8085_ | ~new_n8084_;
  assign po013 = ~new_n8092_ | ~new_n8091_;
  assign po014 = ~new_n8099_ | ~new_n8098_;
  assign po015 = ~new_n8106_ | ~new_n8105_;
  assign po016 = ~new_n8113_ | ~new_n8112_;
  assign po017 = ~new_n8120_ | ~new_n8119_;
  assign po001 = ~new_n8137_ | ~new_n8136_;
  assign po002 = ~new_n8144_ | ~new_n8143_;
  assign po003 = ~new_n8151_ | ~new_n8150_;
  assign po004 = ~new_n8158_ | ~new_n8157_;
  assign po005 = ~new_n8165_ | ~new_n8164_;
  assign po006 = ~new_n8172_ | ~new_n8171_;
  assign po007 = ~new_n8179_ | ~new_n8178_;
  assign po008 = ~new_n8186_ | ~new_n8185_;
  assign po009 = ~new_n8193_ | ~new_n8192_;
  assign new_n7968_ = ~new_n8018_ | ~new_n8017_;
  assign new_n7969_ = ~new_n8014_ | ~new_n8013_;
  assign new_n7970_ = ~new_n8010_ | ~new_n8009_;
  assign new_n7971_ = ~new_n8006_ | ~new_n8005_;
  assign new_n7972_ = ~new_n8002_ | ~new_n8001_;
  assign new_n7973_ = ~new_n7998_ | ~new_n7997_;
  assign new_n7974_ = ~new_n7994_ | ~new_n7993_;
  assign new_n7975_ = ~new_n7976_ | ~new_n7990_;
  assign new_n7976_ = ~pi211 | ~new_n7988_;
  assign new_n7977_ = ~pi438;
  assign new_n7978_ = ~pi193;
  assign new_n7979_ = ~new_n8050_ | ~new_n8049_;
  assign new_n7980_ = ~new_n8046_ | ~new_n8045_;
  assign new_n7981_ = ~new_n8042_ | ~new_n8041_;
  assign new_n7982_ = ~new_n8038_ | ~new_n8037_;
  assign new_n7983_ = ~new_n8034_ | ~new_n8033_;
  assign new_n7984_ = ~new_n8030_ | ~new_n8029_;
  assign new_n7985_ = ~new_n8026_ | ~new_n8025_;
  assign new_n7986_ = ~new_n8022_ | ~new_n8021_;
  assign new_n7987_ = ~new_n7976_;
  assign new_n7988_ = ~new_n7913_;
  assign new_n7989_ = ~new_n7914_ | ~new_n7913_;
  assign new_n7990_ = ~pi456 | ~new_n7989_;
  assign new_n7991_ = ~new_n7975_;
  assign new_n7992_ = pi210 | pi455;
  assign new_n7993_ = ~new_n7992_ | ~new_n7975_;
  assign new_n7994_ = ~pi455 | ~pi210;
  assign new_n7995_ = ~new_n7974_;
  assign new_n7996_ = pi209 | pi454;
  assign new_n7997_ = ~new_n7996_ | ~new_n7974_;
  assign new_n7998_ = ~pi454 | ~pi209;
  assign new_n7999_ = ~new_n7973_;
  assign new_n8000_ = pi208 | pi453;
  assign new_n8001_ = ~new_n8000_ | ~new_n7973_;
  assign new_n8002_ = ~pi453 | ~pi208;
  assign new_n8003_ = ~new_n7972_;
  assign new_n8004_ = pi207 | pi452;
  assign new_n8005_ = ~new_n8004_ | ~new_n7972_;
  assign new_n8006_ = ~pi452 | ~pi207;
  assign new_n8007_ = ~new_n7971_;
  assign new_n8008_ = pi206 | pi451;
  assign new_n8009_ = ~new_n8008_ | ~new_n7971_;
  assign new_n8010_ = ~pi451 | ~pi206;
  assign new_n8011_ = ~new_n7970_;
  assign new_n8012_ = pi205 | pi450;
  assign new_n8013_ = ~new_n8012_ | ~new_n7970_;
  assign new_n8014_ = ~pi450 | ~pi205;
  assign new_n8015_ = ~new_n7969_;
  assign new_n8016_ = pi204 | pi449;
  assign new_n8017_ = ~new_n8016_ | ~new_n7969_;
  assign new_n8018_ = ~pi449 | ~pi204;
  assign new_n8019_ = ~new_n7968_;
  assign new_n8020_ = pi203 | pi448;
  assign new_n8021_ = ~new_n8020_ | ~new_n7968_;
  assign new_n8022_ = ~pi203 | ~pi448;
  assign new_n8023_ = ~new_n7986_;
  assign new_n8024_ = pi202 | pi447;
  assign new_n8025_ = ~new_n8024_ | ~new_n7986_;
  assign new_n8026_ = ~pi447 | ~pi202;
  assign new_n8027_ = ~new_n7985_;
  assign new_n8028_ = pi201 | pi446;
  assign new_n8029_ = ~new_n8028_ | ~new_n7985_;
  assign new_n8030_ = ~pi446 | ~pi201;
  assign new_n8031_ = ~new_n7984_;
  assign new_n8032_ = pi200 | pi445;
  assign new_n8033_ = ~new_n8032_ | ~new_n7984_;
  assign new_n8034_ = ~pi445 | ~pi200;
  assign new_n8035_ = ~new_n7983_;
  assign new_n8036_ = pi199 | pi444;
  assign new_n8037_ = ~new_n8036_ | ~new_n7983_;
  assign new_n8038_ = ~pi444 | ~pi199;
  assign new_n8039_ = ~new_n7982_;
  assign new_n8040_ = pi198 | pi443;
  assign new_n8041_ = ~new_n8040_ | ~new_n7982_;
  assign new_n8042_ = ~pi443 | ~pi198;
  assign new_n8043_ = ~new_n7981_;
  assign new_n8044_ = pi197 | pi442;
  assign new_n8045_ = ~new_n8044_ | ~new_n7981_;
  assign new_n8046_ = ~pi442 | ~pi197;
  assign new_n8047_ = ~new_n7980_;
  assign new_n8048_ = pi196 | pi441;
  assign new_n8049_ = ~new_n8048_ | ~new_n7980_;
  assign new_n8050_ = ~pi441 | ~pi196;
  assign new_n8051_ = ~new_n7979_;
  assign new_n8052_ = pi195 | pi440;
  assign new_n8053_ = ~new_n8052_ | ~new_n7979_;
  assign new_n8054_ = ~pi440 | ~pi195;
  assign new_n8055_ = ~new_n7949_;
  assign new_n8056_ = pi194 | pi439;
  assign new_n8057_ = ~new_n8056_ | ~new_n7949_;
  assign new_n8058_ = ~pi439 | ~pi194;
  assign new_n8059_ = ~new_n8057_ | ~new_n8058_ | ~new_n8127_ | ~new_n8126_;
  assign new_n8060_ = ~pi439 | ~pi194;
  assign new_n8061_ = ~new_n8055_ | ~new_n8060_;
  assign new_n8062_ = pi439 | pi194;
  assign new_n8063_ = ~new_n8061_ | ~new_n8062_ | ~new_n8130_;
  assign new_n8064_ = ~new_n8123_ | ~new_n7914_;
  assign new_n8065_ = ~pi448 | ~new_n7930_;
  assign new_n8066_ = ~pi203 | ~new_n7929_;
  assign new_n8067_ = ~pi448 | ~new_n7930_;
  assign new_n8068_ = ~pi203 | ~new_n7929_;
  assign new_n8069_ = ~new_n8068_ | ~new_n8067_;
  assign new_n8070_ = ~new_n7968_ | ~new_n8066_ | ~new_n8065_;
  assign new_n8071_ = ~new_n8019_ | ~new_n8069_;
  assign new_n8072_ = ~pi449 | ~new_n7927_;
  assign new_n8073_ = ~pi204 | ~new_n7928_;
  assign new_n8074_ = ~pi449 | ~new_n7927_;
  assign new_n8075_ = ~pi204 | ~new_n7928_;
  assign new_n8076_ = ~new_n8075_ | ~new_n8074_;
  assign new_n8077_ = ~new_n7969_ | ~new_n8073_ | ~new_n8072_;
  assign new_n8078_ = ~new_n8015_ | ~new_n8076_;
  assign new_n8079_ = ~pi450 | ~new_n7925_;
  assign new_n8080_ = ~pi205 | ~new_n7926_;
  assign new_n8081_ = ~pi450 | ~new_n7925_;
  assign new_n8082_ = ~pi205 | ~new_n7926_;
  assign new_n8083_ = ~new_n8082_ | ~new_n8081_;
  assign new_n8084_ = ~new_n7970_ | ~new_n8080_ | ~new_n8079_;
  assign new_n8085_ = ~new_n8011_ | ~new_n8083_;
  assign new_n8086_ = ~pi451 | ~new_n7923_;
  assign new_n8087_ = ~pi206 | ~new_n7924_;
  assign new_n8088_ = ~pi451 | ~new_n7923_;
  assign new_n8089_ = ~pi206 | ~new_n7924_;
  assign new_n8090_ = ~new_n8089_ | ~new_n8088_;
  assign new_n8091_ = ~new_n7971_ | ~new_n8087_ | ~new_n8086_;
  assign new_n8092_ = ~new_n8007_ | ~new_n8090_;
  assign new_n8093_ = ~pi452 | ~new_n7921_;
  assign new_n8094_ = ~pi207 | ~new_n7922_;
  assign new_n8095_ = ~pi452 | ~new_n7921_;
  assign new_n8096_ = ~pi207 | ~new_n7922_;
  assign new_n8097_ = ~new_n8096_ | ~new_n8095_;
  assign new_n8098_ = ~new_n7972_ | ~new_n8094_ | ~new_n8093_;
  assign new_n8099_ = ~new_n8003_ | ~new_n8097_;
  assign new_n8100_ = ~pi453 | ~new_n7919_;
  assign new_n8101_ = ~pi208 | ~new_n7920_;
  assign new_n8102_ = ~pi453 | ~new_n7919_;
  assign new_n8103_ = ~pi208 | ~new_n7920_;
  assign new_n8104_ = ~new_n8103_ | ~new_n8102_;
  assign new_n8105_ = ~new_n7973_ | ~new_n8101_ | ~new_n8100_;
  assign new_n8106_ = ~new_n7999_ | ~new_n8104_;
  assign new_n8107_ = ~pi454 | ~new_n7917_;
  assign new_n8108_ = ~pi209 | ~new_n7918_;
  assign new_n8109_ = ~pi454 | ~new_n7917_;
  assign new_n8110_ = ~pi209 | ~new_n7918_;
  assign new_n8111_ = ~new_n8110_ | ~new_n8109_;
  assign new_n8112_ = ~new_n7974_ | ~new_n8108_ | ~new_n8107_;
  assign new_n8113_ = ~new_n7995_ | ~new_n8111_;
  assign new_n8114_ = ~pi455 | ~new_n7915_;
  assign new_n8115_ = ~pi210 | ~new_n7916_;
  assign new_n8116_ = ~pi455 | ~new_n7915_;
  assign new_n8117_ = ~pi210 | ~new_n7916_;
  assign new_n8118_ = ~new_n8117_ | ~new_n8116_;
  assign new_n8119_ = ~new_n7975_ | ~new_n8115_ | ~new_n8114_;
  assign new_n8120_ = ~new_n7991_ | ~new_n8118_;
  assign new_n8121_ = ~pi456 | ~new_n7913_;
  assign new_n8122_ = ~new_n7988_ | ~new_n7912_;
  assign new_n8123_ = ~new_n8122_ | ~new_n8121_;
  assign new_n8124_ = ~new_n7912_ | ~pi211 | ~new_n7913_;
  assign new_n8125_ = ~new_n7987_ | ~pi456;
  assign new_n8126_ = ~pi438 | ~new_n7978_;
  assign new_n8127_ = ~pi193 | ~new_n7977_;
  assign new_n8128_ = ~pi438 | ~new_n7978_;
  assign new_n8129_ = ~pi193 | ~new_n7977_;
  assign new_n8130_ = ~new_n8129_ | ~new_n8128_;
  assign new_n8131_ = ~pi439 | ~new_n7947_;
  assign new_n8132_ = ~pi194 | ~new_n7948_;
  assign new_n8133_ = ~pi439 | ~new_n7947_;
  assign new_n8134_ = ~pi194 | ~new_n7948_;
  assign new_n8135_ = ~new_n8134_ | ~new_n8133_;
  assign new_n8136_ = ~new_n7949_ | ~new_n8132_ | ~new_n8131_;
  assign new_n8137_ = ~new_n8135_ | ~new_n8055_;
  assign new_n8138_ = ~pi440 | ~new_n7945_;
  assign new_n8139_ = ~pi195 | ~new_n7946_;
  assign new_n8140_ = ~pi440 | ~new_n7945_;
  assign new_n8141_ = ~pi195 | ~new_n7946_;
  assign new_n8142_ = ~new_n8141_ | ~new_n8140_;
  assign new_n8143_ = ~new_n7979_ | ~new_n8139_ | ~new_n8138_;
  assign new_n8144_ = ~new_n8051_ | ~new_n8142_;
  assign new_n8145_ = ~pi441 | ~new_n7943_;
  assign new_n8146_ = ~pi196 | ~new_n7944_;
  assign new_n8147_ = ~pi441 | ~new_n7943_;
  assign new_n8148_ = ~pi196 | ~new_n7944_;
  assign new_n8149_ = ~new_n8148_ | ~new_n8147_;
  assign new_n8150_ = ~new_n7980_ | ~new_n8146_ | ~new_n8145_;
  assign new_n8151_ = ~new_n8047_ | ~new_n8149_;
  assign new_n8152_ = ~pi442 | ~new_n7941_;
  assign new_n8153_ = ~pi197 | ~new_n7942_;
  assign new_n8154_ = ~pi442 | ~new_n7941_;
  assign new_n8155_ = ~pi197 | ~new_n7942_;
  assign new_n8156_ = ~new_n8155_ | ~new_n8154_;
  assign new_n8157_ = ~new_n7981_ | ~new_n8153_ | ~new_n8152_;
  assign new_n8158_ = ~new_n8043_ | ~new_n8156_;
  assign new_n8159_ = ~pi443 | ~new_n7939_;
  assign new_n8160_ = ~pi198 | ~new_n7940_;
  assign new_n8161_ = ~pi443 | ~new_n7939_;
  assign new_n8162_ = ~pi198 | ~new_n7940_;
  assign new_n8163_ = ~new_n8162_ | ~new_n8161_;
  assign new_n8164_ = ~new_n7982_ | ~new_n8160_ | ~new_n8159_;
  assign new_n8165_ = ~new_n8039_ | ~new_n8163_;
  assign new_n8166_ = ~pi444 | ~new_n7937_;
  assign new_n8167_ = ~pi199 | ~new_n7938_;
  assign new_n8168_ = ~pi444 | ~new_n7937_;
  assign new_n8169_ = ~pi199 | ~new_n7938_;
  assign new_n8170_ = ~new_n8169_ | ~new_n8168_;
  assign new_n8171_ = ~new_n7983_ | ~new_n8167_ | ~new_n8166_;
  assign new_n8172_ = ~new_n8035_ | ~new_n8170_;
  assign new_n8173_ = ~pi445 | ~new_n7935_;
  assign new_n8174_ = ~pi200 | ~new_n7936_;
  assign new_n8175_ = ~pi445 | ~new_n7935_;
  assign new_n8176_ = ~pi200 | ~new_n7936_;
  assign new_n8177_ = ~new_n8176_ | ~new_n8175_;
  assign new_n8178_ = ~new_n7984_ | ~new_n8174_ | ~new_n8173_;
  assign new_n8179_ = ~new_n8031_ | ~new_n8177_;
  assign new_n8180_ = ~pi446 | ~new_n7933_;
  assign new_n8181_ = ~pi201 | ~new_n7934_;
  assign new_n8182_ = ~pi446 | ~new_n7933_;
  assign new_n8183_ = ~pi201 | ~new_n7934_;
  assign new_n8184_ = ~new_n8183_ | ~new_n8182_;
  assign new_n8185_ = ~new_n7985_ | ~new_n8181_ | ~new_n8180_;
  assign new_n8186_ = ~new_n8027_ | ~new_n8184_;
  assign new_n8187_ = ~pi447 | ~new_n7931_;
  assign new_n8188_ = ~pi202 | ~new_n7932_;
  assign new_n8189_ = ~pi447 | ~new_n7931_;
  assign new_n8190_ = ~pi202 | ~new_n7932_;
  assign new_n8191_ = ~new_n8190_ | ~new_n8189_;
  assign new_n8192_ = ~new_n7986_ | ~new_n8188_ | ~new_n8187_;
  assign new_n8193_ = ~new_n8023_ | ~new_n8191_;
  assign new_n8194_ = ~pi457 | ~new_n7910_;
  assign new_n8195_ = ~pi212 | ~new_n7911_;
  assign new_n8196_ = new_n8389_ & new_n8387_;
  assign new_n8197_ = new_n8395_ & new_n8393_;
  assign new_n8198_ = new_n8197_ & new_n8397_;
  assign new_n8199_ = new_n8405_ & new_n8401_;
  assign new_n8200_ = new_n8199_ & new_n8408_;
  assign new_n8201_ = new_n8570_ & new_n8569_;
  assign new_n8202_ = ~new_n8516_ | ~new_n8661_ | ~new_n8660_;
  assign new_n8203_ = new_n8316_ & new_n8515_;
  assign new_n8204_ = ~pi024;
  assign new_n8205_ = ~new_n1104_;
  assign new_n8206_ = ~pi025;
  assign new_n8207_ = ~new_n1105_;
  assign new_n8208_ = ~new_n1105_ | ~pi025;
  assign new_n8209_ = ~pi026;
  assign new_n8210_ = ~new_n1106_;
  assign new_n8211_ = ~pi027;
  assign new_n8212_ = ~new_n1107_;
  assign new_n8213_ = ~pi028;
  assign new_n8214_ = ~new_n1108_;
  assign new_n8215_ = ~new_n1108_ | ~pi028;
  assign new_n8216_ = ~pi029;
  assign new_n8217_ = ~new_n1111_;
  assign new_n8218_ = ~pi030;
  assign new_n8219_ = ~new_n1122_;
  assign new_n8220_ = ~new_n1122_ | ~pi030;
  assign new_n8221_ = ~pi031;
  assign new_n8222_ = ~pi032;
  assign new_n8223_ = ~new_n1134_;
  assign new_n8224_ = ~new_n1133_;
  assign new_n8225_ = ~new_n1103_;
  assign new_n8226_ = ~pi023;
  assign new_n8227_ = ~new_n8480_ | ~new_n8390_;
  assign new_n8228_ = ~pi018;
  assign new_n8229_ = ~new_n1128_;
  assign new_n8230_ = ~pi022;
  assign new_n8231_ = ~new_n1132_;
  assign new_n8232_ = ~pi019;
  assign new_n8233_ = ~new_n1129_;
  assign new_n8234_ = ~pi020;
  assign new_n8235_ = ~new_n1130_;
  assign new_n8236_ = ~pi021;
  assign new_n8237_ = ~new_n1131_;
  assign new_n8238_ = ~new_n1131_ | ~pi021;
  assign new_n8239_ = ~pi017;
  assign new_n8240_ = ~new_n1127_;
  assign new_n8241_ = ~pi016;
  assign new_n8242_ = ~new_n1126_;
  assign new_n8243_ = ~pi015;
  assign new_n8244_ = ~new_n1125_;
  assign new_n8245_ = ~pi014;
  assign new_n8246_ = ~new_n1124_;
  assign new_n8247_ = ~pi013;
  assign new_n8248_ = ~new_n1123_;
  assign new_n8249_ = ~pi012;
  assign new_n8250_ = ~new_n1121_;
  assign new_n8251_ = ~pi011;
  assign new_n8252_ = ~new_n1120_;
  assign new_n8253_ = ~pi010;
  assign new_n8254_ = ~new_n1119_;
  assign new_n8255_ = ~pi009;
  assign new_n8256_ = ~new_n1118_;
  assign new_n8257_ = ~pi008;
  assign new_n8258_ = ~new_n1117_;
  assign new_n8259_ = ~pi007;
  assign new_n8260_ = ~new_n1116_;
  assign new_n8261_ = ~pi006;
  assign new_n8262_ = ~new_n1115_;
  assign new_n8263_ = ~pi005;
  assign new_n8264_ = ~new_n1114_;
  assign new_n8265_ = ~pi004;
  assign new_n8266_ = ~new_n1113_;
  assign new_n8267_ = ~pi003;
  assign new_n8268_ = ~new_n1112_;
  assign new_n8269_ = ~pi002;
  assign new_n8270_ = ~new_n1110_;
  assign new_n8271_ = ~new_n1134_ | ~pi032 | ~pi031;
  assign new_n8272_ = ~new_n8492_ | ~new_n8409_;
  assign new_n8273_ = ~new_n8489_ | ~new_n8406_;
  assign new_n8274_ = ~new_n8485_ | ~new_n8398_;
  assign new_n8275_ = ~new_n8733_ | ~new_n8732_;
  assign new_n8276_ = ~new_n8523_ | ~new_n8522_;
  assign new_n8277_ = ~new_n8530_ | ~new_n8529_;
  assign new_n8278_ = ~new_n8537_ | ~new_n8536_;
  assign new_n8279_ = ~new_n8544_ | ~new_n8543_;
  assign new_n8280_ = ~new_n8551_ | ~new_n8550_;
  assign new_n8281_ = ~new_n8558_ | ~new_n8557_;
  assign new_n8282_ = ~new_n8565_ | ~new_n8564_;
  assign new_n8283_ = ~new_n8579_ | ~new_n8578_;
  assign new_n8284_ = ~new_n8586_ | ~new_n8585_;
  assign new_n8285_ = ~new_n8593_ | ~new_n8592_;
  assign new_n8286_ = ~new_n8600_ | ~new_n8599_;
  assign new_n8287_ = ~new_n8607_ | ~new_n8606_;
  assign new_n8288_ = ~new_n8614_ | ~new_n8613_;
  assign new_n8289_ = ~new_n8621_ | ~new_n8620_;
  assign new_n8290_ = ~new_n8628_ | ~new_n8627_;
  assign new_n8291_ = ~new_n8635_ | ~new_n8634_;
  assign new_n8292_ = ~new_n8642_ | ~new_n8641_;
  assign new_n8293_ = ~new_n8649_ | ~new_n8648_;
  assign new_n8294_ = ~new_n8656_ | ~new_n8655_;
  assign new_n8295_ = ~new_n8668_ | ~new_n8667_;
  assign new_n8296_ = ~new_n8675_ | ~new_n8674_;
  assign new_n8297_ = ~new_n8682_ | ~new_n8681_;
  assign new_n8298_ = ~new_n8689_ | ~new_n8688_;
  assign new_n8299_ = ~new_n8696_ | ~new_n8695_;
  assign new_n8300_ = ~new_n8703_ | ~new_n8702_;
  assign new_n8301_ = ~new_n8710_ | ~new_n8709_;
  assign new_n8302_ = ~new_n8717_ | ~new_n8716_;
  assign new_n8303_ = ~new_n8724_ | ~new_n8723_;
  assign new_n8304_ = ~new_n8731_ | ~new_n8730_;
  assign new_n8305_ = new_n8381_ & new_n8385_;
  assign new_n8306_ = new_n8479_ & new_n8386_;
  assign new_n8307_ = new_n8196_ & new_n8391_;
  assign new_n8308_ = new_n8482_ & new_n8392_;
  assign new_n8309_ = new_n8483_ & new_n8396_;
  assign new_n8310_ = new_n8198_ & new_n8399_;
  assign new_n8311_ = new_n8487_ & new_n8400_;
  assign new_n8312_ = new_n8200_ & new_n8411_;
  assign new_n8313_ = new_n8495_ & new_n8412_;
  assign new_n8314_ = new_n8472_ & new_n8201_ & new_n8474_;
  assign new_n8315_ = new_n8475_ & new_n8568_;
  assign new_n8316_ = new_n8333_ & new_n8476_;
  assign new_n8317_ = new_n8518_ & new_n8517_;
  assign new_n8318_ = ~new_n8309_ | ~new_n8501_;
  assign new_n8319_ = new_n8525_ & new_n8524_;
  assign new_n8320_ = ~new_n8499_ | ~new_n8208_;
  assign new_n8321_ = new_n8532_ & new_n8531_;
  assign new_n8322_ = ~new_n8308_ | ~new_n8511_;
  assign new_n8323_ = new_n8539_ & new_n8538_;
  assign new_n8324_ = ~new_n8481_ | ~new_n8509_;
  assign new_n8325_ = new_n8546_ & new_n8545_;
  assign new_n8326_ = ~new_n8507_ | ~new_n8215_;
  assign new_n8327_ = new_n8553_ & new_n8552_;
  assign new_n8328_ = ~new_n8306_ | ~new_n8513_;
  assign new_n8329_ = new_n8560_ & new_n8559_;
  assign new_n8330_ = ~new_n8220_ | ~new_n8382_;
  assign new_n8331_ = ~new_n1109_;
  assign new_n8332_ = ~pi001;
  assign new_n8333_ = new_n8572_ & new_n8571_;
  assign new_n8334_ = new_n8574_ & new_n8573_;
  assign new_n8335_ = ~new_n8472_ | ~new_n8471_;
  assign new_n8336_ = ~new_n8477_ | ~new_n8478_ | ~new_n8271_;
  assign new_n8337_ = new_n8588_ & new_n8587_;
  assign new_n8338_ = ~new_n8468_ | ~new_n8467_;
  assign new_n8339_ = new_n8595_ & new_n8594_;
  assign new_n8340_ = ~new_n8464_ | ~new_n8463_;
  assign new_n8341_ = new_n8602_ & new_n8601_;
  assign new_n8342_ = ~new_n8460_ | ~new_n8459_;
  assign new_n8343_ = new_n8609_ & new_n8608_;
  assign new_n8344_ = ~new_n8456_ | ~new_n8455_;
  assign new_n8345_ = new_n8616_ & new_n8615_;
  assign new_n8346_ = ~new_n8452_ | ~new_n8451_;
  assign new_n8347_ = new_n8623_ & new_n8622_;
  assign new_n8348_ = ~new_n8448_ | ~new_n8447_;
  assign new_n8349_ = new_n8630_ & new_n8629_;
  assign new_n8350_ = ~new_n8444_ | ~new_n8443_;
  assign new_n8351_ = new_n8637_ & new_n8636_;
  assign new_n8352_ = ~new_n8440_ | ~new_n8439_;
  assign new_n8353_ = new_n8644_ & new_n8643_;
  assign new_n8354_ = ~new_n8436_ | ~new_n8435_;
  assign new_n8355_ = new_n8651_ & new_n8650_;
  assign new_n8356_ = ~new_n8432_ | ~new_n8431_;
  assign new_n8357_ = ~new_n1134_ | ~pi032;
  assign new_n8358_ = new_n8663_ & new_n8662_;
  assign new_n8359_ = ~new_n8428_ | ~new_n8427_;
  assign new_n8360_ = new_n8670_ & new_n8669_;
  assign new_n8361_ = ~new_n8424_ | ~new_n8423_;
  assign new_n8362_ = new_n8677_ & new_n8676_;
  assign new_n8363_ = ~new_n8420_ | ~new_n8419_;
  assign new_n8364_ = new_n8684_ & new_n8683_;
  assign new_n8365_ = ~new_n8416_ | ~new_n8415_;
  assign new_n8366_ = new_n8691_ & new_n8690_;
  assign new_n8367_ = ~new_n8313_ | ~new_n8494_;
  assign new_n8368_ = new_n8698_ & new_n8697_;
  assign new_n8369_ = ~new_n8493_ | ~new_n8491_;
  assign new_n8370_ = new_n8705_ & new_n8704_;
  assign new_n8371_ = ~new_n8490_ | ~new_n8488_;
  assign new_n8372_ = new_n8712_ & new_n8711_;
  assign new_n8373_ = ~new_n8238_ | ~new_n8402_;
  assign new_n8374_ = new_n8719_ & new_n8718_;
  assign new_n8375_ = ~new_n8311_ | ~new_n8505_;
  assign new_n8376_ = new_n8726_ & new_n8725_;
  assign new_n8377_ = ~new_n8486_ | ~new_n8503_;
  assign new_n8378_ = ~new_n8271_;
  assign new_n8379_ = ~new_n8357_;
  assign new_n8380_ = ~new_n8336_;
  assign new_n8381_ = pi030 | new_n1122_;
  assign new_n8382_ = ~new_n8496_ | ~new_n8381_;
  assign new_n8383_ = ~new_n8220_;
  assign new_n8384_ = ~new_n8330_;
  assign new_n8385_ = pi029 | new_n1111_;
  assign new_n8386_ = ~new_n1111_ | ~pi029;
  assign new_n8387_ = pi028 | new_n1108_;
  assign new_n8388_ = ~new_n8215_;
  assign new_n8389_ = pi027 | new_n1107_;
  assign new_n8390_ = ~new_n1107_ | ~pi027;
  assign new_n8391_ = pi026 | new_n1106_;
  assign new_n8392_ = ~new_n1106_ | ~pi026;
  assign new_n8393_ = pi025 | new_n1105_;
  assign new_n8394_ = ~new_n8208_;
  assign new_n8395_ = pi024 | new_n1104_;
  assign new_n8396_ = ~new_n1104_ | ~pi024;
  assign new_n8397_ = pi023 | new_n1103_;
  assign new_n8398_ = ~pi023 | ~new_n1103_;
  assign new_n8399_ = pi022 | new_n1132_;
  assign new_n8400_ = ~new_n1132_ | ~pi022;
  assign new_n8401_ = pi021 | new_n1131_;
  assign new_n8402_ = ~new_n8401_ | ~new_n8375_;
  assign new_n8403_ = ~new_n8238_;
  assign new_n8404_ = ~new_n8373_;
  assign new_n8405_ = pi020 | new_n1130_;
  assign new_n8406_ = ~new_n1130_ | ~pi020;
  assign new_n8407_ = ~new_n8371_;
  assign new_n8408_ = pi019 | new_n1129_;
  assign new_n8409_ = ~new_n1129_ | ~pi019;
  assign new_n8410_ = ~new_n8369_;
  assign new_n8411_ = pi018 | new_n1128_;
  assign new_n8412_ = ~new_n1128_ | ~pi018;
  assign new_n8413_ = ~new_n8367_;
  assign new_n8414_ = pi017 | new_n1127_;
  assign new_n8415_ = ~new_n8414_ | ~new_n8367_;
  assign new_n8416_ = ~new_n1127_ | ~pi017;
  assign new_n8417_ = ~new_n8365_;
  assign new_n8418_ = pi016 | new_n1126_;
  assign new_n8419_ = ~new_n8418_ | ~new_n8365_;
  assign new_n8420_ = ~new_n1126_ | ~pi016;
  assign new_n8421_ = ~new_n8363_;
  assign new_n8422_ = pi015 | new_n1125_;
  assign new_n8423_ = ~new_n8422_ | ~new_n8363_;
  assign new_n8424_ = ~new_n1125_ | ~pi015;
  assign new_n8425_ = ~new_n8361_;
  assign new_n8426_ = pi014 | new_n1124_;
  assign new_n8427_ = ~new_n8426_ | ~new_n8361_;
  assign new_n8428_ = ~new_n1124_ | ~pi014;
  assign new_n8429_ = ~new_n8359_;
  assign new_n8430_ = pi013 | new_n1123_;
  assign new_n8431_ = ~new_n8430_ | ~new_n8359_;
  assign new_n8432_ = ~new_n1123_ | ~pi013;
  assign new_n8433_ = ~new_n8356_;
  assign new_n8434_ = pi012 | new_n1121_;
  assign new_n8435_ = ~new_n8434_ | ~new_n8356_;
  assign new_n8436_ = ~new_n1121_ | ~pi012;
  assign new_n8437_ = ~new_n8354_;
  assign new_n8438_ = pi011 | new_n1120_;
  assign new_n8439_ = ~new_n8438_ | ~new_n8354_;
  assign new_n8440_ = ~new_n1120_ | ~pi011;
  assign new_n8441_ = ~new_n8352_;
  assign new_n8442_ = pi010 | new_n1119_;
  assign new_n8443_ = ~new_n8442_ | ~new_n8352_;
  assign new_n8444_ = ~new_n1119_ | ~pi010;
  assign new_n8445_ = ~new_n8350_;
  assign new_n8446_ = pi009 | new_n1118_;
  assign new_n8447_ = ~new_n8446_ | ~new_n8350_;
  assign new_n8448_ = ~new_n1118_ | ~pi009;
  assign new_n8449_ = ~new_n8348_;
  assign new_n8450_ = pi008 | new_n1117_;
  assign new_n8451_ = ~new_n8450_ | ~new_n8348_;
  assign new_n8452_ = ~new_n1117_ | ~pi008;
  assign new_n8453_ = ~new_n8346_;
  assign new_n8454_ = pi007 | new_n1116_;
  assign new_n8455_ = ~new_n8454_ | ~new_n8346_;
  assign new_n8456_ = ~new_n1116_ | ~pi007;
  assign new_n8457_ = ~new_n8344_;
  assign new_n8458_ = pi006 | new_n1115_;
  assign new_n8459_ = ~new_n8458_ | ~new_n8344_;
  assign new_n8460_ = ~new_n1115_ | ~pi006;
  assign new_n8461_ = ~new_n8342_;
  assign new_n8462_ = pi005 | new_n1114_;
  assign new_n8463_ = ~new_n8462_ | ~new_n8342_;
  assign new_n8464_ = ~new_n1114_ | ~pi005;
  assign new_n8465_ = ~new_n8340_;
  assign new_n8466_ = pi004 | new_n1113_;
  assign new_n8467_ = ~new_n8466_ | ~new_n8340_;
  assign new_n8468_ = ~new_n1113_ | ~pi004;
  assign new_n8469_ = ~new_n8338_;
  assign new_n8470_ = pi003 | new_n1112_;
  assign new_n8471_ = ~new_n8470_ | ~new_n8338_;
  assign new_n8472_ = ~new_n1112_ | ~pi003;
  assign new_n8473_ = ~new_n8335_;
  assign new_n8474_ = ~new_n1110_ | ~pi002;
  assign new_n8475_ = new_n1110_ | pi002;
  assign new_n8476_ = ~new_n8471_ | ~new_n8314_;
  assign new_n8477_ = ~new_n1133_ | ~new_n1134_ | ~pi032;
  assign new_n8478_ = ~new_n1133_ | ~pi031;
  assign new_n8479_ = ~new_n8383_ | ~new_n8385_;
  assign new_n8480_ = ~new_n8388_ | ~new_n8389_;
  assign new_n8481_ = ~new_n8227_;
  assign new_n8482_ = ~new_n8227_ | ~new_n8391_;
  assign new_n8483_ = ~new_n8394_ | ~new_n8395_;
  assign new_n8484_ = ~new_n8483_ | ~new_n8396_;
  assign new_n8485_ = ~new_n8484_ | ~new_n8397_;
  assign new_n8486_ = ~new_n8274_;
  assign new_n8487_ = ~new_n8274_ | ~new_n8399_;
  assign new_n8488_ = ~new_n8199_ | ~new_n8375_;
  assign new_n8489_ = ~new_n8403_ | ~new_n8405_;
  assign new_n8490_ = ~new_n8273_;
  assign new_n8491_ = ~new_n8200_ | ~new_n8375_;
  assign new_n8492_ = ~new_n8273_ | ~new_n8408_;
  assign new_n8493_ = ~new_n8272_;
  assign new_n8494_ = ~new_n8312_ | ~new_n8375_;
  assign new_n8495_ = ~new_n8272_ | ~new_n8411_;
  assign new_n8496_ = ~new_n8497_ | ~new_n8498_ | ~new_n8478_;
  assign new_n8497_ = ~new_n1133_ | ~new_n1134_ | ~pi032;
  assign new_n8498_ = ~new_n1134_ | ~pi032 | ~pi031;
  assign new_n8499_ = ~new_n8393_ | ~new_n8322_;
  assign new_n8500_ = ~new_n8320_;
  assign new_n8501_ = ~new_n8197_ | ~new_n8322_;
  assign new_n8502_ = ~new_n8318_;
  assign new_n8503_ = ~new_n8198_ | ~new_n8322_;
  assign new_n8504_ = ~new_n8377_;
  assign new_n8505_ = ~new_n8310_ | ~new_n8322_;
  assign new_n8506_ = ~new_n8375_;
  assign new_n8507_ = ~new_n8387_ | ~new_n8328_;
  assign new_n8508_ = ~new_n8326_;
  assign new_n8509_ = ~new_n8196_ | ~new_n8328_;
  assign new_n8510_ = ~new_n8324_;
  assign new_n8511_ = ~new_n8307_ | ~new_n8328_;
  assign new_n8512_ = ~new_n8322_;
  assign new_n8513_ = ~new_n8305_ | ~new_n8336_;
  assign new_n8514_ = ~new_n8328_;
  assign new_n8515_ = ~new_n8315_ | ~new_n8335_;
  assign new_n8516_ = ~new_n8378_ | ~new_n1133_;
  assign new_n8517_ = ~new_n1103_ | ~new_n8226_;
  assign new_n8518_ = ~pi023 | ~new_n8225_;
  assign new_n8519_ = ~new_n1103_ | ~new_n8226_;
  assign new_n8520_ = ~pi023 | ~new_n8225_;
  assign new_n8521_ = ~new_n8520_ | ~new_n8519_;
  assign new_n8522_ = ~new_n8317_ | ~new_n8318_;
  assign new_n8523_ = ~new_n8502_ | ~new_n8521_;
  assign new_n8524_ = ~new_n1104_ | ~new_n8204_;
  assign new_n8525_ = ~pi024 | ~new_n8205_;
  assign new_n8526_ = ~new_n1104_ | ~new_n8204_;
  assign new_n8527_ = ~pi024 | ~new_n8205_;
  assign new_n8528_ = ~new_n8527_ | ~new_n8526_;
  assign new_n8529_ = ~new_n8319_ | ~new_n8320_;
  assign new_n8530_ = ~new_n8500_ | ~new_n8528_;
  assign new_n8531_ = ~new_n1105_ | ~new_n8206_;
  assign new_n8532_ = ~pi025 | ~new_n8207_;
  assign new_n8533_ = ~new_n1105_ | ~new_n8206_;
  assign new_n8534_ = ~pi025 | ~new_n8207_;
  assign new_n8535_ = ~new_n8534_ | ~new_n8533_;
  assign new_n8536_ = ~new_n8321_ | ~new_n8322_;
  assign new_n8537_ = ~new_n8512_ | ~new_n8535_;
  assign new_n8538_ = ~new_n1106_ | ~new_n8209_;
  assign new_n8539_ = ~pi026 | ~new_n8210_;
  assign new_n8540_ = ~new_n1106_ | ~new_n8209_;
  assign new_n8541_ = ~pi026 | ~new_n8210_;
  assign new_n8542_ = ~new_n8541_ | ~new_n8540_;
  assign new_n8543_ = ~new_n8323_ | ~new_n8324_;
  assign new_n8544_ = ~new_n8510_ | ~new_n8542_;
  assign new_n8545_ = ~new_n1107_ | ~new_n8211_;
  assign new_n8546_ = ~pi027 | ~new_n8212_;
  assign new_n8547_ = ~new_n1107_ | ~new_n8211_;
  assign new_n8548_ = ~pi027 | ~new_n8212_;
  assign new_n8549_ = ~new_n8548_ | ~new_n8547_;
  assign new_n8550_ = ~new_n8325_ | ~new_n8326_;
  assign new_n8551_ = ~new_n8508_ | ~new_n8549_;
  assign new_n8552_ = ~new_n1108_ | ~new_n8213_;
  assign new_n8553_ = ~pi028 | ~new_n8214_;
  assign new_n8554_ = ~new_n1108_ | ~new_n8213_;
  assign new_n8555_ = ~pi028 | ~new_n8214_;
  assign new_n8556_ = ~new_n8555_ | ~new_n8554_;
  assign new_n8557_ = ~new_n8327_ | ~new_n8328_;
  assign new_n8558_ = ~new_n8514_ | ~new_n8556_;
  assign new_n8559_ = ~new_n1111_ | ~new_n8216_;
  assign new_n8560_ = ~pi029 | ~new_n8217_;
  assign new_n8561_ = ~new_n1111_ | ~new_n8216_;
  assign new_n8562_ = ~pi029 | ~new_n8217_;
  assign new_n8563_ = ~new_n8562_ | ~new_n8561_;
  assign new_n8564_ = ~new_n8329_ | ~new_n8330_;
  assign new_n8565_ = ~new_n8384_ | ~new_n8563_;
  assign new_n8566_ = ~new_n1109_ | ~new_n8332_;
  assign new_n8567_ = ~pi001 | ~new_n8331_;
  assign new_n8568_ = ~new_n8567_ | ~new_n8566_;
  assign new_n8569_ = ~new_n1109_ | ~new_n8332_;
  assign new_n8570_ = ~pi001 | ~new_n8331_;
  assign new_n8571_ = ~new_n8270_ | ~new_n8201_ | ~new_n8269_;
  assign new_n8572_ = ~new_n1110_ | ~pi002 | ~new_n8568_;
  assign new_n8573_ = ~new_n1110_ | ~new_n8269_;
  assign new_n8574_ = ~pi002 | ~new_n8270_;
  assign new_n8575_ = ~new_n1110_ | ~new_n8269_;
  assign new_n8576_ = ~pi002 | ~new_n8270_;
  assign new_n8577_ = ~new_n8576_ | ~new_n8575_;
  assign new_n8578_ = ~new_n8334_ | ~new_n8335_;
  assign new_n8579_ = ~new_n8473_ | ~new_n8577_;
  assign new_n8580_ = ~new_n1122_ | ~new_n8218_;
  assign new_n8581_ = ~pi030 | ~new_n8219_;
  assign new_n8582_ = ~new_n1122_ | ~new_n8218_;
  assign new_n8583_ = ~pi030 | ~new_n8219_;
  assign new_n8584_ = ~new_n8583_ | ~new_n8582_;
  assign new_n8585_ = ~new_n8336_ | ~new_n8581_ | ~new_n8580_;
  assign new_n8586_ = ~new_n8380_ | ~new_n8584_;
  assign new_n8587_ = ~new_n1112_ | ~new_n8267_;
  assign new_n8588_ = ~pi003 | ~new_n8268_;
  assign new_n8589_ = ~new_n1112_ | ~new_n8267_;
  assign new_n8590_ = ~pi003 | ~new_n8268_;
  assign new_n8591_ = ~new_n8590_ | ~new_n8589_;
  assign new_n8592_ = ~new_n8337_ | ~new_n8338_;
  assign new_n8593_ = ~new_n8469_ | ~new_n8591_;
  assign new_n8594_ = ~new_n1113_ | ~new_n8265_;
  assign new_n8595_ = ~pi004 | ~new_n8266_;
  assign new_n8596_ = ~new_n1113_ | ~new_n8265_;
  assign new_n8597_ = ~pi004 | ~new_n8266_;
  assign new_n8598_ = ~new_n8597_ | ~new_n8596_;
  assign new_n8599_ = ~new_n8339_ | ~new_n8340_;
  assign new_n8600_ = ~new_n8465_ | ~new_n8598_;
  assign new_n8601_ = ~new_n1114_ | ~new_n8263_;
  assign new_n8602_ = ~pi005 | ~new_n8264_;
  assign new_n8603_ = ~new_n1114_ | ~new_n8263_;
  assign new_n8604_ = ~pi005 | ~new_n8264_;
  assign new_n8605_ = ~new_n8604_ | ~new_n8603_;
  assign new_n8606_ = ~new_n8341_ | ~new_n8342_;
  assign new_n8607_ = ~new_n8461_ | ~new_n8605_;
  assign new_n8608_ = ~new_n1115_ | ~new_n8261_;
  assign new_n8609_ = ~pi006 | ~new_n8262_;
  assign new_n8610_ = ~new_n1115_ | ~new_n8261_;
  assign new_n8611_ = ~pi006 | ~new_n8262_;
  assign new_n8612_ = ~new_n8611_ | ~new_n8610_;
  assign new_n8613_ = ~new_n8343_ | ~new_n8344_;
  assign new_n8614_ = ~new_n8457_ | ~new_n8612_;
  assign new_n8615_ = ~new_n1116_ | ~new_n8259_;
  assign new_n8616_ = ~pi007 | ~new_n8260_;
  assign new_n8617_ = ~new_n1116_ | ~new_n8259_;
  assign new_n8618_ = ~pi007 | ~new_n8260_;
  assign new_n8619_ = ~new_n8618_ | ~new_n8617_;
  assign new_n8620_ = ~new_n8345_ | ~new_n8346_;
  assign new_n8621_ = ~new_n8453_ | ~new_n8619_;
  assign new_n8622_ = ~new_n1117_ | ~new_n8257_;
  assign new_n8623_ = ~pi008 | ~new_n8258_;
  assign new_n8624_ = ~new_n1117_ | ~new_n8257_;
  assign new_n8625_ = ~pi008 | ~new_n8258_;
  assign new_n8626_ = ~new_n8625_ | ~new_n8624_;
  assign new_n8627_ = ~new_n8347_ | ~new_n8348_;
  assign new_n8628_ = ~new_n8449_ | ~new_n8626_;
  assign new_n8629_ = ~new_n1118_ | ~new_n8255_;
  assign new_n8630_ = ~pi009 | ~new_n8256_;
  assign new_n8631_ = ~new_n1118_ | ~new_n8255_;
  assign new_n8632_ = ~pi009 | ~new_n8256_;
  assign new_n8633_ = ~new_n8632_ | ~new_n8631_;
  assign new_n8634_ = ~new_n8349_ | ~new_n8350_;
  assign new_n8635_ = ~new_n8445_ | ~new_n8633_;
  assign new_n8636_ = ~new_n1119_ | ~new_n8253_;
  assign new_n8637_ = ~pi010 | ~new_n8254_;
  assign new_n8638_ = ~new_n1119_ | ~new_n8253_;
  assign new_n8639_ = ~pi010 | ~new_n8254_;
  assign new_n8640_ = ~new_n8639_ | ~new_n8638_;
  assign new_n8641_ = ~new_n8351_ | ~new_n8352_;
  assign new_n8642_ = ~new_n8441_ | ~new_n8640_;
  assign new_n8643_ = ~new_n1120_ | ~new_n8251_;
  assign new_n8644_ = ~pi011 | ~new_n8252_;
  assign new_n8645_ = ~new_n1120_ | ~new_n8251_;
  assign new_n8646_ = ~pi011 | ~new_n8252_;
  assign new_n8647_ = ~new_n8646_ | ~new_n8645_;
  assign new_n8648_ = ~new_n8353_ | ~new_n8354_;
  assign new_n8649_ = ~new_n8437_ | ~new_n8647_;
  assign new_n8650_ = ~new_n1121_ | ~new_n8249_;
  assign new_n8651_ = ~pi012 | ~new_n8250_;
  assign new_n8652_ = ~new_n1121_ | ~new_n8249_;
  assign new_n8653_ = ~pi012 | ~new_n8250_;
  assign new_n8654_ = ~new_n8653_ | ~new_n8652_;
  assign new_n8655_ = ~new_n8355_ | ~new_n8356_;
  assign new_n8656_ = ~new_n8433_ | ~new_n8654_;
  assign new_n8657_ = ~new_n1133_ | ~new_n8357_;
  assign new_n8658_ = ~new_n8379_ | ~new_n8224_;
  assign new_n8659_ = ~new_n8658_ | ~new_n8657_;
  assign new_n8660_ = ~pi031 | ~new_n8357_ | ~new_n8224_;
  assign new_n8661_ = ~new_n8659_ | ~new_n8221_;
  assign new_n8662_ = ~new_n1123_ | ~new_n8247_;
  assign new_n8663_ = ~pi013 | ~new_n8248_;
  assign new_n8664_ = ~new_n1123_ | ~new_n8247_;
  assign new_n8665_ = ~pi013 | ~new_n8248_;
  assign new_n8666_ = ~new_n8665_ | ~new_n8664_;
  assign new_n8667_ = ~new_n8358_ | ~new_n8359_;
  assign new_n8668_ = ~new_n8429_ | ~new_n8666_;
  assign new_n8669_ = ~new_n1124_ | ~new_n8245_;
  assign new_n8670_ = ~pi014 | ~new_n8246_;
  assign new_n8671_ = ~new_n1124_ | ~new_n8245_;
  assign new_n8672_ = ~pi014 | ~new_n8246_;
  assign new_n8673_ = ~new_n8672_ | ~new_n8671_;
  assign new_n8674_ = ~new_n8360_ | ~new_n8361_;
  assign new_n8675_ = ~new_n8425_ | ~new_n8673_;
  assign new_n8676_ = ~new_n1125_ | ~new_n8243_;
  assign new_n8677_ = ~pi015 | ~new_n8244_;
  assign new_n8678_ = ~new_n1125_ | ~new_n8243_;
  assign new_n8679_ = ~pi015 | ~new_n8244_;
  assign new_n8680_ = ~new_n8679_ | ~new_n8678_;
  assign new_n8681_ = ~new_n8362_ | ~new_n8363_;
  assign new_n8682_ = ~new_n8421_ | ~new_n8680_;
  assign new_n8683_ = ~new_n1126_ | ~new_n8241_;
  assign new_n8684_ = ~pi016 | ~new_n8242_;
  assign new_n8685_ = ~new_n1126_ | ~new_n8241_;
  assign new_n8686_ = ~pi016 | ~new_n8242_;
  assign new_n8687_ = ~new_n8686_ | ~new_n8685_;
  assign new_n8688_ = ~new_n8364_ | ~new_n8365_;
  assign new_n8689_ = ~new_n8417_ | ~new_n8687_;
  assign new_n8690_ = ~new_n1127_ | ~new_n8239_;
  assign new_n8691_ = ~pi017 | ~new_n8240_;
  assign new_n8692_ = ~new_n1127_ | ~new_n8239_;
  assign new_n8693_ = ~pi017 | ~new_n8240_;
  assign new_n8694_ = ~new_n8693_ | ~new_n8692_;
  assign new_n8695_ = ~new_n8366_ | ~new_n8367_;
  assign new_n8696_ = ~new_n8413_ | ~new_n8694_;
  assign new_n8697_ = ~new_n1128_ | ~new_n8228_;
  assign new_n8698_ = ~pi018 | ~new_n8229_;
  assign new_n8699_ = ~new_n1128_ | ~new_n8228_;
  assign new_n8700_ = ~pi018 | ~new_n8229_;
  assign new_n8701_ = ~new_n8700_ | ~new_n8699_;
  assign new_n8702_ = ~new_n8368_ | ~new_n8369_;
  assign new_n8703_ = ~new_n8410_ | ~new_n8701_;
  assign new_n8704_ = ~new_n1129_ | ~new_n8232_;
  assign new_n8705_ = ~pi019 | ~new_n8233_;
  assign new_n8706_ = ~new_n1129_ | ~new_n8232_;
  assign new_n8707_ = ~pi019 | ~new_n8233_;
  assign new_n8708_ = ~new_n8707_ | ~new_n8706_;
  assign new_n8709_ = ~new_n8370_ | ~new_n8371_;
  assign new_n8710_ = ~new_n8407_ | ~new_n8708_;
  assign new_n8711_ = ~new_n1130_ | ~new_n8234_;
  assign new_n8712_ = ~pi020 | ~new_n8235_;
  assign new_n8713_ = ~new_n1130_ | ~new_n8234_;
  assign new_n8714_ = ~pi020 | ~new_n8235_;
  assign new_n8715_ = ~new_n8714_ | ~new_n8713_;
  assign new_n8716_ = ~new_n8372_ | ~new_n8373_;
  assign new_n8717_ = ~new_n8404_ | ~new_n8715_;
  assign new_n8718_ = ~new_n1131_ | ~new_n8236_;
  assign new_n8719_ = ~pi021 | ~new_n8237_;
  assign new_n8720_ = ~new_n1131_ | ~new_n8236_;
  assign new_n8721_ = ~pi021 | ~new_n8237_;
  assign new_n8722_ = ~new_n8721_ | ~new_n8720_;
  assign new_n8723_ = ~new_n8374_ | ~new_n8375_;
  assign new_n8724_ = ~new_n8506_ | ~new_n8722_;
  assign new_n8725_ = ~new_n1132_ | ~new_n8230_;
  assign new_n8726_ = ~pi022 | ~new_n8231_;
  assign new_n8727_ = ~new_n1132_ | ~new_n8230_;
  assign new_n8728_ = ~pi022 | ~new_n8231_;
  assign new_n8729_ = ~new_n8728_ | ~new_n8727_;
  assign new_n8730_ = ~new_n8376_ | ~new_n8377_;
  assign new_n8731_ = ~new_n8504_ | ~new_n8729_;
  assign new_n8732_ = ~new_n1134_ | ~new_n8222_;
  assign new_n8733_ = ~pi032 | ~new_n8223_;
  assign new_n8734_ = ~pi438;
  assign new_n8735_ = ~pi269;
  assign new_n8736_ = new_n8833_ & pi267 & pi273;
  assign new_n8737_ = ~pi257;
  assign new_n8738_ = ~pi257 | ~pi269;
  assign new_n8739_ = ~pi260;
  assign new_n8740_ = ~pi260 | ~new_n8811_;
  assign new_n8741_ = ~pi248;
  assign new_n8742_ = ~pi248 | ~new_n8812_;
  assign new_n8743_ = ~pi274;
  assign new_n8744_ = ~pi274 | ~new_n8813_;
  assign new_n8745_ = ~pi266;
  assign new_n8746_ = ~pi256;
  assign new_n8747_ = ~pi266 | ~new_n8814_;
  assign new_n8748_ = ~new_n8815_ | ~pi256;
  assign new_n8749_ = ~pi270;
  assign new_n8750_ = ~pi270 | ~new_n8816_;
  assign new_n8751_ = ~pi251;
  assign new_n8752_ = ~pi251 | ~new_n8817_;
  assign new_n8753_ = ~pi263;
  assign new_n8754_ = ~pi263 | ~new_n8818_;
  assign new_n8755_ = ~pi253;
  assign new_n8756_ = ~pi253 | ~new_n8819_;
  assign new_n8757_ = ~pi272;
  assign new_n8758_ = ~pi272 | ~new_n8820_;
  assign new_n8759_ = ~pi246;
  assign new_n8760_ = ~pi246 | ~new_n8821_;
  assign new_n8761_ = ~pi261;
  assign new_n8762_ = ~pi261 | ~new_n8822_;
  assign new_n8763_ = ~pi259;
  assign new_n8764_ = ~pi259 | ~new_n8823_;
  assign new_n8765_ = ~pi249;
  assign new_n8766_ = ~pi249 | ~new_n8824_;
  assign new_n8767_ = ~pi268;
  assign new_n8768_ = ~pi268 | ~new_n8825_;
  assign new_n8769_ = ~pi254;
  assign new_n8770_ = ~pi254 | ~new_n8826_;
  assign new_n8771_ = ~pi264;
  assign new_n8772_ = ~pi264 | ~new_n8827_;
  assign new_n8773_ = ~pi252;
  assign new_n8774_ = ~pi252 | ~new_n8828_;
  assign new_n8775_ = ~pi271;
  assign new_n8776_ = ~pi271 | ~new_n8829_;
  assign new_n8777_ = ~pi258;
  assign new_n8778_ = ~pi258 | ~new_n8830_;
  assign new_n8779_ = ~pi262;
  assign new_n8780_ = ~pi262 | ~new_n8831_;
  assign new_n8781_ = ~pi247;
  assign new_n8782_ = ~pi247 | ~new_n8832_;
  assign new_n8783_ = ~pi267;
  assign new_n8784_ = ~pi273;
  assign new_n8785_ = ~new_n8836_ | ~new_n8835_;
  assign new_n8786_ = ~new_n8838_ | ~new_n8837_;
  assign new_n8787_ = ~new_n8840_ | ~new_n8839_;
  assign new_n8788_ = ~new_n8842_ | ~new_n8841_;
  assign new_n8789_ = ~new_n8844_ | ~new_n8843_;
  assign new_n8790_ = ~new_n8846_ | ~new_n8845_;
  assign new_n8791_ = ~new_n8848_ | ~new_n8847_;
  assign new_n8792_ = ~new_n8850_ | ~new_n8849_;
  assign new_n8793_ = ~new_n8852_ | ~new_n8851_;
  assign new_n8794_ = ~new_n8854_ | ~new_n8853_;
  assign new_n8795_ = ~new_n8856_ | ~new_n8855_;
  assign new_n8796_ = ~new_n8858_ | ~new_n8857_;
  assign new_n8797_ = ~new_n8860_ | ~new_n8859_;
  assign new_n8798_ = ~new_n8862_ | ~new_n8861_;
  assign new_n8799_ = ~new_n8864_ | ~new_n8863_;
  assign new_n8800_ = ~new_n8866_ | ~new_n8865_;
  assign new_n8801_ = ~new_n8868_ | ~new_n8867_;
  assign new_n8802_ = ~new_n8870_ | ~new_n8869_;
  assign new_n8803_ = ~new_n8872_ | ~new_n8871_;
  assign new_n8804_ = ~new_n8874_ | ~new_n8873_;
  assign new_n8805_ = ~new_n8876_ | ~new_n8875_;
  assign new_n8806_ = ~new_n8878_ | ~new_n8877_;
  assign new_n8807_ = ~new_n8880_ | ~new_n8879_;
  assign new_n8808_ = ~new_n8882_ | ~new_n8881_;
  assign new_n8809_ = ~new_n8884_ | ~new_n8883_;
  assign new_n8810_ = ~pi273 | ~new_n8833_;
  assign new_n8811_ = ~new_n8738_;
  assign new_n8812_ = ~new_n8740_;
  assign new_n8813_ = ~new_n8742_;
  assign new_n8814_ = ~new_n8744_;
  assign new_n8815_ = ~new_n8747_;
  assign new_n8816_ = ~new_n8748_;
  assign new_n8817_ = ~new_n8750_;
  assign new_n8818_ = ~new_n8752_;
  assign new_n8819_ = ~new_n8754_;
  assign new_n8820_ = ~new_n8756_;
  assign new_n8821_ = ~new_n8758_;
  assign new_n8822_ = ~new_n8760_;
  assign new_n8823_ = ~new_n8762_;
  assign new_n8824_ = ~new_n8764_;
  assign new_n8825_ = ~new_n8766_;
  assign new_n8826_ = ~new_n8768_;
  assign new_n8827_ = ~new_n8770_;
  assign new_n8828_ = ~new_n8772_;
  assign new_n8829_ = ~new_n8774_;
  assign new_n8830_ = ~new_n8776_;
  assign new_n8831_ = ~new_n8778_;
  assign new_n8832_ = ~new_n8780_;
  assign new_n8833_ = ~new_n8782_;
  assign new_n8834_ = ~new_n8810_;
  assign new_n8835_ = ~pi256 | ~new_n8747_;
  assign new_n8836_ = ~new_n8815_ | ~new_n8746_;
  assign new_n8837_ = ~pi266 | ~new_n8744_;
  assign new_n8838_ = ~new_n8814_ | ~new_n8745_;
  assign new_n8839_ = ~pi274 | ~new_n8742_;
  assign new_n8840_ = ~new_n8813_ | ~new_n8743_;
  assign new_n8841_ = ~pi248 | ~new_n8740_;
  assign new_n8842_ = ~new_n8812_ | ~new_n8741_;
  assign new_n8843_ = ~pi260 | ~new_n8738_;
  assign new_n8844_ = ~new_n8811_ | ~new_n8739_;
  assign new_n8845_ = ~pi257 | ~new_n8735_;
  assign new_n8846_ = ~pi269 | ~new_n8737_;
  assign new_n8847_ = ~pi267 | ~new_n8810_;
  assign new_n8848_ = ~new_n8834_ | ~new_n8783_;
  assign new_n8849_ = ~pi273 | ~new_n8782_;
  assign new_n8850_ = ~new_n8833_ | ~new_n8784_;
  assign new_n8851_ = ~pi247 | ~new_n8780_;
  assign new_n8852_ = ~new_n8832_ | ~new_n8781_;
  assign new_n8853_ = ~pi262 | ~new_n8778_;
  assign new_n8854_ = ~new_n8831_ | ~new_n8779_;
  assign new_n8855_ = ~pi258 | ~new_n8776_;
  assign new_n8856_ = ~new_n8830_ | ~new_n8777_;
  assign new_n8857_ = ~pi271 | ~new_n8774_;
  assign new_n8858_ = ~new_n8829_ | ~new_n8775_;
  assign new_n8859_ = ~pi252 | ~new_n8772_;
  assign new_n8860_ = ~new_n8828_ | ~new_n8773_;
  assign new_n8861_ = ~pi264 | ~new_n8770_;
  assign new_n8862_ = ~new_n8827_ | ~new_n8771_;
  assign new_n8863_ = ~pi254 | ~new_n8768_;
  assign new_n8864_ = ~new_n8826_ | ~new_n8769_;
  assign new_n8865_ = ~pi268 | ~new_n8766_;
  assign new_n8866_ = ~new_n8825_ | ~new_n8767_;
  assign new_n8867_ = ~pi249 | ~new_n8764_;
  assign new_n8868_ = ~new_n8824_ | ~new_n8765_;
  assign new_n8869_ = ~pi259 | ~new_n8762_;
  assign new_n8870_ = ~new_n8823_ | ~new_n8763_;
  assign new_n8871_ = ~pi261 | ~new_n8760_;
  assign new_n8872_ = ~new_n8822_ | ~new_n8761_;
  assign new_n8873_ = ~pi246 | ~new_n8758_;
  assign new_n8874_ = ~new_n8821_ | ~new_n8759_;
  assign new_n8875_ = ~pi272 | ~new_n8756_;
  assign new_n8876_ = ~new_n8820_ | ~new_n8757_;
  assign new_n8877_ = ~pi253 | ~new_n8754_;
  assign new_n8878_ = ~new_n8819_ | ~new_n8755_;
  assign new_n8879_ = ~pi263 | ~new_n8752_;
  assign new_n8880_ = ~new_n8818_ | ~new_n8753_;
  assign new_n8881_ = ~pi251 | ~new_n8750_;
  assign new_n8882_ = ~new_n8817_ | ~new_n8751_;
  assign new_n8883_ = ~pi270 | ~new_n8748_;
  assign new_n8884_ = ~new_n8816_ | ~new_n8749_;
  assign new_n8885_ = new_n8976_ & new_n8975_;
  assign new_n8886_ = new_n8977_ & new_n8978_;
  assign new_n8887_ = new_n8994_ & new_n8993_;
  assign new_n8888_ = new_n9036_ & new_n9035_;
  assign new_n8889_ = new_n9045_ & new_n9044_;
  assign new_n8890_ = new_n9063_ & new_n9062_;
  assign new_n8891_ = new_n9099_ & new_n9096_;
  assign new_n8892_ = new_n9092_ & new_n9089_;
  assign new_n8893_ = new_n9083_ & new_n9080_;
  assign new_n8894_ = new_n9077_ & new_n9073_;
  assign new_n8895_ = new_n9032_ & new_n9029_;
  assign new_n8896_ = new_n9024_ & new_n9021_;
  assign new_n8897_ = new_n9010_ & new_n9007_;
  assign new_n8898_ = ~pi167;
  assign new_n8899_ = ~new_n1809_;
  assign new_n8900_ = ~new_n1812_;
  assign new_n8901_ = ~new_n1809_ | ~pi167;
  assign new_n8902_ = ~pi168;
  assign new_n8903_ = ~pi165;
  assign new_n8904_ = ~new_n1803_;
  assign new_n8905_ = ~new_n1806_;
  assign new_n8906_ = ~pi163;
  assign new_n8907_ = ~new_n1797_;
  assign new_n8908_ = ~pi161;
  assign new_n8909_ = ~new_n1788_;
  assign new_n8910_ = ~new_n1788_ | ~pi161;
  assign new_n8911_ = ~pi164;
  assign new_n8912_ = ~new_n1800_;
  assign new_n8913_ = ~new_n1803_ | ~pi165;
  assign new_n8914_ = ~pi166;
  assign new_n8915_ = ~pi169;
  assign new_n8916_ = ~new_n1815_;
  assign new_n8917_ = ~new_n1818_;
  assign new_n8918_ = ~pi170;
  assign new_n8919_ = ~new_n8930_ | ~new_n9002_;
  assign new_n8920_ = ~new_n8990_ | ~new_n8991_ | ~new_n8989_;
  assign new_n8921_ = ~new_n8979_ | ~new_n8980_;
  assign new_n8922_ = ~pi162 | ~new_n1794_;
  assign new_n8923_ = ~new_n9016_ | ~new_n9017_ | ~new_n9015_;
  assign new_n8924_ = ~new_n9013_ | ~new_n9012_;
  assign new_n8925_ = ~pi177;
  assign new_n8926_ = ~new_n1839_;
  assign new_n8927_ = ~new_n1842_;
  assign new_n8928_ = ~new_n1839_ | ~pi177;
  assign new_n8929_ = ~pi178;
  assign new_n8930_ = ~new_n1815_ | ~pi169;
  assign new_n8931_ = ~pi171;
  assign new_n8932_ = ~new_n1821_;
  assign new_n8933_ = ~pi173;
  assign new_n8934_ = ~new_n1827_;
  assign new_n8935_ = ~pi172;
  assign new_n8936_ = ~new_n1824_;
  assign new_n8937_ = ~new_n1824_ | ~pi172;
  assign new_n8938_ = ~pi174;
  assign new_n8939_ = ~new_n1830_;
  assign new_n8940_ = ~pi175;
  assign new_n8941_ = ~new_n1833_;
  assign new_n8942_ = ~pi176;
  assign new_n8943_ = ~new_n1836_;
  assign new_n8944_ = ~pi179;
  assign new_n8945_ = ~new_n1845_;
  assign new_n8946_ = ~new_n9068_ | ~new_n9067_ | ~new_n9066_;
  assign new_n8947_ = ~new_n9060_ | ~new_n9059_;
  assign new_n8948_ = ~new_n8937_ | ~new_n9085_;
  assign new_n8949_ = ~new_n9140_ | ~new_n9139_;
  assign new_n8950_ = ~new_n9189_ | ~new_n9188_;
  assign new_n8951_ = ~new_n9112_ | ~new_n9111_;
  assign new_n8952_ = ~new_n9117_ | ~new_n9116_;
  assign new_n8953_ = ~new_n9124_ | ~new_n9123_;
  assign new_n8954_ = ~new_n9131_ | ~new_n9130_;
  assign new_n8955_ = ~new_n9136_ | ~new_n9135_;
  assign new_n8956_ = ~new_n9152_ | ~new_n9151_;
  assign new_n8957_ = ~new_n9159_ | ~new_n9158_;
  assign new_n8958_ = ~new_n9166_ | ~new_n9165_;
  assign new_n8959_ = ~new_n9173_ | ~new_n9172_;
  assign new_n8960_ = ~new_n9180_ | ~new_n9179_;
  assign new_n8961_ = ~new_n9185_ | ~new_n9184_;
  assign new_n8962_ = ~new_n8999_ | ~new_n8998_ | ~new_n8997_;
  assign new_n8963_ = ~new_n9014_ | ~new_n9026_;
  assign new_n8964_ = ~new_n8922_ | ~new_n9033_;
  assign new_n8965_ = ~new_n1782_;
  assign new_n8966_ = ~pi180;
  assign new_n8967_ = ~new_n9056_ | ~new_n9055_;
  assign new_n8968_ = ~new_n9052_ | ~new_n9051_;
  assign new_n8969_ = ~new_n9042_ | ~new_n9041_;
  assign new_n8970_ = ~new_n8913_;
  assign new_n8971_ = ~pi170 | ~new_n1818_;
  assign new_n8972_ = ~new_n1827_ | ~pi173;
  assign new_n8973_ = ~new_n8937_;
  assign new_n8974_ = ~new_n8930_;
  assign new_n8975_ = new_n1806_ | pi166;
  assign new_n8976_ = new_n1803_ | pi165;
  assign new_n8977_ = pi164 | new_n1800_;
  assign new_n8978_ = pi163 | new_n1797_;
  assign new_n8979_ = ~new_n8910_;
  assign new_n8980_ = pi162 | new_n1794_;
  assign new_n8981_ = ~new_n8921_;
  assign new_n8982_ = ~new_n8922_;
  assign new_n8983_ = ~new_n8921_ | ~new_n8922_;
  assign new_n8984_ = ~new_n8977_ | ~pi163 | ~new_n1797_;
  assign new_n8985_ = ~new_n8886_ | ~new_n8983_;
  assign new_n8986_ = ~new_n1800_ | ~pi164;
  assign new_n8987_ = ~new_n8985_ | ~new_n8986_ | ~new_n8984_;
  assign new_n8988_ = ~new_n8914_ | ~new_n8913_;
  assign new_n8989_ = ~new_n1806_ | ~new_n8988_;
  assign new_n8990_ = ~new_n8885_ | ~new_n8987_;
  assign new_n8991_ = ~pi166 | ~new_n8970_;
  assign new_n8992_ = ~new_n8920_;
  assign new_n8993_ = new_n1812_ | pi168;
  assign new_n8994_ = new_n1809_ | pi167;
  assign new_n8995_ = ~new_n8901_;
  assign new_n8996_ = ~new_n8902_ | ~new_n8901_;
  assign new_n8997_ = ~new_n1812_ | ~new_n8996_;
  assign new_n8998_ = ~pi168 | ~new_n8995_;
  assign new_n8999_ = ~new_n8887_ | ~new_n8920_;
  assign new_n9000_ = ~new_n8962_;
  assign new_n9001_ = pi169 | new_n1815_;
  assign new_n9002_ = ~new_n9001_ | ~new_n8962_;
  assign new_n9003_ = ~new_n8919_;
  assign new_n9004_ = new_n1818_ | pi170;
  assign new_n9005_ = pi167 | new_n1809_;
  assign new_n9006_ = ~new_n9005_ | ~new_n8920_;
  assign new_n9007_ = ~new_n9006_ | ~new_n8901_ | ~new_n9119_ | ~new_n9118_;
  assign new_n9008_ = ~new_n8992_ | ~new_n8901_;
  assign new_n9009_ = ~pi168 | ~new_n1812_;
  assign new_n9010_ = ~new_n9008_ | ~new_n9009_ | ~new_n8887_;
  assign new_n9011_ = new_n1809_ | pi167;
  assign new_n9012_ = ~new_n8982_ | ~new_n8978_;
  assign new_n9013_ = ~new_n1797_ | ~pi163;
  assign new_n9014_ = ~new_n8924_;
  assign new_n9015_ = ~new_n8981_ | ~new_n8886_;
  assign new_n9016_ = ~new_n8924_ | ~new_n8977_;
  assign new_n9017_ = ~new_n1800_ | ~pi164;
  assign new_n9018_ = ~new_n8923_;
  assign new_n9019_ = pi165 | new_n1803_;
  assign new_n9020_ = ~new_n9019_ | ~new_n8923_;
  assign new_n9021_ = ~new_n9020_ | ~new_n8913_ | ~new_n9126_ | ~new_n9125_;
  assign new_n9022_ = ~new_n9018_ | ~new_n8913_;
  assign new_n9023_ = ~pi166 | ~new_n1806_;
  assign new_n9024_ = ~new_n9022_ | ~new_n9023_ | ~new_n8885_;
  assign new_n9025_ = new_n1803_ | pi165;
  assign new_n9026_ = ~new_n8981_ | ~new_n8978_;
  assign new_n9027_ = ~new_n8963_;
  assign new_n9028_ = ~new_n1800_ | ~pi164;
  assign new_n9029_ = ~new_n9137_ | ~new_n9138_ | ~new_n8922_ | ~new_n8921_;
  assign new_n9030_ = ~new_n8922_ | ~new_n8921_;
  assign new_n9031_ = ~new_n1797_ | ~pi163;
  assign new_n9032_ = ~new_n9030_ | ~new_n9031_ | ~new_n8978_;
  assign new_n9033_ = pi162 | new_n1794_;
  assign new_n9034_ = ~new_n8964_;
  assign new_n9035_ = new_n1818_ | pi170;
  assign new_n9036_ = new_n1821_ | pi171;
  assign new_n9037_ = ~new_n8974_ | ~new_n8888_;
  assign new_n9038_ = ~new_n1821_ | ~pi171;
  assign new_n9039_ = ~new_n9037_ | ~new_n9038_ | ~new_n8971_;
  assign new_n9040_ = pi171 | new_n1821_;
  assign new_n9041_ = ~new_n8962_ | ~new_n9001_ | ~new_n8888_;
  assign new_n9042_ = ~new_n9040_ | ~new_n9039_;
  assign new_n9043_ = ~new_n8969_;
  assign new_n9044_ = new_n1830_ | pi174;
  assign new_n9045_ = new_n1827_ | pi173;
  assign new_n9046_ = ~new_n8973_ | ~new_n8889_;
  assign new_n9047_ = ~new_n1830_ | ~pi174;
  assign new_n9048_ = ~new_n9046_ | ~new_n9047_ | ~new_n8972_;
  assign new_n9049_ = pi172 | new_n1824_;
  assign new_n9050_ = pi174 | new_n1830_;
  assign new_n9051_ = ~new_n8969_ | ~new_n9049_ | ~new_n8889_;
  assign new_n9052_ = ~new_n9050_ | ~new_n9048_;
  assign new_n9053_ = ~new_n8968_;
  assign new_n9054_ = pi175 | new_n1833_;
  assign new_n9055_ = ~new_n9054_ | ~new_n8968_;
  assign new_n9056_ = ~new_n1833_ | ~pi175;
  assign new_n9057_ = ~new_n8967_;
  assign new_n9058_ = pi176 | new_n1836_;
  assign new_n9059_ = ~new_n9058_ | ~new_n8967_;
  assign new_n9060_ = ~new_n1836_ | ~pi176;
  assign new_n9061_ = ~new_n8947_;
  assign new_n9062_ = new_n1842_ | pi178;
  assign new_n9063_ = new_n1839_ | pi177;
  assign new_n9064_ = ~new_n8928_;
  assign new_n9065_ = ~new_n8929_ | ~new_n8928_;
  assign new_n9066_ = ~new_n1842_ | ~new_n9065_;
  assign new_n9067_ = ~pi178 | ~new_n9064_;
  assign new_n9068_ = ~new_n8890_ | ~new_n8947_;
  assign new_n9069_ = ~new_n8946_;
  assign new_n9070_ = pi179 | new_n1845_;
  assign new_n9071_ = ~new_n9070_ | ~new_n8946_;
  assign new_n9072_ = ~new_n1845_ | ~pi179;
  assign new_n9073_ = ~new_n9071_ | ~new_n9072_ | ~new_n9142_ | ~new_n9141_;
  assign new_n9074_ = ~new_n1845_ | ~pi179;
  assign new_n9075_ = ~new_n9069_ | ~new_n9074_;
  assign new_n9076_ = new_n1845_ | pi179;
  assign new_n9077_ = ~new_n9075_ | ~new_n9076_ | ~new_n9145_;
  assign new_n9078_ = pi177 | new_n1839_;
  assign new_n9079_ = ~new_n9078_ | ~new_n8947_;
  assign new_n9080_ = ~new_n9079_ | ~new_n8928_ | ~new_n9154_ | ~new_n9153_;
  assign new_n9081_ = ~new_n9061_ | ~new_n8928_;
  assign new_n9082_ = ~pi178 | ~new_n1842_;
  assign new_n9083_ = ~new_n9081_ | ~new_n9082_ | ~new_n8890_;
  assign new_n9084_ = new_n1839_ | pi177;
  assign new_n9085_ = ~new_n9049_ | ~new_n8969_;
  assign new_n9086_ = ~new_n8948_;
  assign new_n9087_ = pi173 | new_n1827_;
  assign new_n9088_ = ~new_n9087_ | ~new_n8948_;
  assign new_n9089_ = ~new_n9088_ | ~new_n8972_ | ~new_n9175_ | ~new_n9174_;
  assign new_n9090_ = ~new_n9086_ | ~new_n8972_;
  assign new_n9091_ = ~new_n1830_ | ~pi174;
  assign new_n9092_ = ~new_n9090_ | ~new_n9091_ | ~new_n8889_;
  assign new_n9093_ = new_n1827_ | pi173;
  assign new_n9094_ = pi170 | new_n1818_;
  assign new_n9095_ = ~new_n9094_ | ~new_n8919_;
  assign new_n9096_ = ~new_n9095_ | ~new_n8971_ | ~new_n9187_ | ~new_n9186_;
  assign new_n9097_ = ~new_n9003_ | ~new_n8971_;
  assign new_n9098_ = ~new_n1821_ | ~pi171;
  assign new_n9099_ = ~new_n9097_ | ~new_n9098_ | ~new_n8888_;
  assign new_n9100_ = ~new_n9004_ | ~new_n8971_;
  assign new_n9101_ = ~new_n9001_ | ~new_n8930_;
  assign new_n9102_ = ~new_n9011_ | ~new_n8901_;
  assign new_n9103_ = ~new_n9025_ | ~new_n8913_;
  assign new_n9104_ = ~new_n9028_ | ~new_n8977_;
  assign new_n9105_ = ~new_n9084_ | ~new_n8928_;
  assign new_n9106_ = ~new_n9093_ | ~new_n8972_;
  assign new_n9107_ = ~new_n9049_ | ~new_n8937_;
  assign new_n9108_ = ~new_n1818_ | ~new_n8918_;
  assign new_n9109_ = ~pi170 | ~new_n8917_;
  assign new_n9110_ = ~new_n9109_ | ~new_n9108_;
  assign new_n9111_ = ~new_n9100_ | ~new_n8919_;
  assign new_n9112_ = ~new_n9110_ | ~new_n9003_;
  assign new_n9113_ = ~new_n1815_ | ~new_n8915_;
  assign new_n9114_ = ~pi169 | ~new_n8916_;
  assign new_n9115_ = ~new_n9114_ | ~new_n9113_;
  assign new_n9116_ = ~new_n9101_ | ~new_n8962_;
  assign new_n9117_ = ~new_n9000_ | ~new_n9115_;
  assign new_n9118_ = ~new_n1812_ | ~new_n8902_;
  assign new_n9119_ = ~pi168 | ~new_n8900_;
  assign new_n9120_ = ~new_n1809_ | ~new_n8898_;
  assign new_n9121_ = ~pi167 | ~new_n8899_;
  assign new_n9122_ = ~new_n9121_ | ~new_n9120_;
  assign new_n9123_ = ~new_n9102_ | ~new_n8920_;
  assign new_n9124_ = ~new_n9122_ | ~new_n8992_;
  assign new_n9125_ = ~new_n1806_ | ~new_n8914_;
  assign new_n9126_ = ~pi166 | ~new_n8905_;
  assign new_n9127_ = ~new_n1803_ | ~new_n8903_;
  assign new_n9128_ = ~pi165 | ~new_n8904_;
  assign new_n9129_ = ~new_n9128_ | ~new_n9127_;
  assign new_n9130_ = ~new_n9103_ | ~new_n8923_;
  assign new_n9131_ = ~new_n9129_ | ~new_n9018_;
  assign new_n9132_ = ~new_n1800_ | ~new_n8911_;
  assign new_n9133_ = ~pi164 | ~new_n8912_;
  assign new_n9134_ = ~new_n9133_ | ~new_n9132_;
  assign new_n9135_ = ~new_n9104_ | ~new_n8963_;
  assign new_n9136_ = ~new_n9027_ | ~new_n9134_;
  assign new_n9137_ = ~new_n1797_ | ~new_n8906_;
  assign new_n9138_ = ~pi163 | ~new_n8907_;
  assign new_n9139_ = ~new_n8979_ | ~new_n8964_;
  assign new_n9140_ = ~new_n9034_ | ~new_n8910_;
  assign new_n9141_ = ~new_n1782_ | ~new_n8966_;
  assign new_n9142_ = ~pi180 | ~new_n8965_;
  assign new_n9143_ = ~new_n1782_ | ~new_n8966_;
  assign new_n9144_ = ~pi180 | ~new_n8965_;
  assign new_n9145_ = ~new_n9144_ | ~new_n9143_;
  assign new_n9146_ = ~new_n1845_ | ~new_n8944_;
  assign new_n9147_ = ~pi179 | ~new_n8945_;
  assign new_n9148_ = ~new_n1845_ | ~new_n8944_;
  assign new_n9149_ = ~pi179 | ~new_n8945_;
  assign new_n9150_ = ~new_n9149_ | ~new_n9148_;
  assign new_n9151_ = ~new_n8946_ | ~new_n9147_ | ~new_n9146_;
  assign new_n9152_ = ~new_n9150_ | ~new_n9069_;
  assign new_n9153_ = ~new_n1842_ | ~new_n8929_;
  assign new_n9154_ = ~pi178 | ~new_n8927_;
  assign new_n9155_ = ~new_n1839_ | ~new_n8925_;
  assign new_n9156_ = ~pi177 | ~new_n8926_;
  assign new_n9157_ = ~new_n9156_ | ~new_n9155_;
  assign new_n9158_ = ~new_n9105_ | ~new_n8947_;
  assign new_n9159_ = ~new_n9157_ | ~new_n9061_;
  assign new_n9160_ = ~new_n1836_ | ~new_n8942_;
  assign new_n9161_ = ~pi176 | ~new_n8943_;
  assign new_n9162_ = ~new_n1836_ | ~new_n8942_;
  assign new_n9163_ = ~pi176 | ~new_n8943_;
  assign new_n9164_ = ~new_n9163_ | ~new_n9162_;
  assign new_n9165_ = ~new_n8967_ | ~new_n9161_ | ~new_n9160_;
  assign new_n9166_ = ~new_n9057_ | ~new_n9164_;
  assign new_n9167_ = ~new_n1833_ | ~new_n8940_;
  assign new_n9168_ = ~pi175 | ~new_n8941_;
  assign new_n9169_ = ~new_n1833_ | ~new_n8940_;
  assign new_n9170_ = ~pi175 | ~new_n8941_;
  assign new_n9171_ = ~new_n9170_ | ~new_n9169_;
  assign new_n9172_ = ~new_n8968_ | ~new_n9168_ | ~new_n9167_;
  assign new_n9173_ = ~new_n9053_ | ~new_n9171_;
  assign new_n9174_ = ~new_n1830_ | ~new_n8938_;
  assign new_n9175_ = ~pi174 | ~new_n8939_;
  assign new_n9176_ = ~new_n1827_ | ~new_n8933_;
  assign new_n9177_ = ~pi173 | ~new_n8934_;
  assign new_n9178_ = ~new_n9177_ | ~new_n9176_;
  assign new_n9179_ = ~new_n9106_ | ~new_n8948_;
  assign new_n9180_ = ~new_n9178_ | ~new_n9086_;
  assign new_n9181_ = ~new_n1824_ | ~new_n8935_;
  assign new_n9182_ = ~pi172 | ~new_n8936_;
  assign new_n9183_ = ~new_n9182_ | ~new_n9181_;
  assign new_n9184_ = ~new_n9107_ | ~new_n8969_;
  assign new_n9185_ = ~new_n9043_ | ~new_n9183_;
  assign new_n9186_ = ~new_n1821_ | ~new_n8931_;
  assign new_n9187_ = ~pi171 | ~new_n8932_;
  assign new_n9188_ = ~new_n1788_ | ~new_n8908_;
  assign new_n9189_ = ~pi161 | ~new_n8909_;
  assign new_n9190_ = new_n9411_ & new_n9222_;
  assign new_n9191_ = new_n9409_ & new_n9376_;
  assign new_n9192_ = new_n9408_ & new_n9219_;
  assign new_n9193_ = new_n9407_ & new_n9220_;
  assign new_n9194_ = new_n9405_ & new_n9379_;
  assign new_n9195_ = new_n9404_ & new_n9218_;
  assign new_n9196_ = new_n9403_ & new_n9381_;
  assign new_n9197_ = new_n9401_ & new_n9382_;
  assign new_n9198_ = new_n9400_ & new_n9356_;
  assign new_n9199_ = new_n9399_ & new_n9384_;
  assign new_n9200_ = new_n9397_ & new_n9385_;
  assign new_n9201_ = new_n9396_ & new_n9353_;
  assign new_n9202_ = new_n9395_ & new_n9351_;
  assign new_n9203_ = new_n9393_ & new_n9388_;
  assign new_n9204_ = new_n9392_ & new_n9217_;
  assign new_n9205_ = new_n9391_ & new_n9211_;
  assign new_n9206_ = new_n9374_ & new_n9364_;
  assign new_n9207_ = new_n9373_ & new_n9213_;
  assign new_n9208_ = new_n9372_ & new_n9214_;
  assign new_n9209_ = new_n9370_ & new_n9367_;
  assign new_n9210_ = new_n9369_ & new_n9212_;
  assign new_n9211_ = pi033 | pi035 | pi034;
  assign new_n9212_ = ~new_n9227_ | ~new_n9228_ | ~new_n9414_;
  assign new_n9213_ = ~new_n9229_ | ~new_n9414_;
  assign new_n9214_ = ~new_n9230_ | ~new_n9365_;
  assign new_n9215_ = ~pi040;
  assign new_n9216_ = ~pi036;
  assign new_n9217_ = ~new_n9240_ | ~new_n9235_;
  assign new_n9218_ = ~new_n9311_ | ~new_n9312_ | ~new_n9314_ | ~new_n9313_;
  assign new_n9219_ = ~new_n9340_ | ~new_n9368_;
  assign new_n9220_ = ~new_n9341_ | ~new_n9377_;
  assign new_n9221_ = ~pi048;
  assign new_n9222_ = ~new_n9342_ | ~new_n9368_;
  assign new_n9223_ = ~pi044;
  assign new_n9224_ = ~new_n9431_ | ~new_n9430_;
  assign new_n9225_ = ~new_n9421_ | ~new_n9420_;
  assign new_n9226_ = ~new_n9425_ | ~new_n9424_;
  assign new_n9227_ = ~pi037 & ~pi036 & ~pi039 & ~pi038;
  assign new_n9228_ = ~pi040 & ~pi041;
  assign new_n9229_ = ~pi036 & ~pi037;
  assign new_n9230_ = ~pi038 & ~pi039;
  assign new_n9231_ = ~pi044 & ~pi043 & ~pi046 & ~pi045;
  assign new_n9232_ = ~pi048 & ~pi047 & ~pi050 & ~pi049;
  assign new_n9233_ = ~pi052 & ~pi051 & ~pi033 & ~pi034;
  assign new_n9234_ = ~pi053 & ~pi054 & ~pi055;
  assign new_n9235_ = new_n9231_ & new_n9232_ & new_n9234_ & new_n9233_;
  assign new_n9236_ = ~pi057 & ~pi056 & ~pi059 & ~pi058;
  assign new_n9237_ = ~pi061 & ~pi060 & ~pi035 & ~pi062;
  assign new_n9238_ = ~pi037 & ~pi036 & ~pi039 & ~pi038;
  assign new_n9239_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9240_ = new_n9236_ & new_n9237_ & new_n9239_ & new_n9238_;
  assign new_n9241_ = ~pi044 & ~pi043 & ~pi046 & ~pi045;
  assign new_n9242_ = ~pi048 & ~pi047 & ~pi050 & ~pi049;
  assign new_n9243_ = ~pi052 & ~pi051 & ~pi033 & ~pi034;
  assign new_n9244_ = ~pi053 & ~pi054 & ~pi055;
  assign new_n9245_ = new_n9241_ & new_n9242_ & new_n9244_ & new_n9243_;
  assign new_n9246_ = ~pi057 & ~pi056 & ~pi059 & ~pi058;
  assign new_n9247_ = ~pi060 & ~pi061 & ~pi035;
  assign new_n9248_ = ~pi037 & ~pi036 & ~pi039 & ~pi038;
  assign new_n9249_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9250_ = new_n9246_ & new_n9247_ & new_n9249_ & new_n9248_;
  assign new_n9251_ = ~pi044 & ~pi043 & ~pi046 & ~pi045;
  assign new_n9252_ = ~pi047 & ~pi048 & ~pi049;
  assign new_n9253_ = ~pi051 & ~pi050 & ~pi034 & ~pi052;
  assign new_n9254_ = ~pi033 & ~pi053 & ~pi054;
  assign new_n9255_ = new_n9251_ & new_n9252_ & new_n9254_ & new_n9253_;
  assign new_n9256_ = ~pi056 & ~pi055 & ~pi058 & ~pi057;
  assign new_n9257_ = ~pi059 & ~pi060 & ~pi035;
  assign new_n9258_ = ~pi037 & ~pi036 & ~pi039 & ~pi038;
  assign new_n9259_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9260_ = new_n9256_ & new_n9257_ & new_n9259_ & new_n9258_;
  assign new_n9261_ = ~pi044 & ~pi043 & ~pi046 & ~pi045;
  assign new_n9262_ = ~pi047 & ~pi048 & ~pi049;
  assign new_n9263_ = ~pi051 & ~pi050 & ~pi034 & ~pi052;
  assign new_n9264_ = ~pi033 & ~pi053 & ~pi054;
  assign new_n9265_ = new_n9261_ & new_n9262_ & new_n9264_ & new_n9263_;
  assign new_n9266_ = ~pi056 & ~pi055 & ~pi058 & ~pi057;
  assign new_n9267_ = ~pi059 & ~pi035 & ~pi036;
  assign new_n9268_ = ~pi037 & ~pi038 & ~pi039;
  assign new_n9269_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9270_ = new_n9266_ & new_n9267_ & new_n9269_ & new_n9268_;
  assign new_n9271_ = ~pi044 & ~pi043 & ~pi046 & ~pi045;
  assign new_n9272_ = ~pi047 & ~pi048 & ~pi049;
  assign new_n9273_ = ~pi051 & ~pi050 & ~pi034 & ~pi052;
  assign new_n9274_ = ~pi033 & ~pi053 & ~pi054;
  assign new_n9275_ = new_n9271_ & new_n9272_ & new_n9274_ & new_n9273_;
  assign new_n9276_ = ~pi056 & ~pi055 & ~pi058 & ~pi057;
  assign new_n9277_ = ~pi059 & ~pi035 & ~pi036;
  assign new_n9278_ = ~pi037 & ~pi038 & ~pi039;
  assign new_n9279_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9280_ = new_n9276_ & new_n9277_ & new_n9279_ & new_n9278_;
  assign new_n9281_ = ~pi044 & ~pi043 & ~pi046 & ~pi045;
  assign new_n9282_ = ~pi047 & ~pi048 & ~pi049;
  assign new_n9283_ = ~pi050 & ~pi051 & ~pi052;
  assign new_n9284_ = ~pi034 & ~pi033 & ~pi053;
  assign new_n9285_ = new_n9281_ & new_n9282_ & new_n9284_ & new_n9283_;
  assign new_n9286_ = ~pi055 & ~pi054 & ~pi057 & ~pi056;
  assign new_n9287_ = ~pi058 & ~pi035 & ~pi036;
  assign new_n9288_ = ~pi037 & ~pi038 & ~pi039;
  assign new_n9289_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9290_ = new_n9286_ & new_n9287_ & new_n9289_ & new_n9288_;
  assign new_n9291_ = ~pi044 & ~pi043 & ~pi046 & ~pi045;
  assign new_n9292_ = ~pi047 & ~pi048 & ~pi049;
  assign new_n9293_ = ~pi050 & ~pi051 & ~pi052;
  assign new_n9294_ = ~pi034 & ~pi033 & ~pi053;
  assign new_n9295_ = new_n9291_ & new_n9292_ & new_n9294_ & new_n9293_;
  assign new_n9296_ = ~pi054 & ~pi055 & ~pi056;
  assign new_n9297_ = ~pi057 & ~pi035 & ~pi036;
  assign new_n9298_ = ~pi037 & ~pi038 & ~pi039;
  assign new_n9299_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9300_ = new_n9296_ & new_n9297_ & new_n9299_ & new_n9298_;
  assign new_n9301_ = ~pi043 & ~pi044 & ~pi045;
  assign new_n9302_ = ~pi046 & ~pi047 & ~pi048;
  assign new_n9303_ = ~pi049 & ~pi050 & ~pi051;
  assign new_n9304_ = ~pi052 & ~pi034 & ~pi033;
  assign new_n9305_ = new_n9301_ & new_n9302_ & new_n9304_ & new_n9303_;
  assign new_n9306_ = ~pi053 & ~pi054 & ~pi055;
  assign new_n9307_ = ~pi056 & ~pi035 & ~pi036;
  assign new_n9308_ = ~pi037 & ~pi038 & ~pi039;
  assign new_n9309_ = ~pi040 & ~pi041 & ~pi042;
  assign new_n9310_ = new_n9306_ & new_n9307_ & new_n9309_ & new_n9308_;
  assign new_n9311_ = ~pi047 & ~pi046 & ~pi045 & ~pi044 & ~pi043;
  assign new_n9312_ = ~pi049 & ~pi048 & ~pi033 & ~pi034;
  assign new_n9313_ = ~pi036 & ~pi035 & ~pi038 & ~pi037;
  assign new_n9314_ = ~pi040 & ~pi039 & ~pi042 & ~pi041;
  assign new_n9315_ = ~pi050 & ~pi051;
  assign new_n9316_ = ~pi052 & ~pi053;
  assign new_n9317_ = ~pi054 & ~pi055;
  assign new_n9318_ = new_n9317_ & new_n9316_ & new_n9315_;
  assign new_n9319_ = ~pi043 & ~pi044 & ~pi045;
  assign new_n9320_ = ~pi046 & ~pi047 & ~pi048;
  assign new_n9321_ = new_n9320_ & new_n9319_;
  assign new_n9322_ = ~pi034 & ~pi052 & ~pi051 & ~pi050 & ~pi049;
  assign new_n9323_ = ~pi033 & ~pi053 & ~pi054;
  assign new_n9324_ = ~pi035 & ~pi036 & ~pi037;
  assign new_n9325_ = new_n9324_ & new_n9323_;
  assign new_n9326_ = ~pi042 & ~pi041 & ~pi040 & ~pi039 & ~pi038;
  assign new_n9327_ = ~pi043 & ~pi044 & ~pi045;
  assign new_n9328_ = ~pi046 & ~pi047 & ~pi048;
  assign new_n9329_ = ~pi034 & ~pi052 & ~pi051 & ~pi050 & ~pi049;
  assign new_n9330_ = ~pi037 & ~pi036 & ~pi035 & ~pi053 & ~pi033;
  assign new_n9331_ = ~pi042 & ~pi041 & ~pi040 & ~pi039 & ~pi038;
  assign new_n9332_ = ~pi047 & ~pi046 & ~pi045 & ~pi044 & ~pi043;
  assign new_n9333_ = ~pi052 & ~pi051 & ~pi050 & ~pi049 & ~pi048;
  assign new_n9334_ = ~pi037 & ~pi036 & ~pi035 & ~pi033 & ~pi034;
  assign new_n9335_ = ~pi042 & ~pi041 & ~pi040 & ~pi039 & ~pi038;
  assign new_n9336_ = ~pi047 & ~pi046 & ~pi045 & ~pi044 & ~pi043;
  assign new_n9337_ = ~pi034 & ~pi051 & ~pi050 & ~pi049 & ~pi048;
  assign new_n9338_ = ~pi038 & ~pi037 & ~pi036 & ~pi035 & ~pi033;
  assign new_n9339_ = ~pi040 & ~pi039 & ~pi042 & ~pi041;
  assign new_n9340_ = ~pi044 & ~pi043 & ~pi042 & ~pi045;
  assign new_n9341_ = ~pi046 & ~pi047;
  assign new_n9342_ = ~pi043 & ~pi042;
  assign new_n9343_ = ~pi042;
  assign new_n9344_ = new_n9417_ & new_n9416_;
  assign new_n9345_ = ~pi038;
  assign new_n9346_ = new_n9419_ & new_n9418_;
  assign new_n9347_ = ~pi064;
  assign new_n9348_ = ~pi063;
  assign new_n9349_ = new_n9423_ & new_n9422_;
  assign new_n9350_ = ~pi060;
  assign new_n9351_ = ~new_n9280_ | ~new_n9275_;
  assign new_n9352_ = ~pi058;
  assign new_n9353_ = ~new_n9300_ | ~new_n9295_;
  assign new_n9354_ = new_n9427_ & new_n9426_;
  assign new_n9355_ = ~pi054;
  assign new_n9356_ = ~new_n9330_ | ~new_n9331_ | ~new_n9329_ | ~new_n9328_ | ~new_n9327_;
  assign new_n9357_ = new_n9429_ & new_n9428_;
  assign new_n9358_ = ~pi034;
  assign new_n9359_ = ~pi033;
  assign new_n9360_ = ~pi050;
  assign new_n9361_ = new_n9433_ & new_n9432_;
  assign new_n9362_ = ~pi046;
  assign new_n9363_ = new_n9435_ & new_n9434_;
  assign new_n9364_ = ~new_n9414_ | ~new_n9216_;
  assign new_n9365_ = ~new_n9213_;
  assign new_n9366_ = ~new_n9214_;
  assign new_n9367_ = ~new_n9366_ | ~new_n9215_;
  assign new_n9368_ = ~new_n9212_;
  assign new_n9369_ = ~pi041 | ~new_n9367_;
  assign new_n9370_ = ~pi040 | ~new_n9214_;
  assign new_n9371_ = ~new_n9365_ | ~new_n9345_;
  assign new_n9372_ = ~pi039 | ~new_n9371_;
  assign new_n9373_ = ~pi037 | ~new_n9364_;
  assign new_n9374_ = ~pi036 | ~new_n9211_;
  assign new_n9375_ = ~new_n9222_;
  assign new_n9376_ = ~new_n9375_ | ~new_n9223_;
  assign new_n9377_ = ~new_n9219_;
  assign new_n9378_ = ~new_n9220_;
  assign new_n9379_ = ~new_n9378_ | ~new_n9221_;
  assign new_n9380_ = ~new_n9218_;
  assign new_n9381_ = ~new_n9336_ | ~new_n9337_ | ~new_n9339_ | ~new_n9338_;
  assign new_n9382_ = ~new_n9332_ | ~new_n9333_ | ~new_n9335_ | ~new_n9334_;
  assign new_n9383_ = ~new_n9356_;
  assign new_n9384_ = ~new_n9318_ | ~new_n9380_;
  assign new_n9385_ = ~new_n9310_ | ~new_n9305_;
  assign new_n9386_ = ~new_n9353_;
  assign new_n9387_ = ~new_n9351_;
  assign new_n9388_ = ~new_n9250_ | ~new_n9245_;
  assign new_n9389_ = ~new_n9217_;
  assign new_n9390_ = pi034 | pi033;
  assign new_n9391_ = ~pi035 | ~new_n9390_;
  assign new_n9392_ = ~pi062 | ~new_n9388_;
  assign new_n9393_ = ~pi061 | ~new_n9413_;
  assign new_n9394_ = ~new_n9290_ | ~new_n9285_;
  assign new_n9395_ = ~pi059 | ~new_n9394_;
  assign new_n9396_ = ~pi057 | ~new_n9385_;
  assign new_n9397_ = ~pi056 | ~new_n9384_;
  assign new_n9398_ = ~new_n9321_ | ~new_n9322_ | ~new_n9326_ | ~new_n9325_;
  assign new_n9399_ = ~pi055 | ~new_n9398_;
  assign new_n9400_ = ~pi053 | ~new_n9382_;
  assign new_n9401_ = ~pi052 | ~new_n9381_;
  assign new_n9402_ = ~new_n9380_ | ~new_n9360_;
  assign new_n9403_ = ~pi051 | ~new_n9402_;
  assign new_n9404_ = ~pi049 | ~new_n9379_;
  assign new_n9405_ = ~pi048 | ~new_n9220_;
  assign new_n9406_ = ~new_n9377_ | ~new_n9362_;
  assign new_n9407_ = ~pi047 | ~new_n9406_;
  assign new_n9408_ = ~pi045 | ~new_n9376_;
  assign new_n9409_ = ~pi044 | ~new_n9222_;
  assign new_n9410_ = ~new_n9368_ | ~new_n9343_;
  assign new_n9411_ = ~pi043 | ~new_n9410_;
  assign new_n9412_ = ~new_n9389_ | ~new_n9348_;
  assign new_n9413_ = ~new_n9260_ | ~new_n9255_;
  assign new_n9414_ = ~new_n9211_;
  assign new_n9415_ = ~new_n9270_ | ~new_n9265_;
  assign new_n9416_ = ~pi042 | ~new_n9212_;
  assign new_n9417_ = ~new_n9368_ | ~new_n9343_;
  assign new_n9418_ = ~pi038 | ~new_n9213_;
  assign new_n9419_ = ~new_n9365_ | ~new_n9345_;
  assign new_n9420_ = ~new_n9412_ | ~new_n9347_;
  assign new_n9421_ = ~pi064 | ~new_n9389_ | ~new_n9348_;
  assign new_n9422_ = ~pi063 | ~new_n9217_;
  assign new_n9423_ = ~new_n9389_ | ~new_n9348_;
  assign new_n9424_ = ~new_n9387_ | ~pi060;
  assign new_n9425_ = ~new_n9415_ | ~new_n9350_;
  assign new_n9426_ = ~pi058 | ~new_n9353_;
  assign new_n9427_ = ~new_n9386_ | ~new_n9352_;
  assign new_n9428_ = ~pi054 | ~new_n9356_;
  assign new_n9429_ = ~new_n9383_ | ~new_n9355_;
  assign new_n9430_ = ~pi034 | ~new_n9359_;
  assign new_n9431_ = ~pi033 | ~new_n9358_;
  assign new_n9432_ = ~pi050 | ~new_n9218_;
  assign new_n9433_ = ~new_n9380_ | ~new_n9360_;
  assign new_n9434_ = ~pi046 | ~new_n9219_;
  assign new_n9435_ = ~new_n9377_ | ~new_n9362_;
  assign new_n9436_ = ~new_n1396_;
  assign new_n9437_ = ~new_n1393_;
  assign new_n9438_ = new_n9440_ & new_n9439_;
  assign new_n9439_ = ~new_n1393_ | ~new_n9436_;
  assign new_n9440_ = ~new_n1396_ | ~new_n9437_;
  assign new_n9441_ = new_n9570_ & new_n9470_;
  assign new_n9442_ = new_n9568_ & new_n9471_;
  assign new_n9443_ = new_n9567_ & new_n9472_;
  assign new_n9444_ = new_n9566_ & new_n9473_;
  assign new_n9445_ = new_n9564_ & new_n9474_;
  assign new_n9446_ = new_n9563_ & new_n9475_;
  assign new_n9447_ = new_n9562_ & new_n9476_;
  assign new_n9448_ = new_n9560_ & new_n9477_;
  assign new_n9449_ = new_n9558_ & new_n9478_;
  assign new_n9450_ = new_n9556_ & new_n9479_;
  assign new_n9451_ = new_n9554_ & new_n9480_;
  assign new_n9452_ = new_n9552_ & new_n9481_;
  assign new_n9453_ = new_n9550_ & new_n9460_;
  assign new_n9454_ = new_n9548_ & new_n9502_;
  assign new_n9455_ = new_n9533_ & new_n9461_;
  assign new_n9456_ = new_n9532_ & new_n9462_;
  assign new_n9457_ = new_n9531_ & new_n9463_;
  assign new_n9458_ = new_n9529_ & new_n9464_;
  assign new_n9459_ = new_n9528_ & new_n9465_;
  assign new_n9460_ = new_n1790_ | new_n1798_ | new_n1795_;
  assign new_n9461_ = ~new_n9522_ | ~new_n9469_;
  assign new_n9462_ = ~new_n9523_ | ~new_n9468_;
  assign new_n9463_ = ~new_n9493_ | ~new_n9524_;
  assign new_n9464_ = ~new_n9525_ | ~new_n9467_;
  assign new_n9465_ = ~new_n9526_ | ~new_n9466_;
  assign new_n9466_ = ~new_n1816_;
  assign new_n9467_ = ~new_n1813_;
  assign new_n9468_ = ~new_n1804_;
  assign new_n9469_ = ~new_n1801_;
  assign new_n9470_ = ~new_n9494_ | ~new_n9527_;
  assign new_n9471_ = ~new_n9534_ | ~new_n9491_;
  assign new_n9472_ = ~new_n9535_ | ~new_n9490_;
  assign new_n9473_ = ~new_n9495_ | ~new_n9536_;
  assign new_n9474_ = ~new_n9537_ | ~new_n9489_;
  assign new_n9475_ = ~new_n9538_ | ~new_n9488_;
  assign new_n9476_ = ~new_n9496_ | ~new_n9539_;
  assign new_n9477_ = ~new_n9487_ | ~new_n9540_ | ~new_n9516_;
  assign new_n9478_ = ~new_n9486_ | ~new_n9541_ | ~new_n9512_;
  assign new_n9479_ = ~new_n9485_ | ~new_n9542_ | ~new_n9510_;
  assign new_n9480_ = ~new_n9484_ | ~new_n9543_ | ~new_n9508_;
  assign new_n9481_ = ~new_n9483_ | ~new_n9544_ | ~new_n9506_;
  assign new_n9482_ = ~new_n2356_;
  assign new_n9483_ = ~new_n2346_;
  assign new_n9484_ = ~new_n2348_;
  assign new_n9485_ = ~new_n2350_;
  assign new_n9486_ = ~new_n2352_;
  assign new_n9487_ = ~new_n2354_;
  assign new_n9488_ = ~new_n1840_;
  assign new_n9489_ = ~new_n1837_;
  assign new_n9490_ = ~new_n1828_;
  assign new_n9491_ = ~new_n1825_;
  assign new_n9492_ = ~new_n9588_ | ~new_n9587_;
  assign new_n9493_ = ~new_n1807_ & ~new_n1810_;
  assign new_n9494_ = ~new_n1822_ & ~new_n1819_;
  assign new_n9495_ = ~new_n1831_ & ~new_n1834_;
  assign new_n9496_ = ~new_n1843_ & ~new_n1846_;
  assign new_n9497_ = ~new_n1819_;
  assign new_n9498_ = new_n9572_ & new_n9571_;
  assign new_n9499_ = ~new_n1807_;
  assign new_n9500_ = new_n9574_ & new_n9573_;
  assign new_n9501_ = ~new_n2355_;
  assign new_n9502_ = ~new_n9482_ | ~new_n9545_ | ~new_n9504_;
  assign new_n9503_ = new_n9576_ & new_n9575_;
  assign new_n9504_ = ~new_n2357_;
  assign new_n9505_ = new_n9578_ & new_n9577_;
  assign new_n9506_ = ~new_n2347_;
  assign new_n9507_ = new_n9580_ & new_n9579_;
  assign new_n9508_ = ~new_n2349_;
  assign new_n9509_ = new_n9582_ & new_n9581_;
  assign new_n9510_ = ~new_n2351_;
  assign new_n9511_ = new_n9584_ & new_n9583_;
  assign new_n9512_ = ~new_n2353_;
  assign new_n9513_ = new_n9586_ & new_n9585_;
  assign new_n9514_ = ~new_n1795_;
  assign new_n9515_ = ~new_n1790_;
  assign new_n9516_ = ~new_n1848_;
  assign new_n9517_ = new_n9590_ & new_n9589_;
  assign new_n9518_ = ~new_n1843_;
  assign new_n9519_ = new_n9592_ & new_n9591_;
  assign new_n9520_ = ~new_n1831_;
  assign new_n9521_ = new_n9594_ & new_n9593_;
  assign new_n9522_ = ~new_n9460_;
  assign new_n9523_ = ~new_n9461_;
  assign new_n9524_ = ~new_n9462_;
  assign new_n9525_ = ~new_n9463_;
  assign new_n9526_ = ~new_n9464_;
  assign new_n9527_ = ~new_n9465_;
  assign new_n9528_ = ~new_n1816_ | ~new_n9464_;
  assign new_n9529_ = ~new_n1813_ | ~new_n9463_;
  assign new_n9530_ = ~new_n9524_ | ~new_n9499_;
  assign new_n9531_ = ~new_n1810_ | ~new_n9530_;
  assign new_n9532_ = ~new_n1804_ | ~new_n9461_;
  assign new_n9533_ = ~new_n1801_ | ~new_n9460_;
  assign new_n9534_ = ~new_n9470_;
  assign new_n9535_ = ~new_n9471_;
  assign new_n9536_ = ~new_n9472_;
  assign new_n9537_ = ~new_n9473_;
  assign new_n9538_ = ~new_n9474_;
  assign new_n9539_ = ~new_n9475_;
  assign new_n9540_ = ~new_n9476_;
  assign new_n9541_ = ~new_n9477_;
  assign new_n9542_ = ~new_n9478_;
  assign new_n9543_ = ~new_n9479_;
  assign new_n9544_ = ~new_n9480_;
  assign new_n9545_ = ~new_n9481_;
  assign new_n9546_ = ~new_n9502_;
  assign new_n9547_ = ~new_n9545_ | ~new_n9504_;
  assign new_n9548_ = ~new_n2356_ | ~new_n9547_;
  assign new_n9549_ = new_n1795_ | new_n1790_;
  assign new_n9550_ = ~new_n1798_ | ~new_n9549_;
  assign new_n9551_ = ~new_n9544_ | ~new_n9506_;
  assign new_n9552_ = ~new_n2346_ | ~new_n9551_;
  assign new_n9553_ = ~new_n9543_ | ~new_n9508_;
  assign new_n9554_ = ~new_n2348_ | ~new_n9553_;
  assign new_n9555_ = ~new_n9542_ | ~new_n9510_;
  assign new_n9556_ = ~new_n2350_ | ~new_n9555_;
  assign new_n9557_ = ~new_n9541_ | ~new_n9512_;
  assign new_n9558_ = ~new_n2352_ | ~new_n9557_;
  assign new_n9559_ = ~new_n9540_ | ~new_n9516_;
  assign new_n9560_ = ~new_n2354_ | ~new_n9559_;
  assign new_n9561_ = ~new_n9539_ | ~new_n9518_;
  assign new_n9562_ = ~new_n1846_ | ~new_n9561_;
  assign new_n9563_ = ~new_n1840_ | ~new_n9474_;
  assign new_n9564_ = ~new_n1837_ | ~new_n9473_;
  assign new_n9565_ = ~new_n9536_ | ~new_n9520_;
  assign new_n9566_ = ~new_n1834_ | ~new_n9565_;
  assign new_n9567_ = ~new_n1828_ | ~new_n9471_;
  assign new_n9568_ = ~new_n1825_ | ~new_n9470_;
  assign new_n9569_ = ~new_n9527_ | ~new_n9497_;
  assign new_n9570_ = ~new_n1822_ | ~new_n9569_;
  assign new_n9571_ = ~new_n1819_ | ~new_n9465_;
  assign new_n9572_ = ~new_n9527_ | ~new_n9497_;
  assign new_n9573_ = ~new_n1807_ | ~new_n9462_;
  assign new_n9574_ = ~new_n9524_ | ~new_n9499_;
  assign new_n9575_ = ~new_n2355_ | ~new_n9502_;
  assign new_n9576_ = ~new_n9546_ | ~new_n9501_;
  assign new_n9577_ = ~new_n2357_ | ~new_n9481_;
  assign new_n9578_ = ~new_n9545_ | ~new_n9504_;
  assign new_n9579_ = ~new_n2347_ | ~new_n9480_;
  assign new_n9580_ = ~new_n9544_ | ~new_n9506_;
  assign new_n9581_ = ~new_n2349_ | ~new_n9479_;
  assign new_n9582_ = ~new_n9543_ | ~new_n9508_;
  assign new_n9583_ = ~new_n2351_ | ~new_n9478_;
  assign new_n9584_ = ~new_n9542_ | ~new_n9510_;
  assign new_n9585_ = ~new_n2353_ | ~new_n9477_;
  assign new_n9586_ = ~new_n9541_ | ~new_n9512_;
  assign new_n9587_ = ~new_n1795_ | ~new_n9515_;
  assign new_n9588_ = ~new_n1790_ | ~new_n9514_;
  assign new_n9589_ = ~new_n1848_ | ~new_n9476_;
  assign new_n9590_ = ~new_n9540_ | ~new_n9516_;
  assign new_n9591_ = ~new_n1843_ | ~new_n9475_;
  assign new_n9592_ = ~new_n9539_ | ~new_n9518_;
  assign new_n9593_ = ~new_n1831_ | ~new_n9472_;
  assign new_n9594_ = ~new_n9536_ | ~new_n9520_;
  assign new_n9595_ = new_n9767_ & new_n9766_;
  assign new_n9596_ = new_n9768_ & new_n9769_;
  assign new_n9597_ = new_n9785_ & new_n9784_;
  assign new_n9598_ = new_n9825_ & new_n9824_;
  assign new_n9599_ = new_n9834_ & new_n9833_;
  assign new_n9600_ = new_n9852_ & new_n9851_;
  assign new_n9601_ = new_n9860_ & new_n9859_;
  assign new_n9602_ = new_n9939_ & new_n9936_;
  assign new_n9603_ = new_n9932_ & new_n9929_;
  assign new_n9604_ = new_n9923_ & new_n9920_;
  assign new_n9605_ = new_n9914_ & new_n9911_;
  assign new_n9606_ = new_n9908_ & new_n9906_;
  assign new_n9607_ = new_n9901_ & new_n9898_;
  assign new_n9608_ = new_n9823_ & new_n9820_;
  assign new_n9609_ = new_n9815_ & new_n9812_;
  assign new_n9610_ = new_n9801_ & new_n9798_;
  assign new_n9611_ = ~new_n1810_;
  assign new_n9612_ = ~new_n1408_;
  assign new_n9613_ = ~new_n1407_;
  assign new_n9614_ = ~new_n1408_ | ~new_n1810_;
  assign new_n9615_ = ~new_n1813_;
  assign new_n9616_ = ~new_n1804_;
  assign new_n9617_ = ~new_n1397_;
  assign new_n9618_ = ~new_n1404_;
  assign new_n9619_ = ~new_n1798_;
  assign new_n9620_ = ~new_n1405_;
  assign new_n9621_ = ~new_n1790_;
  assign new_n9622_ = ~new_n1414_;
  assign new_n9623_ = ~new_n1414_ | ~new_n1790_;
  assign new_n9624_ = ~new_n1801_;
  assign new_n9625_ = ~new_n1401_;
  assign new_n9626_ = ~new_n1397_ | ~new_n1804_;
  assign new_n9627_ = ~new_n1807_;
  assign new_n9628_ = ~new_n1816_;
  assign new_n9629_ = ~new_n1421_;
  assign new_n9630_ = ~new_n1420_;
  assign new_n9631_ = ~new_n1819_;
  assign new_n9632_ = ~new_n9653_ | ~new_n9793_;
  assign new_n9633_ = ~new_n9709_ | ~new_n9781_;
  assign new_n9634_ = ~new_n9770_ | ~new_n9771_;
  assign new_n9635_ = ~new_n1795_ | ~new_n1415_;
  assign new_n9636_ = ~new_n9713_ | ~new_n9807_;
  assign new_n9637_ = ~new_n9804_ | ~new_n9803_;
  assign new_n9638_ = ~new_n2347_;
  assign new_n9639_ = ~new_n1390_;
  assign new_n9640_ = ~new_n1394_;
  assign new_n9641_ = ~new_n2348_;
  assign new_n9642_ = ~new_n2349_;
  assign new_n9643_ = ~new_n1395_;
  assign new_n9644_ = ~new_n2350_;
  assign new_n9645_ = ~new_n1402_;
  assign new_n9646_ = ~new_n2353_;
  assign new_n9647_ = ~new_n1412_;
  assign new_n9648_ = ~new_n1840_;
  assign new_n9649_ = ~new_n1410_;
  assign new_n9650_ = ~new_n1406_;
  assign new_n9651_ = ~new_n1410_ | ~new_n1840_;
  assign new_n9652_ = ~new_n1843_;
  assign new_n9653_ = ~new_n1421_ | ~new_n1816_;
  assign new_n9654_ = ~new_n1822_;
  assign new_n9655_ = ~new_n1399_;
  assign new_n9656_ = ~new_n1828_;
  assign new_n9657_ = ~new_n1409_;
  assign new_n9658_ = ~new_n1825_;
  assign new_n9659_ = ~new_n1400_;
  assign new_n9660_ = ~new_n1400_ | ~new_n1825_;
  assign new_n9661_ = ~new_n1831_;
  assign new_n9662_ = ~new_n1417_;
  assign new_n9663_ = ~new_n1834_;
  assign new_n9664_ = ~new_n1416_;
  assign new_n9665_ = ~new_n1837_;
  assign new_n9666_ = ~new_n1411_;
  assign new_n9667_ = ~new_n1846_;
  assign new_n9668_ = ~new_n1419_;
  assign new_n9669_ = ~new_n1419_ | ~new_n1846_;
  assign new_n9670_ = ~new_n1848_;
  assign new_n9671_ = ~new_n1418_;
  assign new_n9672_ = ~new_n1418_ | ~new_n1848_;
  assign new_n9673_ = ~new_n2354_;
  assign new_n9674_ = ~new_n2352_;
  assign new_n9675_ = ~new_n1398_;
  assign new_n9676_ = ~new_n2351_;
  assign new_n9677_ = ~new_n1403_;
  assign new_n9678_ = ~new_n2348_ | ~new_n1394_;
  assign new_n9679_ = ~new_n1391_;
  assign new_n9680_ = ~new_n2346_;
  assign new_n9681_ = ~new_n9894_ | ~new_n9764_;
  assign new_n9682_ = ~new_n1413_;
  assign new_n9683_ = ~new_n9669_ | ~new_n9903_;
  assign new_n9684_ = ~new_n9849_ | ~new_n9848_;
  assign new_n9685_ = ~new_n9660_ | ~new_n9925_;
  assign new_n9686_ = ~new_n10045_ | ~new_n10044_;
  assign new_n9687_ = ~new_n10092_ | ~new_n10091_;
  assign new_n9688_ = ~new_n9963_ | ~new_n9962_;
  assign new_n9689_ = ~new_n9968_ | ~new_n9967_;
  assign new_n9690_ = ~new_n9975_ | ~new_n9974_;
  assign new_n9691_ = ~new_n9982_ | ~new_n9981_;
  assign new_n9692_ = ~new_n9987_ | ~new_n9986_;
  assign new_n9693_ = ~new_n9996_ | ~new_n9995_;
  assign new_n9694_ = ~new_n10003_ | ~new_n10002_;
  assign new_n9695_ = ~new_n10010_ | ~new_n10009_;
  assign new_n9696_ = ~new_n10017_ | ~new_n10016_;
  assign new_n9697_ = ~new_n10022_ | ~new_n10021_;
  assign new_n9698_ = ~new_n10029_ | ~new_n10028_;
  assign new_n9699_ = ~new_n10036_ | ~new_n10035_;
  assign new_n9700_ = ~new_n10050_ | ~new_n10049_;
  assign new_n9701_ = ~new_n10055_ | ~new_n10054_;
  assign new_n9702_ = ~new_n10062_ | ~new_n10061_;
  assign new_n9703_ = ~new_n10069_ | ~new_n10068_;
  assign new_n9704_ = ~new_n10076_ | ~new_n10075_;
  assign new_n9705_ = ~new_n10083_ | ~new_n10082_;
  assign new_n9706_ = ~new_n10088_ | ~new_n10087_;
  assign new_n9707_ = new_n1798_ & new_n1405_;
  assign new_n9708_ = new_n9777_ & new_n9775_;
  assign new_n9709_ = new_n9782_ & new_n9780_;
  assign new_n9710_ = new_n9789_ & new_n9788_;
  assign new_n9711_ = new_n9614_ & new_n9970_ & new_n9969_;
  assign new_n9712_ = new_n9800_ & new_n9597_;
  assign new_n9713_ = new_n9808_ & new_n9806_;
  assign new_n9714_ = new_n9626_ & new_n9977_ & new_n9976_;
  assign new_n9715_ = new_n9814_ & new_n9595_;
  assign new_n9716_ = new_n9822_ & new_n9769_;
  assign new_n9717_ = new_n9792_ & new_n9598_;
  assign new_n9718_ = new_n9827_ & new_n9759_;
  assign new_n9719_ = new_n9836_ & new_n9760_;
  assign new_n9720_ = new_n9856_ & new_n9855_;
  assign new_n9721_ = new_n9601_ & new_n9870_;
  assign new_n9722_ = new_n9873_ & new_n9868_;
  assign new_n9723_ = new_n9889_ & new_n9886_;
  assign new_n9724_ = new_n9956_ & new_n9890_;
  assign new_n9725_ = new_n9747_ & new_n9866_;
  assign new_n9726_ = new_n9651_ & new_n10057_ & new_n10056_;
  assign new_n9727_ = new_n9760_ & new_n10078_ & new_n10077_;
  assign new_n9728_ = new_n9931_ & new_n9599_;
  assign new_n9729_ = new_n9759_ & new_n10090_ & new_n10089_;
  assign new_n9730_ = new_n9938_ & new_n9598_;
  assign new_n9731_ = ~new_n9710_ | ~new_n9790_;
  assign new_n9732_ = ~new_n9805_ | ~new_n9817_;
  assign new_n9733_ = ~new_n1392_;
  assign new_n9734_ = ~new_n2357_;
  assign new_n9735_ = new_n9991_ & new_n9990_;
  assign new_n9736_ = ~new_n9952_ | ~new_n9892_ | ~new_n9757_;
  assign new_n9737_ = new_n9998_ & new_n9997_;
  assign new_n9738_ = ~new_n9724_ | ~new_n9958_ | ~new_n9957_;
  assign new_n9739_ = new_n10005_ & new_n10004_;
  assign new_n9740_ = ~new_n9678_ | ~new_n9953_ | ~new_n9887_;
  assign new_n9741_ = new_n10012_ & new_n10011_;
  assign new_n9742_ = ~new_n9881_ | ~new_n9880_;
  assign new_n9743_ = new_n10024_ & new_n10023_;
  assign new_n9744_ = ~new_n9877_ | ~new_n9876_;
  assign new_n9745_ = new_n10031_ & new_n10030_;
  assign new_n9746_ = ~new_n9722_ | ~new_n9872_;
  assign new_n9747_ = new_n10038_ & new_n10037_;
  assign new_n9748_ = new_n10043_ & new_n10042_;
  assign new_n9749_ = ~new_n9635_ | ~new_n9915_;
  assign new_n9750_ = ~new_n9720_ | ~new_n9857_;
  assign new_n9751_ = new_n10064_ & new_n10063_;
  assign new_n9752_ = ~new_n9845_ | ~new_n9844_;
  assign new_n9753_ = new_n10071_ & new_n10070_;
  assign new_n9754_ = ~new_n9841_ | ~new_n9840_;
  assign new_n9755_ = ~new_n9831_ | ~new_n9830_;
  assign new_n9756_ = ~new_n9955_ | ~new_n9954_;
  assign new_n9757_ = ~new_n1391_ | ~new_n9738_;
  assign new_n9758_ = ~new_n9626_;
  assign new_n9759_ = ~new_n1819_ | ~new_n1420_;
  assign new_n9760_ = ~new_n1409_ | ~new_n1828_;
  assign new_n9761_ = ~new_n1395_ | ~new_n2349_;
  assign new_n9762_ = ~new_n9660_;
  assign new_n9763_ = ~new_n9669_;
  assign new_n9764_ = ~new_n1402_ | ~new_n2350_;
  assign new_n9765_ = ~new_n9653_;
  assign new_n9766_ = new_n1404_ | new_n1807_;
  assign new_n9767_ = new_n1397_ | new_n1804_;
  assign new_n9768_ = new_n1801_ | new_n1401_;
  assign new_n9769_ = new_n1798_ | new_n1405_;
  assign new_n9770_ = ~new_n9623_;
  assign new_n9771_ = new_n1795_ | new_n1415_;
  assign new_n9772_ = ~new_n9634_;
  assign new_n9773_ = ~new_n9635_;
  assign new_n9774_ = ~new_n9634_ | ~new_n9635_;
  assign new_n9775_ = ~new_n9707_ | ~new_n9768_;
  assign new_n9776_ = ~new_n9596_ | ~new_n9774_;
  assign new_n9777_ = ~new_n1401_ | ~new_n1801_;
  assign new_n9778_ = ~new_n9708_ | ~new_n9776_;
  assign new_n9779_ = ~new_n9627_ | ~new_n9626_;
  assign new_n9780_ = ~new_n1404_ | ~new_n9779_;
  assign new_n9781_ = ~new_n9595_ | ~new_n9778_;
  assign new_n9782_ = ~new_n1807_ | ~new_n9758_;
  assign new_n9783_ = ~new_n9633_;
  assign new_n9784_ = new_n1407_ | new_n1813_;
  assign new_n9785_ = new_n1408_ | new_n1810_;
  assign new_n9786_ = ~new_n9614_;
  assign new_n9787_ = ~new_n9615_ | ~new_n9614_;
  assign new_n9788_ = ~new_n1407_ | ~new_n9787_;
  assign new_n9789_ = ~new_n1813_ | ~new_n9786_;
  assign new_n9790_ = ~new_n9597_ | ~new_n9633_;
  assign new_n9791_ = ~new_n9731_;
  assign new_n9792_ = new_n1816_ | new_n1421_;
  assign new_n9793_ = ~new_n9792_ | ~new_n9731_;
  assign new_n9794_ = ~new_n9632_;
  assign new_n9795_ = new_n1420_ | new_n1819_;
  assign new_n9796_ = new_n1810_ | new_n1408_;
  assign new_n9797_ = ~new_n9796_ | ~new_n9633_;
  assign new_n9798_ = ~new_n9711_ | ~new_n9797_;
  assign new_n9799_ = ~new_n9783_ | ~new_n9614_;
  assign new_n9800_ = ~new_n1813_ | ~new_n1407_;
  assign new_n9801_ = ~new_n9712_ | ~new_n9799_;
  assign new_n9802_ = new_n1408_ | new_n1810_;
  assign new_n9803_ = ~new_n9773_ | ~new_n9769_;
  assign new_n9804_ = ~new_n1405_ | ~new_n1798_;
  assign new_n9805_ = ~new_n9637_;
  assign new_n9806_ = ~new_n9772_ | ~new_n9596_;
  assign new_n9807_ = ~new_n9637_ | ~new_n9768_;
  assign new_n9808_ = ~new_n1401_ | ~new_n1801_;
  assign new_n9809_ = ~new_n9636_;
  assign new_n9810_ = new_n1804_ | new_n1397_;
  assign new_n9811_ = ~new_n9810_ | ~new_n9636_;
  assign new_n9812_ = ~new_n9714_ | ~new_n9811_;
  assign new_n9813_ = ~new_n9809_ | ~new_n9626_;
  assign new_n9814_ = ~new_n1807_ | ~new_n1404_;
  assign new_n9815_ = ~new_n9715_ | ~new_n9813_;
  assign new_n9816_ = new_n1397_ | new_n1804_;
  assign new_n9817_ = ~new_n9772_ | ~new_n9769_;
  assign new_n9818_ = ~new_n9732_;
  assign new_n9819_ = ~new_n1401_ | ~new_n1801_;
  assign new_n9820_ = ~new_n9634_ | ~new_n9635_ | ~new_n9989_ | ~new_n9988_;
  assign new_n9821_ = ~new_n9635_ | ~new_n9634_;
  assign new_n9822_ = ~new_n1405_ | ~new_n1798_;
  assign new_n9823_ = ~new_n9716_ | ~new_n9821_;
  assign new_n9824_ = new_n1420_ | new_n1819_;
  assign new_n9825_ = new_n1399_ | new_n1822_;
  assign new_n9826_ = ~new_n9765_ | ~new_n9598_;
  assign new_n9827_ = ~new_n1399_ | ~new_n1822_;
  assign new_n9828_ = ~new_n9718_ | ~new_n9826_;
  assign new_n9829_ = new_n1822_ | new_n1399_;
  assign new_n9830_ = ~new_n9717_ | ~new_n9731_;
  assign new_n9831_ = ~new_n9829_ | ~new_n9828_;
  assign new_n9832_ = ~new_n9755_;
  assign new_n9833_ = new_n1417_ | new_n1831_;
  assign new_n9834_ = new_n1409_ | new_n1828_;
  assign new_n9835_ = ~new_n9762_ | ~new_n9599_;
  assign new_n9836_ = ~new_n1417_ | ~new_n1831_;
  assign new_n9837_ = ~new_n9719_ | ~new_n9835_;
  assign new_n9838_ = new_n1825_ | new_n1400_;
  assign new_n9839_ = new_n1831_ | new_n1417_;
  assign new_n9840_ = ~new_n9599_ | ~new_n9838_ | ~new_n9755_;
  assign new_n9841_ = ~new_n9839_ | ~new_n9837_;
  assign new_n9842_ = ~new_n9754_;
  assign new_n9843_ = new_n1834_ | new_n1416_;
  assign new_n9844_ = ~new_n9843_ | ~new_n9754_;
  assign new_n9845_ = ~new_n1416_ | ~new_n1834_;
  assign new_n9846_ = ~new_n9752_;
  assign new_n9847_ = new_n1837_ | new_n1411_;
  assign new_n9848_ = ~new_n9847_ | ~new_n9752_;
  assign new_n9849_ = ~new_n1411_ | ~new_n1837_;
  assign new_n9850_ = ~new_n9684_;
  assign new_n9851_ = new_n1406_ | new_n1843_;
  assign new_n9852_ = new_n1410_ | new_n1840_;
  assign new_n9853_ = ~new_n9651_;
  assign new_n9854_ = ~new_n9652_ | ~new_n9651_;
  assign new_n9855_ = ~new_n1406_ | ~new_n9854_;
  assign new_n9856_ = ~new_n1843_ | ~new_n9853_;
  assign new_n9857_ = ~new_n9600_ | ~new_n9684_;
  assign new_n9858_ = ~new_n9750_;
  assign new_n9859_ = new_n1413_ | new_n2354_;
  assign new_n9860_ = new_n1418_ | new_n1848_;
  assign new_n9861_ = new_n1412_ | new_n2353_;
  assign new_n9862_ = ~new_n9672_;
  assign new_n9863_ = ~new_n2354_ | ~new_n9862_;
  assign new_n9864_ = ~new_n9863_ | ~new_n9682_;
  assign new_n9865_ = ~new_n9672_ | ~new_n9673_;
  assign new_n9866_ = ~new_n9865_ | ~new_n9864_;
  assign new_n9867_ = ~new_n9763_ | ~new_n9601_;
  assign new_n9868_ = ~new_n1412_ | ~new_n2353_;
  assign new_n9869_ = ~new_n9866_ | ~new_n9867_;
  assign new_n9870_ = new_n1846_ | new_n1419_;
  assign new_n9871_ = new_n2353_ | new_n1412_;
  assign new_n9872_ = ~new_n9721_ | ~new_n9861_ | ~new_n9750_;
  assign new_n9873_ = ~new_n9871_ | ~new_n9869_;
  assign new_n9874_ = ~new_n9746_;
  assign new_n9875_ = new_n2352_ | new_n1398_;
  assign new_n9876_ = ~new_n9875_ | ~new_n9746_;
  assign new_n9877_ = ~new_n1398_ | ~new_n2352_;
  assign new_n9878_ = ~new_n9744_;
  assign new_n9879_ = new_n2351_ | new_n1403_;
  assign new_n9880_ = ~new_n9879_ | ~new_n9744_;
  assign new_n9881_ = ~new_n1403_ | ~new_n2351_;
  assign new_n9882_ = ~new_n9742_;
  assign new_n9883_ = new_n1395_ | new_n2349_;
  assign new_n9884_ = ~new_n9764_ | ~new_n9761_;
  assign new_n9885_ = ~new_n9678_;
  assign new_n9886_ = new_n2350_ | new_n1402_;
  assign new_n9887_ = ~new_n9756_ | ~new_n9742_ | ~new_n9886_;
  assign new_n9888_ = ~new_n9740_;
  assign new_n9889_ = new_n2347_ | new_n1390_;
  assign new_n9890_ = ~new_n1390_ | ~new_n2347_;
  assign new_n9891_ = ~new_n9738_;
  assign new_n9892_ = ~new_n2346_ | ~new_n9738_;
  assign new_n9893_ = ~new_n9736_;
  assign new_n9894_ = ~new_n9886_ | ~new_n9742_;
  assign new_n9895_ = ~new_n9681_;
  assign new_n9896_ = new_n2349_ | new_n1395_;
  assign new_n9897_ = ~new_n9896_ | ~new_n9681_;
  assign new_n9898_ = ~new_n9741_ | ~new_n9897_ | ~new_n9761_;
  assign new_n9899_ = ~new_n9895_ | ~new_n9761_;
  assign new_n9900_ = ~new_n2348_ | ~new_n1394_;
  assign new_n9901_ = ~new_n9756_ | ~new_n9899_ | ~new_n9900_;
  assign new_n9902_ = new_n1395_ | new_n2349_;
  assign new_n9903_ = ~new_n9870_ | ~new_n9750_;
  assign new_n9904_ = ~new_n9683_;
  assign new_n9905_ = ~new_n9601_ | ~new_n9683_;
  assign new_n9906_ = ~new_n9725_ | ~new_n9905_;
  assign new_n9907_ = ~new_n9905_ | ~new_n9866_;
  assign new_n9908_ = ~new_n10041_ | ~new_n9907_;
  assign new_n9909_ = new_n1848_ | new_n1418_;
  assign new_n9910_ = ~new_n9909_ | ~new_n9683_;
  assign new_n9911_ = ~new_n9748_ | ~new_n9910_ | ~new_n9672_;
  assign new_n9912_ = ~new_n9904_ | ~new_n9672_;
  assign new_n9913_ = ~new_n1413_ | ~new_n2354_;
  assign new_n9914_ = ~new_n9601_ | ~new_n9913_ | ~new_n9912_;
  assign new_n9915_ = new_n1795_ | new_n1415_;
  assign new_n9916_ = ~new_n9749_;
  assign new_n9917_ = new_n1418_ | new_n1848_;
  assign new_n9918_ = new_n1840_ | new_n1410_;
  assign new_n9919_ = ~new_n9918_ | ~new_n9684_;
  assign new_n9920_ = ~new_n9726_ | ~new_n9919_;
  assign new_n9921_ = ~new_n9850_ | ~new_n9651_;
  assign new_n9922_ = ~new_n1843_ | ~new_n1406_;
  assign new_n9923_ = ~new_n9600_ | ~new_n9922_ | ~new_n9921_;
  assign new_n9924_ = new_n1410_ | new_n1840_;
  assign new_n9925_ = ~new_n9838_ | ~new_n9755_;
  assign new_n9926_ = ~new_n9685_;
  assign new_n9927_ = new_n1828_ | new_n1409_;
  assign new_n9928_ = ~new_n9927_ | ~new_n9685_;
  assign new_n9929_ = ~new_n9727_ | ~new_n9928_;
  assign new_n9930_ = ~new_n9926_ | ~new_n9760_;
  assign new_n9931_ = ~new_n1417_ | ~new_n1831_;
  assign new_n9932_ = ~new_n9728_ | ~new_n9930_;
  assign new_n9933_ = new_n1409_ | new_n1828_;
  assign new_n9934_ = new_n1819_ | new_n1420_;
  assign new_n9935_ = ~new_n9934_ | ~new_n9632_;
  assign new_n9936_ = ~new_n9729_ | ~new_n9935_;
  assign new_n9937_ = ~new_n9794_ | ~new_n9759_;
  assign new_n9938_ = ~new_n1399_ | ~new_n1822_;
  assign new_n9939_ = ~new_n9730_ | ~new_n9937_;
  assign new_n9940_ = ~new_n9795_ | ~new_n9759_;
  assign new_n9941_ = ~new_n9792_ | ~new_n9653_;
  assign new_n9942_ = ~new_n9802_ | ~new_n9614_;
  assign new_n9943_ = ~new_n9816_ | ~new_n9626_;
  assign new_n9944_ = ~new_n9819_ | ~new_n9768_;
  assign new_n9945_ = ~new_n9902_ | ~new_n9761_;
  assign new_n9946_ = ~new_n9886_ | ~new_n9764_;
  assign new_n9947_ = ~new_n9917_ | ~new_n9672_;
  assign new_n9948_ = ~new_n9870_ | ~new_n9669_;
  assign new_n9949_ = ~new_n9924_ | ~new_n9651_;
  assign new_n9950_ = ~new_n9933_ | ~new_n9760_;
  assign new_n9951_ = ~new_n9838_ | ~new_n9660_;
  assign new_n9952_ = ~new_n2346_ | ~new_n1391_;
  assign new_n9953_ = ~new_n9884_ | ~new_n9756_;
  assign new_n9954_ = ~new_n1394_ | ~new_n9883_;
  assign new_n9955_ = ~new_n2348_ | ~new_n9883_;
  assign new_n9956_ = ~new_n9889_ | ~new_n9884_ | ~new_n9756_;
  assign new_n9957_ = ~new_n9723_ | ~new_n9742_ | ~new_n9756_;
  assign new_n9958_ = ~new_n9885_ | ~new_n9889_;
  assign new_n9959_ = ~new_n1420_ | ~new_n9631_;
  assign new_n9960_ = ~new_n1819_ | ~new_n9630_;
  assign new_n9961_ = ~new_n9960_ | ~new_n9959_;
  assign new_n9962_ = ~new_n9940_ | ~new_n9632_;
  assign new_n9963_ = ~new_n9961_ | ~new_n9794_;
  assign new_n9964_ = ~new_n1421_ | ~new_n9628_;
  assign new_n9965_ = ~new_n1816_ | ~new_n9629_;
  assign new_n9966_ = ~new_n9965_ | ~new_n9964_;
  assign new_n9967_ = ~new_n9941_ | ~new_n9731_;
  assign new_n9968_ = ~new_n9791_ | ~new_n9966_;
  assign new_n9969_ = ~new_n1407_ | ~new_n9615_;
  assign new_n9970_ = ~new_n1813_ | ~new_n9613_;
  assign new_n9971_ = ~new_n1408_ | ~new_n9611_;
  assign new_n9972_ = ~new_n1810_ | ~new_n9612_;
  assign new_n9973_ = ~new_n9972_ | ~new_n9971_;
  assign new_n9974_ = ~new_n9942_ | ~new_n9633_;
  assign new_n9975_ = ~new_n9973_ | ~new_n9783_;
  assign new_n9976_ = ~new_n1404_ | ~new_n9627_;
  assign new_n9977_ = ~new_n1807_ | ~new_n9618_;
  assign new_n9978_ = ~new_n1397_ | ~new_n9616_;
  assign new_n9979_ = ~new_n1804_ | ~new_n9617_;
  assign new_n9980_ = ~new_n9979_ | ~new_n9978_;
  assign new_n9981_ = ~new_n9943_ | ~new_n9636_;
  assign new_n9982_ = ~new_n9980_ | ~new_n9809_;
  assign new_n9983_ = ~new_n1401_ | ~new_n9624_;
  assign new_n9984_ = ~new_n1801_ | ~new_n9625_;
  assign new_n9985_ = ~new_n9984_ | ~new_n9983_;
  assign new_n9986_ = ~new_n9944_ | ~new_n9732_;
  assign new_n9987_ = ~new_n9818_ | ~new_n9985_;
  assign new_n9988_ = ~new_n1405_ | ~new_n9619_;
  assign new_n9989_ = ~new_n1798_ | ~new_n9620_;
  assign new_n9990_ = ~new_n1392_ | ~new_n9734_;
  assign new_n9991_ = ~new_n2357_ | ~new_n9733_;
  assign new_n9992_ = ~new_n1392_ | ~new_n9734_;
  assign new_n9993_ = ~new_n2357_ | ~new_n9733_;
  assign new_n9994_ = ~new_n9993_ | ~new_n9992_;
  assign new_n9995_ = ~new_n9735_ | ~new_n9736_;
  assign new_n9996_ = ~new_n9893_ | ~new_n9994_;
  assign new_n9997_ = ~new_n1391_ | ~new_n9680_;
  assign new_n9998_ = ~new_n2346_ | ~new_n9679_;
  assign new_n9999_ = ~new_n1391_ | ~new_n9680_;
  assign new_n10000_ = ~new_n2346_ | ~new_n9679_;
  assign new_n10001_ = ~new_n10000_ | ~new_n9999_;
  assign new_n10002_ = ~new_n9737_ | ~new_n9738_;
  assign new_n10003_ = ~new_n9891_ | ~new_n10001_;
  assign new_n10004_ = ~new_n1390_ | ~new_n9638_;
  assign new_n10005_ = ~new_n2347_ | ~new_n9639_;
  assign new_n10006_ = ~new_n1390_ | ~new_n9638_;
  assign new_n10007_ = ~new_n2347_ | ~new_n9639_;
  assign new_n10008_ = ~new_n10007_ | ~new_n10006_;
  assign new_n10009_ = ~new_n9739_ | ~new_n9740_;
  assign new_n10010_ = ~new_n9888_ | ~new_n10008_;
  assign new_n10011_ = ~new_n1394_ | ~new_n9641_;
  assign new_n10012_ = ~new_n2348_ | ~new_n9640_;
  assign new_n10013_ = ~new_n1395_ | ~new_n9642_;
  assign new_n10014_ = ~new_n2349_ | ~new_n9643_;
  assign new_n10015_ = ~new_n10014_ | ~new_n10013_;
  assign new_n10016_ = ~new_n9945_ | ~new_n9681_;
  assign new_n10017_ = ~new_n10015_ | ~new_n9895_;
  assign new_n10018_ = ~new_n1402_ | ~new_n9644_;
  assign new_n10019_ = ~new_n2350_ | ~new_n9645_;
  assign new_n10020_ = ~new_n10019_ | ~new_n10018_;
  assign new_n10021_ = ~new_n9946_ | ~new_n9742_;
  assign new_n10022_ = ~new_n9882_ | ~new_n10020_;
  assign new_n10023_ = ~new_n1403_ | ~new_n9676_;
  assign new_n10024_ = ~new_n2351_ | ~new_n9677_;
  assign new_n10025_ = ~new_n1403_ | ~new_n9676_;
  assign new_n10026_ = ~new_n2351_ | ~new_n9677_;
  assign new_n10027_ = ~new_n10026_ | ~new_n10025_;
  assign new_n10028_ = ~new_n9743_ | ~new_n9744_;
  assign new_n10029_ = ~new_n9878_ | ~new_n10027_;
  assign new_n10030_ = ~new_n1398_ | ~new_n9674_;
  assign new_n10031_ = ~new_n2352_ | ~new_n9675_;
  assign new_n10032_ = ~new_n1398_ | ~new_n9674_;
  assign new_n10033_ = ~new_n2352_ | ~new_n9675_;
  assign new_n10034_ = ~new_n10033_ | ~new_n10032_;
  assign new_n10035_ = ~new_n9745_ | ~new_n9746_;
  assign new_n10036_ = ~new_n9874_ | ~new_n10034_;
  assign new_n10037_ = ~new_n1412_ | ~new_n9646_;
  assign new_n10038_ = ~new_n2353_ | ~new_n9647_;
  assign new_n10039_ = ~new_n1412_ | ~new_n9646_;
  assign new_n10040_ = ~new_n2353_ | ~new_n9647_;
  assign new_n10041_ = ~new_n10040_ | ~new_n10039_;
  assign new_n10042_ = ~new_n1413_ | ~new_n9673_;
  assign new_n10043_ = ~new_n2354_ | ~new_n9682_;
  assign new_n10044_ = ~new_n9770_ | ~new_n9749_;
  assign new_n10045_ = ~new_n9916_ | ~new_n9623_;
  assign new_n10046_ = ~new_n1418_ | ~new_n9670_;
  assign new_n10047_ = ~new_n1848_ | ~new_n9671_;
  assign new_n10048_ = ~new_n10047_ | ~new_n10046_;
  assign new_n10049_ = ~new_n9947_ | ~new_n9683_;
  assign new_n10050_ = ~new_n10048_ | ~new_n9904_;
  assign new_n10051_ = ~new_n1419_ | ~new_n9667_;
  assign new_n10052_ = ~new_n1846_ | ~new_n9668_;
  assign new_n10053_ = ~new_n10052_ | ~new_n10051_;
  assign new_n10054_ = ~new_n9948_ | ~new_n9750_;
  assign new_n10055_ = ~new_n9858_ | ~new_n10053_;
  assign new_n10056_ = ~new_n1406_ | ~new_n9652_;
  assign new_n10057_ = ~new_n1843_ | ~new_n9650_;
  assign new_n10058_ = ~new_n1410_ | ~new_n9648_;
  assign new_n10059_ = ~new_n1840_ | ~new_n9649_;
  assign new_n10060_ = ~new_n10059_ | ~new_n10058_;
  assign new_n10061_ = ~new_n9949_ | ~new_n9684_;
  assign new_n10062_ = ~new_n10060_ | ~new_n9850_;
  assign new_n10063_ = ~new_n1411_ | ~new_n9665_;
  assign new_n10064_ = ~new_n1837_ | ~new_n9666_;
  assign new_n10065_ = ~new_n1411_ | ~new_n9665_;
  assign new_n10066_ = ~new_n1837_ | ~new_n9666_;
  assign new_n10067_ = ~new_n10066_ | ~new_n10065_;
  assign new_n10068_ = ~new_n9751_ | ~new_n9752_;
  assign new_n10069_ = ~new_n9846_ | ~new_n10067_;
  assign new_n10070_ = ~new_n1416_ | ~new_n9663_;
  assign new_n10071_ = ~new_n1834_ | ~new_n9664_;
  assign new_n10072_ = ~new_n1416_ | ~new_n9663_;
  assign new_n10073_ = ~new_n1834_ | ~new_n9664_;
  assign new_n10074_ = ~new_n10073_ | ~new_n10072_;
  assign new_n10075_ = ~new_n9753_ | ~new_n9754_;
  assign new_n10076_ = ~new_n9842_ | ~new_n10074_;
  assign new_n10077_ = ~new_n1417_ | ~new_n9661_;
  assign new_n10078_ = ~new_n1831_ | ~new_n9662_;
  assign new_n10079_ = ~new_n1409_ | ~new_n9656_;
  assign new_n10080_ = ~new_n1828_ | ~new_n9657_;
  assign new_n10081_ = ~new_n10080_ | ~new_n10079_;
  assign new_n10082_ = ~new_n9950_ | ~new_n9685_;
  assign new_n10083_ = ~new_n10081_ | ~new_n9926_;
  assign new_n10084_ = ~new_n1400_ | ~new_n9658_;
  assign new_n10085_ = ~new_n1825_ | ~new_n9659_;
  assign new_n10086_ = ~new_n10085_ | ~new_n10084_;
  assign new_n10087_ = ~new_n9951_ | ~new_n9755_;
  assign new_n10088_ = ~new_n9832_ | ~new_n10086_;
  assign new_n10089_ = ~new_n1399_ | ~new_n9654_;
  assign new_n10090_ = ~new_n1822_ | ~new_n9655_;
  assign new_n10091_ = ~new_n1414_ | ~new_n9621_;
  assign new_n10092_ = ~new_n1790_ | ~new_n9622_;
  assign new_n10093_ = new_n10184_ & new_n10183_;
  assign new_n10094_ = new_n10185_ & new_n10186_;
  assign new_n10095_ = new_n10202_ & new_n10201_;
  assign new_n10096_ = new_n10244_ & new_n10243_;
  assign new_n10097_ = new_n10253_ & new_n10252_;
  assign new_n10098_ = new_n10271_ & new_n10270_;
  assign new_n10099_ = new_n10307_ & new_n10304_;
  assign new_n10100_ = new_n10300_ & new_n10297_;
  assign new_n10101_ = new_n10291_ & new_n10288_;
  assign new_n10102_ = new_n10285_ & new_n10281_;
  assign new_n10103_ = new_n10240_ & new_n10237_;
  assign new_n10104_ = new_n10232_ & new_n10229_;
  assign new_n10105_ = new_n10218_ & new_n10215_;
  assign new_n10106_ = ~pi135;
  assign new_n10107_ = ~new_n1809_;
  assign new_n10108_ = ~new_n1812_;
  assign new_n10109_ = ~new_n1809_ | ~pi135;
  assign new_n10110_ = ~pi136;
  assign new_n10111_ = ~pi133;
  assign new_n10112_ = ~new_n1803_;
  assign new_n10113_ = ~new_n1806_;
  assign new_n10114_ = ~pi131;
  assign new_n10115_ = ~new_n1797_;
  assign new_n10116_ = ~pi129;
  assign new_n10117_ = ~new_n1788_;
  assign new_n10118_ = ~new_n1788_ | ~pi129;
  assign new_n10119_ = ~pi132;
  assign new_n10120_ = ~new_n1800_;
  assign new_n10121_ = ~new_n1803_ | ~pi133;
  assign new_n10122_ = ~pi134;
  assign new_n10123_ = ~pi137;
  assign new_n10124_ = ~new_n1815_;
  assign new_n10125_ = ~new_n1818_;
  assign new_n10126_ = ~pi138;
  assign new_n10127_ = ~new_n10138_ | ~new_n10210_;
  assign new_n10128_ = ~new_n10198_ | ~new_n10199_ | ~new_n10197_;
  assign new_n10129_ = ~new_n10187_ | ~new_n10188_;
  assign new_n10130_ = ~pi130 | ~new_n1794_;
  assign new_n10131_ = ~new_n10224_ | ~new_n10225_ | ~new_n10223_;
  assign new_n10132_ = ~new_n10221_ | ~new_n10220_;
  assign new_n10133_ = ~pi145;
  assign new_n10134_ = ~new_n1839_;
  assign new_n10135_ = ~new_n1842_;
  assign new_n10136_ = ~new_n1839_ | ~pi145;
  assign new_n10137_ = ~pi146;
  assign new_n10138_ = ~new_n1815_ | ~pi137;
  assign new_n10139_ = ~pi139;
  assign new_n10140_ = ~new_n1821_;
  assign new_n10141_ = ~pi141;
  assign new_n10142_ = ~new_n1827_;
  assign new_n10143_ = ~pi140;
  assign new_n10144_ = ~new_n1824_;
  assign new_n10145_ = ~new_n1824_ | ~pi140;
  assign new_n10146_ = ~pi142;
  assign new_n10147_ = ~new_n1830_;
  assign new_n10148_ = ~pi143;
  assign new_n10149_ = ~new_n1833_;
  assign new_n10150_ = ~pi144;
  assign new_n10151_ = ~new_n1836_;
  assign new_n10152_ = ~pi147;
  assign new_n10153_ = ~new_n1845_;
  assign new_n10154_ = ~new_n10276_ | ~new_n10275_ | ~new_n10274_;
  assign new_n10155_ = ~new_n10268_ | ~new_n10267_;
  assign new_n10156_ = ~new_n10145_ | ~new_n10293_;
  assign new_n10157_ = ~new_n10348_ | ~new_n10347_;
  assign new_n10158_ = ~new_n10397_ | ~new_n10396_;
  assign new_n10159_ = ~new_n10320_ | ~new_n10319_;
  assign new_n10160_ = ~new_n10325_ | ~new_n10324_;
  assign new_n10161_ = ~new_n10332_ | ~new_n10331_;
  assign new_n10162_ = ~new_n10339_ | ~new_n10338_;
  assign new_n10163_ = ~new_n10344_ | ~new_n10343_;
  assign new_n10164_ = ~new_n10360_ | ~new_n10359_;
  assign new_n10165_ = ~new_n10367_ | ~new_n10366_;
  assign new_n10166_ = ~new_n10374_ | ~new_n10373_;
  assign new_n10167_ = ~new_n10381_ | ~new_n10380_;
  assign new_n10168_ = ~new_n10388_ | ~new_n10387_;
  assign new_n10169_ = ~new_n10393_ | ~new_n10392_;
  assign new_n10170_ = ~new_n10207_ | ~new_n10206_ | ~new_n10205_;
  assign new_n10171_ = ~new_n10222_ | ~new_n10234_;
  assign new_n10172_ = ~new_n10130_ | ~new_n10241_;
  assign new_n10173_ = ~new_n1782_;
  assign new_n10174_ = ~pi148;
  assign new_n10175_ = ~new_n10264_ | ~new_n10263_;
  assign new_n10176_ = ~new_n10260_ | ~new_n10259_;
  assign new_n10177_ = ~new_n10250_ | ~new_n10249_;
  assign new_n10178_ = ~new_n10121_;
  assign new_n10179_ = ~pi138 | ~new_n1818_;
  assign new_n10180_ = ~new_n1827_ | ~pi141;
  assign new_n10181_ = ~new_n10145_;
  assign new_n10182_ = ~new_n10138_;
  assign new_n10183_ = new_n1806_ | pi134;
  assign new_n10184_ = new_n1803_ | pi133;
  assign new_n10185_ = pi132 | new_n1800_;
  assign new_n10186_ = pi131 | new_n1797_;
  assign new_n10187_ = ~new_n10118_;
  assign new_n10188_ = pi130 | new_n1794_;
  assign new_n10189_ = ~new_n10129_;
  assign new_n10190_ = ~new_n10130_;
  assign new_n10191_ = ~new_n10129_ | ~new_n10130_;
  assign new_n10192_ = ~new_n10185_ | ~pi131 | ~new_n1797_;
  assign new_n10193_ = ~new_n10094_ | ~new_n10191_;
  assign new_n10194_ = ~new_n1800_ | ~pi132;
  assign new_n10195_ = ~new_n10193_ | ~new_n10194_ | ~new_n10192_;
  assign new_n10196_ = ~new_n10122_ | ~new_n10121_;
  assign new_n10197_ = ~new_n1806_ | ~new_n10196_;
  assign new_n10198_ = ~new_n10093_ | ~new_n10195_;
  assign new_n10199_ = ~pi134 | ~new_n10178_;
  assign new_n10200_ = ~new_n10128_;
  assign new_n10201_ = new_n1812_ | pi136;
  assign new_n10202_ = new_n1809_ | pi135;
  assign new_n10203_ = ~new_n10109_;
  assign new_n10204_ = ~new_n10110_ | ~new_n10109_;
  assign new_n10205_ = ~new_n1812_ | ~new_n10204_;
  assign new_n10206_ = ~pi136 | ~new_n10203_;
  assign new_n10207_ = ~new_n10095_ | ~new_n10128_;
  assign new_n10208_ = ~new_n10170_;
  assign new_n10209_ = pi137 | new_n1815_;
  assign new_n10210_ = ~new_n10209_ | ~new_n10170_;
  assign new_n10211_ = ~new_n10127_;
  assign new_n10212_ = new_n1818_ | pi138;
  assign new_n10213_ = pi135 | new_n1809_;
  assign new_n10214_ = ~new_n10213_ | ~new_n10128_;
  assign new_n10215_ = ~new_n10214_ | ~new_n10109_ | ~new_n10327_ | ~new_n10326_;
  assign new_n10216_ = ~new_n10200_ | ~new_n10109_;
  assign new_n10217_ = ~pi136 | ~new_n1812_;
  assign new_n10218_ = ~new_n10216_ | ~new_n10217_ | ~new_n10095_;
  assign new_n10219_ = new_n1809_ | pi135;
  assign new_n10220_ = ~new_n10190_ | ~new_n10186_;
  assign new_n10221_ = ~new_n1797_ | ~pi131;
  assign new_n10222_ = ~new_n10132_;
  assign new_n10223_ = ~new_n10189_ | ~new_n10094_;
  assign new_n10224_ = ~new_n10132_ | ~new_n10185_;
  assign new_n10225_ = ~new_n1800_ | ~pi132;
  assign new_n10226_ = ~new_n10131_;
  assign new_n10227_ = pi133 | new_n1803_;
  assign new_n10228_ = ~new_n10227_ | ~new_n10131_;
  assign new_n10229_ = ~new_n10228_ | ~new_n10121_ | ~new_n10334_ | ~new_n10333_;
  assign new_n10230_ = ~new_n10226_ | ~new_n10121_;
  assign new_n10231_ = ~pi134 | ~new_n1806_;
  assign new_n10232_ = ~new_n10230_ | ~new_n10231_ | ~new_n10093_;
  assign new_n10233_ = new_n1803_ | pi133;
  assign new_n10234_ = ~new_n10189_ | ~new_n10186_;
  assign new_n10235_ = ~new_n10171_;
  assign new_n10236_ = ~new_n1800_ | ~pi132;
  assign new_n10237_ = ~new_n10129_ | ~new_n10130_ | ~new_n10346_ | ~new_n10345_;
  assign new_n10238_ = ~new_n10130_ | ~new_n10129_;
  assign new_n10239_ = ~new_n1797_ | ~pi131;
  assign new_n10240_ = ~new_n10238_ | ~new_n10239_ | ~new_n10186_;
  assign new_n10241_ = pi130 | new_n1794_;
  assign new_n10242_ = ~new_n10172_;
  assign new_n10243_ = new_n1818_ | pi138;
  assign new_n10244_ = new_n1821_ | pi139;
  assign new_n10245_ = ~new_n10182_ | ~new_n10096_;
  assign new_n10246_ = ~new_n1821_ | ~pi139;
  assign new_n10247_ = ~new_n10245_ | ~new_n10246_ | ~new_n10179_;
  assign new_n10248_ = pi139 | new_n1821_;
  assign new_n10249_ = ~new_n10170_ | ~new_n10209_ | ~new_n10096_;
  assign new_n10250_ = ~new_n10248_ | ~new_n10247_;
  assign new_n10251_ = ~new_n10177_;
  assign new_n10252_ = new_n1830_ | pi142;
  assign new_n10253_ = new_n1827_ | pi141;
  assign new_n10254_ = ~new_n10181_ | ~new_n10097_;
  assign new_n10255_ = ~new_n1830_ | ~pi142;
  assign new_n10256_ = ~new_n10254_ | ~new_n10255_ | ~new_n10180_;
  assign new_n10257_ = pi140 | new_n1824_;
  assign new_n10258_ = pi142 | new_n1830_;
  assign new_n10259_ = ~new_n10177_ | ~new_n10257_ | ~new_n10097_;
  assign new_n10260_ = ~new_n10258_ | ~new_n10256_;
  assign new_n10261_ = ~new_n10176_;
  assign new_n10262_ = pi143 | new_n1833_;
  assign new_n10263_ = ~new_n10262_ | ~new_n10176_;
  assign new_n10264_ = ~new_n1833_ | ~pi143;
  assign new_n10265_ = ~new_n10175_;
  assign new_n10266_ = pi144 | new_n1836_;
  assign new_n10267_ = ~new_n10266_ | ~new_n10175_;
  assign new_n10268_ = ~new_n1836_ | ~pi144;
  assign new_n10269_ = ~new_n10155_;
  assign new_n10270_ = new_n1842_ | pi146;
  assign new_n10271_ = new_n1839_ | pi145;
  assign new_n10272_ = ~new_n10136_;
  assign new_n10273_ = ~new_n10137_ | ~new_n10136_;
  assign new_n10274_ = ~new_n1842_ | ~new_n10273_;
  assign new_n10275_ = ~pi146 | ~new_n10272_;
  assign new_n10276_ = ~new_n10098_ | ~new_n10155_;
  assign new_n10277_ = ~new_n10154_;
  assign new_n10278_ = pi147 | new_n1845_;
  assign new_n10279_ = ~new_n10278_ | ~new_n10154_;
  assign new_n10280_ = ~new_n1845_ | ~pi147;
  assign new_n10281_ = ~new_n10279_ | ~new_n10280_ | ~new_n10350_ | ~new_n10349_;
  assign new_n10282_ = ~new_n1845_ | ~pi147;
  assign new_n10283_ = ~new_n10277_ | ~new_n10282_;
  assign new_n10284_ = new_n1845_ | pi147;
  assign new_n10285_ = ~new_n10283_ | ~new_n10284_ | ~new_n10353_;
  assign new_n10286_ = pi145 | new_n1839_;
  assign new_n10287_ = ~new_n10286_ | ~new_n10155_;
  assign new_n10288_ = ~new_n10287_ | ~new_n10136_ | ~new_n10362_ | ~new_n10361_;
  assign new_n10289_ = ~new_n10269_ | ~new_n10136_;
  assign new_n10290_ = ~pi146 | ~new_n1842_;
  assign new_n10291_ = ~new_n10289_ | ~new_n10290_ | ~new_n10098_;
  assign new_n10292_ = new_n1839_ | pi145;
  assign new_n10293_ = ~new_n10257_ | ~new_n10177_;
  assign new_n10294_ = ~new_n10156_;
  assign new_n10295_ = pi141 | new_n1827_;
  assign new_n10296_ = ~new_n10295_ | ~new_n10156_;
  assign new_n10297_ = ~new_n10296_ | ~new_n10180_ | ~new_n10383_ | ~new_n10382_;
  assign new_n10298_ = ~new_n10294_ | ~new_n10180_;
  assign new_n10299_ = ~new_n1830_ | ~pi142;
  assign new_n10300_ = ~new_n10298_ | ~new_n10299_ | ~new_n10097_;
  assign new_n10301_ = new_n1827_ | pi141;
  assign new_n10302_ = pi138 | new_n1818_;
  assign new_n10303_ = ~new_n10302_ | ~new_n10127_;
  assign new_n10304_ = ~new_n10303_ | ~new_n10179_ | ~new_n10395_ | ~new_n10394_;
  assign new_n10305_ = ~new_n10211_ | ~new_n10179_;
  assign new_n10306_ = ~new_n1821_ | ~pi139;
  assign new_n10307_ = ~new_n10305_ | ~new_n10306_ | ~new_n10096_;
  assign new_n10308_ = ~new_n10212_ | ~new_n10179_;
  assign new_n10309_ = ~new_n10209_ | ~new_n10138_;
  assign new_n10310_ = ~new_n10219_ | ~new_n10109_;
  assign new_n10311_ = ~new_n10233_ | ~new_n10121_;
  assign new_n10312_ = ~new_n10236_ | ~new_n10185_;
  assign new_n10313_ = ~new_n10292_ | ~new_n10136_;
  assign new_n10314_ = ~new_n10301_ | ~new_n10180_;
  assign new_n10315_ = ~new_n10257_ | ~new_n10145_;
  assign new_n10316_ = ~new_n1818_ | ~new_n10126_;
  assign new_n10317_ = ~pi138 | ~new_n10125_;
  assign new_n10318_ = ~new_n10317_ | ~new_n10316_;
  assign new_n10319_ = ~new_n10308_ | ~new_n10127_;
  assign new_n10320_ = ~new_n10318_ | ~new_n10211_;
  assign new_n10321_ = ~new_n1815_ | ~new_n10123_;
  assign new_n10322_ = ~pi137 | ~new_n10124_;
  assign new_n10323_ = ~new_n10322_ | ~new_n10321_;
  assign new_n10324_ = ~new_n10309_ | ~new_n10170_;
  assign new_n10325_ = ~new_n10208_ | ~new_n10323_;
  assign new_n10326_ = ~new_n1812_ | ~new_n10110_;
  assign new_n10327_ = ~pi136 | ~new_n10108_;
  assign new_n10328_ = ~new_n1809_ | ~new_n10106_;
  assign new_n10329_ = ~pi135 | ~new_n10107_;
  assign new_n10330_ = ~new_n10329_ | ~new_n10328_;
  assign new_n10331_ = ~new_n10310_ | ~new_n10128_;
  assign new_n10332_ = ~new_n10330_ | ~new_n10200_;
  assign new_n10333_ = ~new_n1806_ | ~new_n10122_;
  assign new_n10334_ = ~pi134 | ~new_n10113_;
  assign new_n10335_ = ~new_n1803_ | ~new_n10111_;
  assign new_n10336_ = ~pi133 | ~new_n10112_;
  assign new_n10337_ = ~new_n10336_ | ~new_n10335_;
  assign new_n10338_ = ~new_n10311_ | ~new_n10131_;
  assign new_n10339_ = ~new_n10337_ | ~new_n10226_;
  assign new_n10340_ = ~new_n1800_ | ~new_n10119_;
  assign new_n10341_ = ~pi132 | ~new_n10120_;
  assign new_n10342_ = ~new_n10341_ | ~new_n10340_;
  assign new_n10343_ = ~new_n10312_ | ~new_n10171_;
  assign new_n10344_ = ~new_n10235_ | ~new_n10342_;
  assign new_n10345_ = ~new_n1797_ | ~new_n10114_;
  assign new_n10346_ = ~pi131 | ~new_n10115_;
  assign new_n10347_ = ~new_n10187_ | ~new_n10172_;
  assign new_n10348_ = ~new_n10242_ | ~new_n10118_;
  assign new_n10349_ = ~new_n1782_ | ~new_n10174_;
  assign new_n10350_ = ~pi148 | ~new_n10173_;
  assign new_n10351_ = ~new_n1782_ | ~new_n10174_;
  assign new_n10352_ = ~pi148 | ~new_n10173_;
  assign new_n10353_ = ~new_n10352_ | ~new_n10351_;
  assign new_n10354_ = ~new_n1845_ | ~new_n10152_;
  assign new_n10355_ = ~pi147 | ~new_n10153_;
  assign new_n10356_ = ~new_n1845_ | ~new_n10152_;
  assign new_n10357_ = ~pi147 | ~new_n10153_;
  assign new_n10358_ = ~new_n10357_ | ~new_n10356_;
  assign new_n10359_ = ~new_n10154_ | ~new_n10355_ | ~new_n10354_;
  assign new_n10360_ = ~new_n10358_ | ~new_n10277_;
  assign new_n10361_ = ~new_n1842_ | ~new_n10137_;
  assign new_n10362_ = ~pi146 | ~new_n10135_;
  assign new_n10363_ = ~new_n1839_ | ~new_n10133_;
  assign new_n10364_ = ~pi145 | ~new_n10134_;
  assign new_n10365_ = ~new_n10364_ | ~new_n10363_;
  assign new_n10366_ = ~new_n10313_ | ~new_n10155_;
  assign new_n10367_ = ~new_n10365_ | ~new_n10269_;
  assign new_n10368_ = ~new_n1836_ | ~new_n10150_;
  assign new_n10369_ = ~pi144 | ~new_n10151_;
  assign new_n10370_ = ~new_n1836_ | ~new_n10150_;
  assign new_n10371_ = ~pi144 | ~new_n10151_;
  assign new_n10372_ = ~new_n10371_ | ~new_n10370_;
  assign new_n10373_ = ~new_n10175_ | ~new_n10369_ | ~new_n10368_;
  assign new_n10374_ = ~new_n10265_ | ~new_n10372_;
  assign new_n10375_ = ~new_n1833_ | ~new_n10148_;
  assign new_n10376_ = ~pi143 | ~new_n10149_;
  assign new_n10377_ = ~new_n1833_ | ~new_n10148_;
  assign new_n10378_ = ~pi143 | ~new_n10149_;
  assign new_n10379_ = ~new_n10378_ | ~new_n10377_;
  assign new_n10380_ = ~new_n10176_ | ~new_n10376_ | ~new_n10375_;
  assign new_n10381_ = ~new_n10261_ | ~new_n10379_;
  assign new_n10382_ = ~new_n1830_ | ~new_n10146_;
  assign new_n10383_ = ~pi142 | ~new_n10147_;
  assign new_n10384_ = ~new_n1827_ | ~new_n10141_;
  assign new_n10385_ = ~pi141 | ~new_n10142_;
  assign new_n10386_ = ~new_n10385_ | ~new_n10384_;
  assign new_n10387_ = ~new_n10314_ | ~new_n10156_;
  assign new_n10388_ = ~new_n10386_ | ~new_n10294_;
  assign new_n10389_ = ~new_n1824_ | ~new_n10143_;
  assign new_n10390_ = ~pi140 | ~new_n10144_;
  assign new_n10391_ = ~new_n10390_ | ~new_n10389_;
  assign new_n10392_ = ~new_n10315_ | ~new_n10177_;
  assign new_n10393_ = ~new_n10251_ | ~new_n10391_;
  assign new_n10394_ = ~new_n1821_ | ~new_n10139_;
  assign new_n10395_ = ~pi139 | ~new_n10140_;
  assign new_n10396_ = ~new_n1788_ | ~new_n10116_;
  assign new_n10397_ = ~pi129 | ~new_n10117_;
  assign new_n10398_ = new_n10576_ & new_n10593_;
  assign new_n10399_ = new_n10595_ & new_n10594_;
  assign new_n10400_ = new_n10571_ & new_n10632_;
  assign new_n10401_ = new_n10634_ & new_n10633_;
  assign new_n10402_ = new_n10651_ & new_n10650_;
  assign new_n10403_ = new_n10677_ & new_n10676_;
  assign new_n10404_ = new_n10775_ & new_n10774_;
  assign new_n10405_ = ~new_n10732_ | ~new_n10735_;
  assign new_n10406_ = ~new_n10721_ | ~new_n10724_;
  assign new_n10407_ = ~new_n10710_ | ~new_n10713_;
  assign new_n10408_ = ~new_n10702_ | ~new_n10704_;
  assign new_n10409_ = ~new_n10740_ | ~new_n10548_ | ~new_n10567_;
  assign new_n10410_ = ~new_n10628_ | ~new_n10630_;
  assign new_n10411_ = ~new_n10620_ | ~new_n10623_;
  assign new_n10412_ = ~new_n10612_ | ~new_n10614_;
  assign new_n10413_ = ~new_n10417_ | ~new_n10738_;
  assign new_n10414_ = ~new_n1813_;
  assign new_n10415_ = ~new_n1798_;
  assign new_n10416_ = ~new_n1790_;
  assign new_n10417_ = ~new_n1790_ | ~new_n10485_;
  assign new_n10418_ = ~new_n1415_;
  assign new_n10419_ = ~new_n1801_;
  assign new_n10420_ = ~new_n1405_;
  assign new_n10421_ = ~new_n1405_ | ~new_n10415_;
  assign new_n10422_ = ~new_n1401_;
  assign new_n10423_ = ~new_n1810_;
  assign new_n10424_ = ~new_n1807_;
  assign new_n10425_ = ~new_n1804_;
  assign new_n10426_ = ~new_n1408_;
  assign new_n10427_ = ~new_n1404_;
  assign new_n10428_ = ~new_n1397_;
  assign new_n10429_ = ~new_n1397_ | ~new_n10425_;
  assign new_n10430_ = ~new_n1816_;
  assign new_n10431_ = ~new_n1407_;
  assign new_n10432_ = ~new_n1407_ | ~new_n10414_;
  assign new_n10433_ = ~new_n1421_;
  assign new_n10434_ = ~new_n1819_;
  assign new_n10435_ = ~new_n1420_;
  assign new_n10436_ = ~new_n10601_ | ~new_n10600_;
  assign new_n10437_ = ~new_n10429_ | ~new_n10616_;
  assign new_n10438_ = ~new_n10585_ | ~new_n10584_;
  assign new_n10439_ = ~new_n2348_;
  assign new_n10440_ = ~new_n2352_;
  assign new_n10441_ = ~new_n1837_;
  assign new_n10442_ = ~new_n1825_;
  assign new_n10443_ = ~new_n1822_;
  assign new_n10444_ = ~new_n1400_;
  assign new_n10445_ = ~new_n1399_;
  assign new_n10446_ = ~new_n1420_ | ~new_n10434_;
  assign new_n10447_ = ~new_n1828_;
  assign new_n10448_ = ~new_n1409_;
  assign new_n10449_ = ~new_n1831_;
  assign new_n10450_ = ~new_n1417_;
  assign new_n10451_ = ~new_n1840_;
  assign new_n10452_ = ~new_n1834_;
  assign new_n10453_ = ~new_n1410_;
  assign new_n10454_ = ~new_n1411_;
  assign new_n10455_ = ~new_n1416_;
  assign new_n10456_ = ~new_n1416_ | ~new_n10452_;
  assign new_n10457_ = ~new_n1843_;
  assign new_n10458_ = ~new_n1406_;
  assign new_n10459_ = ~new_n10661_ | ~new_n10660_;
  assign new_n10460_ = ~new_n1419_;
  assign new_n10461_ = ~new_n1848_;
  assign new_n10462_ = ~new_n1418_;
  assign new_n10463_ = ~new_n2354_;
  assign new_n10464_ = ~new_n1413_;
  assign new_n10465_ = ~new_n2351_;
  assign new_n10466_ = ~new_n2353_;
  assign new_n10467_ = ~new_n1403_;
  assign new_n10468_ = ~new_n1398_;
  assign new_n10469_ = ~new_n1412_;
  assign new_n10470_ = ~new_n1412_ | ~new_n10466_;
  assign new_n10471_ = ~new_n2350_;
  assign new_n10472_ = ~new_n1402_;
  assign new_n10473_ = ~new_n2349_;
  assign new_n10474_ = ~new_n1395_;
  assign new_n10475_ = ~new_n2347_;
  assign new_n10476_ = ~new_n1394_;
  assign new_n10477_ = ~new_n1394_ | ~new_n10439_;
  assign new_n10478_ = ~new_n1390_;
  assign new_n10479_ = ~new_n2346_;
  assign new_n10480_ = ~new_n1391_;
  assign new_n10481_ = ~new_n10691_ | ~new_n10690_;
  assign new_n10482_ = ~new_n10470_ | ~new_n10706_;
  assign new_n10483_ = ~new_n10456_ | ~new_n10717_;
  assign new_n10484_ = ~new_n10446_ | ~new_n10728_;
  assign new_n10485_ = ~new_n1414_;
  assign new_n10486_ = ~new_n10785_ | ~new_n10784_;
  assign new_n10487_ = ~new_n10799_ | ~new_n10798_;
  assign new_n10488_ = ~new_n10804_ | ~new_n10803_;
  assign new_n10489_ = ~new_n10820_ | ~new_n10819_;
  assign new_n10490_ = ~new_n10825_ | ~new_n10824_;
  assign new_n10491_ = ~new_n10830_ | ~new_n10829_;
  assign new_n10492_ = ~new_n10835_ | ~new_n10834_;
  assign new_n10493_ = ~new_n10840_ | ~new_n10839_;
  assign new_n10494_ = ~new_n10856_ | ~new_n10855_;
  assign new_n10495_ = ~new_n10861_ | ~new_n10860_;
  assign new_n10496_ = ~new_n10744_ | ~new_n10743_;
  assign new_n10497_ = ~new_n10753_ | ~new_n10752_;
  assign new_n10498_ = ~new_n10760_ | ~new_n10759_;
  assign new_n10499_ = ~new_n10764_ | ~new_n10763_;
  assign new_n10500_ = ~new_n10773_ | ~new_n10772_;
  assign new_n10501_ = ~new_n10794_ | ~new_n10793_;
  assign new_n10502_ = ~new_n10811_ | ~new_n10810_;
  assign new_n10503_ = ~new_n10815_ | ~new_n10814_;
  assign new_n10504_ = ~new_n10847_ | ~new_n10846_;
  assign new_n10505_ = ~new_n10851_ | ~new_n10850_;
  assign new_n10506_ = ~new_n10868_ | ~new_n10867_;
  assign new_n10507_ = new_n10587_ & new_n10575_;
  assign new_n10508_ = new_n10590_ & new_n10591_;
  assign new_n10509_ = new_n10603_ & new_n10577_;
  assign new_n10510_ = new_n10606_ & new_n10607_;
  assign new_n10511_ = new_n10432_ & new_n10746_ & new_n10745_;
  assign new_n10512_ = new_n10749_ & new_n10577_;
  assign new_n10513_ = new_n10622_ & new_n10399_;
  assign new_n10514_ = new_n10756_ & new_n10576_;
  assign new_n10515_ = new_n10421_ & new_n10766_ & new_n10765_;
  assign new_n10516_ = new_n10769_ & new_n10575_;
  assign new_n10517_ = new_n10609_ & new_n10400_;
  assign new_n10518_ = new_n10654_ & new_n10572_;
  assign new_n10519_ = new_n10680_ & new_n10573_;
  assign new_n10520_ = new_n10696_ & new_n10697_;
  assign new_n10521_ = new_n10699_ & new_n10778_;
  assign new_n10522_ = new_n10700_ & new_n10697_ & new_n10696_;
  assign new_n10523_ = ~new_n10782_ | ~new_n10781_;
  assign new_n10524_ = new_n10477_ & new_n10787_ & new_n10786_;
  assign new_n10525_ = new_n10790_ & new_n10574_;
  assign new_n10526_ = ~new_n10796_ | ~new_n10795_;
  assign new_n10527_ = ~new_n10801_ | ~new_n10800_;
  assign new_n10528_ = new_n10807_ & new_n10573_;
  assign new_n10529_ = ~new_n10817_ | ~new_n10816_;
  assign new_n10530_ = ~new_n10822_ | ~new_n10821_;
  assign new_n10531_ = ~new_n10827_ | ~new_n10826_;
  assign new_n10532_ = ~new_n10832_ | ~new_n10831_;
  assign new_n10533_ = ~new_n10837_ | ~new_n10836_;
  assign new_n10534_ = new_n10843_ & new_n10572_;
  assign new_n10535_ = ~new_n10853_ | ~new_n10852_;
  assign new_n10536_ = ~new_n10858_ | ~new_n10857_;
  assign new_n10537_ = new_n10734_ & new_n10401_;
  assign new_n10538_ = new_n10864_ & new_n10571_;
  assign new_n10539_ = new_n10742_ & new_n10741_;
  assign new_n10540_ = ~new_n10510_ | ~new_n10604_;
  assign new_n10541_ = new_n10751_ & new_n10750_;
  assign new_n10542_ = new_n10758_ & new_n10757_;
  assign new_n10543_ = new_n10762_ & new_n10761_;
  assign new_n10544_ = ~new_n10508_ | ~new_n10588_;
  assign new_n10545_ = new_n10771_ & new_n10770_;
  assign new_n10546_ = ~new_n2357_;
  assign new_n10547_ = ~new_n1392_;
  assign new_n10548_ = new_n10780_ & new_n10779_;
  assign new_n10549_ = ~new_n10520_ | ~new_n10694_;
  assign new_n10550_ = new_n10792_ & new_n10791_;
  assign new_n10551_ = ~new_n10687_ | ~new_n10686_;
  assign new_n10552_ = ~new_n10683_ | ~new_n10682_;
  assign new_n10553_ = new_n10809_ & new_n10808_;
  assign new_n10554_ = new_n10813_ & new_n10812_;
  assign new_n10555_ = ~new_n10673_ | ~new_n10672_;
  assign new_n10556_ = ~new_n10669_ | ~new_n10668_;
  assign new_n10557_ = ~new_n1795_;
  assign new_n10558_ = ~new_n10665_ | ~new_n10664_;
  assign new_n10559_ = ~new_n1846_;
  assign new_n10560_ = ~new_n10657_ | ~new_n10656_;
  assign new_n10561_ = new_n10845_ & new_n10844_;
  assign new_n10562_ = new_n10849_ & new_n10848_;
  assign new_n10563_ = ~new_n10647_ | ~new_n10646_;
  assign new_n10564_ = ~new_n10643_ | ~new_n10642_;
  assign new_n10565_ = ~new_n10639_ | ~new_n10638_;
  assign new_n10566_ = new_n10866_ & new_n10865_;
  assign new_n10567_ = ~new_n10521_ | ~new_n10549_;
  assign new_n10568_ = ~new_n10477_;
  assign new_n10569_ = ~new_n10421_;
  assign new_n10570_ = ~new_n10432_;
  assign new_n10571_ = ~new_n1822_ | ~new_n10445_;
  assign new_n10572_ = ~new_n1837_ | ~new_n10454_;
  assign new_n10573_ = ~new_n2352_ | ~new_n10468_;
  assign new_n10574_ = ~new_n2348_ | ~new_n10476_;
  assign new_n10575_ = ~new_n1798_ | ~new_n10420_;
  assign new_n10576_ = ~new_n1807_ | ~new_n10427_;
  assign new_n10577_ = ~new_n1813_ | ~new_n10431_;
  assign new_n10578_ = ~new_n10456_;
  assign new_n10579_ = ~new_n10470_;
  assign new_n10580_ = ~new_n10429_;
  assign new_n10581_ = ~new_n10446_;
  assign new_n10582_ = ~new_n10417_;
  assign new_n10583_ = ~new_n10582_ | ~new_n10418_;
  assign new_n10584_ = ~new_n10583_ | ~new_n10557_;
  assign new_n10585_ = ~new_n1415_ | ~new_n10417_;
  assign new_n10586_ = ~new_n10438_;
  assign new_n10587_ = ~new_n1801_ | ~new_n10422_;
  assign new_n10588_ = ~new_n10507_ | ~new_n10438_;
  assign new_n10589_ = ~new_n10422_ | ~new_n10421_;
  assign new_n10590_ = ~new_n10589_ | ~new_n10419_;
  assign new_n10591_ = ~new_n1401_ | ~new_n10569_;
  assign new_n10592_ = ~new_n10544_;
  assign new_n10593_ = ~new_n1810_ | ~new_n10426_;
  assign new_n10594_ = ~new_n1408_ | ~new_n10423_;
  assign new_n10595_ = ~new_n1404_ | ~new_n10424_;
  assign new_n10596_ = ~new_n10580_ | ~new_n10398_;
  assign new_n10597_ = ~new_n10399_ | ~new_n10596_;
  assign new_n10598_ = ~new_n1804_ | ~new_n10428_;
  assign new_n10599_ = ~new_n1810_ | ~new_n10426_;
  assign new_n10600_ = ~new_n10398_ | ~new_n10598_ | ~new_n10544_;
  assign new_n10601_ = ~new_n10599_ | ~new_n10597_;
  assign new_n10602_ = ~new_n10436_;
  assign new_n10603_ = ~new_n1816_ | ~new_n10433_;
  assign new_n10604_ = ~new_n10509_ | ~new_n10436_;
  assign new_n10605_ = ~new_n10433_ | ~new_n10432_;
  assign new_n10606_ = ~new_n10605_ | ~new_n10430_;
  assign new_n10607_ = ~new_n1421_ | ~new_n10570_;
  assign new_n10608_ = ~new_n10540_;
  assign new_n10609_ = ~new_n1819_ | ~new_n10435_;
  assign new_n10610_ = ~new_n10609_ | ~new_n10446_;
  assign new_n10611_ = ~new_n10602_ | ~new_n10432_;
  assign new_n10612_ = ~new_n10512_ | ~new_n10611_;
  assign new_n10613_ = ~new_n10436_ | ~new_n10577_;
  assign new_n10614_ = ~new_n10511_ | ~new_n10613_;
  assign new_n10615_ = ~new_n10432_ | ~new_n10577_;
  assign new_n10616_ = ~new_n10598_ | ~new_n10544_;
  assign new_n10617_ = ~new_n10437_;
  assign new_n10618_ = ~new_n1404_ | ~new_n10424_;
  assign new_n10619_ = ~new_n10617_ | ~new_n10618_;
  assign new_n10620_ = ~new_n10514_ | ~new_n10619_;
  assign new_n10621_ = ~new_n10437_ | ~new_n10576_;
  assign new_n10622_ = ~new_n1810_ | ~new_n10426_;
  assign new_n10623_ = ~new_n10513_ | ~new_n10621_;
  assign new_n10624_ = ~new_n1404_ | ~new_n10424_;
  assign new_n10625_ = ~new_n10576_ | ~new_n10624_;
  assign new_n10626_ = ~new_n10598_ | ~new_n10429_;
  assign new_n10627_ = ~new_n10586_ | ~new_n10421_;
  assign new_n10628_ = ~new_n10516_ | ~new_n10627_;
  assign new_n10629_ = ~new_n10438_ | ~new_n10575_;
  assign new_n10630_ = ~new_n10515_ | ~new_n10629_;
  assign new_n10631_ = ~new_n10421_ | ~new_n10575_;
  assign new_n10632_ = ~new_n1825_ | ~new_n10444_;
  assign new_n10633_ = ~new_n1400_ | ~new_n10442_;
  assign new_n10634_ = ~new_n1399_ | ~new_n10443_;
  assign new_n10635_ = ~new_n10581_ | ~new_n10400_;
  assign new_n10636_ = ~new_n10401_ | ~new_n10635_;
  assign new_n10637_ = ~new_n1825_ | ~new_n10444_;
  assign new_n10638_ = ~new_n10517_ | ~new_n10540_;
  assign new_n10639_ = ~new_n10637_ | ~new_n10636_;
  assign new_n10640_ = ~new_n10565_;
  assign new_n10641_ = ~new_n1828_ | ~new_n10448_;
  assign new_n10642_ = ~new_n10641_ | ~new_n10565_;
  assign new_n10643_ = ~new_n1409_ | ~new_n10447_;
  assign new_n10644_ = ~new_n10564_;
  assign new_n10645_ = ~new_n1831_ | ~new_n10450_;
  assign new_n10646_ = ~new_n10645_ | ~new_n10564_;
  assign new_n10647_ = ~new_n1417_ | ~new_n10449_;
  assign new_n10648_ = ~new_n10563_;
  assign new_n10649_ = ~new_n1840_ | ~new_n10453_;
  assign new_n10650_ = ~new_n1410_ | ~new_n10451_;
  assign new_n10651_ = ~new_n1411_ | ~new_n10441_;
  assign new_n10652_ = ~new_n10578_ | ~new_n10572_;
  assign new_n10653_ = ~new_n10402_ | ~new_n10652_;
  assign new_n10654_ = ~new_n1834_ | ~new_n10455_;
  assign new_n10655_ = ~new_n1840_ | ~new_n10453_;
  assign new_n10656_ = ~new_n10649_ | ~new_n10563_ | ~new_n10518_;
  assign new_n10657_ = ~new_n10655_ | ~new_n10653_;
  assign new_n10658_ = ~new_n10560_;
  assign new_n10659_ = ~new_n1843_ | ~new_n10458_;
  assign new_n10660_ = ~new_n10659_ | ~new_n10560_;
  assign new_n10661_ = ~new_n1406_ | ~new_n10457_;
  assign new_n10662_ = ~new_n10459_;
  assign new_n10663_ = ~new_n10662_ | ~new_n10460_;
  assign new_n10664_ = ~new_n10663_ | ~new_n10559_;
  assign new_n10665_ = ~new_n1419_ | ~new_n10459_;
  assign new_n10666_ = ~new_n10558_;
  assign new_n10667_ = ~new_n1848_ | ~new_n10462_;
  assign new_n10668_ = ~new_n10667_ | ~new_n10558_;
  assign new_n10669_ = ~new_n1418_ | ~new_n10461_;
  assign new_n10670_ = ~new_n10556_;
  assign new_n10671_ = ~new_n2354_ | ~new_n10464_;
  assign new_n10672_ = ~new_n10671_ | ~new_n10556_;
  assign new_n10673_ = ~new_n1413_ | ~new_n10463_;
  assign new_n10674_ = ~new_n10555_;
  assign new_n10675_ = ~new_n2351_ | ~new_n10467_;
  assign new_n10676_ = ~new_n1403_ | ~new_n10465_;
  assign new_n10677_ = ~new_n1398_ | ~new_n10440_;
  assign new_n10678_ = ~new_n10579_ | ~new_n10573_;
  assign new_n10679_ = ~new_n10403_ | ~new_n10678_;
  assign new_n10680_ = ~new_n2353_ | ~new_n10469_;
  assign new_n10681_ = ~new_n2351_ | ~new_n10467_;
  assign new_n10682_ = ~new_n10675_ | ~new_n10555_ | ~new_n10519_;
  assign new_n10683_ = ~new_n10681_ | ~new_n10679_;
  assign new_n10684_ = ~new_n10552_;
  assign new_n10685_ = ~new_n2350_ | ~new_n10472_;
  assign new_n10686_ = ~new_n10685_ | ~new_n10552_;
  assign new_n10687_ = ~new_n1402_ | ~new_n10471_;
  assign new_n10688_ = ~new_n10551_;
  assign new_n10689_ = ~new_n2349_ | ~new_n10474_;
  assign new_n10690_ = ~new_n10689_ | ~new_n10551_;
  assign new_n10691_ = ~new_n1395_ | ~new_n10473_;
  assign new_n10692_ = ~new_n10481_;
  assign new_n10693_ = ~new_n2347_ | ~new_n10478_;
  assign new_n10694_ = ~new_n10693_ | ~new_n10481_ | ~new_n10574_;
  assign new_n10695_ = ~new_n10478_ | ~new_n10477_;
  assign new_n10696_ = ~new_n10695_ | ~new_n10475_;
  assign new_n10697_ = ~new_n1390_ | ~new_n10568_;
  assign new_n10698_ = ~new_n10549_;
  assign new_n10699_ = ~new_n2346_ | ~new_n10480_;
  assign new_n10700_ = ~new_n1391_ | ~new_n10479_;
  assign new_n10701_ = ~new_n10692_ | ~new_n10477_;
  assign new_n10702_ = ~new_n10525_ | ~new_n10701_;
  assign new_n10703_ = ~new_n10481_ | ~new_n10574_;
  assign new_n10704_ = ~new_n10524_ | ~new_n10703_;
  assign new_n10705_ = ~new_n10477_ | ~new_n10574_;
  assign new_n10706_ = ~new_n10680_ | ~new_n10555_;
  assign new_n10707_ = ~new_n10482_;
  assign new_n10708_ = ~new_n1398_ | ~new_n10440_;
  assign new_n10709_ = ~new_n10707_ | ~new_n10708_;
  assign new_n10710_ = ~new_n10528_ | ~new_n10709_;
  assign new_n10711_ = ~new_n10482_ | ~new_n10573_;
  assign new_n10712_ = ~new_n2351_ | ~new_n10467_;
  assign new_n10713_ = ~new_n10403_ | ~new_n10712_ | ~new_n10711_;
  assign new_n10714_ = ~new_n1398_ | ~new_n10440_;
  assign new_n10715_ = ~new_n10573_ | ~new_n10714_;
  assign new_n10716_ = ~new_n10680_ | ~new_n10470_;
  assign new_n10717_ = ~new_n10654_ | ~new_n10563_;
  assign new_n10718_ = ~new_n10483_;
  assign new_n10719_ = ~new_n1411_ | ~new_n10441_;
  assign new_n10720_ = ~new_n10718_ | ~new_n10719_;
  assign new_n10721_ = ~new_n10534_ | ~new_n10720_;
  assign new_n10722_ = ~new_n10483_ | ~new_n10572_;
  assign new_n10723_ = ~new_n1840_ | ~new_n10453_;
  assign new_n10724_ = ~new_n10402_ | ~new_n10723_ | ~new_n10722_;
  assign new_n10725_ = ~new_n1411_ | ~new_n10441_;
  assign new_n10726_ = ~new_n10572_ | ~new_n10725_;
  assign new_n10727_ = ~new_n10654_ | ~new_n10456_;
  assign new_n10728_ = ~new_n10609_ | ~new_n10540_;
  assign new_n10729_ = ~new_n10484_;
  assign new_n10730_ = ~new_n1399_ | ~new_n10443_;
  assign new_n10731_ = ~new_n10729_ | ~new_n10730_;
  assign new_n10732_ = ~new_n10538_ | ~new_n10731_;
  assign new_n10733_ = ~new_n10484_ | ~new_n10571_;
  assign new_n10734_ = ~new_n1825_ | ~new_n10444_;
  assign new_n10735_ = ~new_n10537_ | ~new_n10733_;
  assign new_n10736_ = ~new_n1399_ | ~new_n10443_;
  assign new_n10737_ = ~new_n10571_ | ~new_n10736_;
  assign new_n10738_ = ~new_n1414_ | ~new_n10416_;
  assign new_n10739_ = ~new_n10693_ | ~new_n10481_ | ~new_n10574_;
  assign new_n10740_ = ~new_n10522_ | ~new_n10404_ | ~new_n10739_;
  assign new_n10741_ = ~new_n1819_ | ~new_n10435_;
  assign new_n10742_ = ~new_n1420_ | ~new_n10434_;
  assign new_n10743_ = ~new_n10610_ | ~new_n10540_;
  assign new_n10744_ = ~new_n10608_ | ~new_n10539_;
  assign new_n10745_ = ~new_n1816_ | ~new_n10433_;
  assign new_n10746_ = ~new_n1421_ | ~new_n10430_;
  assign new_n10747_ = ~new_n1816_ | ~new_n10433_;
  assign new_n10748_ = ~new_n1421_ | ~new_n10430_;
  assign new_n10749_ = ~new_n10748_ | ~new_n10747_;
  assign new_n10750_ = ~new_n1813_ | ~new_n10431_;
  assign new_n10751_ = ~new_n1407_ | ~new_n10414_;
  assign new_n10752_ = ~new_n10615_ | ~new_n10436_;
  assign new_n10753_ = ~new_n10541_ | ~new_n10602_;
  assign new_n10754_ = ~new_n1810_ | ~new_n10426_;
  assign new_n10755_ = ~new_n1408_ | ~new_n10423_;
  assign new_n10756_ = ~new_n10755_ | ~new_n10754_;
  assign new_n10757_ = ~new_n1807_ | ~new_n10427_;
  assign new_n10758_ = ~new_n1404_ | ~new_n10424_;
  assign new_n10759_ = ~new_n10625_ | ~new_n10437_;
  assign new_n10760_ = ~new_n10542_ | ~new_n10617_;
  assign new_n10761_ = ~new_n1804_ | ~new_n10428_;
  assign new_n10762_ = ~new_n1397_ | ~new_n10425_;
  assign new_n10763_ = ~new_n10626_ | ~new_n10544_;
  assign new_n10764_ = ~new_n10592_ | ~new_n10543_;
  assign new_n10765_ = ~new_n1801_ | ~new_n10422_;
  assign new_n10766_ = ~new_n1401_ | ~new_n10419_;
  assign new_n10767_ = ~new_n1801_ | ~new_n10422_;
  assign new_n10768_ = ~new_n1401_ | ~new_n10419_;
  assign new_n10769_ = ~new_n10768_ | ~new_n10767_;
  assign new_n10770_ = ~new_n1798_ | ~new_n10420_;
  assign new_n10771_ = ~new_n1405_ | ~new_n10415_;
  assign new_n10772_ = ~new_n10631_ | ~new_n10438_;
  assign new_n10773_ = ~new_n10545_ | ~new_n10586_;
  assign new_n10774_ = ~new_n2357_ | ~new_n10547_;
  assign new_n10775_ = ~new_n1392_ | ~new_n10546_;
  assign new_n10776_ = ~new_n2357_ | ~new_n10547_;
  assign new_n10777_ = ~new_n1392_ | ~new_n10546_;
  assign new_n10778_ = ~new_n10777_ | ~new_n10776_;
  assign new_n10779_ = ~new_n10479_ | ~new_n1391_ | ~new_n10778_;
  assign new_n10780_ = ~new_n2346_ | ~new_n10404_ | ~new_n10480_;
  assign new_n10781_ = ~new_n2346_ | ~new_n10480_;
  assign new_n10782_ = ~new_n1391_ | ~new_n10479_;
  assign new_n10783_ = ~new_n10523_;
  assign new_n10784_ = ~new_n10698_ | ~new_n10783_;
  assign new_n10785_ = ~new_n10523_ | ~new_n10549_;
  assign new_n10786_ = ~new_n2347_ | ~new_n10478_;
  assign new_n10787_ = ~new_n1390_ | ~new_n10475_;
  assign new_n10788_ = ~new_n2347_ | ~new_n10478_;
  assign new_n10789_ = ~new_n1390_ | ~new_n10475_;
  assign new_n10790_ = ~new_n10789_ | ~new_n10788_;
  assign new_n10791_ = ~new_n2348_ | ~new_n10476_;
  assign new_n10792_ = ~new_n1394_ | ~new_n10439_;
  assign new_n10793_ = ~new_n10705_ | ~new_n10481_;
  assign new_n10794_ = ~new_n10550_ | ~new_n10692_;
  assign new_n10795_ = ~new_n2349_ | ~new_n10474_;
  assign new_n10796_ = ~new_n1395_ | ~new_n10473_;
  assign new_n10797_ = ~new_n10526_;
  assign new_n10798_ = ~new_n10688_ | ~new_n10797_;
  assign new_n10799_ = ~new_n10526_ | ~new_n10551_;
  assign new_n10800_ = ~new_n2350_ | ~new_n10472_;
  assign new_n10801_ = ~new_n1402_ | ~new_n10471_;
  assign new_n10802_ = ~new_n10527_;
  assign new_n10803_ = ~new_n10684_ | ~new_n10802_;
  assign new_n10804_ = ~new_n10527_ | ~new_n10552_;
  assign new_n10805_ = ~new_n2351_ | ~new_n10467_;
  assign new_n10806_ = ~new_n1403_ | ~new_n10465_;
  assign new_n10807_ = ~new_n10806_ | ~new_n10805_;
  assign new_n10808_ = ~new_n2352_ | ~new_n10468_;
  assign new_n10809_ = ~new_n1398_ | ~new_n10440_;
  assign new_n10810_ = ~new_n10715_ | ~new_n10482_;
  assign new_n10811_ = ~new_n10553_ | ~new_n10707_;
  assign new_n10812_ = ~new_n2353_ | ~new_n10469_;
  assign new_n10813_ = ~new_n1412_ | ~new_n10466_;
  assign new_n10814_ = ~new_n10716_ | ~new_n10555_;
  assign new_n10815_ = ~new_n10674_ | ~new_n10554_;
  assign new_n10816_ = ~new_n2354_ | ~new_n10464_;
  assign new_n10817_ = ~new_n1413_ | ~new_n10463_;
  assign new_n10818_ = ~new_n10529_;
  assign new_n10819_ = ~new_n10670_ | ~new_n10818_;
  assign new_n10820_ = ~new_n10529_ | ~new_n10556_;
  assign new_n10821_ = ~new_n1795_ | ~new_n10418_;
  assign new_n10822_ = ~new_n1415_ | ~new_n10557_;
  assign new_n10823_ = ~new_n10530_;
  assign new_n10824_ = ~new_n10823_ | ~new_n10582_;
  assign new_n10825_ = ~new_n10530_ | ~new_n10417_;
  assign new_n10826_ = ~new_n1848_ | ~new_n10462_;
  assign new_n10827_ = ~new_n1418_ | ~new_n10461_;
  assign new_n10828_ = ~new_n10531_;
  assign new_n10829_ = ~new_n10666_ | ~new_n10828_;
  assign new_n10830_ = ~new_n10531_ | ~new_n10558_;
  assign new_n10831_ = ~new_n1846_ | ~new_n10460_;
  assign new_n10832_ = ~new_n1419_ | ~new_n10559_;
  assign new_n10833_ = ~new_n10532_;
  assign new_n10834_ = ~new_n10833_ | ~new_n10662_;
  assign new_n10835_ = ~new_n10532_ | ~new_n10459_;
  assign new_n10836_ = ~new_n1843_ | ~new_n10458_;
  assign new_n10837_ = ~new_n1406_ | ~new_n10457_;
  assign new_n10838_ = ~new_n10533_;
  assign new_n10839_ = ~new_n10658_ | ~new_n10838_;
  assign new_n10840_ = ~new_n10533_ | ~new_n10560_;
  assign new_n10841_ = ~new_n1840_ | ~new_n10453_;
  assign new_n10842_ = ~new_n1410_ | ~new_n10451_;
  assign new_n10843_ = ~new_n10842_ | ~new_n10841_;
  assign new_n10844_ = ~new_n1837_ | ~new_n10454_;
  assign new_n10845_ = ~new_n1411_ | ~new_n10441_;
  assign new_n10846_ = ~new_n10726_ | ~new_n10483_;
  assign new_n10847_ = ~new_n10561_ | ~new_n10718_;
  assign new_n10848_ = ~new_n1834_ | ~new_n10455_;
  assign new_n10849_ = ~new_n1416_ | ~new_n10452_;
  assign new_n10850_ = ~new_n10727_ | ~new_n10563_;
  assign new_n10851_ = ~new_n10648_ | ~new_n10562_;
  assign new_n10852_ = ~new_n1831_ | ~new_n10450_;
  assign new_n10853_ = ~new_n1417_ | ~new_n10449_;
  assign new_n10854_ = ~new_n10535_;
  assign new_n10855_ = ~new_n10644_ | ~new_n10854_;
  assign new_n10856_ = ~new_n10535_ | ~new_n10564_;
  assign new_n10857_ = ~new_n1828_ | ~new_n10448_;
  assign new_n10858_ = ~new_n1409_ | ~new_n10447_;
  assign new_n10859_ = ~new_n10536_;
  assign new_n10860_ = ~new_n10640_ | ~new_n10859_;
  assign new_n10861_ = ~new_n10536_ | ~new_n10565_;
  assign new_n10862_ = ~new_n1825_ | ~new_n10444_;
  assign new_n10863_ = ~new_n1400_ | ~new_n10442_;
  assign new_n10864_ = ~new_n10863_ | ~new_n10862_;
  assign new_n10865_ = ~new_n1822_ | ~new_n10445_;
  assign new_n10866_ = ~new_n1399_ | ~new_n10443_;
  assign new_n10867_ = ~new_n10737_ | ~new_n10484_;
  assign new_n10868_ = ~new_n10566_ | ~new_n10729_;
  assign new_n10869_ = new_n10982_ & new_n10983_;
  assign new_n10870_ = new_n11000_ & new_n10999_;
  assign new_n10871_ = new_n11004_ & new_n11005_ & new_n11007_ & new_n11006_;
  assign new_n10872_ = new_n11027_ & new_n11026_;
  assign new_n10873_ = new_n10869_ & new_n11061_ & new_n11060_ & new_n11059_;
  assign new_n10874_ = new_n2357_ & new_n10883_;
  assign new_n10875_ = new_n10980_ & new_n10981_ & new_n11070_ & new_n11069_;
  assign new_n10876_ = new_n1790_ & new_n10911_;
  assign new_n10877_ = new_n11067_ & new_n11068_ & new_n10978_;
  assign new_n10878_ = ~new_n2355_;
  assign new_n10879_ = ~new_n2356_;
  assign new_n10880_ = ~new_n1393_;
  assign new_n10881_ = ~new_n2357_;
  assign new_n10882_ = ~new_n1396_;
  assign new_n10883_ = ~new_n1392_;
  assign new_n10884_ = ~new_n1391_;
  assign new_n10885_ = ~new_n2347_;
  assign new_n10886_ = ~new_n1394_;
  assign new_n10887_ = ~new_n2349_;
  assign new_n10888_ = ~new_n2346_;
  assign new_n10889_ = ~new_n2348_;
  assign new_n10890_ = ~new_n2350_;
  assign new_n10891_ = ~new_n1403_;
  assign new_n10892_ = ~new_n2351_;
  assign new_n10893_ = ~new_n1398_;
  assign new_n10894_ = ~new_n1395_;
  assign new_n10895_ = ~new_n1402_;
  assign new_n10896_ = ~new_n1412_;
  assign new_n10897_ = ~new_n1413_;
  assign new_n10898_ = ~new_n1843_;
  assign new_n10899_ = ~new_n1846_;
  assign new_n10900_ = ~new_n1411_;
  assign new_n10901_ = ~new_n1416_;
  assign new_n10902_ = ~new_n1810_;
  assign new_n10903_ = ~new_n1404_;
  assign new_n10904_ = ~new_n1420_;
  assign new_n10905_ = ~new_n1421_;
  assign new_n10906_ = ~new_n1408_;
  assign new_n10907_ = ~new_n1407_;
  assign new_n10908_ = ~new_n1397_;
  assign new_n10909_ = ~new_n1401_;
  assign new_n10910_ = ~new_n1790_;
  assign new_n10911_ = ~new_n1414_;
  assign new_n10912_ = ~new_n11010_ | ~new_n11009_;
  assign new_n10913_ = ~new_n1795_;
  assign new_n10914_ = ~new_n1405_;
  assign new_n10915_ = ~new_n1825_;
  assign new_n10916_ = ~new_n1828_;
  assign new_n10917_ = ~new_n1798_;
  assign new_n10918_ = ~new_n1801_;
  assign new_n10919_ = ~new_n1807_;
  assign new_n10920_ = ~new_n1804_;
  assign new_n10921_ = ~new_n1813_;
  assign new_n10922_ = ~new_n1816_;
  assign new_n10923_ = ~new_n1819_;
  assign new_n10924_ = ~new_n1822_;
  assign new_n10925_ = ~new_n1399_;
  assign new_n10926_ = ~new_n1409_;
  assign new_n10927_ = ~new_n1400_;
  assign new_n10928_ = ~new_n1417_;
  assign new_n10929_ = ~new_n1831_;
  assign new_n10930_ = ~new_n1834_;
  assign new_n10931_ = ~new_n1837_;
  assign new_n10932_ = ~new_n1840_;
  assign new_n10933_ = ~new_n1410_;
  assign new_n10934_ = ~new_n1406_;
  assign new_n10935_ = ~new_n1419_;
  assign new_n10936_ = ~new_n1418_;
  assign new_n10937_ = ~new_n1848_;
  assign new_n10938_ = ~new_n2354_;
  assign new_n10939_ = ~new_n2353_;
  assign new_n10940_ = ~new_n2352_;
  assign new_n10941_ = ~new_n10874_ | ~new_n10988_;
  assign new_n10942_ = ~new_n10875_ | ~new_n10950_ | ~new_n10987_ | ~new_n10985_;
  assign new_n10943_ = ~new_n10972_ | ~new_n11058_;
  assign new_n10944_ = new_n2347_ & new_n10976_;
  assign new_n10945_ = new_n2349_ & new_n10894_;
  assign new_n10946_ = new_n2346_ & new_n10884_;
  assign new_n10947_ = new_n2348_ & new_n10886_;
  assign new_n10948_ = new_n1403_ & new_n10892_;
  assign new_n10949_ = new_n1398_ & new_n10940_;
  assign new_n10950_ = new_n10986_ & new_n10984_;
  assign new_n10951_ = new_n10992_ & new_n10989_;
  assign new_n10952_ = new_n10991_ & new_n10994_ & new_n11064_;
  assign new_n10953_ = new_n1404_ & new_n10919_;
  assign new_n10954_ = new_n11008_ & new_n11012_;
  assign new_n10955_ = new_n10954_ & new_n11003_;
  assign new_n10956_ = new_n10871_ & new_n11016_ & new_n11015_;
  assign new_n10957_ = new_n1798_ & new_n10914_;
  assign new_n10958_ = new_n11022_ & new_n11024_ & new_n11023_;
  assign new_n10959_ = new_n1813_ & new_n10907_;
  assign new_n10960_ = new_n11034_ & new_n11033_;
  assign new_n10961_ = new_n10960_ & new_n10872_;
  assign new_n10962_ = new_n1399_ & new_n10924_;
  assign new_n10963_ = new_n1400_ & new_n10915_;
  assign new_n10964_ = new_n10965_ & new_n11036_ & new_n11037_;
  assign new_n10965_ = new_n11040_ & new_n11039_;
  assign new_n10966_ = new_n10870_ & new_n10967_;
  assign new_n10967_ = new_n11048_ & new_n11049_;
  assign new_n10968_ = new_n1410_ & new_n10932_;
  assign new_n10969_ = new_n1406_ & new_n10898_;
  assign new_n10970_ = new_n10971_ & new_n11051_ & new_n11053_;
  assign new_n10971_ = new_n11055_ & new_n11054_;
  assign new_n10972_ = new_n10997_ & new_n10996_;
  assign new_n10973_ = new_n2354_ & new_n10897_;
  assign new_n10974_ = new_n10991_ & new_n10990_;
  assign new_n10975_ = new_n10993_ & new_n10992_ & new_n10873_ & new_n10994_;
  assign new_n10976_ = ~new_n1390_;
  assign new_n10977_ = ~new_n11063_ | ~new_n11062_;
  assign new_n10978_ = ~new_n2355_ | ~new_n10880_;
  assign new_n10979_ = ~new_n1392_ | ~new_n10881_;
  assign new_n10980_ = ~new_n1391_ | ~new_n10888_;
  assign new_n10981_ = ~new_n1394_ | ~new_n10889_;
  assign new_n10982_ = ~new_n2350_ | ~new_n10895_;
  assign new_n10983_ = ~new_n2351_ | ~new_n10891_;
  assign new_n10984_ = ~new_n10948_ | ~new_n10982_;
  assign new_n10985_ = ~new_n10949_ | ~new_n10869_;
  assign new_n10986_ = ~new_n1395_ | ~new_n10887_;
  assign new_n10987_ = ~new_n1402_ | ~new_n10890_;
  assign new_n10988_ = ~new_n1396_ | ~new_n10879_;
  assign new_n10989_ = ~new_n10978_ | ~new_n10944_ | ~new_n10980_;
  assign new_n10990_ = ~new_n10978_ | ~new_n10945_ | ~new_n10875_;
  assign new_n10991_ = ~new_n2356_ | ~new_n10978_ | ~new_n10882_;
  assign new_n10992_ = ~new_n10946_ | ~new_n10978_;
  assign new_n10993_ = ~new_n10978_ | ~new_n10947_ | ~new_n10875_;
  assign new_n10994_ = ~new_n1393_ | ~new_n10878_;
  assign new_n10995_ = ~new_n10990_ | ~new_n10951_ | ~new_n10942_ | ~new_n10993_;
  assign new_n10996_ = ~new_n1412_ | ~new_n10939_;
  assign new_n10997_ = ~new_n1413_ | ~new_n10938_;
  assign new_n10998_ = ~new_n1411_ | ~new_n10931_;
  assign new_n10999_ = ~new_n1843_ | ~new_n10934_;
  assign new_n11000_ = ~new_n1846_ | ~new_n10935_;
  assign new_n11001_ = ~new_n1416_ | ~new_n10930_;
  assign new_n11002_ = ~new_n1810_ | ~new_n10906_;
  assign new_n11003_ = ~new_n10953_ | ~new_n11002_;
  assign new_n11004_ = ~new_n1420_ | ~new_n10923_;
  assign new_n11005_ = ~new_n1421_ | ~new_n10922_;
  assign new_n11006_ = ~new_n1408_ | ~new_n10902_;
  assign new_n11007_ = ~new_n1407_ | ~new_n10921_;
  assign new_n11008_ = ~new_n1397_ | ~new_n10920_;
  assign new_n11009_ = new_n1787_ | new_n10876_;
  assign new_n11010_ = ~new_n1414_ | ~new_n10910_;
  assign new_n11011_ = ~new_n10912_;
  assign new_n11012_ = ~new_n1401_ | ~new_n10918_;
  assign new_n11013_ = ~new_n1795_ | ~new_n11011_;
  assign new_n11014_ = ~new_n1415_ | ~new_n11013_;
  assign new_n11015_ = ~new_n10912_ | ~new_n10913_;
  assign new_n11016_ = ~new_n1405_ | ~new_n10917_;
  assign new_n11017_ = ~new_n10956_ | ~new_n10955_ | ~new_n11014_;
  assign new_n11018_ = ~new_n10957_ | ~new_n11012_;
  assign new_n11019_ = ~new_n1801_ | ~new_n10909_;
  assign new_n11020_ = ~new_n11019_ | ~new_n11018_;
  assign new_n11021_ = ~new_n11020_ | ~new_n11008_;
  assign new_n11022_ = ~new_n1807_ | ~new_n10903_;
  assign new_n11023_ = ~new_n1804_ | ~new_n10908_;
  assign new_n11024_ = ~new_n1810_ | ~new_n10906_;
  assign new_n11025_ = ~new_n11021_ | ~new_n10958_;
  assign new_n11026_ = ~new_n1825_ | ~new_n10927_;
  assign new_n11027_ = ~new_n1828_ | ~new_n10926_;
  assign new_n11028_ = ~new_n10959_ | ~new_n11005_;
  assign new_n11029_ = ~new_n1816_ | ~new_n10905_;
  assign new_n11030_ = ~new_n11029_ | ~new_n11028_;
  assign new_n11031_ = ~new_n10871_ | ~new_n11025_ | ~new_n11003_;
  assign new_n11032_ = ~new_n11030_ | ~new_n11004_;
  assign new_n11033_ = ~new_n1819_ | ~new_n10904_;
  assign new_n11034_ = ~new_n1822_ | ~new_n10925_;
  assign new_n11035_ = ~new_n11017_ | ~new_n10961_ | ~new_n11031_ | ~new_n11032_;
  assign new_n11036_ = ~new_n10962_ | ~new_n10872_;
  assign new_n11037_ = ~new_n1409_ | ~new_n10916_;
  assign new_n11038_ = ~new_n1828_ | ~new_n10926_;
  assign new_n11039_ = ~new_n10963_ | ~new_n11038_;
  assign new_n11040_ = ~new_n1417_ | ~new_n10929_;
  assign new_n11041_ = ~new_n11035_ | ~new_n10964_;
  assign new_n11042_ = ~new_n1831_ | ~new_n10928_;
  assign new_n11043_ = ~new_n11042_ | ~new_n11041_;
  assign new_n11044_ = ~new_n11043_ | ~new_n11001_;
  assign new_n11045_ = ~new_n1834_ | ~new_n10901_;
  assign new_n11046_ = ~new_n11045_ | ~new_n11044_;
  assign new_n11047_ = ~new_n11046_ | ~new_n10998_;
  assign new_n11048_ = ~new_n1837_ | ~new_n10900_;
  assign new_n11049_ = ~new_n1840_ | ~new_n10933_;
  assign new_n11050_ = ~new_n11047_ | ~new_n10966_;
  assign new_n11051_ = ~new_n10968_ | ~new_n10870_;
  assign new_n11052_ = ~new_n1846_ | ~new_n10935_;
  assign new_n11053_ = ~new_n10969_ | ~new_n11052_;
  assign new_n11054_ = ~new_n1419_ | ~new_n10899_;
  assign new_n11055_ = ~new_n1418_ | ~new_n10937_;
  assign new_n11056_ = ~new_n11050_ | ~new_n10970_;
  assign new_n11057_ = ~new_n1848_ | ~new_n10936_;
  assign new_n11058_ = ~new_n11057_ | ~new_n11056_;
  assign new_n11059_ = ~new_n10973_ | ~new_n10996_;
  assign new_n11060_ = ~new_n2353_ | ~new_n10896_;
  assign new_n11061_ = ~new_n2352_ | ~new_n10893_;
  assign new_n11062_ = ~new_n2356_ | ~new_n10979_;
  assign new_n11063_ = ~new_n10882_ | ~new_n10979_;
  assign new_n11064_ = ~new_n10874_ | ~new_n11065_;
  assign new_n11065_ = ~new_n1396_ | ~new_n10879_;
  assign new_n11066_ = ~new_n10995_ | ~new_n10977_;
  assign new_n11067_ = ~new_n10952_ | ~new_n11066_;
  assign new_n11068_ = ~new_n10975_ | ~new_n10974_ | ~new_n10941_ | ~new_n10989_ | ~new_n10943_;
  assign new_n11069_ = ~new_n1390_ | ~new_n10885_;
  assign new_n11070_ = ~new_n2347_ | ~new_n10976_;
  assign new_n11071_ = new_n1396_ & new_n11072_;
  assign new_n11072_ = ~new_n1393_;
  assign new_n11073_ = new_n11251_ & new_n11268_;
  assign new_n11074_ = new_n11270_ & new_n11269_;
  assign new_n11075_ = new_n11246_ & new_n11307_;
  assign new_n11076_ = new_n11309_ & new_n11308_;
  assign new_n11077_ = new_n11326_ & new_n11325_;
  assign new_n11078_ = new_n11352_ & new_n11351_;
  assign new_n11079_ = new_n11450_ & new_n11449_;
  assign new_n11080_ = ~new_n11407_ | ~new_n11410_;
  assign new_n11081_ = ~new_n11396_ | ~new_n11399_;
  assign new_n11082_ = ~new_n11385_ | ~new_n11388_;
  assign new_n11083_ = ~new_n11377_ | ~new_n11379_;
  assign new_n11084_ = ~new_n11415_ | ~new_n11223_ | ~new_n11242_;
  assign new_n11085_ = ~new_n11303_ | ~new_n11305_;
  assign new_n11086_ = ~new_n11295_ | ~new_n11298_;
  assign new_n11087_ = ~new_n11287_ | ~new_n11289_;
  assign new_n11088_ = ~new_n11092_ | ~new_n11413_;
  assign new_n11089_ = ~new_n1813_;
  assign new_n11090_ = ~new_n1798_;
  assign new_n11091_ = ~new_n1790_;
  assign new_n11092_ = ~new_n1790_ | ~new_n11160_;
  assign new_n11093_ = ~new_n1415_;
  assign new_n11094_ = ~new_n1801_;
  assign new_n11095_ = ~new_n1405_;
  assign new_n11096_ = ~new_n1405_ | ~new_n11090_;
  assign new_n11097_ = ~new_n1401_;
  assign new_n11098_ = ~new_n1810_;
  assign new_n11099_ = ~new_n1807_;
  assign new_n11100_ = ~new_n1804_;
  assign new_n11101_ = ~new_n1408_;
  assign new_n11102_ = ~new_n1404_;
  assign new_n11103_ = ~new_n1397_;
  assign new_n11104_ = ~new_n1397_ | ~new_n11100_;
  assign new_n11105_ = ~new_n1816_;
  assign new_n11106_ = ~new_n1407_;
  assign new_n11107_ = ~new_n1407_ | ~new_n11089_;
  assign new_n11108_ = ~new_n1421_;
  assign new_n11109_ = ~new_n1819_;
  assign new_n11110_ = ~new_n1420_;
  assign new_n11111_ = ~new_n11276_ | ~new_n11275_;
  assign new_n11112_ = ~new_n11104_ | ~new_n11291_;
  assign new_n11113_ = ~new_n11260_ | ~new_n11259_;
  assign new_n11114_ = ~new_n2348_;
  assign new_n11115_ = ~new_n2352_;
  assign new_n11116_ = ~new_n1837_;
  assign new_n11117_ = ~new_n1825_;
  assign new_n11118_ = ~new_n1822_;
  assign new_n11119_ = ~new_n1400_;
  assign new_n11120_ = ~new_n1399_;
  assign new_n11121_ = ~new_n1420_ | ~new_n11109_;
  assign new_n11122_ = ~new_n1828_;
  assign new_n11123_ = ~new_n1409_;
  assign new_n11124_ = ~new_n1831_;
  assign new_n11125_ = ~new_n1417_;
  assign new_n11126_ = ~new_n1840_;
  assign new_n11127_ = ~new_n1834_;
  assign new_n11128_ = ~new_n1410_;
  assign new_n11129_ = ~new_n1411_;
  assign new_n11130_ = ~new_n1416_;
  assign new_n11131_ = ~new_n1416_ | ~new_n11127_;
  assign new_n11132_ = ~new_n1843_;
  assign new_n11133_ = ~new_n1406_;
  assign new_n11134_ = ~new_n11336_ | ~new_n11335_;
  assign new_n11135_ = ~new_n1419_;
  assign new_n11136_ = ~new_n1848_;
  assign new_n11137_ = ~new_n1418_;
  assign new_n11138_ = ~new_n2354_;
  assign new_n11139_ = ~new_n1413_;
  assign new_n11140_ = ~new_n2351_;
  assign new_n11141_ = ~new_n2353_;
  assign new_n11142_ = ~new_n1403_;
  assign new_n11143_ = ~new_n1398_;
  assign new_n11144_ = ~new_n1412_;
  assign new_n11145_ = ~new_n1412_ | ~new_n11141_;
  assign new_n11146_ = ~new_n2350_;
  assign new_n11147_ = ~new_n1402_;
  assign new_n11148_ = ~new_n2349_;
  assign new_n11149_ = ~new_n1395_;
  assign new_n11150_ = ~new_n2347_;
  assign new_n11151_ = ~new_n1394_;
  assign new_n11152_ = ~new_n1394_ | ~new_n11114_;
  assign new_n11153_ = ~new_n1390_;
  assign new_n11154_ = ~new_n2346_;
  assign new_n11155_ = ~new_n1391_;
  assign new_n11156_ = ~new_n11366_ | ~new_n11365_;
  assign new_n11157_ = ~new_n11145_ | ~new_n11381_;
  assign new_n11158_ = ~new_n11131_ | ~new_n11392_;
  assign new_n11159_ = ~new_n11121_ | ~new_n11403_;
  assign new_n11160_ = ~new_n1414_;
  assign new_n11161_ = ~new_n11460_ | ~new_n11459_;
  assign new_n11162_ = ~new_n11474_ | ~new_n11473_;
  assign new_n11163_ = ~new_n11479_ | ~new_n11478_;
  assign new_n11164_ = ~new_n11495_ | ~new_n11494_;
  assign new_n11165_ = ~new_n11500_ | ~new_n11499_;
  assign new_n11166_ = ~new_n11505_ | ~new_n11504_;
  assign new_n11167_ = ~new_n11510_ | ~new_n11509_;
  assign new_n11168_ = ~new_n11515_ | ~new_n11514_;
  assign new_n11169_ = ~new_n11531_ | ~new_n11530_;
  assign new_n11170_ = ~new_n11536_ | ~new_n11535_;
  assign new_n11171_ = ~new_n11419_ | ~new_n11418_;
  assign new_n11172_ = ~new_n11428_ | ~new_n11427_;
  assign new_n11173_ = ~new_n11435_ | ~new_n11434_;
  assign new_n11174_ = ~new_n11439_ | ~new_n11438_;
  assign new_n11175_ = ~new_n11448_ | ~new_n11447_;
  assign new_n11176_ = ~new_n11469_ | ~new_n11468_;
  assign new_n11177_ = ~new_n11486_ | ~new_n11485_;
  assign new_n11178_ = ~new_n11490_ | ~new_n11489_;
  assign new_n11179_ = ~new_n11522_ | ~new_n11521_;
  assign new_n11180_ = ~new_n11526_ | ~new_n11525_;
  assign new_n11181_ = ~new_n11543_ | ~new_n11542_;
  assign new_n11182_ = new_n11262_ & new_n11250_;
  assign new_n11183_ = new_n11265_ & new_n11266_;
  assign new_n11184_ = new_n11278_ & new_n11252_;
  assign new_n11185_ = new_n11281_ & new_n11282_;
  assign new_n11186_ = new_n11107_ & new_n11421_ & new_n11420_;
  assign new_n11187_ = new_n11424_ & new_n11252_;
  assign new_n11188_ = new_n11297_ & new_n11074_;
  assign new_n11189_ = new_n11431_ & new_n11251_;
  assign new_n11190_ = new_n11096_ & new_n11441_ & new_n11440_;
  assign new_n11191_ = new_n11444_ & new_n11250_;
  assign new_n11192_ = new_n11284_ & new_n11075_;
  assign new_n11193_ = new_n11329_ & new_n11247_;
  assign new_n11194_ = new_n11355_ & new_n11248_;
  assign new_n11195_ = new_n11371_ & new_n11372_;
  assign new_n11196_ = new_n11374_ & new_n11453_;
  assign new_n11197_ = new_n11375_ & new_n11372_ & new_n11371_;
  assign new_n11198_ = ~new_n11457_ | ~new_n11456_;
  assign new_n11199_ = new_n11152_ & new_n11462_ & new_n11461_;
  assign new_n11200_ = new_n11465_ & new_n11249_;
  assign new_n11201_ = ~new_n11471_ | ~new_n11470_;
  assign new_n11202_ = ~new_n11476_ | ~new_n11475_;
  assign new_n11203_ = new_n11482_ & new_n11248_;
  assign new_n11204_ = ~new_n11492_ | ~new_n11491_;
  assign new_n11205_ = ~new_n11497_ | ~new_n11496_;
  assign new_n11206_ = ~new_n11502_ | ~new_n11501_;
  assign new_n11207_ = ~new_n11507_ | ~new_n11506_;
  assign new_n11208_ = ~new_n11512_ | ~new_n11511_;
  assign new_n11209_ = new_n11518_ & new_n11247_;
  assign new_n11210_ = ~new_n11528_ | ~new_n11527_;
  assign new_n11211_ = ~new_n11533_ | ~new_n11532_;
  assign new_n11212_ = new_n11409_ & new_n11076_;
  assign new_n11213_ = new_n11539_ & new_n11246_;
  assign new_n11214_ = new_n11417_ & new_n11416_;
  assign new_n11215_ = ~new_n11185_ | ~new_n11279_;
  assign new_n11216_ = new_n11426_ & new_n11425_;
  assign new_n11217_ = new_n11433_ & new_n11432_;
  assign new_n11218_ = new_n11437_ & new_n11436_;
  assign new_n11219_ = ~new_n11183_ | ~new_n11263_;
  assign new_n11220_ = new_n11446_ & new_n11445_;
  assign new_n11221_ = ~new_n2357_;
  assign new_n11222_ = ~new_n1392_;
  assign new_n11223_ = new_n11455_ & new_n11454_;
  assign new_n11224_ = ~new_n11195_ | ~new_n11369_;
  assign new_n11225_ = new_n11467_ & new_n11466_;
  assign new_n11226_ = ~new_n11362_ | ~new_n11361_;
  assign new_n11227_ = ~new_n11358_ | ~new_n11357_;
  assign new_n11228_ = new_n11484_ & new_n11483_;
  assign new_n11229_ = new_n11488_ & new_n11487_;
  assign new_n11230_ = ~new_n11348_ | ~new_n11347_;
  assign new_n11231_ = ~new_n11344_ | ~new_n11343_;
  assign new_n11232_ = ~new_n1795_;
  assign new_n11233_ = ~new_n11340_ | ~new_n11339_;
  assign new_n11234_ = ~new_n1846_;
  assign new_n11235_ = ~new_n11332_ | ~new_n11331_;
  assign new_n11236_ = new_n11520_ & new_n11519_;
  assign new_n11237_ = new_n11524_ & new_n11523_;
  assign new_n11238_ = ~new_n11322_ | ~new_n11321_;
  assign new_n11239_ = ~new_n11318_ | ~new_n11317_;
  assign new_n11240_ = ~new_n11314_ | ~new_n11313_;
  assign new_n11241_ = new_n11541_ & new_n11540_;
  assign new_n11242_ = ~new_n11196_ | ~new_n11224_;
  assign new_n11243_ = ~new_n11152_;
  assign new_n11244_ = ~new_n11096_;
  assign new_n11245_ = ~new_n11107_;
  assign new_n11246_ = ~new_n1822_ | ~new_n11120_;
  assign new_n11247_ = ~new_n1837_ | ~new_n11129_;
  assign new_n11248_ = ~new_n2352_ | ~new_n11143_;
  assign new_n11249_ = ~new_n2348_ | ~new_n11151_;
  assign new_n11250_ = ~new_n1798_ | ~new_n11095_;
  assign new_n11251_ = ~new_n1807_ | ~new_n11102_;
  assign new_n11252_ = ~new_n1813_ | ~new_n11106_;
  assign new_n11253_ = ~new_n11131_;
  assign new_n11254_ = ~new_n11145_;
  assign new_n11255_ = ~new_n11104_;
  assign new_n11256_ = ~new_n11121_;
  assign new_n11257_ = ~new_n11092_;
  assign new_n11258_ = ~new_n11257_ | ~new_n11093_;
  assign new_n11259_ = ~new_n11258_ | ~new_n11232_;
  assign new_n11260_ = ~new_n1415_ | ~new_n11092_;
  assign new_n11261_ = ~new_n11113_;
  assign new_n11262_ = ~new_n1801_ | ~new_n11097_;
  assign new_n11263_ = ~new_n11182_ | ~new_n11113_;
  assign new_n11264_ = ~new_n11097_ | ~new_n11096_;
  assign new_n11265_ = ~new_n11264_ | ~new_n11094_;
  assign new_n11266_ = ~new_n1401_ | ~new_n11244_;
  assign new_n11267_ = ~new_n11219_;
  assign new_n11268_ = ~new_n1810_ | ~new_n11101_;
  assign new_n11269_ = ~new_n1408_ | ~new_n11098_;
  assign new_n11270_ = ~new_n1404_ | ~new_n11099_;
  assign new_n11271_ = ~new_n11255_ | ~new_n11073_;
  assign new_n11272_ = ~new_n11074_ | ~new_n11271_;
  assign new_n11273_ = ~new_n1804_ | ~new_n11103_;
  assign new_n11274_ = ~new_n1810_ | ~new_n11101_;
  assign new_n11275_ = ~new_n11073_ | ~new_n11273_ | ~new_n11219_;
  assign new_n11276_ = ~new_n11274_ | ~new_n11272_;
  assign new_n11277_ = ~new_n11111_;
  assign new_n11278_ = ~new_n1816_ | ~new_n11108_;
  assign new_n11279_ = ~new_n11184_ | ~new_n11111_;
  assign new_n11280_ = ~new_n11108_ | ~new_n11107_;
  assign new_n11281_ = ~new_n11280_ | ~new_n11105_;
  assign new_n11282_ = ~new_n1421_ | ~new_n11245_;
  assign new_n11283_ = ~new_n11215_;
  assign new_n11284_ = ~new_n1819_ | ~new_n11110_;
  assign new_n11285_ = ~new_n11284_ | ~new_n11121_;
  assign new_n11286_ = ~new_n11277_ | ~new_n11107_;
  assign new_n11287_ = ~new_n11187_ | ~new_n11286_;
  assign new_n11288_ = ~new_n11111_ | ~new_n11252_;
  assign new_n11289_ = ~new_n11186_ | ~new_n11288_;
  assign new_n11290_ = ~new_n11107_ | ~new_n11252_;
  assign new_n11291_ = ~new_n11273_ | ~new_n11219_;
  assign new_n11292_ = ~new_n11112_;
  assign new_n11293_ = ~new_n1404_ | ~new_n11099_;
  assign new_n11294_ = ~new_n11292_ | ~new_n11293_;
  assign new_n11295_ = ~new_n11189_ | ~new_n11294_;
  assign new_n11296_ = ~new_n11112_ | ~new_n11251_;
  assign new_n11297_ = ~new_n1810_ | ~new_n11101_;
  assign new_n11298_ = ~new_n11188_ | ~new_n11296_;
  assign new_n11299_ = ~new_n1404_ | ~new_n11099_;
  assign new_n11300_ = ~new_n11251_ | ~new_n11299_;
  assign new_n11301_ = ~new_n11273_ | ~new_n11104_;
  assign new_n11302_ = ~new_n11261_ | ~new_n11096_;
  assign new_n11303_ = ~new_n11191_ | ~new_n11302_;
  assign new_n11304_ = ~new_n11113_ | ~new_n11250_;
  assign new_n11305_ = ~new_n11190_ | ~new_n11304_;
  assign new_n11306_ = ~new_n11096_ | ~new_n11250_;
  assign new_n11307_ = ~new_n1825_ | ~new_n11119_;
  assign new_n11308_ = ~new_n1400_ | ~new_n11117_;
  assign new_n11309_ = ~new_n1399_ | ~new_n11118_;
  assign new_n11310_ = ~new_n11256_ | ~new_n11075_;
  assign new_n11311_ = ~new_n11076_ | ~new_n11310_;
  assign new_n11312_ = ~new_n1825_ | ~new_n11119_;
  assign new_n11313_ = ~new_n11192_ | ~new_n11215_;
  assign new_n11314_ = ~new_n11312_ | ~new_n11311_;
  assign new_n11315_ = ~new_n11240_;
  assign new_n11316_ = ~new_n1828_ | ~new_n11123_;
  assign new_n11317_ = ~new_n11316_ | ~new_n11240_;
  assign new_n11318_ = ~new_n1409_ | ~new_n11122_;
  assign new_n11319_ = ~new_n11239_;
  assign new_n11320_ = ~new_n1831_ | ~new_n11125_;
  assign new_n11321_ = ~new_n11320_ | ~new_n11239_;
  assign new_n11322_ = ~new_n1417_ | ~new_n11124_;
  assign new_n11323_ = ~new_n11238_;
  assign new_n11324_ = ~new_n1840_ | ~new_n11128_;
  assign new_n11325_ = ~new_n1410_ | ~new_n11126_;
  assign new_n11326_ = ~new_n1411_ | ~new_n11116_;
  assign new_n11327_ = ~new_n11253_ | ~new_n11247_;
  assign new_n11328_ = ~new_n11077_ | ~new_n11327_;
  assign new_n11329_ = ~new_n1834_ | ~new_n11130_;
  assign new_n11330_ = ~new_n1840_ | ~new_n11128_;
  assign new_n11331_ = ~new_n11324_ | ~new_n11238_ | ~new_n11193_;
  assign new_n11332_ = ~new_n11330_ | ~new_n11328_;
  assign new_n11333_ = ~new_n11235_;
  assign new_n11334_ = ~new_n1843_ | ~new_n11133_;
  assign new_n11335_ = ~new_n11334_ | ~new_n11235_;
  assign new_n11336_ = ~new_n1406_ | ~new_n11132_;
  assign new_n11337_ = ~new_n11134_;
  assign new_n11338_ = ~new_n11337_ | ~new_n11135_;
  assign new_n11339_ = ~new_n11338_ | ~new_n11234_;
  assign new_n11340_ = ~new_n1419_ | ~new_n11134_;
  assign new_n11341_ = ~new_n11233_;
  assign new_n11342_ = ~new_n1848_ | ~new_n11137_;
  assign new_n11343_ = ~new_n11342_ | ~new_n11233_;
  assign new_n11344_ = ~new_n1418_ | ~new_n11136_;
  assign new_n11345_ = ~new_n11231_;
  assign new_n11346_ = ~new_n2354_ | ~new_n11139_;
  assign new_n11347_ = ~new_n11346_ | ~new_n11231_;
  assign new_n11348_ = ~new_n1413_ | ~new_n11138_;
  assign new_n11349_ = ~new_n11230_;
  assign new_n11350_ = ~new_n2351_ | ~new_n11142_;
  assign new_n11351_ = ~new_n1403_ | ~new_n11140_;
  assign new_n11352_ = ~new_n1398_ | ~new_n11115_;
  assign new_n11353_ = ~new_n11254_ | ~new_n11248_;
  assign new_n11354_ = ~new_n11078_ | ~new_n11353_;
  assign new_n11355_ = ~new_n2353_ | ~new_n11144_;
  assign new_n11356_ = ~new_n2351_ | ~new_n11142_;
  assign new_n11357_ = ~new_n11350_ | ~new_n11230_ | ~new_n11194_;
  assign new_n11358_ = ~new_n11356_ | ~new_n11354_;
  assign new_n11359_ = ~new_n11227_;
  assign new_n11360_ = ~new_n2350_ | ~new_n11147_;
  assign new_n11361_ = ~new_n11360_ | ~new_n11227_;
  assign new_n11362_ = ~new_n1402_ | ~new_n11146_;
  assign new_n11363_ = ~new_n11226_;
  assign new_n11364_ = ~new_n2349_ | ~new_n11149_;
  assign new_n11365_ = ~new_n11364_ | ~new_n11226_;
  assign new_n11366_ = ~new_n1395_ | ~new_n11148_;
  assign new_n11367_ = ~new_n11156_;
  assign new_n11368_ = ~new_n2347_ | ~new_n11153_;
  assign new_n11369_ = ~new_n11368_ | ~new_n11156_ | ~new_n11249_;
  assign new_n11370_ = ~new_n11153_ | ~new_n11152_;
  assign new_n11371_ = ~new_n11370_ | ~new_n11150_;
  assign new_n11372_ = ~new_n1390_ | ~new_n11243_;
  assign new_n11373_ = ~new_n11224_;
  assign new_n11374_ = ~new_n2346_ | ~new_n11155_;
  assign new_n11375_ = ~new_n1391_ | ~new_n11154_;
  assign new_n11376_ = ~new_n11367_ | ~new_n11152_;
  assign new_n11377_ = ~new_n11200_ | ~new_n11376_;
  assign new_n11378_ = ~new_n11156_ | ~new_n11249_;
  assign new_n11379_ = ~new_n11199_ | ~new_n11378_;
  assign new_n11380_ = ~new_n11152_ | ~new_n11249_;
  assign new_n11381_ = ~new_n11355_ | ~new_n11230_;
  assign new_n11382_ = ~new_n11157_;
  assign new_n11383_ = ~new_n1398_ | ~new_n11115_;
  assign new_n11384_ = ~new_n11382_ | ~new_n11383_;
  assign new_n11385_ = ~new_n11203_ | ~new_n11384_;
  assign new_n11386_ = ~new_n11157_ | ~new_n11248_;
  assign new_n11387_ = ~new_n2351_ | ~new_n11142_;
  assign new_n11388_ = ~new_n11078_ | ~new_n11387_ | ~new_n11386_;
  assign new_n11389_ = ~new_n1398_ | ~new_n11115_;
  assign new_n11390_ = ~new_n11248_ | ~new_n11389_;
  assign new_n11391_ = ~new_n11355_ | ~new_n11145_;
  assign new_n11392_ = ~new_n11329_ | ~new_n11238_;
  assign new_n11393_ = ~new_n11158_;
  assign new_n11394_ = ~new_n1411_ | ~new_n11116_;
  assign new_n11395_ = ~new_n11393_ | ~new_n11394_;
  assign new_n11396_ = ~new_n11209_ | ~new_n11395_;
  assign new_n11397_ = ~new_n11158_ | ~new_n11247_;
  assign new_n11398_ = ~new_n1840_ | ~new_n11128_;
  assign new_n11399_ = ~new_n11077_ | ~new_n11398_ | ~new_n11397_;
  assign new_n11400_ = ~new_n1411_ | ~new_n11116_;
  assign new_n11401_ = ~new_n11247_ | ~new_n11400_;
  assign new_n11402_ = ~new_n11329_ | ~new_n11131_;
  assign new_n11403_ = ~new_n11284_ | ~new_n11215_;
  assign new_n11404_ = ~new_n11159_;
  assign new_n11405_ = ~new_n1399_ | ~new_n11118_;
  assign new_n11406_ = ~new_n11404_ | ~new_n11405_;
  assign new_n11407_ = ~new_n11213_ | ~new_n11406_;
  assign new_n11408_ = ~new_n11159_ | ~new_n11246_;
  assign new_n11409_ = ~new_n1825_ | ~new_n11119_;
  assign new_n11410_ = ~new_n11212_ | ~new_n11408_;
  assign new_n11411_ = ~new_n1399_ | ~new_n11118_;
  assign new_n11412_ = ~new_n11246_ | ~new_n11411_;
  assign new_n11413_ = ~new_n1414_ | ~new_n11091_;
  assign new_n11414_ = ~new_n11368_ | ~new_n11156_ | ~new_n11249_;
  assign new_n11415_ = ~new_n11197_ | ~new_n11079_ | ~new_n11414_;
  assign new_n11416_ = ~new_n1819_ | ~new_n11110_;
  assign new_n11417_ = ~new_n1420_ | ~new_n11109_;
  assign new_n11418_ = ~new_n11285_ | ~new_n11215_;
  assign new_n11419_ = ~new_n11283_ | ~new_n11214_;
  assign new_n11420_ = ~new_n1816_ | ~new_n11108_;
  assign new_n11421_ = ~new_n1421_ | ~new_n11105_;
  assign new_n11422_ = ~new_n1816_ | ~new_n11108_;
  assign new_n11423_ = ~new_n1421_ | ~new_n11105_;
  assign new_n11424_ = ~new_n11423_ | ~new_n11422_;
  assign new_n11425_ = ~new_n1813_ | ~new_n11106_;
  assign new_n11426_ = ~new_n1407_ | ~new_n11089_;
  assign new_n11427_ = ~new_n11290_ | ~new_n11111_;
  assign new_n11428_ = ~new_n11216_ | ~new_n11277_;
  assign new_n11429_ = ~new_n1810_ | ~new_n11101_;
  assign new_n11430_ = ~new_n1408_ | ~new_n11098_;
  assign new_n11431_ = ~new_n11430_ | ~new_n11429_;
  assign new_n11432_ = ~new_n1807_ | ~new_n11102_;
  assign new_n11433_ = ~new_n1404_ | ~new_n11099_;
  assign new_n11434_ = ~new_n11300_ | ~new_n11112_;
  assign new_n11435_ = ~new_n11217_ | ~new_n11292_;
  assign new_n11436_ = ~new_n1804_ | ~new_n11103_;
  assign new_n11437_ = ~new_n1397_ | ~new_n11100_;
  assign new_n11438_ = ~new_n11301_ | ~new_n11219_;
  assign new_n11439_ = ~new_n11267_ | ~new_n11218_;
  assign new_n11440_ = ~new_n1801_ | ~new_n11097_;
  assign new_n11441_ = ~new_n1401_ | ~new_n11094_;
  assign new_n11442_ = ~new_n1801_ | ~new_n11097_;
  assign new_n11443_ = ~new_n1401_ | ~new_n11094_;
  assign new_n11444_ = ~new_n11443_ | ~new_n11442_;
  assign new_n11445_ = ~new_n1798_ | ~new_n11095_;
  assign new_n11446_ = ~new_n1405_ | ~new_n11090_;
  assign new_n11447_ = ~new_n11306_ | ~new_n11113_;
  assign new_n11448_ = ~new_n11220_ | ~new_n11261_;
  assign new_n11449_ = ~new_n2357_ | ~new_n11222_;
  assign new_n11450_ = ~new_n1392_ | ~new_n11221_;
  assign new_n11451_ = ~new_n2357_ | ~new_n11222_;
  assign new_n11452_ = ~new_n1392_ | ~new_n11221_;
  assign new_n11453_ = ~new_n11452_ | ~new_n11451_;
  assign new_n11454_ = ~new_n11154_ | ~new_n1391_ | ~new_n11453_;
  assign new_n11455_ = ~new_n2346_ | ~new_n11079_ | ~new_n11155_;
  assign new_n11456_ = ~new_n2346_ | ~new_n11155_;
  assign new_n11457_ = ~new_n1391_ | ~new_n11154_;
  assign new_n11458_ = ~new_n11198_;
  assign new_n11459_ = ~new_n11373_ | ~new_n11458_;
  assign new_n11460_ = ~new_n11198_ | ~new_n11224_;
  assign new_n11461_ = ~new_n2347_ | ~new_n11153_;
  assign new_n11462_ = ~new_n1390_ | ~new_n11150_;
  assign new_n11463_ = ~new_n2347_ | ~new_n11153_;
  assign new_n11464_ = ~new_n1390_ | ~new_n11150_;
  assign new_n11465_ = ~new_n11464_ | ~new_n11463_;
  assign new_n11466_ = ~new_n2348_ | ~new_n11151_;
  assign new_n11467_ = ~new_n1394_ | ~new_n11114_;
  assign new_n11468_ = ~new_n11380_ | ~new_n11156_;
  assign new_n11469_ = ~new_n11225_ | ~new_n11367_;
  assign new_n11470_ = ~new_n2349_ | ~new_n11149_;
  assign new_n11471_ = ~new_n1395_ | ~new_n11148_;
  assign new_n11472_ = ~new_n11201_;
  assign new_n11473_ = ~new_n11363_ | ~new_n11472_;
  assign new_n11474_ = ~new_n11201_ | ~new_n11226_;
  assign new_n11475_ = ~new_n2350_ | ~new_n11147_;
  assign new_n11476_ = ~new_n1402_ | ~new_n11146_;
  assign new_n11477_ = ~new_n11202_;
  assign new_n11478_ = ~new_n11359_ | ~new_n11477_;
  assign new_n11479_ = ~new_n11202_ | ~new_n11227_;
  assign new_n11480_ = ~new_n2351_ | ~new_n11142_;
  assign new_n11481_ = ~new_n1403_ | ~new_n11140_;
  assign new_n11482_ = ~new_n11481_ | ~new_n11480_;
  assign new_n11483_ = ~new_n2352_ | ~new_n11143_;
  assign new_n11484_ = ~new_n1398_ | ~new_n11115_;
  assign new_n11485_ = ~new_n11390_ | ~new_n11157_;
  assign new_n11486_ = ~new_n11228_ | ~new_n11382_;
  assign new_n11487_ = ~new_n2353_ | ~new_n11144_;
  assign new_n11488_ = ~new_n1412_ | ~new_n11141_;
  assign new_n11489_ = ~new_n11391_ | ~new_n11230_;
  assign new_n11490_ = ~new_n11349_ | ~new_n11229_;
  assign new_n11491_ = ~new_n2354_ | ~new_n11139_;
  assign new_n11492_ = ~new_n1413_ | ~new_n11138_;
  assign new_n11493_ = ~new_n11204_;
  assign new_n11494_ = ~new_n11345_ | ~new_n11493_;
  assign new_n11495_ = ~new_n11204_ | ~new_n11231_;
  assign new_n11496_ = ~new_n1795_ | ~new_n11093_;
  assign new_n11497_ = ~new_n1415_ | ~new_n11232_;
  assign new_n11498_ = ~new_n11205_;
  assign new_n11499_ = ~new_n11498_ | ~new_n11257_;
  assign new_n11500_ = ~new_n11205_ | ~new_n11092_;
  assign new_n11501_ = ~new_n1848_ | ~new_n11137_;
  assign new_n11502_ = ~new_n1418_ | ~new_n11136_;
  assign new_n11503_ = ~new_n11206_;
  assign new_n11504_ = ~new_n11341_ | ~new_n11503_;
  assign new_n11505_ = ~new_n11206_ | ~new_n11233_;
  assign new_n11506_ = ~new_n1846_ | ~new_n11135_;
  assign new_n11507_ = ~new_n1419_ | ~new_n11234_;
  assign new_n11508_ = ~new_n11207_;
  assign new_n11509_ = ~new_n11508_ | ~new_n11337_;
  assign new_n11510_ = ~new_n11207_ | ~new_n11134_;
  assign new_n11511_ = ~new_n1843_ | ~new_n11133_;
  assign new_n11512_ = ~new_n1406_ | ~new_n11132_;
  assign new_n11513_ = ~new_n11208_;
  assign new_n11514_ = ~new_n11333_ | ~new_n11513_;
  assign new_n11515_ = ~new_n11208_ | ~new_n11235_;
  assign new_n11516_ = ~new_n1840_ | ~new_n11128_;
  assign new_n11517_ = ~new_n1410_ | ~new_n11126_;
  assign new_n11518_ = ~new_n11517_ | ~new_n11516_;
  assign new_n11519_ = ~new_n1837_ | ~new_n11129_;
  assign new_n11520_ = ~new_n1411_ | ~new_n11116_;
  assign new_n11521_ = ~new_n11401_ | ~new_n11158_;
  assign new_n11522_ = ~new_n11236_ | ~new_n11393_;
  assign new_n11523_ = ~new_n1834_ | ~new_n11130_;
  assign new_n11524_ = ~new_n1416_ | ~new_n11127_;
  assign new_n11525_ = ~new_n11402_ | ~new_n11238_;
  assign new_n11526_ = ~new_n11323_ | ~new_n11237_;
  assign new_n11527_ = ~new_n1831_ | ~new_n11125_;
  assign new_n11528_ = ~new_n1417_ | ~new_n11124_;
  assign new_n11529_ = ~new_n11210_;
  assign new_n11530_ = ~new_n11319_ | ~new_n11529_;
  assign new_n11531_ = ~new_n11210_ | ~new_n11239_;
  assign new_n11532_ = ~new_n1828_ | ~new_n11123_;
  assign new_n11533_ = ~new_n1409_ | ~new_n11122_;
  assign new_n11534_ = ~new_n11211_;
  assign new_n11535_ = ~new_n11315_ | ~new_n11534_;
  assign new_n11536_ = ~new_n11211_ | ~new_n11240_;
  assign new_n11537_ = ~new_n1825_ | ~new_n11119_;
  assign new_n11538_ = ~new_n1400_ | ~new_n11117_;
  assign new_n11539_ = ~new_n11538_ | ~new_n11537_;
  assign new_n11540_ = ~new_n1822_ | ~new_n11120_;
  assign new_n11541_ = ~new_n1399_ | ~new_n11118_;
  assign new_n11542_ = ~new_n11412_ | ~new_n11159_;
  assign new_n11543_ = ~new_n11241_ | ~new_n11404_;
  assign new_n11544_ = new_n11750_ & new_n11749_;
  assign new_n11545_ = new_n11762_ & new_n11761_;
  assign new_n11546_ = new_n11793_ & new_n11792_;
  assign new_n11547_ = new_n11811_ & new_n11810_;
  assign new_n11548_ = new_n11823_ & new_n11822_;
  assign new_n11549_ = new_n12047_ & new_n12046_;
  assign new_n11550_ = new_n11879_ & new_n11876_;
  assign new_n11551_ = new_n11870_ & new_n11867_;
  assign new_n11552_ = new_n11863_ & new_n11860_;
  assign new_n11553_ = new_n11854_ & new_n11900_ & new_n11851_;
  assign new_n11554_ = new_n11785_ & new_n11782_;
  assign new_n11555_ = new_n11778_ & new_n11775_;
  assign new_n11556_ = ~new_n1548_;
  assign new_n11557_ = ~new_n1512_;
  assign new_n11558_ = ~new_n1512_ | ~new_n11598_;
  assign new_n11559_ = ~new_n1511_;
  assign new_n11560_ = ~new_n1514_;
  assign new_n11561_ = ~new_n1516_;
  assign new_n11562_ = ~new_n1516_ | ~new_n11601_;
  assign new_n11563_ = ~new_n1515_;
  assign new_n11564_ = ~new_n1518_;
  assign new_n11565_ = ~new_n1517_;
  assign new_n11566_ = ~new_n1513_;
  assign new_n11567_ = ~new_n1510_;
  assign new_n11568_ = ~new_n1509_;
  assign new_n11569_ = ~new_n11759_ | ~new_n11758_;
  assign new_n11570_ = ~new_n11747_ | ~new_n11746_;
  assign new_n11571_ = ~new_n1491_;
  assign new_n11572_ = ~new_n1492_;
  assign new_n11573_ = ~new_n1493_;
  assign new_n11574_ = ~new_n1494_;
  assign new_n11575_ = ~new_n1502_;
  assign new_n11576_ = ~new_n1502_ | ~new_n11611_;
  assign new_n11577_ = ~new_n1501_;
  assign new_n11578_ = ~new_n1508_;
  assign new_n11579_ = ~new_n1506_;
  assign new_n11580_ = ~new_n1507_;
  assign new_n11581_ = ~new_n1507_ | ~new_n11614_;
  assign new_n11582_ = ~new_n1505_;
  assign new_n11583_ = ~new_n1504_;
  assign new_n11584_ = ~new_n1503_;
  assign new_n11585_ = ~new_n1500_;
  assign new_n11586_ = ~new_n1498_;
  assign new_n11587_ = ~new_n1499_;
  assign new_n11588_ = ~new_n1499_ | ~new_n11620_;
  assign new_n11589_ = ~new_n1497_;
  assign new_n11590_ = ~new_n1496_;
  assign new_n11591_ = ~new_n1495_;
  assign new_n11592_ = ~new_n1492_ | ~new_n11609_;
  assign new_n11593_ = ~new_n11740_ | ~new_n11849_;
  assign new_n11594_ = ~new_n11588_ | ~new_n11856_;
  assign new_n11595_ = ~new_n11808_ | ~new_n11807_;
  assign new_n11596_ = ~new_n11581_ | ~new_n11872_;
  assign new_n11597_ = ~new_n11906_ | ~new_n11905_;
  assign new_n11598_ = ~new_n11935_ | ~new_n11934_;
  assign new_n11599_ = ~new_n11932_ | ~new_n11931_;
  assign new_n11600_ = ~new_n11914_ | ~new_n11913_;
  assign new_n11601_ = ~new_n11926_ | ~new_n11925_;
  assign new_n11602_ = ~new_n11923_ | ~new_n11922_;
  assign new_n11603_ = ~new_n11917_ | ~new_n11916_;
  assign new_n11604_ = ~new_n11920_ | ~new_n11919_;
  assign new_n11605_ = ~new_n11929_ | ~new_n11928_;
  assign new_n11606_ = ~new_n11938_ | ~new_n11937_;
  assign new_n11607_ = ~new_n11978_ | ~new_n11977_;
  assign new_n11608_ = ~new_n11981_ | ~new_n11980_;
  assign new_n11609_ = ~new_n11984_ | ~new_n11983_;
  assign new_n11610_ = ~new_n11987_ | ~new_n11986_;
  assign new_n11611_ = ~new_n12011_ | ~new_n12010_;
  assign new_n11612_ = ~new_n12008_ | ~new_n12007_;
  assign new_n11613_ = ~new_n11990_ | ~new_n11989_;
  assign new_n11614_ = ~new_n11999_ | ~new_n11998_;
  assign new_n11615_ = ~new_n11993_ | ~new_n11992_;
  assign new_n11616_ = ~new_n11996_ | ~new_n11995_;
  assign new_n11617_ = ~new_n12002_ | ~new_n12001_;
  assign new_n11618_ = ~new_n12005_ | ~new_n12004_;
  assign new_n11619_ = ~new_n12014_ | ~new_n12013_;
  assign new_n11620_ = ~new_n12023_ | ~new_n12022_;
  assign new_n11621_ = ~new_n12017_ | ~new_n12016_;
  assign new_n11622_ = ~new_n12020_ | ~new_n12019_;
  assign new_n11623_ = ~new_n12026_ | ~new_n12025_;
  assign new_n11624_ = ~new_n12029_ | ~new_n12028_;
  assign new_n11625_ = ~new_n12035_ | ~new_n12034_;
  assign new_n11626_ = ~new_n12142_ | ~new_n12141_;
  assign new_n11627_ = ~new_n11941_ | ~new_n11940_;
  assign new_n11628_ = ~new_n11948_ | ~new_n11947_;
  assign new_n11629_ = ~new_n11955_ | ~new_n11954_;
  assign new_n11630_ = ~new_n11962_ | ~new_n11961_;
  assign new_n11631_ = ~new_n11969_ | ~new_n11968_;
  assign new_n11632_ = ~new_n11976_ | ~new_n11975_;
  assign new_n11633_ = ~new_n12038_ | ~new_n12037_;
  assign new_n11634_ = ~new_n12045_ | ~new_n12044_;
  assign new_n11635_ = ~new_n12052_ | ~new_n12051_;
  assign new_n11636_ = ~new_n12057_ | ~new_n12056_;
  assign new_n11637_ = ~new_n12064_ | ~new_n12063_;
  assign new_n11638_ = ~new_n12071_ | ~new_n12070_;
  assign new_n11639_ = ~new_n12078_ | ~new_n12077_;
  assign new_n11640_ = ~new_n12085_ | ~new_n12084_;
  assign new_n11641_ = ~new_n12090_ | ~new_n12089_;
  assign new_n11642_ = ~new_n12097_ | ~new_n12096_;
  assign new_n11643_ = ~new_n12104_ | ~new_n12103_;
  assign new_n11644_ = ~new_n12111_ | ~new_n12110_;
  assign new_n11645_ = ~new_n12118_ | ~new_n12117_;
  assign new_n11646_ = ~new_n12125_ | ~new_n12124_;
  assign new_n11647_ = ~new_n12130_ | ~new_n12129_;
  assign new_n11648_ = ~new_n12137_ | ~new_n12136_;
  assign new_n11649_ = new_n11753_ & new_n11752_;
  assign new_n11650_ = new_n11766_ & new_n11765_;
  assign new_n11651_ = new_n11558_ & new_n11950_ & new_n11949_;
  assign new_n11652_ = new_n11777_ & new_n11545_;
  assign new_n11653_ = new_n11562_ & new_n11971_ & new_n11970_;
  assign new_n11654_ = new_n11784_ & new_n11544_;
  assign new_n11655_ = new_n11797_ & new_n11546_;
  assign new_n11656_ = new_n11795_ & new_n11735_;
  assign new_n11657_ = new_n11815_ & new_n11814_;
  assign new_n11658_ = new_n11827_ & new_n11548_;
  assign new_n11659_ = new_n11825_ & new_n11736_;
  assign new_n11660_ = new_n11899_ & new_n11592_;
  assign new_n11661_ = new_n11848_ & new_n11843_;
  assign new_n11662_ = new_n11896_ & new_n11847_;
  assign new_n11663_ = ~new_n12032_ | ~new_n12031_;
  assign new_n11664_ = new_n11892_ & new_n11592_;
  assign new_n11665_ = new_n11982_ & new_n11573_;
  assign new_n11666_ = new_n11740_ & new_n11737_;
  assign new_n11667_ = new_n11853_ & new_n11733_;
  assign new_n11668_ = new_n11549_ & new_n11737_;
  assign new_n11669_ = new_n11736_ & new_n12073_ & new_n12072_;
  assign new_n11670_ = new_n11862_ & new_n11548_;
  assign new_n11671_ = new_n11576_ & new_n12099_ & new_n12098_;
  assign new_n11672_ = new_n11869_ & new_n11547_;
  assign new_n11673_ = new_n11735_ & new_n12120_ & new_n12119_;
  assign new_n11674_ = new_n11878_ & new_n11546_;
  assign new_n11675_ = ~new_n12139_ | ~new_n12138_;
  assign new_n11676_ = ~new_n1538_;
  assign new_n11677_ = new_n11909_ & new_n11908_;
  assign new_n11678_ = ~new_n1543_;
  assign new_n11679_ = ~new_n1547_;
  assign new_n11680_ = ~new_n1546_;
  assign new_n11681_ = ~new_n1544_;
  assign new_n11682_ = ~new_n1545_;
  assign new_n11683_ = ~new_n1542_;
  assign new_n11684_ = ~new_n1540_;
  assign new_n11685_ = ~new_n1541_;
  assign new_n11686_ = ~new_n1539_;
  assign new_n11687_ = ~new_n11771_ | ~new_n11770_;
  assign new_n11688_ = new_n11943_ & new_n11942_;
  assign new_n11689_ = ~new_n11650_ | ~new_n11767_;
  assign new_n11690_ = new_n11957_ & new_n11956_;
  assign new_n11691_ = ~new_n11901_ | ~new_n11890_;
  assign new_n11692_ = new_n11964_ & new_n11963_;
  assign new_n11693_ = ~new_n11649_ | ~new_n11754_;
  assign new_n11694_ = ~new_n1520_;
  assign new_n11695_ = ~new_n1522_;
  assign new_n11696_ = ~new_n1521_;
  assign new_n11697_ = ~new_n1523_;
  assign new_n11698_ = ~new_n1537_;
  assign new_n11699_ = ~new_n1534_;
  assign new_n11700_ = ~new_n1535_;
  assign new_n11701_ = ~new_n1536_;
  assign new_n11702_ = ~new_n1533_;
  assign new_n11703_ = ~new_n1532_;
  assign new_n11704_ = ~new_n1530_;
  assign new_n11705_ = ~new_n1531_;
  assign new_n11706_ = ~new_n1529_;
  assign new_n11707_ = ~new_n1526_;
  assign new_n11708_ = ~new_n1527_;
  assign new_n11709_ = ~new_n1528_;
  assign new_n11710_ = ~new_n1525_;
  assign new_n11711_ = ~new_n1524_;
  assign new_n11712_ = ~new_n1490_;
  assign new_n11713_ = ~new_n1519_;
  assign new_n11714_ = new_n12040_ & new_n12039_;
  assign new_n11715_ = ~new_n11664_ | ~new_n11844_;
  assign new_n11716_ = ~new_n11838_ | ~new_n11837_;
  assign new_n11717_ = new_n12059_ & new_n12058_;
  assign new_n11718_ = ~new_n11834_ | ~new_n11833_;
  assign new_n11719_ = new_n12066_ & new_n12065_;
  assign new_n11720_ = ~new_n11830_ | ~new_n11829_;
  assign new_n11721_ = new_n12080_ & new_n12079_;
  assign new_n11722_ = ~new_n11743_ | ~new_n11742_;
  assign new_n11723_ = ~new_n11820_ | ~new_n11819_;
  assign new_n11724_ = new_n12092_ & new_n12091_;
  assign new_n11725_ = ~new_n11657_ | ~new_n11816_;
  assign new_n11726_ = new_n12106_ & new_n12105_;
  assign new_n11727_ = ~new_n11804_ | ~new_n11803_;
  assign new_n11728_ = new_n12113_ & new_n12112_;
  assign new_n11729_ = ~new_n11800_ | ~new_n11799_;
  assign new_n11730_ = ~new_n11790_ | ~new_n11789_;
  assign new_n11731_ = new_n12132_ & new_n12131_;
  assign new_n11732_ = ~new_n11903_ | ~new_n11893_;
  assign new_n11733_ = ~new_n11895_ | ~new_n11894_;
  assign new_n11734_ = ~new_n11562_;
  assign new_n11735_ = ~new_n1506_ | ~new_n11616_;
  assign new_n11736_ = ~new_n1498_ | ~new_n11622_;
  assign new_n11737_ = ~new_n1493_ | ~new_n11608_;
  assign new_n11738_ = ~new_n11581_;
  assign new_n11739_ = ~new_n11588_;
  assign new_n11740_ = ~new_n1494_ | ~new_n11610_;
  assign new_n11741_ = new_n1548_ | new_n1518_;
  assign new_n11742_ = ~new_n11603_ | ~new_n11741_;
  assign new_n11743_ = ~new_n1518_ | ~new_n1548_;
  assign new_n11744_ = ~new_n11722_;
  assign new_n11745_ = ~new_n11921_ | ~new_n11565_;
  assign new_n11746_ = ~new_n11745_ | ~new_n11722_;
  assign new_n11747_ = ~new_n1517_ | ~new_n11604_;
  assign new_n11748_ = ~new_n11570_;
  assign new_n11749_ = ~new_n11924_ | ~new_n11563_;
  assign new_n11750_ = ~new_n11927_ | ~new_n11561_;
  assign new_n11751_ = ~new_n11563_ | ~new_n11562_;
  assign new_n11752_ = ~new_n11602_ | ~new_n11751_;
  assign new_n11753_ = ~new_n1515_ | ~new_n11734_;
  assign new_n11754_ = ~new_n11544_ | ~new_n11570_;
  assign new_n11755_ = ~new_n11693_;
  assign new_n11756_ = ~new_n11915_ | ~new_n11560_;
  assign new_n11757_ = ~new_n11930_ | ~new_n11566_;
  assign new_n11758_ = ~new_n11757_ | ~new_n11691_;
  assign new_n11759_ = ~new_n1513_ | ~new_n11605_;
  assign new_n11760_ = ~new_n11569_;
  assign new_n11761_ = ~new_n11933_ | ~new_n11559_;
  assign new_n11762_ = ~new_n11936_ | ~new_n11557_;
  assign new_n11763_ = ~new_n11558_;
  assign new_n11764_ = ~new_n11559_ | ~new_n11558_;
  assign new_n11765_ = ~new_n11599_ | ~new_n11764_;
  assign new_n11766_ = ~new_n1511_ | ~new_n11763_;
  assign new_n11767_ = ~new_n11545_ | ~new_n11569_;
  assign new_n11768_ = ~new_n11689_;
  assign new_n11769_ = ~new_n11939_ | ~new_n11567_;
  assign new_n11770_ = ~new_n11769_ | ~new_n11689_;
  assign new_n11771_ = ~new_n1510_ | ~new_n11606_;
  assign new_n11772_ = ~new_n11687_;
  assign new_n11773_ = ~new_n11936_ | ~new_n11557_;
  assign new_n11774_ = ~new_n11773_ | ~new_n11569_;
  assign new_n11775_ = ~new_n11651_ | ~new_n11774_;
  assign new_n11776_ = ~new_n11760_ | ~new_n11558_;
  assign new_n11777_ = ~new_n1511_ | ~new_n11599_;
  assign new_n11778_ = ~new_n11652_ | ~new_n11776_;
  assign new_n11779_ = ~new_n11936_ | ~new_n11557_;
  assign new_n11780_ = ~new_n11927_ | ~new_n11561_;
  assign new_n11781_ = ~new_n11780_ | ~new_n11570_;
  assign new_n11782_ = ~new_n11653_ | ~new_n11781_;
  assign new_n11783_ = ~new_n11748_ | ~new_n11562_;
  assign new_n11784_ = ~new_n1515_ | ~new_n11602_;
  assign new_n11785_ = ~new_n11654_ | ~new_n11783_;
  assign new_n11786_ = ~new_n11927_ | ~new_n11561_;
  assign new_n11787_ = ~new_n11907_ | ~new_n11568_;
  assign new_n11788_ = ~new_n11991_ | ~new_n11578_;
  assign new_n11789_ = ~new_n11788_ | ~new_n11732_;
  assign new_n11790_ = ~new_n1508_ | ~new_n11613_;
  assign new_n11791_ = ~new_n11730_;
  assign new_n11792_ = ~new_n11994_ | ~new_n11582_;
  assign new_n11793_ = ~new_n11997_ | ~new_n11579_;
  assign new_n11794_ = ~new_n11738_ | ~new_n11546_;
  assign new_n11795_ = ~new_n1505_ | ~new_n11615_;
  assign new_n11796_ = ~new_n11656_ | ~new_n11794_;
  assign new_n11797_ = ~new_n12000_ | ~new_n11580_;
  assign new_n11798_ = ~new_n11994_ | ~new_n11582_;
  assign new_n11799_ = ~new_n11655_ | ~new_n11730_;
  assign new_n11800_ = ~new_n11798_ | ~new_n11796_;
  assign new_n11801_ = ~new_n11729_;
  assign new_n11802_ = ~new_n12003_ | ~new_n11583_;
  assign new_n11803_ = ~new_n11802_ | ~new_n11729_;
  assign new_n11804_ = ~new_n1504_ | ~new_n11617_;
  assign new_n11805_ = ~new_n11727_;
  assign new_n11806_ = ~new_n12006_ | ~new_n11584_;
  assign new_n11807_ = ~new_n11806_ | ~new_n11727_;
  assign new_n11808_ = ~new_n1503_ | ~new_n11618_;
  assign new_n11809_ = ~new_n11595_;
  assign new_n11810_ = ~new_n12009_ | ~new_n11577_;
  assign new_n11811_ = ~new_n12012_ | ~new_n11575_;
  assign new_n11812_ = ~new_n11576_;
  assign new_n11813_ = ~new_n11577_ | ~new_n11576_;
  assign new_n11814_ = ~new_n11612_ | ~new_n11813_;
  assign new_n11815_ = ~new_n1501_ | ~new_n11812_;
  assign new_n11816_ = ~new_n11547_ | ~new_n11595_;
  assign new_n11817_ = ~new_n11725_;
  assign new_n11818_ = ~new_n12015_ | ~new_n11585_;
  assign new_n11819_ = ~new_n11818_ | ~new_n11725_;
  assign new_n11820_ = ~new_n1500_ | ~new_n11619_;
  assign new_n11821_ = ~new_n11723_;
  assign new_n11822_ = ~new_n12018_ | ~new_n11589_;
  assign new_n11823_ = ~new_n12021_ | ~new_n11586_;
  assign new_n11824_ = ~new_n11739_ | ~new_n11548_;
  assign new_n11825_ = ~new_n1497_ | ~new_n11621_;
  assign new_n11826_ = ~new_n11659_ | ~new_n11824_;
  assign new_n11827_ = ~new_n12024_ | ~new_n11587_;
  assign new_n11828_ = ~new_n12018_ | ~new_n11589_;
  assign new_n11829_ = ~new_n11658_ | ~new_n11723_;
  assign new_n11830_ = ~new_n11828_ | ~new_n11826_;
  assign new_n11831_ = ~new_n11720_;
  assign new_n11832_ = ~new_n12027_ | ~new_n11590_;
  assign new_n11833_ = ~new_n11832_ | ~new_n11720_;
  assign new_n11834_ = ~new_n1496_ | ~new_n11623_;
  assign new_n11835_ = ~new_n11718_;
  assign new_n11836_ = ~new_n12030_ | ~new_n11591_;
  assign new_n11837_ = ~new_n11836_ | ~new_n11718_;
  assign new_n11838_ = ~new_n1495_ | ~new_n11624_;
  assign new_n11839_ = ~new_n11716_;
  assign new_n11840_ = ~new_n11982_ | ~new_n11573_;
  assign new_n11841_ = ~new_n11740_ | ~new_n11737_;
  assign new_n11842_ = ~new_n11592_;
  assign new_n11843_ = ~new_n11988_ | ~new_n11574_;
  assign new_n11844_ = ~new_n11733_ | ~new_n11716_ | ~new_n11843_;
  assign new_n11845_ = ~new_n11715_;
  assign new_n11846_ = ~new_n11979_ | ~new_n11571_;
  assign new_n11847_ = ~new_n1491_ | ~new_n11607_;
  assign new_n11848_ = ~new_n11979_ | ~new_n11571_;
  assign new_n11849_ = ~new_n11843_ | ~new_n11716_;
  assign new_n11850_ = ~new_n11593_;
  assign new_n11851_ = ~new_n11665_ | ~new_n11549_;
  assign new_n11852_ = ~new_n11666_ | ~new_n11849_;
  assign new_n11853_ = ~new_n1492_ | ~new_n11609_;
  assign new_n11854_ = ~new_n11667_ | ~new_n11852_;
  assign new_n11855_ = ~new_n11982_ | ~new_n11573_;
  assign new_n11856_ = ~new_n11827_ | ~new_n11723_;
  assign new_n11857_ = ~new_n11594_;
  assign new_n11858_ = ~new_n12021_ | ~new_n11586_;
  assign new_n11859_ = ~new_n11858_ | ~new_n11594_;
  assign new_n11860_ = ~new_n11669_ | ~new_n11859_;
  assign new_n11861_ = ~new_n11857_ | ~new_n11736_;
  assign new_n11862_ = ~new_n1497_ | ~new_n11621_;
  assign new_n11863_ = ~new_n11670_ | ~new_n11861_;
  assign new_n11864_ = ~new_n12021_ | ~new_n11586_;
  assign new_n11865_ = ~new_n12012_ | ~new_n11575_;
  assign new_n11866_ = ~new_n11865_ | ~new_n11595_;
  assign new_n11867_ = ~new_n11671_ | ~new_n11866_;
  assign new_n11868_ = ~new_n11809_ | ~new_n11576_;
  assign new_n11869_ = ~new_n1501_ | ~new_n11612_;
  assign new_n11870_ = ~new_n11672_ | ~new_n11868_;
  assign new_n11871_ = ~new_n12012_ | ~new_n11575_;
  assign new_n11872_ = ~new_n11797_ | ~new_n11730_;
  assign new_n11873_ = ~new_n11596_;
  assign new_n11874_ = ~new_n11997_ | ~new_n11579_;
  assign new_n11875_ = ~new_n11874_ | ~new_n11596_;
  assign new_n11876_ = ~new_n11673_ | ~new_n11875_;
  assign new_n11877_ = ~new_n11873_ | ~new_n11735_;
  assign new_n11878_ = ~new_n1505_ | ~new_n11615_;
  assign new_n11879_ = ~new_n11674_ | ~new_n11877_;
  assign new_n11880_ = ~new_n11997_ | ~new_n11579_;
  assign new_n11881_ = ~new_n11779_ | ~new_n11558_;
  assign new_n11882_ = ~new_n11786_ | ~new_n11562_;
  assign new_n11883_ = ~new_n11855_ | ~new_n11737_;
  assign new_n11884_ = ~new_n11843_ | ~new_n11740_;
  assign new_n11885_ = ~new_n11864_ | ~new_n11736_;
  assign new_n11886_ = ~new_n11827_ | ~new_n11588_;
  assign new_n11887_ = ~new_n11871_ | ~new_n11576_;
  assign new_n11888_ = ~new_n11880_ | ~new_n11735_;
  assign new_n11889_ = ~new_n11797_ | ~new_n11581_;
  assign new_n11890_ = ~new_n1514_ | ~new_n11600_;
  assign new_n11891_ = ~new_n11660_ | ~new_n11892_ | ~new_n11844_;
  assign new_n11892_ = ~new_n11841_ | ~new_n11733_;
  assign new_n11893_ = ~new_n1509_ | ~new_n11597_;
  assign new_n11894_ = ~new_n11609_ | ~new_n11840_;
  assign new_n11895_ = ~new_n1492_ | ~new_n11840_;
  assign new_n11896_ = ~new_n11848_ | ~new_n11841_ | ~new_n11733_;
  assign new_n11897_ = ~new_n11661_ | ~new_n11716_ | ~new_n11733_;
  assign new_n11898_ = ~new_n11842_ | ~new_n11848_;
  assign new_n11899_ = ~new_n1491_ | ~new_n11607_;
  assign new_n11900_ = ~new_n11668_ | ~new_n11850_;
  assign new_n11901_ = ~new_n11756_ | ~new_n11693_;
  assign new_n11902_ = ~new_n11691_;
  assign new_n11903_ = ~new_n11787_ | ~new_n11687_;
  assign new_n11904_ = ~new_n11732_;
  assign new_n11905_ = ~new_n1548_ | ~new_n11676_;
  assign new_n11906_ = ~new_n1538_ | ~new_n11556_;
  assign new_n11907_ = ~new_n11597_;
  assign new_n11908_ = ~new_n11907_ | ~new_n1509_;
  assign new_n11909_ = ~new_n11597_ | ~new_n11568_;
  assign new_n11910_ = ~new_n11907_ | ~new_n1509_;
  assign new_n11911_ = ~new_n11597_ | ~new_n11568_;
  assign new_n11912_ = ~new_n11911_ | ~new_n11910_;
  assign new_n11913_ = ~new_n1548_ | ~new_n11678_;
  assign new_n11914_ = ~new_n1543_ | ~new_n11556_;
  assign new_n11915_ = ~new_n11600_;
  assign new_n11916_ = ~new_n1548_ | ~new_n11679_;
  assign new_n11917_ = ~new_n1547_ | ~new_n11556_;
  assign new_n11918_ = ~new_n11603_;
  assign new_n11919_ = ~new_n1548_ | ~new_n11680_;
  assign new_n11920_ = ~new_n1546_ | ~new_n11556_;
  assign new_n11921_ = ~new_n11604_;
  assign new_n11922_ = ~new_n1548_ | ~new_n11681_;
  assign new_n11923_ = ~new_n1544_ | ~new_n11556_;
  assign new_n11924_ = ~new_n11602_;
  assign new_n11925_ = ~new_n1548_ | ~new_n11682_;
  assign new_n11926_ = ~new_n1545_ | ~new_n11556_;
  assign new_n11927_ = ~new_n11601_;
  assign new_n11928_ = ~new_n1548_ | ~new_n11683_;
  assign new_n11929_ = ~new_n1542_ | ~new_n11556_;
  assign new_n11930_ = ~new_n11605_;
  assign new_n11931_ = ~new_n1548_ | ~new_n11684_;
  assign new_n11932_ = ~new_n1540_ | ~new_n11556_;
  assign new_n11933_ = ~new_n11599_;
  assign new_n11934_ = ~new_n1548_ | ~new_n11685_;
  assign new_n11935_ = ~new_n1541_ | ~new_n11556_;
  assign new_n11936_ = ~new_n11598_;
  assign new_n11937_ = ~new_n1548_ | ~new_n11686_;
  assign new_n11938_ = ~new_n1539_ | ~new_n11556_;
  assign new_n11939_ = ~new_n11606_;
  assign new_n11940_ = ~new_n11677_ | ~new_n11687_;
  assign new_n11941_ = ~new_n11772_ | ~new_n11912_;
  assign new_n11942_ = ~new_n11939_ | ~new_n1510_;
  assign new_n11943_ = ~new_n11606_ | ~new_n11567_;
  assign new_n11944_ = ~new_n11939_ | ~new_n1510_;
  assign new_n11945_ = ~new_n11606_ | ~new_n11567_;
  assign new_n11946_ = ~new_n11945_ | ~new_n11944_;
  assign new_n11947_ = ~new_n11688_ | ~new_n11689_;
  assign new_n11948_ = ~new_n11768_ | ~new_n11946_;
  assign new_n11949_ = ~new_n11933_ | ~new_n1511_;
  assign new_n11950_ = ~new_n11599_ | ~new_n11559_;
  assign new_n11951_ = ~new_n11936_ | ~new_n1512_;
  assign new_n11952_ = ~new_n11598_ | ~new_n11557_;
  assign new_n11953_ = ~new_n11952_ | ~new_n11951_;
  assign new_n11954_ = ~new_n11881_ | ~new_n11569_;
  assign new_n11955_ = ~new_n11953_ | ~new_n11760_;
  assign new_n11956_ = ~new_n11930_ | ~new_n1513_;
  assign new_n11957_ = ~new_n11605_ | ~new_n11566_;
  assign new_n11958_ = ~new_n11930_ | ~new_n1513_;
  assign new_n11959_ = ~new_n11605_ | ~new_n11566_;
  assign new_n11960_ = ~new_n11959_ | ~new_n11958_;
  assign new_n11961_ = ~new_n11690_ | ~new_n11691_;
  assign new_n11962_ = ~new_n11902_ | ~new_n11960_;
  assign new_n11963_ = ~new_n11915_ | ~new_n1514_;
  assign new_n11964_ = ~new_n11600_ | ~new_n11560_;
  assign new_n11965_ = ~new_n11915_ | ~new_n1514_;
  assign new_n11966_ = ~new_n11600_ | ~new_n11560_;
  assign new_n11967_ = ~new_n11966_ | ~new_n11965_;
  assign new_n11968_ = ~new_n11692_ | ~new_n11693_;
  assign new_n11969_ = ~new_n11755_ | ~new_n11967_;
  assign new_n11970_ = ~new_n11924_ | ~new_n1515_;
  assign new_n11971_ = ~new_n11602_ | ~new_n11563_;
  assign new_n11972_ = ~new_n11927_ | ~new_n1516_;
  assign new_n11973_ = ~new_n11601_ | ~new_n11561_;
  assign new_n11974_ = ~new_n11973_ | ~new_n11972_;
  assign new_n11975_ = ~new_n11882_ | ~new_n11570_;
  assign new_n11976_ = ~new_n11974_ | ~new_n11748_;
  assign new_n11977_ = ~new_n1548_ | ~new_n11694_;
  assign new_n11978_ = ~new_n1520_ | ~new_n11556_;
  assign new_n11979_ = ~new_n11607_;
  assign new_n11980_ = ~new_n1548_ | ~new_n11695_;
  assign new_n11981_ = ~new_n1522_ | ~new_n11556_;
  assign new_n11982_ = ~new_n11608_;
  assign new_n11983_ = ~new_n1548_ | ~new_n11696_;
  assign new_n11984_ = ~new_n1521_ | ~new_n11556_;
  assign new_n11985_ = ~new_n11609_;
  assign new_n11986_ = ~new_n1548_ | ~new_n11697_;
  assign new_n11987_ = ~new_n1523_ | ~new_n11556_;
  assign new_n11988_ = ~new_n11610_;
  assign new_n11989_ = ~new_n1548_ | ~new_n11698_;
  assign new_n11990_ = ~new_n1537_ | ~new_n11556_;
  assign new_n11991_ = ~new_n11613_;
  assign new_n11992_ = ~new_n1548_ | ~new_n11699_;
  assign new_n11993_ = ~new_n1534_ | ~new_n11556_;
  assign new_n11994_ = ~new_n11615_;
  assign new_n11995_ = ~new_n1548_ | ~new_n11700_;
  assign new_n11996_ = ~new_n1535_ | ~new_n11556_;
  assign new_n11997_ = ~new_n11616_;
  assign new_n11998_ = ~new_n1548_ | ~new_n11701_;
  assign new_n11999_ = ~new_n1536_ | ~new_n11556_;
  assign new_n12000_ = ~new_n11614_;
  assign new_n12001_ = ~new_n1548_ | ~new_n11702_;
  assign new_n12002_ = ~new_n1533_ | ~new_n11556_;
  assign new_n12003_ = ~new_n11617_;
  assign new_n12004_ = ~new_n1548_ | ~new_n11703_;
  assign new_n12005_ = ~new_n1532_ | ~new_n11556_;
  assign new_n12006_ = ~new_n11618_;
  assign new_n12007_ = ~new_n1548_ | ~new_n11704_;
  assign new_n12008_ = ~new_n1530_ | ~new_n11556_;
  assign new_n12009_ = ~new_n11612_;
  assign new_n12010_ = ~new_n1548_ | ~new_n11705_;
  assign new_n12011_ = ~new_n1531_ | ~new_n11556_;
  assign new_n12012_ = ~new_n11611_;
  assign new_n12013_ = ~new_n1548_ | ~new_n11706_;
  assign new_n12014_ = ~new_n1529_ | ~new_n11556_;
  assign new_n12015_ = ~new_n11619_;
  assign new_n12016_ = ~new_n1548_ | ~new_n11707_;
  assign new_n12017_ = ~new_n1526_ | ~new_n11556_;
  assign new_n12018_ = ~new_n11621_;
  assign new_n12019_ = ~new_n1548_ | ~new_n11708_;
  assign new_n12020_ = ~new_n1527_ | ~new_n11556_;
  assign new_n12021_ = ~new_n11622_;
  assign new_n12022_ = ~new_n1548_ | ~new_n11709_;
  assign new_n12023_ = ~new_n1528_ | ~new_n11556_;
  assign new_n12024_ = ~new_n11620_;
  assign new_n12025_ = ~new_n1548_ | ~new_n11710_;
  assign new_n12026_ = ~new_n1525_ | ~new_n11556_;
  assign new_n12027_ = ~new_n11623_;
  assign new_n12028_ = ~new_n1548_ | ~new_n11711_;
  assign new_n12029_ = ~new_n1524_ | ~new_n11556_;
  assign new_n12030_ = ~new_n11624_;
  assign new_n12031_ = ~new_n1548_ | ~new_n11712_;
  assign new_n12032_ = ~new_n1490_ | ~new_n11556_;
  assign new_n12033_ = ~new_n11663_;
  assign new_n12034_ = ~new_n1519_ | ~new_n12033_;
  assign new_n12035_ = ~new_n11663_ | ~new_n11713_;
  assign new_n12036_ = ~new_n11625_;
  assign new_n12037_ = ~new_n12036_ | ~new_n11891_ | ~new_n11846_;
  assign new_n12038_ = ~new_n11625_ | ~new_n11662_ | ~new_n11898_ | ~new_n11897_;
  assign new_n12039_ = ~new_n11979_ | ~new_n1491_;
  assign new_n12040_ = ~new_n11607_ | ~new_n11571_;
  assign new_n12041_ = ~new_n11979_ | ~new_n1491_;
  assign new_n12042_ = ~new_n11607_ | ~new_n11571_;
  assign new_n12043_ = ~new_n12042_ | ~new_n12041_;
  assign new_n12044_ = ~new_n11714_ | ~new_n11715_;
  assign new_n12045_ = ~new_n11845_ | ~new_n12043_;
  assign new_n12046_ = ~new_n11985_ | ~new_n1492_;
  assign new_n12047_ = ~new_n11609_ | ~new_n11572_;
  assign new_n12048_ = ~new_n11982_ | ~new_n1493_;
  assign new_n12049_ = ~new_n11608_ | ~new_n11573_;
  assign new_n12050_ = ~new_n12049_ | ~new_n12048_;
  assign new_n12051_ = ~new_n11883_ | ~new_n11593_;
  assign new_n12052_ = ~new_n12050_ | ~new_n11850_;
  assign new_n12053_ = ~new_n11988_ | ~new_n1494_;
  assign new_n12054_ = ~new_n11610_ | ~new_n11574_;
  assign new_n12055_ = ~new_n12054_ | ~new_n12053_;
  assign new_n12056_ = ~new_n11884_ | ~new_n11716_;
  assign new_n12057_ = ~new_n11839_ | ~new_n12055_;
  assign new_n12058_ = ~new_n12030_ | ~new_n1495_;
  assign new_n12059_ = ~new_n11624_ | ~new_n11591_;
  assign new_n12060_ = ~new_n12030_ | ~new_n1495_;
  assign new_n12061_ = ~new_n11624_ | ~new_n11591_;
  assign new_n12062_ = ~new_n12061_ | ~new_n12060_;
  assign new_n12063_ = ~new_n11717_ | ~new_n11718_;
  assign new_n12064_ = ~new_n11835_ | ~new_n12062_;
  assign new_n12065_ = ~new_n12027_ | ~new_n1496_;
  assign new_n12066_ = ~new_n11623_ | ~new_n11590_;
  assign new_n12067_ = ~new_n12027_ | ~new_n1496_;
  assign new_n12068_ = ~new_n11623_ | ~new_n11590_;
  assign new_n12069_ = ~new_n12068_ | ~new_n12067_;
  assign new_n12070_ = ~new_n11719_ | ~new_n11720_;
  assign new_n12071_ = ~new_n11831_ | ~new_n12069_;
  assign new_n12072_ = ~new_n12018_ | ~new_n1497_;
  assign new_n12073_ = ~new_n11621_ | ~new_n11589_;
  assign new_n12074_ = ~new_n12021_ | ~new_n1498_;
  assign new_n12075_ = ~new_n11622_ | ~new_n11586_;
  assign new_n12076_ = ~new_n12075_ | ~new_n12074_;
  assign new_n12077_ = ~new_n11885_ | ~new_n11594_;
  assign new_n12078_ = ~new_n12076_ | ~new_n11857_;
  assign new_n12079_ = ~new_n11921_ | ~new_n1517_;
  assign new_n12080_ = ~new_n11604_ | ~new_n11565_;
  assign new_n12081_ = ~new_n11921_ | ~new_n1517_;
  assign new_n12082_ = ~new_n11604_ | ~new_n11565_;
  assign new_n12083_ = ~new_n12082_ | ~new_n12081_;
  assign new_n12084_ = ~new_n11721_ | ~new_n11722_;
  assign new_n12085_ = ~new_n11744_ | ~new_n12083_;
  assign new_n12086_ = ~new_n12024_ | ~new_n1499_;
  assign new_n12087_ = ~new_n11620_ | ~new_n11587_;
  assign new_n12088_ = ~new_n12087_ | ~new_n12086_;
  assign new_n12089_ = ~new_n11886_ | ~new_n11723_;
  assign new_n12090_ = ~new_n11821_ | ~new_n12088_;
  assign new_n12091_ = ~new_n12015_ | ~new_n1500_;
  assign new_n12092_ = ~new_n11619_ | ~new_n11585_;
  assign new_n12093_ = ~new_n12015_ | ~new_n1500_;
  assign new_n12094_ = ~new_n11619_ | ~new_n11585_;
  assign new_n12095_ = ~new_n12094_ | ~new_n12093_;
  assign new_n12096_ = ~new_n11724_ | ~new_n11725_;
  assign new_n12097_ = ~new_n11817_ | ~new_n12095_;
  assign new_n12098_ = ~new_n12009_ | ~new_n1501_;
  assign new_n12099_ = ~new_n11612_ | ~new_n11577_;
  assign new_n12100_ = ~new_n12012_ | ~new_n1502_;
  assign new_n12101_ = ~new_n11611_ | ~new_n11575_;
  assign new_n12102_ = ~new_n12101_ | ~new_n12100_;
  assign new_n12103_ = ~new_n11887_ | ~new_n11595_;
  assign new_n12104_ = ~new_n12102_ | ~new_n11809_;
  assign new_n12105_ = ~new_n12006_ | ~new_n1503_;
  assign new_n12106_ = ~new_n11618_ | ~new_n11584_;
  assign new_n12107_ = ~new_n12006_ | ~new_n1503_;
  assign new_n12108_ = ~new_n11618_ | ~new_n11584_;
  assign new_n12109_ = ~new_n12108_ | ~new_n12107_;
  assign new_n12110_ = ~new_n11726_ | ~new_n11727_;
  assign new_n12111_ = ~new_n11805_ | ~new_n12109_;
  assign new_n12112_ = ~new_n12003_ | ~new_n1504_;
  assign new_n12113_ = ~new_n11617_ | ~new_n11583_;
  assign new_n12114_ = ~new_n12003_ | ~new_n1504_;
  assign new_n12115_ = ~new_n11617_ | ~new_n11583_;
  assign new_n12116_ = ~new_n12115_ | ~new_n12114_;
  assign new_n12117_ = ~new_n11728_ | ~new_n11729_;
  assign new_n12118_ = ~new_n11801_ | ~new_n12116_;
  assign new_n12119_ = ~new_n11994_ | ~new_n1505_;
  assign new_n12120_ = ~new_n11615_ | ~new_n11582_;
  assign new_n12121_ = ~new_n11997_ | ~new_n1506_;
  assign new_n12122_ = ~new_n11616_ | ~new_n11579_;
  assign new_n12123_ = ~new_n12122_ | ~new_n12121_;
  assign new_n12124_ = ~new_n11888_ | ~new_n11596_;
  assign new_n12125_ = ~new_n12123_ | ~new_n11873_;
  assign new_n12126_ = ~new_n12000_ | ~new_n1507_;
  assign new_n12127_ = ~new_n11614_ | ~new_n11580_;
  assign new_n12128_ = ~new_n12127_ | ~new_n12126_;
  assign new_n12129_ = ~new_n11889_ | ~new_n11730_;
  assign new_n12130_ = ~new_n11791_ | ~new_n12128_;
  assign new_n12131_ = ~new_n11991_ | ~new_n1508_;
  assign new_n12132_ = ~new_n11613_ | ~new_n11578_;
  assign new_n12133_ = ~new_n11991_ | ~new_n1508_;
  assign new_n12134_ = ~new_n11613_ | ~new_n11578_;
  assign new_n12135_ = ~new_n12134_ | ~new_n12133_;
  assign new_n12136_ = ~new_n11731_ | ~new_n11732_;
  assign new_n12137_ = ~new_n11904_ | ~new_n12135_;
  assign new_n12138_ = ~new_n1518_ | ~new_n11556_;
  assign new_n12139_ = ~new_n1548_ | ~new_n11564_;
  assign new_n12140_ = ~new_n11675_;
  assign new_n12141_ = ~new_n11603_ | ~new_n12140_;
  assign new_n12142_ = ~new_n11675_ | ~new_n11918_;
  assign new_n12143_ = new_n12321_ & new_n12338_;
  assign new_n12144_ = new_n12340_ & new_n12339_;
  assign new_n12145_ = new_n12316_ & new_n12377_;
  assign new_n12146_ = new_n12379_ & new_n12378_;
  assign new_n12147_ = new_n12396_ & new_n12395_;
  assign new_n12148_ = new_n12422_ & new_n12421_;
  assign new_n12149_ = new_n12520_ & new_n12519_;
  assign new_n12150_ = ~new_n12477_ | ~new_n12480_;
  assign new_n12151_ = ~new_n12466_ | ~new_n12469_;
  assign new_n12152_ = ~new_n12455_ | ~new_n12458_;
  assign new_n12153_ = ~new_n12447_ | ~new_n12449_;
  assign new_n12154_ = ~new_n12485_ | ~new_n12293_ | ~new_n12312_;
  assign new_n12155_ = ~new_n12373_ | ~new_n12375_;
  assign new_n12156_ = ~new_n12365_ | ~new_n12368_;
  assign new_n12157_ = ~new_n12357_ | ~new_n12359_;
  assign new_n12158_ = ~new_n12162_ | ~new_n12483_;
  assign new_n12159_ = ~new_n1813_;
  assign new_n12160_ = ~new_n1798_;
  assign new_n12161_ = ~new_n1790_;
  assign new_n12162_ = ~new_n1790_ | ~new_n12230_;
  assign new_n12163_ = ~new_n1415_;
  assign new_n12164_ = ~new_n1801_;
  assign new_n12165_ = ~new_n1405_;
  assign new_n12166_ = ~new_n1405_ | ~new_n12160_;
  assign new_n12167_ = ~new_n1401_;
  assign new_n12168_ = ~new_n1810_;
  assign new_n12169_ = ~new_n1807_;
  assign new_n12170_ = ~new_n1804_;
  assign new_n12171_ = ~new_n1408_;
  assign new_n12172_ = ~new_n1404_;
  assign new_n12173_ = ~new_n1397_;
  assign new_n12174_ = ~new_n1397_ | ~new_n12170_;
  assign new_n12175_ = ~new_n1816_;
  assign new_n12176_ = ~new_n1407_;
  assign new_n12177_ = ~new_n1407_ | ~new_n12159_;
  assign new_n12178_ = ~new_n1421_;
  assign new_n12179_ = ~new_n1819_;
  assign new_n12180_ = ~new_n1420_;
  assign new_n12181_ = ~new_n12346_ | ~new_n12345_;
  assign new_n12182_ = ~new_n12174_ | ~new_n12361_;
  assign new_n12183_ = ~new_n12330_ | ~new_n12329_;
  assign new_n12184_ = ~new_n2348_;
  assign new_n12185_ = ~new_n2352_;
  assign new_n12186_ = ~new_n1837_;
  assign new_n12187_ = ~new_n1825_;
  assign new_n12188_ = ~new_n1822_;
  assign new_n12189_ = ~new_n1400_;
  assign new_n12190_ = ~new_n1399_;
  assign new_n12191_ = ~new_n1420_ | ~new_n12179_;
  assign new_n12192_ = ~new_n1828_;
  assign new_n12193_ = ~new_n1409_;
  assign new_n12194_ = ~new_n1831_;
  assign new_n12195_ = ~new_n1417_;
  assign new_n12196_ = ~new_n1840_;
  assign new_n12197_ = ~new_n1834_;
  assign new_n12198_ = ~new_n1410_;
  assign new_n12199_ = ~new_n1411_;
  assign new_n12200_ = ~new_n1416_;
  assign new_n12201_ = ~new_n1416_ | ~new_n12197_;
  assign new_n12202_ = ~new_n1843_;
  assign new_n12203_ = ~new_n1406_;
  assign new_n12204_ = ~new_n12406_ | ~new_n12405_;
  assign new_n12205_ = ~new_n1419_;
  assign new_n12206_ = ~new_n1848_;
  assign new_n12207_ = ~new_n1418_;
  assign new_n12208_ = ~new_n2354_;
  assign new_n12209_ = ~new_n1413_;
  assign new_n12210_ = ~new_n2351_;
  assign new_n12211_ = ~new_n2353_;
  assign new_n12212_ = ~new_n1403_;
  assign new_n12213_ = ~new_n1398_;
  assign new_n12214_ = ~new_n1412_;
  assign new_n12215_ = ~new_n1412_ | ~new_n12211_;
  assign new_n12216_ = ~new_n2350_;
  assign new_n12217_ = ~new_n1402_;
  assign new_n12218_ = ~new_n2349_;
  assign new_n12219_ = ~new_n1395_;
  assign new_n12220_ = ~new_n2347_;
  assign new_n12221_ = ~new_n1394_;
  assign new_n12222_ = ~new_n1394_ | ~new_n12184_;
  assign new_n12223_ = ~new_n1390_;
  assign new_n12224_ = ~new_n2346_;
  assign new_n12225_ = ~new_n1391_;
  assign new_n12226_ = ~new_n12436_ | ~new_n12435_;
  assign new_n12227_ = ~new_n12215_ | ~new_n12451_;
  assign new_n12228_ = ~new_n12201_ | ~new_n12462_;
  assign new_n12229_ = ~new_n12191_ | ~new_n12473_;
  assign new_n12230_ = ~new_n1414_;
  assign new_n12231_ = ~new_n12530_ | ~new_n12529_;
  assign new_n12232_ = ~new_n12544_ | ~new_n12543_;
  assign new_n12233_ = ~new_n12549_ | ~new_n12548_;
  assign new_n12234_ = ~new_n12565_ | ~new_n12564_;
  assign new_n12235_ = ~new_n12570_ | ~new_n12569_;
  assign new_n12236_ = ~new_n12575_ | ~new_n12574_;
  assign new_n12237_ = ~new_n12580_ | ~new_n12579_;
  assign new_n12238_ = ~new_n12585_ | ~new_n12584_;
  assign new_n12239_ = ~new_n12601_ | ~new_n12600_;
  assign new_n12240_ = ~new_n12606_ | ~new_n12605_;
  assign new_n12241_ = ~new_n12489_ | ~new_n12488_;
  assign new_n12242_ = ~new_n12498_ | ~new_n12497_;
  assign new_n12243_ = ~new_n12505_ | ~new_n12504_;
  assign new_n12244_ = ~new_n12509_ | ~new_n12508_;
  assign new_n12245_ = ~new_n12518_ | ~new_n12517_;
  assign new_n12246_ = ~new_n12539_ | ~new_n12538_;
  assign new_n12247_ = ~new_n12556_ | ~new_n12555_;
  assign new_n12248_ = ~new_n12560_ | ~new_n12559_;
  assign new_n12249_ = ~new_n12592_ | ~new_n12591_;
  assign new_n12250_ = ~new_n12596_ | ~new_n12595_;
  assign new_n12251_ = ~new_n12613_ | ~new_n12612_;
  assign new_n12252_ = new_n12332_ & new_n12320_;
  assign new_n12253_ = new_n12335_ & new_n12336_;
  assign new_n12254_ = new_n12348_ & new_n12322_;
  assign new_n12255_ = new_n12351_ & new_n12352_;
  assign new_n12256_ = new_n12177_ & new_n12491_ & new_n12490_;
  assign new_n12257_ = new_n12494_ & new_n12322_;
  assign new_n12258_ = new_n12367_ & new_n12144_;
  assign new_n12259_ = new_n12501_ & new_n12321_;
  assign new_n12260_ = new_n12166_ & new_n12511_ & new_n12510_;
  assign new_n12261_ = new_n12514_ & new_n12320_;
  assign new_n12262_ = new_n12354_ & new_n12145_;
  assign new_n12263_ = new_n12399_ & new_n12317_;
  assign new_n12264_ = new_n12425_ & new_n12318_;
  assign new_n12265_ = new_n12441_ & new_n12442_;
  assign new_n12266_ = new_n12444_ & new_n12523_;
  assign new_n12267_ = new_n12445_ & new_n12442_ & new_n12441_;
  assign new_n12268_ = ~new_n12527_ | ~new_n12526_;
  assign new_n12269_ = new_n12222_ & new_n12532_ & new_n12531_;
  assign new_n12270_ = new_n12535_ & new_n12319_;
  assign new_n12271_ = ~new_n12541_ | ~new_n12540_;
  assign new_n12272_ = ~new_n12546_ | ~new_n12545_;
  assign new_n12273_ = new_n12552_ & new_n12318_;
  assign new_n12274_ = ~new_n12562_ | ~new_n12561_;
  assign new_n12275_ = ~new_n12567_ | ~new_n12566_;
  assign new_n12276_ = ~new_n12572_ | ~new_n12571_;
  assign new_n12277_ = ~new_n12577_ | ~new_n12576_;
  assign new_n12278_ = ~new_n12582_ | ~new_n12581_;
  assign new_n12279_ = new_n12588_ & new_n12317_;
  assign new_n12280_ = ~new_n12598_ | ~new_n12597_;
  assign new_n12281_ = ~new_n12603_ | ~new_n12602_;
  assign new_n12282_ = new_n12479_ & new_n12146_;
  assign new_n12283_ = new_n12609_ & new_n12316_;
  assign new_n12284_ = new_n12487_ & new_n12486_;
  assign new_n12285_ = ~new_n12255_ | ~new_n12349_;
  assign new_n12286_ = new_n12496_ & new_n12495_;
  assign new_n12287_ = new_n12503_ & new_n12502_;
  assign new_n12288_ = new_n12507_ & new_n12506_;
  assign new_n12289_ = ~new_n12253_ | ~new_n12333_;
  assign new_n12290_ = new_n12516_ & new_n12515_;
  assign new_n12291_ = ~new_n2357_;
  assign new_n12292_ = ~new_n1392_;
  assign new_n12293_ = new_n12525_ & new_n12524_;
  assign new_n12294_ = ~new_n12265_ | ~new_n12439_;
  assign new_n12295_ = new_n12537_ & new_n12536_;
  assign new_n12296_ = ~new_n12432_ | ~new_n12431_;
  assign new_n12297_ = ~new_n12428_ | ~new_n12427_;
  assign new_n12298_ = new_n12554_ & new_n12553_;
  assign new_n12299_ = new_n12558_ & new_n12557_;
  assign new_n12300_ = ~new_n12418_ | ~new_n12417_;
  assign new_n12301_ = ~new_n12414_ | ~new_n12413_;
  assign new_n12302_ = ~new_n1795_;
  assign new_n12303_ = ~new_n12410_ | ~new_n12409_;
  assign new_n12304_ = ~new_n1846_;
  assign new_n12305_ = ~new_n12402_ | ~new_n12401_;
  assign new_n12306_ = new_n12590_ & new_n12589_;
  assign new_n12307_ = new_n12594_ & new_n12593_;
  assign new_n12308_ = ~new_n12392_ | ~new_n12391_;
  assign new_n12309_ = ~new_n12388_ | ~new_n12387_;
  assign new_n12310_ = ~new_n12384_ | ~new_n12383_;
  assign new_n12311_ = new_n12611_ & new_n12610_;
  assign new_n12312_ = ~new_n12266_ | ~new_n12294_;
  assign new_n12313_ = ~new_n12222_;
  assign new_n12314_ = ~new_n12166_;
  assign new_n12315_ = ~new_n12177_;
  assign new_n12316_ = ~new_n1822_ | ~new_n12190_;
  assign new_n12317_ = ~new_n1837_ | ~new_n12199_;
  assign new_n12318_ = ~new_n2352_ | ~new_n12213_;
  assign new_n12319_ = ~new_n2348_ | ~new_n12221_;
  assign new_n12320_ = ~new_n1798_ | ~new_n12165_;
  assign new_n12321_ = ~new_n1807_ | ~new_n12172_;
  assign new_n12322_ = ~new_n1813_ | ~new_n12176_;
  assign new_n12323_ = ~new_n12201_;
  assign new_n12324_ = ~new_n12215_;
  assign new_n12325_ = ~new_n12174_;
  assign new_n12326_ = ~new_n12191_;
  assign new_n12327_ = ~new_n12162_;
  assign new_n12328_ = ~new_n12327_ | ~new_n12163_;
  assign new_n12329_ = ~new_n12328_ | ~new_n12302_;
  assign new_n12330_ = ~new_n1415_ | ~new_n12162_;
  assign new_n12331_ = ~new_n12183_;
  assign new_n12332_ = ~new_n1801_ | ~new_n12167_;
  assign new_n12333_ = ~new_n12252_ | ~new_n12183_;
  assign new_n12334_ = ~new_n12167_ | ~new_n12166_;
  assign new_n12335_ = ~new_n12334_ | ~new_n12164_;
  assign new_n12336_ = ~new_n1401_ | ~new_n12314_;
  assign new_n12337_ = ~new_n12289_;
  assign new_n12338_ = ~new_n1810_ | ~new_n12171_;
  assign new_n12339_ = ~new_n1408_ | ~new_n12168_;
  assign new_n12340_ = ~new_n1404_ | ~new_n12169_;
  assign new_n12341_ = ~new_n12325_ | ~new_n12143_;
  assign new_n12342_ = ~new_n12144_ | ~new_n12341_;
  assign new_n12343_ = ~new_n1804_ | ~new_n12173_;
  assign new_n12344_ = ~new_n1810_ | ~new_n12171_;
  assign new_n12345_ = ~new_n12143_ | ~new_n12343_ | ~new_n12289_;
  assign new_n12346_ = ~new_n12344_ | ~new_n12342_;
  assign new_n12347_ = ~new_n12181_;
  assign new_n12348_ = ~new_n1816_ | ~new_n12178_;
  assign new_n12349_ = ~new_n12254_ | ~new_n12181_;
  assign new_n12350_ = ~new_n12178_ | ~new_n12177_;
  assign new_n12351_ = ~new_n12350_ | ~new_n12175_;
  assign new_n12352_ = ~new_n1421_ | ~new_n12315_;
  assign new_n12353_ = ~new_n12285_;
  assign new_n12354_ = ~new_n1819_ | ~new_n12180_;
  assign new_n12355_ = ~new_n12354_ | ~new_n12191_;
  assign new_n12356_ = ~new_n12347_ | ~new_n12177_;
  assign new_n12357_ = ~new_n12257_ | ~new_n12356_;
  assign new_n12358_ = ~new_n12181_ | ~new_n12322_;
  assign new_n12359_ = ~new_n12256_ | ~new_n12358_;
  assign new_n12360_ = ~new_n12177_ | ~new_n12322_;
  assign new_n12361_ = ~new_n12343_ | ~new_n12289_;
  assign new_n12362_ = ~new_n12182_;
  assign new_n12363_ = ~new_n1404_ | ~new_n12169_;
  assign new_n12364_ = ~new_n12362_ | ~new_n12363_;
  assign new_n12365_ = ~new_n12259_ | ~new_n12364_;
  assign new_n12366_ = ~new_n12182_ | ~new_n12321_;
  assign new_n12367_ = ~new_n1810_ | ~new_n12171_;
  assign new_n12368_ = ~new_n12258_ | ~new_n12366_;
  assign new_n12369_ = ~new_n1404_ | ~new_n12169_;
  assign new_n12370_ = ~new_n12321_ | ~new_n12369_;
  assign new_n12371_ = ~new_n12343_ | ~new_n12174_;
  assign new_n12372_ = ~new_n12331_ | ~new_n12166_;
  assign new_n12373_ = ~new_n12261_ | ~new_n12372_;
  assign new_n12374_ = ~new_n12183_ | ~new_n12320_;
  assign new_n12375_ = ~new_n12260_ | ~new_n12374_;
  assign new_n12376_ = ~new_n12166_ | ~new_n12320_;
  assign new_n12377_ = ~new_n1825_ | ~new_n12189_;
  assign new_n12378_ = ~new_n1400_ | ~new_n12187_;
  assign new_n12379_ = ~new_n1399_ | ~new_n12188_;
  assign new_n12380_ = ~new_n12326_ | ~new_n12145_;
  assign new_n12381_ = ~new_n12146_ | ~new_n12380_;
  assign new_n12382_ = ~new_n1825_ | ~new_n12189_;
  assign new_n12383_ = ~new_n12262_ | ~new_n12285_;
  assign new_n12384_ = ~new_n12382_ | ~new_n12381_;
  assign new_n12385_ = ~new_n12310_;
  assign new_n12386_ = ~new_n1828_ | ~new_n12193_;
  assign new_n12387_ = ~new_n12386_ | ~new_n12310_;
  assign new_n12388_ = ~new_n1409_ | ~new_n12192_;
  assign new_n12389_ = ~new_n12309_;
  assign new_n12390_ = ~new_n1831_ | ~new_n12195_;
  assign new_n12391_ = ~new_n12390_ | ~new_n12309_;
  assign new_n12392_ = ~new_n1417_ | ~new_n12194_;
  assign new_n12393_ = ~new_n12308_;
  assign new_n12394_ = ~new_n1840_ | ~new_n12198_;
  assign new_n12395_ = ~new_n1410_ | ~new_n12196_;
  assign new_n12396_ = ~new_n1411_ | ~new_n12186_;
  assign new_n12397_ = ~new_n12323_ | ~new_n12317_;
  assign new_n12398_ = ~new_n12147_ | ~new_n12397_;
  assign new_n12399_ = ~new_n1834_ | ~new_n12200_;
  assign new_n12400_ = ~new_n1840_ | ~new_n12198_;
  assign new_n12401_ = ~new_n12394_ | ~new_n12308_ | ~new_n12263_;
  assign new_n12402_ = ~new_n12400_ | ~new_n12398_;
  assign new_n12403_ = ~new_n12305_;
  assign new_n12404_ = ~new_n1843_ | ~new_n12203_;
  assign new_n12405_ = ~new_n12404_ | ~new_n12305_;
  assign new_n12406_ = ~new_n1406_ | ~new_n12202_;
  assign new_n12407_ = ~new_n12204_;
  assign new_n12408_ = ~new_n12407_ | ~new_n12205_;
  assign new_n12409_ = ~new_n12408_ | ~new_n12304_;
  assign new_n12410_ = ~new_n1419_ | ~new_n12204_;
  assign new_n12411_ = ~new_n12303_;
  assign new_n12412_ = ~new_n1848_ | ~new_n12207_;
  assign new_n12413_ = ~new_n12412_ | ~new_n12303_;
  assign new_n12414_ = ~new_n1418_ | ~new_n12206_;
  assign new_n12415_ = ~new_n12301_;
  assign new_n12416_ = ~new_n2354_ | ~new_n12209_;
  assign new_n12417_ = ~new_n12416_ | ~new_n12301_;
  assign new_n12418_ = ~new_n1413_ | ~new_n12208_;
  assign new_n12419_ = ~new_n12300_;
  assign new_n12420_ = ~new_n2351_ | ~new_n12212_;
  assign new_n12421_ = ~new_n1403_ | ~new_n12210_;
  assign new_n12422_ = ~new_n1398_ | ~new_n12185_;
  assign new_n12423_ = ~new_n12324_ | ~new_n12318_;
  assign new_n12424_ = ~new_n12148_ | ~new_n12423_;
  assign new_n12425_ = ~new_n2353_ | ~new_n12214_;
  assign new_n12426_ = ~new_n2351_ | ~new_n12212_;
  assign new_n12427_ = ~new_n12420_ | ~new_n12300_ | ~new_n12264_;
  assign new_n12428_ = ~new_n12426_ | ~new_n12424_;
  assign new_n12429_ = ~new_n12297_;
  assign new_n12430_ = ~new_n2350_ | ~new_n12217_;
  assign new_n12431_ = ~new_n12430_ | ~new_n12297_;
  assign new_n12432_ = ~new_n1402_ | ~new_n12216_;
  assign new_n12433_ = ~new_n12296_;
  assign new_n12434_ = ~new_n2349_ | ~new_n12219_;
  assign new_n12435_ = ~new_n12434_ | ~new_n12296_;
  assign new_n12436_ = ~new_n1395_ | ~new_n12218_;
  assign new_n12437_ = ~new_n12226_;
  assign new_n12438_ = ~new_n2347_ | ~new_n12223_;
  assign new_n12439_ = ~new_n12438_ | ~new_n12226_ | ~new_n12319_;
  assign new_n12440_ = ~new_n12223_ | ~new_n12222_;
  assign new_n12441_ = ~new_n12440_ | ~new_n12220_;
  assign new_n12442_ = ~new_n1390_ | ~new_n12313_;
  assign new_n12443_ = ~new_n12294_;
  assign new_n12444_ = ~new_n2346_ | ~new_n12225_;
  assign new_n12445_ = ~new_n1391_ | ~new_n12224_;
  assign new_n12446_ = ~new_n12437_ | ~new_n12222_;
  assign new_n12447_ = ~new_n12270_ | ~new_n12446_;
  assign new_n12448_ = ~new_n12226_ | ~new_n12319_;
  assign new_n12449_ = ~new_n12269_ | ~new_n12448_;
  assign new_n12450_ = ~new_n12222_ | ~new_n12319_;
  assign new_n12451_ = ~new_n12425_ | ~new_n12300_;
  assign new_n12452_ = ~new_n12227_;
  assign new_n12453_ = ~new_n1398_ | ~new_n12185_;
  assign new_n12454_ = ~new_n12452_ | ~new_n12453_;
  assign new_n12455_ = ~new_n12273_ | ~new_n12454_;
  assign new_n12456_ = ~new_n12227_ | ~new_n12318_;
  assign new_n12457_ = ~new_n2351_ | ~new_n12212_;
  assign new_n12458_ = ~new_n12148_ | ~new_n12457_ | ~new_n12456_;
  assign new_n12459_ = ~new_n1398_ | ~new_n12185_;
  assign new_n12460_ = ~new_n12318_ | ~new_n12459_;
  assign new_n12461_ = ~new_n12425_ | ~new_n12215_;
  assign new_n12462_ = ~new_n12399_ | ~new_n12308_;
  assign new_n12463_ = ~new_n12228_;
  assign new_n12464_ = ~new_n1411_ | ~new_n12186_;
  assign new_n12465_ = ~new_n12463_ | ~new_n12464_;
  assign new_n12466_ = ~new_n12279_ | ~new_n12465_;
  assign new_n12467_ = ~new_n12228_ | ~new_n12317_;
  assign new_n12468_ = ~new_n1840_ | ~new_n12198_;
  assign new_n12469_ = ~new_n12147_ | ~new_n12468_ | ~new_n12467_;
  assign new_n12470_ = ~new_n1411_ | ~new_n12186_;
  assign new_n12471_ = ~new_n12317_ | ~new_n12470_;
  assign new_n12472_ = ~new_n12399_ | ~new_n12201_;
  assign new_n12473_ = ~new_n12354_ | ~new_n12285_;
  assign new_n12474_ = ~new_n12229_;
  assign new_n12475_ = ~new_n1399_ | ~new_n12188_;
  assign new_n12476_ = ~new_n12474_ | ~new_n12475_;
  assign new_n12477_ = ~new_n12283_ | ~new_n12476_;
  assign new_n12478_ = ~new_n12229_ | ~new_n12316_;
  assign new_n12479_ = ~new_n1825_ | ~new_n12189_;
  assign new_n12480_ = ~new_n12282_ | ~new_n12478_;
  assign new_n12481_ = ~new_n1399_ | ~new_n12188_;
  assign new_n12482_ = ~new_n12316_ | ~new_n12481_;
  assign new_n12483_ = ~new_n1414_ | ~new_n12161_;
  assign new_n12484_ = ~new_n12438_ | ~new_n12226_ | ~new_n12319_;
  assign new_n12485_ = ~new_n12267_ | ~new_n12149_ | ~new_n12484_;
  assign new_n12486_ = ~new_n1819_ | ~new_n12180_;
  assign new_n12487_ = ~new_n1420_ | ~new_n12179_;
  assign new_n12488_ = ~new_n12355_ | ~new_n12285_;
  assign new_n12489_ = ~new_n12353_ | ~new_n12284_;
  assign new_n12490_ = ~new_n1816_ | ~new_n12178_;
  assign new_n12491_ = ~new_n1421_ | ~new_n12175_;
  assign new_n12492_ = ~new_n1816_ | ~new_n12178_;
  assign new_n12493_ = ~new_n1421_ | ~new_n12175_;
  assign new_n12494_ = ~new_n12493_ | ~new_n12492_;
  assign new_n12495_ = ~new_n1813_ | ~new_n12176_;
  assign new_n12496_ = ~new_n1407_ | ~new_n12159_;
  assign new_n12497_ = ~new_n12360_ | ~new_n12181_;
  assign new_n12498_ = ~new_n12286_ | ~new_n12347_;
  assign new_n12499_ = ~new_n1810_ | ~new_n12171_;
  assign new_n12500_ = ~new_n1408_ | ~new_n12168_;
  assign new_n12501_ = ~new_n12500_ | ~new_n12499_;
  assign new_n12502_ = ~new_n1807_ | ~new_n12172_;
  assign new_n12503_ = ~new_n1404_ | ~new_n12169_;
  assign new_n12504_ = ~new_n12370_ | ~new_n12182_;
  assign new_n12505_ = ~new_n12287_ | ~new_n12362_;
  assign new_n12506_ = ~new_n1804_ | ~new_n12173_;
  assign new_n12507_ = ~new_n1397_ | ~new_n12170_;
  assign new_n12508_ = ~new_n12371_ | ~new_n12289_;
  assign new_n12509_ = ~new_n12337_ | ~new_n12288_;
  assign new_n12510_ = ~new_n1801_ | ~new_n12167_;
  assign new_n12511_ = ~new_n1401_ | ~new_n12164_;
  assign new_n12512_ = ~new_n1801_ | ~new_n12167_;
  assign new_n12513_ = ~new_n1401_ | ~new_n12164_;
  assign new_n12514_ = ~new_n12513_ | ~new_n12512_;
  assign new_n12515_ = ~new_n1798_ | ~new_n12165_;
  assign new_n12516_ = ~new_n1405_ | ~new_n12160_;
  assign new_n12517_ = ~new_n12376_ | ~new_n12183_;
  assign new_n12518_ = ~new_n12290_ | ~new_n12331_;
  assign new_n12519_ = ~new_n2357_ | ~new_n12292_;
  assign new_n12520_ = ~new_n1392_ | ~new_n12291_;
  assign new_n12521_ = ~new_n2357_ | ~new_n12292_;
  assign new_n12522_ = ~new_n1392_ | ~new_n12291_;
  assign new_n12523_ = ~new_n12522_ | ~new_n12521_;
  assign new_n12524_ = ~new_n12224_ | ~new_n1391_ | ~new_n12523_;
  assign new_n12525_ = ~new_n2346_ | ~new_n12149_ | ~new_n12225_;
  assign new_n12526_ = ~new_n2346_ | ~new_n12225_;
  assign new_n12527_ = ~new_n1391_ | ~new_n12224_;
  assign new_n12528_ = ~new_n12268_;
  assign new_n12529_ = ~new_n12443_ | ~new_n12528_;
  assign new_n12530_ = ~new_n12268_ | ~new_n12294_;
  assign new_n12531_ = ~new_n2347_ | ~new_n12223_;
  assign new_n12532_ = ~new_n1390_ | ~new_n12220_;
  assign new_n12533_ = ~new_n2347_ | ~new_n12223_;
  assign new_n12534_ = ~new_n1390_ | ~new_n12220_;
  assign new_n12535_ = ~new_n12534_ | ~new_n12533_;
  assign new_n12536_ = ~new_n2348_ | ~new_n12221_;
  assign new_n12537_ = ~new_n1394_ | ~new_n12184_;
  assign new_n12538_ = ~new_n12450_ | ~new_n12226_;
  assign new_n12539_ = ~new_n12295_ | ~new_n12437_;
  assign new_n12540_ = ~new_n2349_ | ~new_n12219_;
  assign new_n12541_ = ~new_n1395_ | ~new_n12218_;
  assign new_n12542_ = ~new_n12271_;
  assign new_n12543_ = ~new_n12433_ | ~new_n12542_;
  assign new_n12544_ = ~new_n12271_ | ~new_n12296_;
  assign new_n12545_ = ~new_n2350_ | ~new_n12217_;
  assign new_n12546_ = ~new_n1402_ | ~new_n12216_;
  assign new_n12547_ = ~new_n12272_;
  assign new_n12548_ = ~new_n12429_ | ~new_n12547_;
  assign new_n12549_ = ~new_n12272_ | ~new_n12297_;
  assign new_n12550_ = ~new_n2351_ | ~new_n12212_;
  assign new_n12551_ = ~new_n1403_ | ~new_n12210_;
  assign new_n12552_ = ~new_n12551_ | ~new_n12550_;
  assign new_n12553_ = ~new_n2352_ | ~new_n12213_;
  assign new_n12554_ = ~new_n1398_ | ~new_n12185_;
  assign new_n12555_ = ~new_n12460_ | ~new_n12227_;
  assign new_n12556_ = ~new_n12298_ | ~new_n12452_;
  assign new_n12557_ = ~new_n2353_ | ~new_n12214_;
  assign new_n12558_ = ~new_n1412_ | ~new_n12211_;
  assign new_n12559_ = ~new_n12461_ | ~new_n12300_;
  assign new_n12560_ = ~new_n12419_ | ~new_n12299_;
  assign new_n12561_ = ~new_n2354_ | ~new_n12209_;
  assign new_n12562_ = ~new_n1413_ | ~new_n12208_;
  assign new_n12563_ = ~new_n12274_;
  assign new_n12564_ = ~new_n12415_ | ~new_n12563_;
  assign new_n12565_ = ~new_n12274_ | ~new_n12301_;
  assign new_n12566_ = ~new_n1795_ | ~new_n12163_;
  assign new_n12567_ = ~new_n1415_ | ~new_n12302_;
  assign new_n12568_ = ~new_n12275_;
  assign new_n12569_ = ~new_n12568_ | ~new_n12327_;
  assign new_n12570_ = ~new_n12275_ | ~new_n12162_;
  assign new_n12571_ = ~new_n1848_ | ~new_n12207_;
  assign new_n12572_ = ~new_n1418_ | ~new_n12206_;
  assign new_n12573_ = ~new_n12276_;
  assign new_n12574_ = ~new_n12411_ | ~new_n12573_;
  assign new_n12575_ = ~new_n12276_ | ~new_n12303_;
  assign new_n12576_ = ~new_n1846_ | ~new_n12205_;
  assign new_n12577_ = ~new_n1419_ | ~new_n12304_;
  assign new_n12578_ = ~new_n12277_;
  assign new_n12579_ = ~new_n12578_ | ~new_n12407_;
  assign new_n12580_ = ~new_n12277_ | ~new_n12204_;
  assign new_n12581_ = ~new_n1843_ | ~new_n12203_;
  assign new_n12582_ = ~new_n1406_ | ~new_n12202_;
  assign new_n12583_ = ~new_n12278_;
  assign new_n12584_ = ~new_n12403_ | ~new_n12583_;
  assign new_n12585_ = ~new_n12278_ | ~new_n12305_;
  assign new_n12586_ = ~new_n1840_ | ~new_n12198_;
  assign new_n12587_ = ~new_n1410_ | ~new_n12196_;
  assign new_n12588_ = ~new_n12587_ | ~new_n12586_;
  assign new_n12589_ = ~new_n1837_ | ~new_n12199_;
  assign new_n12590_ = ~new_n1411_ | ~new_n12186_;
  assign new_n12591_ = ~new_n12471_ | ~new_n12228_;
  assign new_n12592_ = ~new_n12306_ | ~new_n12463_;
  assign new_n12593_ = ~new_n1834_ | ~new_n12200_;
  assign new_n12594_ = ~new_n1416_ | ~new_n12197_;
  assign new_n12595_ = ~new_n12472_ | ~new_n12308_;
  assign new_n12596_ = ~new_n12393_ | ~new_n12307_;
  assign new_n12597_ = ~new_n1831_ | ~new_n12195_;
  assign new_n12598_ = ~new_n1417_ | ~new_n12194_;
  assign new_n12599_ = ~new_n12280_;
  assign new_n12600_ = ~new_n12389_ | ~new_n12599_;
  assign new_n12601_ = ~new_n12280_ | ~new_n12309_;
  assign new_n12602_ = ~new_n1828_ | ~new_n12193_;
  assign new_n12603_ = ~new_n1409_ | ~new_n12192_;
  assign new_n12604_ = ~new_n12281_;
  assign new_n12605_ = ~new_n12385_ | ~new_n12604_;
  assign new_n12606_ = ~new_n12281_ | ~new_n12310_;
  assign new_n12607_ = ~new_n1825_ | ~new_n12189_;
  assign new_n12608_ = ~new_n1400_ | ~new_n12187_;
  assign new_n12609_ = ~new_n12608_ | ~new_n12607_;
  assign new_n12610_ = ~new_n1822_ | ~new_n12190_;
  assign new_n12611_ = ~new_n1399_ | ~new_n12188_;
  assign new_n12612_ = ~new_n12482_ | ~new_n12229_;
  assign new_n12613_ = ~new_n12311_ | ~new_n12474_;
  assign new_n12614_ = new_n12792_ & new_n12809_;
  assign new_n12615_ = new_n12811_ & new_n12810_;
  assign new_n12616_ = new_n12787_ & new_n12848_;
  assign new_n12617_ = new_n12850_ & new_n12849_;
  assign new_n12618_ = new_n12867_ & new_n12866_;
  assign new_n12619_ = new_n12893_ & new_n12892_;
  assign new_n12620_ = new_n12991_ & new_n12990_;
  assign new_n12621_ = ~new_n12948_ | ~new_n12951_;
  assign new_n12622_ = ~new_n12937_ | ~new_n12940_;
  assign new_n12623_ = ~new_n12926_ | ~new_n12929_;
  assign new_n12624_ = ~new_n12918_ | ~new_n12920_;
  assign new_n12625_ = ~new_n12956_ | ~new_n12764_ | ~new_n12783_;
  assign new_n12626_ = ~new_n12844_ | ~new_n12846_;
  assign new_n12627_ = ~new_n12836_ | ~new_n12839_;
  assign new_n12628_ = ~new_n12828_ | ~new_n12830_;
  assign new_n12629_ = ~new_n12633_ | ~new_n12954_;
  assign new_n12630_ = ~new_n1813_;
  assign new_n12631_ = ~new_n1798_;
  assign new_n12632_ = ~new_n1790_;
  assign new_n12633_ = ~new_n1790_ | ~new_n12701_;
  assign new_n12634_ = ~new_n1415_;
  assign new_n12635_ = ~new_n1801_;
  assign new_n12636_ = ~new_n1405_;
  assign new_n12637_ = ~new_n1405_ | ~new_n12631_;
  assign new_n12638_ = ~new_n1401_;
  assign new_n12639_ = ~new_n1810_;
  assign new_n12640_ = ~new_n1807_;
  assign new_n12641_ = ~new_n1804_;
  assign new_n12642_ = ~new_n1408_;
  assign new_n12643_ = ~new_n1404_;
  assign new_n12644_ = ~new_n1397_;
  assign new_n12645_ = ~new_n1397_ | ~new_n12641_;
  assign new_n12646_ = ~new_n1816_;
  assign new_n12647_ = ~new_n1407_;
  assign new_n12648_ = ~new_n1407_ | ~new_n12630_;
  assign new_n12649_ = ~new_n1421_;
  assign new_n12650_ = ~new_n1819_;
  assign new_n12651_ = ~new_n1420_;
  assign new_n12652_ = ~new_n12817_ | ~new_n12816_;
  assign new_n12653_ = ~new_n12645_ | ~new_n12832_;
  assign new_n12654_ = ~new_n12801_ | ~new_n12800_;
  assign new_n12655_ = ~new_n2348_;
  assign new_n12656_ = ~new_n2352_;
  assign new_n12657_ = ~new_n1837_;
  assign new_n12658_ = ~new_n1825_;
  assign new_n12659_ = ~new_n1822_;
  assign new_n12660_ = ~new_n1400_;
  assign new_n12661_ = ~new_n1399_;
  assign new_n12662_ = ~new_n1420_ | ~new_n12650_;
  assign new_n12663_ = ~new_n1828_;
  assign new_n12664_ = ~new_n1409_;
  assign new_n12665_ = ~new_n1831_;
  assign new_n12666_ = ~new_n1417_;
  assign new_n12667_ = ~new_n1840_;
  assign new_n12668_ = ~new_n1834_;
  assign new_n12669_ = ~new_n1410_;
  assign new_n12670_ = ~new_n1411_;
  assign new_n12671_ = ~new_n1416_;
  assign new_n12672_ = ~new_n1416_ | ~new_n12668_;
  assign new_n12673_ = ~new_n1843_;
  assign new_n12674_ = ~new_n1406_;
  assign new_n12675_ = ~new_n12877_ | ~new_n12876_;
  assign new_n12676_ = ~new_n1419_;
  assign new_n12677_ = ~new_n1848_;
  assign new_n12678_ = ~new_n1418_;
  assign new_n12679_ = ~new_n2354_;
  assign new_n12680_ = ~new_n1413_;
  assign new_n12681_ = ~new_n2351_;
  assign new_n12682_ = ~new_n2353_;
  assign new_n12683_ = ~new_n1403_;
  assign new_n12684_ = ~new_n1398_;
  assign new_n12685_ = ~new_n1412_;
  assign new_n12686_ = ~new_n1412_ | ~new_n12682_;
  assign new_n12687_ = ~new_n2350_;
  assign new_n12688_ = ~new_n1402_;
  assign new_n12689_ = ~new_n2349_;
  assign new_n12690_ = ~new_n1395_;
  assign new_n12691_ = ~new_n2347_;
  assign new_n12692_ = ~new_n1394_;
  assign new_n12693_ = ~new_n1394_ | ~new_n12655_;
  assign new_n12694_ = ~new_n1390_;
  assign new_n12695_ = ~new_n2346_;
  assign new_n12696_ = ~new_n1391_;
  assign new_n12697_ = ~new_n12907_ | ~new_n12906_;
  assign new_n12698_ = ~new_n12686_ | ~new_n12922_;
  assign new_n12699_ = ~new_n12672_ | ~new_n12933_;
  assign new_n12700_ = ~new_n12662_ | ~new_n12944_;
  assign new_n12701_ = ~new_n1414_;
  assign new_n12702_ = ~new_n13001_ | ~new_n13000_;
  assign new_n12703_ = ~new_n13015_ | ~new_n13014_;
  assign new_n12704_ = ~new_n13020_ | ~new_n13019_;
  assign new_n12705_ = ~new_n13036_ | ~new_n13035_;
  assign new_n12706_ = ~new_n13041_ | ~new_n13040_;
  assign new_n12707_ = ~new_n13046_ | ~new_n13045_;
  assign new_n12708_ = ~new_n13051_ | ~new_n13050_;
  assign new_n12709_ = ~new_n13056_ | ~new_n13055_;
  assign new_n12710_ = ~new_n13072_ | ~new_n13071_;
  assign new_n12711_ = ~new_n13077_ | ~new_n13076_;
  assign new_n12712_ = ~new_n12960_ | ~new_n12959_;
  assign new_n12713_ = ~new_n12969_ | ~new_n12968_;
  assign new_n12714_ = ~new_n12976_ | ~new_n12975_;
  assign new_n12715_ = ~new_n12980_ | ~new_n12979_;
  assign new_n12716_ = ~new_n12989_ | ~new_n12988_;
  assign new_n12717_ = ~new_n13010_ | ~new_n13009_;
  assign new_n12718_ = ~new_n13027_ | ~new_n13026_;
  assign new_n12719_ = ~new_n13031_ | ~new_n13030_;
  assign new_n12720_ = ~new_n13063_ | ~new_n13062_;
  assign new_n12721_ = ~new_n13067_ | ~new_n13066_;
  assign new_n12722_ = ~new_n13084_ | ~new_n13083_;
  assign new_n12723_ = new_n12803_ & new_n12791_;
  assign new_n12724_ = new_n12806_ & new_n12807_;
  assign new_n12725_ = new_n12819_ & new_n12793_;
  assign new_n12726_ = new_n12822_ & new_n12823_;
  assign new_n12727_ = new_n12648_ & new_n12962_ & new_n12961_;
  assign new_n12728_ = new_n12965_ & new_n12793_;
  assign new_n12729_ = new_n12838_ & new_n12615_;
  assign new_n12730_ = new_n12972_ & new_n12792_;
  assign new_n12731_ = new_n12637_ & new_n12982_ & new_n12981_;
  assign new_n12732_ = new_n12985_ & new_n12791_;
  assign new_n12733_ = new_n12825_ & new_n12616_;
  assign new_n12734_ = new_n12870_ & new_n12788_;
  assign new_n12735_ = new_n12896_ & new_n12789_;
  assign new_n12736_ = new_n12912_ & new_n12913_;
  assign new_n12737_ = new_n12915_ & new_n12994_;
  assign new_n12738_ = new_n12916_ & new_n12913_ & new_n12912_;
  assign new_n12739_ = ~new_n12998_ | ~new_n12997_;
  assign new_n12740_ = new_n12693_ & new_n13003_ & new_n13002_;
  assign new_n12741_ = new_n13006_ & new_n12790_;
  assign new_n12742_ = ~new_n13012_ | ~new_n13011_;
  assign new_n12743_ = ~new_n13017_ | ~new_n13016_;
  assign new_n12744_ = new_n13023_ & new_n12789_;
  assign new_n12745_ = ~new_n13033_ | ~new_n13032_;
  assign new_n12746_ = ~new_n13038_ | ~new_n13037_;
  assign new_n12747_ = ~new_n13043_ | ~new_n13042_;
  assign new_n12748_ = ~new_n13048_ | ~new_n13047_;
  assign new_n12749_ = ~new_n13053_ | ~new_n13052_;
  assign new_n12750_ = new_n13059_ & new_n12788_;
  assign new_n12751_ = ~new_n13069_ | ~new_n13068_;
  assign new_n12752_ = ~new_n13074_ | ~new_n13073_;
  assign new_n12753_ = new_n12950_ & new_n12617_;
  assign new_n12754_ = new_n13080_ & new_n12787_;
  assign new_n12755_ = new_n12958_ & new_n12957_;
  assign new_n12756_ = ~new_n12726_ | ~new_n12820_;
  assign new_n12757_ = new_n12967_ & new_n12966_;
  assign new_n12758_ = new_n12974_ & new_n12973_;
  assign new_n12759_ = new_n12978_ & new_n12977_;
  assign new_n12760_ = ~new_n12724_ | ~new_n12804_;
  assign new_n12761_ = new_n12987_ & new_n12986_;
  assign new_n12762_ = ~new_n2357_;
  assign new_n12763_ = ~new_n1392_;
  assign new_n12764_ = new_n12996_ & new_n12995_;
  assign new_n12765_ = ~new_n12736_ | ~new_n12910_;
  assign new_n12766_ = new_n13008_ & new_n13007_;
  assign new_n12767_ = ~new_n12903_ | ~new_n12902_;
  assign new_n12768_ = ~new_n12899_ | ~new_n12898_;
  assign new_n12769_ = new_n13025_ & new_n13024_;
  assign new_n12770_ = new_n13029_ & new_n13028_;
  assign new_n12771_ = ~new_n12889_ | ~new_n12888_;
  assign new_n12772_ = ~new_n12885_ | ~new_n12884_;
  assign new_n12773_ = ~new_n1795_;
  assign new_n12774_ = ~new_n12881_ | ~new_n12880_;
  assign new_n12775_ = ~new_n1846_;
  assign new_n12776_ = ~new_n12873_ | ~new_n12872_;
  assign new_n12777_ = new_n13061_ & new_n13060_;
  assign new_n12778_ = new_n13065_ & new_n13064_;
  assign new_n12779_ = ~new_n12863_ | ~new_n12862_;
  assign new_n12780_ = ~new_n12859_ | ~new_n12858_;
  assign new_n12781_ = ~new_n12855_ | ~new_n12854_;
  assign new_n12782_ = new_n13082_ & new_n13081_;
  assign new_n12783_ = ~new_n12737_ | ~new_n12765_;
  assign new_n12784_ = ~new_n12693_;
  assign new_n12785_ = ~new_n12637_;
  assign new_n12786_ = ~new_n12648_;
  assign new_n12787_ = ~new_n1822_ | ~new_n12661_;
  assign new_n12788_ = ~new_n1837_ | ~new_n12670_;
  assign new_n12789_ = ~new_n2352_ | ~new_n12684_;
  assign new_n12790_ = ~new_n2348_ | ~new_n12692_;
  assign new_n12791_ = ~new_n1798_ | ~new_n12636_;
  assign new_n12792_ = ~new_n1807_ | ~new_n12643_;
  assign new_n12793_ = ~new_n1813_ | ~new_n12647_;
  assign new_n12794_ = ~new_n12672_;
  assign new_n12795_ = ~new_n12686_;
  assign new_n12796_ = ~new_n12645_;
  assign new_n12797_ = ~new_n12662_;
  assign new_n12798_ = ~new_n12633_;
  assign new_n12799_ = ~new_n12798_ | ~new_n12634_;
  assign new_n12800_ = ~new_n12799_ | ~new_n12773_;
  assign new_n12801_ = ~new_n1415_ | ~new_n12633_;
  assign new_n12802_ = ~new_n12654_;
  assign new_n12803_ = ~new_n1801_ | ~new_n12638_;
  assign new_n12804_ = ~new_n12723_ | ~new_n12654_;
  assign new_n12805_ = ~new_n12638_ | ~new_n12637_;
  assign new_n12806_ = ~new_n12805_ | ~new_n12635_;
  assign new_n12807_ = ~new_n1401_ | ~new_n12785_;
  assign new_n12808_ = ~new_n12760_;
  assign new_n12809_ = ~new_n1810_ | ~new_n12642_;
  assign new_n12810_ = ~new_n1408_ | ~new_n12639_;
  assign new_n12811_ = ~new_n1404_ | ~new_n12640_;
  assign new_n12812_ = ~new_n12796_ | ~new_n12614_;
  assign new_n12813_ = ~new_n12615_ | ~new_n12812_;
  assign new_n12814_ = ~new_n1804_ | ~new_n12644_;
  assign new_n12815_ = ~new_n1810_ | ~new_n12642_;
  assign new_n12816_ = ~new_n12614_ | ~new_n12814_ | ~new_n12760_;
  assign new_n12817_ = ~new_n12815_ | ~new_n12813_;
  assign new_n12818_ = ~new_n12652_;
  assign new_n12819_ = ~new_n1816_ | ~new_n12649_;
  assign new_n12820_ = ~new_n12725_ | ~new_n12652_;
  assign new_n12821_ = ~new_n12649_ | ~new_n12648_;
  assign new_n12822_ = ~new_n12821_ | ~new_n12646_;
  assign new_n12823_ = ~new_n1421_ | ~new_n12786_;
  assign new_n12824_ = ~new_n12756_;
  assign new_n12825_ = ~new_n1819_ | ~new_n12651_;
  assign new_n12826_ = ~new_n12825_ | ~new_n12662_;
  assign new_n12827_ = ~new_n12818_ | ~new_n12648_;
  assign new_n12828_ = ~new_n12728_ | ~new_n12827_;
  assign new_n12829_ = ~new_n12652_ | ~new_n12793_;
  assign new_n12830_ = ~new_n12727_ | ~new_n12829_;
  assign new_n12831_ = ~new_n12648_ | ~new_n12793_;
  assign new_n12832_ = ~new_n12814_ | ~new_n12760_;
  assign new_n12833_ = ~new_n12653_;
  assign new_n12834_ = ~new_n1404_ | ~new_n12640_;
  assign new_n12835_ = ~new_n12833_ | ~new_n12834_;
  assign new_n12836_ = ~new_n12730_ | ~new_n12835_;
  assign new_n12837_ = ~new_n12653_ | ~new_n12792_;
  assign new_n12838_ = ~new_n1810_ | ~new_n12642_;
  assign new_n12839_ = ~new_n12729_ | ~new_n12837_;
  assign new_n12840_ = ~new_n1404_ | ~new_n12640_;
  assign new_n12841_ = ~new_n12792_ | ~new_n12840_;
  assign new_n12842_ = ~new_n12814_ | ~new_n12645_;
  assign new_n12843_ = ~new_n12802_ | ~new_n12637_;
  assign new_n12844_ = ~new_n12732_ | ~new_n12843_;
  assign new_n12845_ = ~new_n12654_ | ~new_n12791_;
  assign new_n12846_ = ~new_n12731_ | ~new_n12845_;
  assign new_n12847_ = ~new_n12637_ | ~new_n12791_;
  assign new_n12848_ = ~new_n1825_ | ~new_n12660_;
  assign new_n12849_ = ~new_n1400_ | ~new_n12658_;
  assign new_n12850_ = ~new_n1399_ | ~new_n12659_;
  assign new_n12851_ = ~new_n12797_ | ~new_n12616_;
  assign new_n12852_ = ~new_n12617_ | ~new_n12851_;
  assign new_n12853_ = ~new_n1825_ | ~new_n12660_;
  assign new_n12854_ = ~new_n12733_ | ~new_n12756_;
  assign new_n12855_ = ~new_n12853_ | ~new_n12852_;
  assign new_n12856_ = ~new_n12781_;
  assign new_n12857_ = ~new_n1828_ | ~new_n12664_;
  assign new_n12858_ = ~new_n12857_ | ~new_n12781_;
  assign new_n12859_ = ~new_n1409_ | ~new_n12663_;
  assign new_n12860_ = ~new_n12780_;
  assign new_n12861_ = ~new_n1831_ | ~new_n12666_;
  assign new_n12862_ = ~new_n12861_ | ~new_n12780_;
  assign new_n12863_ = ~new_n1417_ | ~new_n12665_;
  assign new_n12864_ = ~new_n12779_;
  assign new_n12865_ = ~new_n1840_ | ~new_n12669_;
  assign new_n12866_ = ~new_n1410_ | ~new_n12667_;
  assign new_n12867_ = ~new_n1411_ | ~new_n12657_;
  assign new_n12868_ = ~new_n12794_ | ~new_n12788_;
  assign new_n12869_ = ~new_n12618_ | ~new_n12868_;
  assign new_n12870_ = ~new_n1834_ | ~new_n12671_;
  assign new_n12871_ = ~new_n1840_ | ~new_n12669_;
  assign new_n12872_ = ~new_n12865_ | ~new_n12779_ | ~new_n12734_;
  assign new_n12873_ = ~new_n12871_ | ~new_n12869_;
  assign new_n12874_ = ~new_n12776_;
  assign new_n12875_ = ~new_n1843_ | ~new_n12674_;
  assign new_n12876_ = ~new_n12875_ | ~new_n12776_;
  assign new_n12877_ = ~new_n1406_ | ~new_n12673_;
  assign new_n12878_ = ~new_n12675_;
  assign new_n12879_ = ~new_n12878_ | ~new_n12676_;
  assign new_n12880_ = ~new_n12879_ | ~new_n12775_;
  assign new_n12881_ = ~new_n1419_ | ~new_n12675_;
  assign new_n12882_ = ~new_n12774_;
  assign new_n12883_ = ~new_n1848_ | ~new_n12678_;
  assign new_n12884_ = ~new_n12883_ | ~new_n12774_;
  assign new_n12885_ = ~new_n1418_ | ~new_n12677_;
  assign new_n12886_ = ~new_n12772_;
  assign new_n12887_ = ~new_n2354_ | ~new_n12680_;
  assign new_n12888_ = ~new_n12887_ | ~new_n12772_;
  assign new_n12889_ = ~new_n1413_ | ~new_n12679_;
  assign new_n12890_ = ~new_n12771_;
  assign new_n12891_ = ~new_n2351_ | ~new_n12683_;
  assign new_n12892_ = ~new_n1403_ | ~new_n12681_;
  assign new_n12893_ = ~new_n1398_ | ~new_n12656_;
  assign new_n12894_ = ~new_n12795_ | ~new_n12789_;
  assign new_n12895_ = ~new_n12619_ | ~new_n12894_;
  assign new_n12896_ = ~new_n2353_ | ~new_n12685_;
  assign new_n12897_ = ~new_n2351_ | ~new_n12683_;
  assign new_n12898_ = ~new_n12891_ | ~new_n12771_ | ~new_n12735_;
  assign new_n12899_ = ~new_n12897_ | ~new_n12895_;
  assign new_n12900_ = ~new_n12768_;
  assign new_n12901_ = ~new_n2350_ | ~new_n12688_;
  assign new_n12902_ = ~new_n12901_ | ~new_n12768_;
  assign new_n12903_ = ~new_n1402_ | ~new_n12687_;
  assign new_n12904_ = ~new_n12767_;
  assign new_n12905_ = ~new_n2349_ | ~new_n12690_;
  assign new_n12906_ = ~new_n12905_ | ~new_n12767_;
  assign new_n12907_ = ~new_n1395_ | ~new_n12689_;
  assign new_n12908_ = ~new_n12697_;
  assign new_n12909_ = ~new_n2347_ | ~new_n12694_;
  assign new_n12910_ = ~new_n12909_ | ~new_n12697_ | ~new_n12790_;
  assign new_n12911_ = ~new_n12694_ | ~new_n12693_;
  assign new_n12912_ = ~new_n12911_ | ~new_n12691_;
  assign new_n12913_ = ~new_n1390_ | ~new_n12784_;
  assign new_n12914_ = ~new_n12765_;
  assign new_n12915_ = ~new_n2346_ | ~new_n12696_;
  assign new_n12916_ = ~new_n1391_ | ~new_n12695_;
  assign new_n12917_ = ~new_n12908_ | ~new_n12693_;
  assign new_n12918_ = ~new_n12741_ | ~new_n12917_;
  assign new_n12919_ = ~new_n12697_ | ~new_n12790_;
  assign new_n12920_ = ~new_n12740_ | ~new_n12919_;
  assign new_n12921_ = ~new_n12693_ | ~new_n12790_;
  assign new_n12922_ = ~new_n12896_ | ~new_n12771_;
  assign new_n12923_ = ~new_n12698_;
  assign new_n12924_ = ~new_n1398_ | ~new_n12656_;
  assign new_n12925_ = ~new_n12923_ | ~new_n12924_;
  assign new_n12926_ = ~new_n12744_ | ~new_n12925_;
  assign new_n12927_ = ~new_n12698_ | ~new_n12789_;
  assign new_n12928_ = ~new_n2351_ | ~new_n12683_;
  assign new_n12929_ = ~new_n12619_ | ~new_n12928_ | ~new_n12927_;
  assign new_n12930_ = ~new_n1398_ | ~new_n12656_;
  assign new_n12931_ = ~new_n12789_ | ~new_n12930_;
  assign new_n12932_ = ~new_n12896_ | ~new_n12686_;
  assign new_n12933_ = ~new_n12870_ | ~new_n12779_;
  assign new_n12934_ = ~new_n12699_;
  assign new_n12935_ = ~new_n1411_ | ~new_n12657_;
  assign new_n12936_ = ~new_n12934_ | ~new_n12935_;
  assign new_n12937_ = ~new_n12750_ | ~new_n12936_;
  assign new_n12938_ = ~new_n12699_ | ~new_n12788_;
  assign new_n12939_ = ~new_n1840_ | ~new_n12669_;
  assign new_n12940_ = ~new_n12618_ | ~new_n12939_ | ~new_n12938_;
  assign new_n12941_ = ~new_n1411_ | ~new_n12657_;
  assign new_n12942_ = ~new_n12788_ | ~new_n12941_;
  assign new_n12943_ = ~new_n12870_ | ~new_n12672_;
  assign new_n12944_ = ~new_n12825_ | ~new_n12756_;
  assign new_n12945_ = ~new_n12700_;
  assign new_n12946_ = ~new_n1399_ | ~new_n12659_;
  assign new_n12947_ = ~new_n12945_ | ~new_n12946_;
  assign new_n12948_ = ~new_n12754_ | ~new_n12947_;
  assign new_n12949_ = ~new_n12700_ | ~new_n12787_;
  assign new_n12950_ = ~new_n1825_ | ~new_n12660_;
  assign new_n12951_ = ~new_n12753_ | ~new_n12949_;
  assign new_n12952_ = ~new_n1399_ | ~new_n12659_;
  assign new_n12953_ = ~new_n12787_ | ~new_n12952_;
  assign new_n12954_ = ~new_n1414_ | ~new_n12632_;
  assign new_n12955_ = ~new_n12909_ | ~new_n12697_ | ~new_n12790_;
  assign new_n12956_ = ~new_n12738_ | ~new_n12620_ | ~new_n12955_;
  assign new_n12957_ = ~new_n1819_ | ~new_n12651_;
  assign new_n12958_ = ~new_n1420_ | ~new_n12650_;
  assign new_n12959_ = ~new_n12826_ | ~new_n12756_;
  assign new_n12960_ = ~new_n12824_ | ~new_n12755_;
  assign new_n12961_ = ~new_n1816_ | ~new_n12649_;
  assign new_n12962_ = ~new_n1421_ | ~new_n12646_;
  assign new_n12963_ = ~new_n1816_ | ~new_n12649_;
  assign new_n12964_ = ~new_n1421_ | ~new_n12646_;
  assign new_n12965_ = ~new_n12964_ | ~new_n12963_;
  assign new_n12966_ = ~new_n1813_ | ~new_n12647_;
  assign new_n12967_ = ~new_n1407_ | ~new_n12630_;
  assign new_n12968_ = ~new_n12831_ | ~new_n12652_;
  assign new_n12969_ = ~new_n12757_ | ~new_n12818_;
  assign new_n12970_ = ~new_n1810_ | ~new_n12642_;
  assign new_n12971_ = ~new_n1408_ | ~new_n12639_;
  assign new_n12972_ = ~new_n12971_ | ~new_n12970_;
  assign new_n12973_ = ~new_n1807_ | ~new_n12643_;
  assign new_n12974_ = ~new_n1404_ | ~new_n12640_;
  assign new_n12975_ = ~new_n12841_ | ~new_n12653_;
  assign new_n12976_ = ~new_n12758_ | ~new_n12833_;
  assign new_n12977_ = ~new_n1804_ | ~new_n12644_;
  assign new_n12978_ = ~new_n1397_ | ~new_n12641_;
  assign new_n12979_ = ~new_n12842_ | ~new_n12760_;
  assign new_n12980_ = ~new_n12808_ | ~new_n12759_;
  assign new_n12981_ = ~new_n1801_ | ~new_n12638_;
  assign new_n12982_ = ~new_n1401_ | ~new_n12635_;
  assign new_n12983_ = ~new_n1801_ | ~new_n12638_;
  assign new_n12984_ = ~new_n1401_ | ~new_n12635_;
  assign new_n12985_ = ~new_n12984_ | ~new_n12983_;
  assign new_n12986_ = ~new_n1798_ | ~new_n12636_;
  assign new_n12987_ = ~new_n1405_ | ~new_n12631_;
  assign new_n12988_ = ~new_n12847_ | ~new_n12654_;
  assign new_n12989_ = ~new_n12761_ | ~new_n12802_;
  assign new_n12990_ = ~new_n2357_ | ~new_n12763_;
  assign new_n12991_ = ~new_n1392_ | ~new_n12762_;
  assign new_n12992_ = ~new_n2357_ | ~new_n12763_;
  assign new_n12993_ = ~new_n1392_ | ~new_n12762_;
  assign new_n12994_ = ~new_n12993_ | ~new_n12992_;
  assign new_n12995_ = ~new_n12695_ | ~new_n1391_ | ~new_n12994_;
  assign new_n12996_ = ~new_n2346_ | ~new_n12620_ | ~new_n12696_;
  assign new_n12997_ = ~new_n2346_ | ~new_n12696_;
  assign new_n12998_ = ~new_n1391_ | ~new_n12695_;
  assign new_n12999_ = ~new_n12739_;
  assign new_n13000_ = ~new_n12914_ | ~new_n12999_;
  assign new_n13001_ = ~new_n12739_ | ~new_n12765_;
  assign new_n13002_ = ~new_n2347_ | ~new_n12694_;
  assign new_n13003_ = ~new_n1390_ | ~new_n12691_;
  assign new_n13004_ = ~new_n2347_ | ~new_n12694_;
  assign new_n13005_ = ~new_n1390_ | ~new_n12691_;
  assign new_n13006_ = ~new_n13005_ | ~new_n13004_;
  assign new_n13007_ = ~new_n2348_ | ~new_n12692_;
  assign new_n13008_ = ~new_n1394_ | ~new_n12655_;
  assign new_n13009_ = ~new_n12921_ | ~new_n12697_;
  assign new_n13010_ = ~new_n12766_ | ~new_n12908_;
  assign new_n13011_ = ~new_n2349_ | ~new_n12690_;
  assign new_n13012_ = ~new_n1395_ | ~new_n12689_;
  assign new_n13013_ = ~new_n12742_;
  assign new_n13014_ = ~new_n12904_ | ~new_n13013_;
  assign new_n13015_ = ~new_n12742_ | ~new_n12767_;
  assign new_n13016_ = ~new_n2350_ | ~new_n12688_;
  assign new_n13017_ = ~new_n1402_ | ~new_n12687_;
  assign new_n13018_ = ~new_n12743_;
  assign new_n13019_ = ~new_n12900_ | ~new_n13018_;
  assign new_n13020_ = ~new_n12743_ | ~new_n12768_;
  assign new_n13021_ = ~new_n2351_ | ~new_n12683_;
  assign new_n13022_ = ~new_n1403_ | ~new_n12681_;
  assign new_n13023_ = ~new_n13022_ | ~new_n13021_;
  assign new_n13024_ = ~new_n2352_ | ~new_n12684_;
  assign new_n13025_ = ~new_n1398_ | ~new_n12656_;
  assign new_n13026_ = ~new_n12931_ | ~new_n12698_;
  assign new_n13027_ = ~new_n12769_ | ~new_n12923_;
  assign new_n13028_ = ~new_n2353_ | ~new_n12685_;
  assign new_n13029_ = ~new_n1412_ | ~new_n12682_;
  assign new_n13030_ = ~new_n12932_ | ~new_n12771_;
  assign new_n13031_ = ~new_n12890_ | ~new_n12770_;
  assign new_n13032_ = ~new_n2354_ | ~new_n12680_;
  assign new_n13033_ = ~new_n1413_ | ~new_n12679_;
  assign new_n13034_ = ~new_n12745_;
  assign new_n13035_ = ~new_n12886_ | ~new_n13034_;
  assign new_n13036_ = ~new_n12745_ | ~new_n12772_;
  assign new_n13037_ = ~new_n1795_ | ~new_n12634_;
  assign new_n13038_ = ~new_n1415_ | ~new_n12773_;
  assign new_n13039_ = ~new_n12746_;
  assign new_n13040_ = ~new_n13039_ | ~new_n12798_;
  assign new_n13041_ = ~new_n12746_ | ~new_n12633_;
  assign new_n13042_ = ~new_n1848_ | ~new_n12678_;
  assign new_n13043_ = ~new_n1418_ | ~new_n12677_;
  assign new_n13044_ = ~new_n12747_;
  assign new_n13045_ = ~new_n12882_ | ~new_n13044_;
  assign new_n13046_ = ~new_n12747_ | ~new_n12774_;
  assign new_n13047_ = ~new_n1846_ | ~new_n12676_;
  assign new_n13048_ = ~new_n1419_ | ~new_n12775_;
  assign new_n13049_ = ~new_n12748_;
  assign new_n13050_ = ~new_n13049_ | ~new_n12878_;
  assign new_n13051_ = ~new_n12748_ | ~new_n12675_;
  assign new_n13052_ = ~new_n1843_ | ~new_n12674_;
  assign new_n13053_ = ~new_n1406_ | ~new_n12673_;
  assign new_n13054_ = ~new_n12749_;
  assign new_n13055_ = ~new_n12874_ | ~new_n13054_;
  assign new_n13056_ = ~new_n12749_ | ~new_n12776_;
  assign new_n13057_ = ~new_n1840_ | ~new_n12669_;
  assign new_n13058_ = ~new_n1410_ | ~new_n12667_;
  assign new_n13059_ = ~new_n13058_ | ~new_n13057_;
  assign new_n13060_ = ~new_n1837_ | ~new_n12670_;
  assign new_n13061_ = ~new_n1411_ | ~new_n12657_;
  assign new_n13062_ = ~new_n12942_ | ~new_n12699_;
  assign new_n13063_ = ~new_n12777_ | ~new_n12934_;
  assign new_n13064_ = ~new_n1834_ | ~new_n12671_;
  assign new_n13065_ = ~new_n1416_ | ~new_n12668_;
  assign new_n13066_ = ~new_n12943_ | ~new_n12779_;
  assign new_n13067_ = ~new_n12864_ | ~new_n12778_;
  assign new_n13068_ = ~new_n1831_ | ~new_n12666_;
  assign new_n13069_ = ~new_n1417_ | ~new_n12665_;
  assign new_n13070_ = ~new_n12751_;
  assign new_n13071_ = ~new_n12860_ | ~new_n13070_;
  assign new_n13072_ = ~new_n12751_ | ~new_n12780_;
  assign new_n13073_ = ~new_n1828_ | ~new_n12664_;
  assign new_n13074_ = ~new_n1409_ | ~new_n12663_;
  assign new_n13075_ = ~new_n12752_;
  assign new_n13076_ = ~new_n12856_ | ~new_n13075_;
  assign new_n13077_ = ~new_n12752_ | ~new_n12781_;
  assign new_n13078_ = ~new_n1825_ | ~new_n12660_;
  assign new_n13079_ = ~new_n1400_ | ~new_n12658_;
  assign new_n13080_ = ~new_n13079_ | ~new_n13078_;
  assign new_n13081_ = ~new_n1822_ | ~new_n12661_;
  assign new_n13082_ = ~new_n1399_ | ~new_n12659_;
  assign new_n13083_ = ~new_n12953_ | ~new_n12700_;
  assign new_n13084_ = ~new_n12782_ | ~new_n12945_;
  assign new_n13085_ = new_n13188_ & new_n13187_;
  assign new_n13086_ = new_n13190_ & new_n13191_;
  assign new_n13087_ = new_n13192_ & new_n13193_;
  assign new_n13088_ = new_n13087_ & new_n13197_ & new_n13160_ & new_n13195_;
  assign new_n13089_ = new_n13205_ & new_n13204_;
  assign new_n13090_ = new_n13164_ & new_n13163_ & new_n13206_ & new_n13203_;
  assign new_n13091_ = new_n13220_ & new_n13219_;
  assign new_n13092_ = new_n13181_ & new_n13272_;
  assign new_n13093_ = new_n13268_ & new_n13183_;
  assign new_n13094_ = ~new_n1933_;
  assign new_n13095_ = ~new_n1934_;
  assign new_n13096_ = ~new_n2356_;
  assign new_n13097_ = ~new_n2357_;
  assign new_n13098_ = ~new_n1938_;
  assign new_n13099_ = ~new_n2350_;
  assign new_n13100_ = ~new_n2349_;
  assign new_n13101_ = ~new_n1943_;
  assign new_n13102_ = ~new_n2353_;
  assign new_n13103_ = ~new_n1944_;
  assign new_n13104_ = ~new_n2354_;
  assign new_n13105_ = ~new_n1848_;
  assign new_n13106_ = ~new_n1948_;
  assign new_n13107_ = ~new_n1846_;
  assign new_n13108_ = ~new_n1949_;
  assign new_n13109_ = ~new_n1947_;
  assign new_n13110_ = ~new_n1945_;
  assign new_n13111_ = ~new_n1843_;
  assign new_n13112_ = ~new_n1840_;
  assign new_n13113_ = ~new_n1950_;
  assign new_n13114_ = ~new_n1951_;
  assign new_n13115_ = ~new_n1813_;
  assign new_n13116_ = ~new_n1929_;
  assign new_n13117_ = ~new_n1810_;
  assign new_n13118_ = ~new_n1930_;
  assign new_n13119_ = ~new_n1926_;
  assign new_n13120_ = ~new_n1956_;
  assign new_n13121_ = ~new_n1927_;
  assign new_n13122_ = ~new_n1928_;
  assign new_n13123_ = ~new_n1931_;
  assign new_n13124_ = ~new_n1932_;
  assign new_n13125_ = ~new_n1790_ | ~new_n13184_;
  assign new_n13126_ = ~new_n1795_;
  assign new_n13127_ = ~new_n1935_;
  assign new_n13128_ = ~new_n1828_;
  assign new_n13129_ = ~new_n1831_;
  assign new_n13130_ = ~new_n1798_;
  assign new_n13131_ = ~new_n1801_;
  assign new_n13132_ = ~new_n1804_;
  assign new_n13133_ = ~new_n1807_;
  assign new_n13134_ = ~new_n1816_;
  assign new_n13135_ = ~new_n1819_;
  assign new_n13136_ = ~new_n1822_;
  assign new_n13137_ = ~new_n1825_;
  assign new_n13138_ = ~new_n1954_;
  assign new_n13139_ = ~new_n1955_;
  assign new_n13140_ = ~new_n1952_;
  assign new_n13141_ = ~new_n1953_;
  assign new_n13142_ = ~new_n1834_;
  assign new_n13143_ = ~new_n1837_;
  assign new_n13144_ = ~new_n2352_;
  assign new_n13145_ = ~new_n2351_;
  assign new_n13146_ = ~new_n1942_;
  assign new_n13147_ = ~new_n1939_;
  assign new_n13148_ = ~new_n1941_;
  assign new_n13149_ = ~new_n1940_;
  assign new_n13150_ = ~new_n2348_;
  assign new_n13151_ = ~new_n2347_;
  assign new_n13152_ = ~new_n2346_;
  assign new_n13153_ = ~new_n1936_;
  assign new_n13154_ = ~new_n2355_;
  assign new_n13155_ = new_n2353_ & new_n13103_;
  assign new_n13156_ = new_n2354_ & new_n13110_;
  assign new_n13157_ = new_n13250_ & new_n13249_;
  assign new_n13158_ = new_n1948_ & new_n13107_;
  assign new_n13159_ = new_n1949_ & new_n13111_;
  assign new_n13160_ = new_n13196_ & new_n13194_;
  assign new_n13161_ = new_n1929_ & new_n13117_;
  assign new_n13162_ = new_n1930_ & new_n13133_;
  assign new_n13163_ = new_n13208_ & new_n13207_;
  assign new_n13164_ = new_n13209_ & new_n13210_ & new_n13212_ & new_n13211_;
  assign new_n13165_ = new_n13216_ & new_n13217_;
  assign new_n13166_ = new_n13165_ & new_n13215_;
  assign new_n13167_ = new_n1798_ & new_n13127_;
  assign new_n13168_ = new_n1801_ & new_n13124_;
  assign new_n13169_ = new_n13209_ & new_n13210_ & new_n13203_;
  assign new_n13170_ = new_n13233_ & new_n13218_;
  assign new_n13171_ = new_n13236_ & new_n13235_;
  assign new_n13172_ = new_n13171_ & new_n13091_;
  assign new_n13173_ = new_n1954_ & new_n13128_;
  assign new_n13174_ = new_n1955_ & new_n13137_;
  assign new_n13175_ = new_n13239_ & new_n13240_;
  assign new_n13176_ = new_n13242_ & new_n13241_;
  assign new_n13177_ = new_n13200_ & new_n13199_ & new_n13253_ & new_n13252_;
  assign new_n13178_ = new_n13257_ & new_n13256_;
  assign new_n13179_ = new_n1942_ & new_n13145_;
  assign new_n13180_ = new_n13274_ & new_n13263_;
  assign new_n13181_ = new_n13266_ & new_n13152_;
  assign new_n13182_ = new_n1936_ & new_n13097_;
  assign new_n13183_ = new_n13269_ & new_n13270_ & new_n13186_;
  assign new_n13184_ = ~new_n1957_;
  assign new_n13185_ = ~new_n1933_ | ~new_n13154_;
  assign new_n13186_ = ~new_n13096_ | ~new_n13185_ | ~new_n1934_;
  assign new_n13187_ = ~new_n2356_ | ~new_n13095_;
  assign new_n13188_ = ~new_n1933_ | ~new_n13154_;
  assign new_n13189_ = ~new_n1938_ | ~new_n13151_;
  assign new_n13190_ = ~new_n1848_ | ~new_n13109_;
  assign new_n13191_ = ~new_n1846_ | ~new_n13106_;
  assign new_n13192_ = ~new_n1943_ | ~new_n13144_;
  assign new_n13193_ = ~new_n1944_ | ~new_n13102_;
  assign new_n13194_ = ~new_n13158_ | ~new_n13190_;
  assign new_n13195_ = ~new_n13159_ | ~new_n13086_;
  assign new_n13196_ = ~new_n1947_ | ~new_n13105_;
  assign new_n13197_ = ~new_n1945_ | ~new_n13104_;
  assign new_n13198_ = ~new_n1950_ | ~new_n13112_;
  assign new_n13199_ = ~new_n2350_ | ~new_n13148_;
  assign new_n13200_ = ~new_n2349_ | ~new_n13149_;
  assign new_n13201_ = ~new_n1951_ | ~new_n13143_;
  assign new_n13202_ = ~new_n1813_ | ~new_n13122_;
  assign new_n13203_ = ~new_n13161_ | ~new_n13202_;
  assign new_n13204_ = ~new_n1810_ | ~new_n13116_;
  assign new_n13205_ = ~new_n1813_ | ~new_n13122_;
  assign new_n13206_ = ~new_n13162_ | ~new_n13089_;
  assign new_n13207_ = ~new_n1926_ | ~new_n13135_;
  assign new_n13208_ = ~new_n1956_ | ~new_n13136_;
  assign new_n13209_ = ~new_n1927_ | ~new_n13134_;
  assign new_n13210_ = ~new_n1928_ | ~new_n13115_;
  assign new_n13211_ = ~new_n1931_ | ~new_n13132_;
  assign new_n13212_ = ~new_n1932_ | ~new_n13131_;
  assign new_n13213_ = ~new_n13125_;
  assign new_n13214_ = ~new_n1795_ | ~new_n13213_;
  assign new_n13215_ = ~new_n1946_ | ~new_n13214_;
  assign new_n13216_ = ~new_n13125_ | ~new_n13126_;
  assign new_n13217_ = ~new_n1935_ | ~new_n13130_;
  assign new_n13218_ = ~new_n13166_ | ~new_n13090_;
  assign new_n13219_ = ~new_n1828_ | ~new_n13138_;
  assign new_n13220_ = ~new_n1831_ | ~new_n13141_;
  assign new_n13221_ = ~new_n13168_ | ~new_n13211_;
  assign new_n13222_ = ~new_n1804_ | ~new_n13123_;
  assign new_n13223_ = ~new_n13089_ | ~new_n13222_ | ~new_n13221_;
  assign new_n13224_ = ~new_n13223_ | ~new_n13206_;
  assign new_n13225_ = ~new_n1807_ | ~new_n13118_;
  assign new_n13226_ = ~new_n13225_ | ~new_n13224_;
  assign new_n13227_ = ~new_n13169_ | ~new_n13226_;
  assign new_n13228_ = ~new_n1816_ | ~new_n13121_;
  assign new_n13229_ = ~new_n13228_ | ~new_n13227_;
  assign new_n13230_ = ~new_n13229_ | ~new_n13207_;
  assign new_n13231_ = ~new_n1819_ | ~new_n13119_;
  assign new_n13232_ = ~new_n13231_ | ~new_n13230_;
  assign new_n13233_ = ~new_n13167_ | ~new_n13090_;
  assign new_n13234_ = ~new_n13232_ | ~new_n13208_;
  assign new_n13235_ = ~new_n1822_ | ~new_n13120_;
  assign new_n13236_ = ~new_n1825_ | ~new_n13139_;
  assign new_n13237_ = ~new_n13172_ | ~new_n13170_ | ~new_n13234_;
  assign new_n13238_ = ~new_n1831_ | ~new_n13141_;
  assign new_n13239_ = ~new_n13173_ | ~new_n13238_;
  assign new_n13240_ = ~new_n13174_ | ~new_n13091_;
  assign new_n13241_ = ~new_n1952_ | ~new_n13142_;
  assign new_n13242_ = ~new_n1953_ | ~new_n13129_;
  assign new_n13243_ = ~new_n13176_ | ~new_n13175_ | ~new_n13237_;
  assign new_n13244_ = ~new_n1834_ | ~new_n13140_;
  assign new_n13245_ = ~new_n13244_ | ~new_n13243_;
  assign new_n13246_ = ~new_n13245_ | ~new_n13201_;
  assign new_n13247_ = ~new_n1837_ | ~new_n13114_;
  assign new_n13248_ = ~new_n13247_ | ~new_n13246_;
  assign new_n13249_ = ~new_n1843_ | ~new_n13108_;
  assign new_n13250_ = ~new_n1840_ | ~new_n13113_;
  assign new_n13251_ = ~new_n13157_ | ~new_n13086_;
  assign new_n13252_ = ~new_n13155_ | ~new_n13192_;
  assign new_n13253_ = ~new_n13156_ | ~new_n13087_;
  assign new_n13254_ = ~new_n13088_ | ~new_n13251_;
  assign new_n13255_ = ~new_n13088_ | ~new_n13248_ | ~new_n13198_;
  assign new_n13256_ = ~new_n2352_ | ~new_n13101_;
  assign new_n13257_ = ~new_n2351_ | ~new_n13146_;
  assign new_n13258_ = ~new_n13177_ | ~new_n13178_ | ~new_n13255_ | ~new_n13254_;
  assign new_n13259_ = ~new_n13200_ | ~new_n13199_ | ~new_n13179_;
  assign new_n13260_ = ~new_n2349_ | ~new_n13149_;
  assign new_n13261_ = ~new_n1941_ | ~new_n13099_;
  assign new_n13262_ = ~new_n1940_ | ~new_n13100_;
  assign new_n13263_ = ~new_n1939_ | ~new_n13150_;
  assign new_n13264_ = ~new_n13180_ | ~new_n13259_ | ~new_n13258_;
  assign new_n13265_ = ~new_n2348_ | ~new_n13147_;
  assign new_n13266_ = ~new_n2347_ | ~new_n13098_;
  assign new_n13267_ = ~new_n2357_ | ~new_n13153_;
  assign new_n13268_ = ~new_n13267_ | ~new_n13275_ | ~new_n13085_ | ~new_n13277_;
  assign new_n13269_ = ~new_n13182_ | ~new_n13085_;
  assign new_n13270_ = ~new_n2355_ | ~new_n13094_;
  assign new_n13271_ = ~new_n13265_ | ~new_n13264_;
  assign new_n13272_ = ~new_n13271_ | ~new_n13189_;
  assign new_n13273_ = ~new_n13262_ | ~new_n13261_;
  assign new_n13274_ = ~new_n13273_ | ~new_n13260_;
  assign new_n13275_ = new_n1937_ | new_n13092_;
  assign new_n13276_ = ~new_n13266_ | ~new_n13272_;
  assign new_n13277_ = ~new_n2346_ | ~new_n13276_;
  assign new_n13278_ = new_n13383_ & new_n13384_;
  assign new_n13279_ = new_n13388_ & new_n13387_;
  assign new_n13280_ = new_n13390_ & new_n13391_;
  assign new_n13281_ = new_n13395_ & new_n13394_;
  assign new_n13282_ = new_n13455_ & new_n13456_ & new_n13458_ & new_n13471_ & new_n13457_;
  assign new_n13283_ = new_n13455_ & new_n13376_;
  assign new_n13284_ = new_n13475_ & new_n13474_;
  assign new_n13285_ = new_n13477_ & new_n13476_;
  assign new_n13286_ = ~new_n13379_ | ~new_n13380_ | ~new_n13472_;
  assign new_n13287_ = ~new_n1425_;
  assign new_n13288_ = ~new_n1424_;
  assign new_n13289_ = ~new_n1458_;
  assign new_n13290_ = ~new_n1426_;
  assign new_n13291_ = ~new_n1427_;
  assign new_n13292_ = ~new_n1460_;
  assign new_n13293_ = ~new_n1459_;
  assign new_n13294_ = ~new_n1457_;
  assign new_n13295_ = ~new_n1464_;
  assign new_n13296_ = ~new_n1463_;
  assign new_n13297_ = ~new_n1434_;
  assign new_n13298_ = ~new_n1435_;
  assign new_n13299_ = ~new_n1470_;
  assign new_n13300_ = ~new_n1469_;
  assign new_n13301_ = ~new_n1440_;
  assign new_n13302_ = ~new_n1441_;
  assign new_n13303_ = ~new_n1476_;
  assign new_n13304_ = ~new_n1475_;
  assign new_n13305_ = ~new_n1446_;
  assign new_n13306_ = ~new_n1479_;
  assign new_n13307_ = ~new_n1447_;
  assign new_n13308_ = ~new_n1480_;
  assign new_n13309_ = ~new_n1449_;
  assign new_n13310_ = ~new_n1448_;
  assign new_n13311_ = ~new_n1451_;
  assign new_n13312_ = ~new_n1450_;
  assign new_n13313_ = ~new_n1453_;
  assign new_n13314_ = ~new_n1452_;
  assign new_n13315_ = ~new_n1454_;
  assign new_n13316_ = ~new_n1486_;
  assign new_n13317_ = ~new_n1485_;
  assign new_n13318_ = ~new_n1484_;
  assign new_n13319_ = ~new_n1483_;
  assign new_n13320_ = ~new_n1482_;
  assign new_n13321_ = ~new_n1481_;
  assign new_n13322_ = ~new_n1478_;
  assign new_n13323_ = ~new_n1477_;
  assign new_n13324_ = ~new_n1445_;
  assign new_n13325_ = ~new_n1443_;
  assign new_n13326_ = ~new_n1444_;
  assign new_n13327_ = ~new_n1442_;
  assign new_n13328_ = ~new_n1474_;
  assign new_n13329_ = ~new_n1473_;
  assign new_n13330_ = ~new_n1472_;
  assign new_n13331_ = ~new_n1471_;
  assign new_n13332_ = ~new_n1439_;
  assign new_n13333_ = ~new_n1438_;
  assign new_n13334_ = ~new_n1437_;
  assign new_n13335_ = ~new_n1436_;
  assign new_n13336_ = ~new_n1468_;
  assign new_n13337_ = ~new_n1467_;
  assign new_n13338_ = ~new_n1466_;
  assign new_n13339_ = ~new_n1465_;
  assign new_n13340_ = ~new_n1429_;
  assign new_n13341_ = ~new_n1428_;
  assign new_n13342_ = ~new_n1432_;
  assign new_n13343_ = ~new_n1433_;
  assign new_n13344_ = ~new_n1430_;
  assign new_n13345_ = ~new_n1431_;
  assign new_n13346_ = ~new_n1461_;
  assign new_n13347_ = ~new_n1462_;
  assign new_n13348_ = ~new_n1489_;
  assign new_n13349_ = new_n13290_ & new_n1458_;
  assign new_n13350_ = new_n13455_ & new_n13456_;
  assign new_n13351_ = new_n1479_ & new_n13307_;
  assign new_n13352_ = new_n1480_ & new_n13310_;
  assign new_n13353_ = new_n13396_ & new_n13397_ & new_n13399_ & new_n13398_;
  assign new_n13354_ = new_n13401_ & new_n13402_ & new_n13403_;
  assign new_n13355_ = new_n1486_ & new_n13315_;
  assign new_n13356_ = new_n13357_ & new_n13404_;
  assign new_n13357_ = new_n13416_ & new_n13415_;
  assign new_n13358_ = new_n13393_ & new_n13392_;
  assign new_n13359_ = new_n13280_ & new_n13358_;
  assign new_n13360_ = new_n13362_ & new_n13419_ & new_n13418_;
  assign new_n13361_ = new_n13422_ & new_n13421_;
  assign new_n13362_ = new_n13361_ & new_n13281_;
  assign new_n13363_ = new_n1445_ & new_n13323_;
  assign new_n13364_ = new_n1444_ & new_n13303_;
  assign new_n13365_ = new_n13366_ & new_n13424_ & new_n13425_;
  assign new_n13366_ = new_n13428_ & new_n13427_;
  assign new_n13367_ = new_n13279_ & new_n13368_;
  assign new_n13368_ = new_n13436_ & new_n13437_;
  assign new_n13369_ = new_n1439_ & new_n13331_;
  assign new_n13370_ = new_n1438_ & new_n13299_;
  assign new_n13371_ = new_n13372_ & new_n13439_ & new_n13441_;
  assign new_n13372_ = new_n13443_ & new_n13442_;
  assign new_n13373_ = new_n13451_ & new_n13452_;
  assign new_n13374_ = new_n1432_ & new_n13295_;
  assign new_n13375_ = new_n1433_ & new_n13339_;
  assign new_n13376_ = new_n13456_ & new_n13378_ & new_n13458_ & new_n13453_ & new_n13457_;
  assign new_n13377_ = new_n13462_ & new_n13461_;
  assign new_n13378_ = new_n13377_ & new_n13460_ & new_n13459_;
  assign new_n13379_ = new_n13467_ & new_n13468_ & new_n13466_;
  assign new_n13380_ = new_n13473_ & new_n13285_;
  assign new_n13381_ = ~new_n1456_;
  assign new_n13382_ = ~new_n1434_ | ~new_n13338_;
  assign new_n13383_ = ~new_n1463_ | ~new_n13345_;
  assign new_n13384_ = ~new_n1464_ | ~new_n13342_;
  assign new_n13385_ = ~new_n1435_ | ~new_n13337_;
  assign new_n13386_ = ~new_n1440_ | ~new_n13330_;
  assign new_n13387_ = ~new_n1470_ | ~new_n13333_;
  assign new_n13388_ = ~new_n1469_ | ~new_n13334_;
  assign new_n13389_ = ~new_n1441_ | ~new_n13329_;
  assign new_n13390_ = ~new_n1446_ | ~new_n13322_;
  assign new_n13391_ = ~new_n1447_ | ~new_n13306_;
  assign new_n13392_ = ~new_n1449_ | ~new_n13321_;
  assign new_n13393_ = ~new_n1448_ | ~new_n13308_;
  assign new_n13394_ = ~new_n1476_ | ~new_n13326_;
  assign new_n13395_ = ~new_n1475_ | ~new_n13325_;
  assign new_n13396_ = ~new_n1451_ | ~new_n13319_;
  assign new_n13397_ = ~new_n1450_ | ~new_n13320_;
  assign new_n13398_ = ~new_n1453_ | ~new_n13317_;
  assign new_n13399_ = ~new_n1452_ | ~new_n13318_;
  assign new_n13400_ = ~new_n1487_ | ~new_n1488_;
  assign new_n13401_ = ~new_n1455_ | ~new_n13400_;
  assign new_n13402_ = new_n1487_ | new_n1488_;
  assign new_n13403_ = ~new_n1454_ | ~new_n13316_;
  assign new_n13404_ = ~new_n13354_ | ~new_n13353_;
  assign new_n13405_ = ~new_n13355_ | ~new_n13398_;
  assign new_n13406_ = ~new_n1485_ | ~new_n13313_;
  assign new_n13407_ = ~new_n13406_ | ~new_n13405_;
  assign new_n13408_ = ~new_n13407_ | ~new_n13399_;
  assign new_n13409_ = ~new_n1484_ | ~new_n13314_;
  assign new_n13410_ = ~new_n13409_ | ~new_n13408_;
  assign new_n13411_ = ~new_n13410_ | ~new_n13396_;
  assign new_n13412_ = ~new_n1483_ | ~new_n13311_;
  assign new_n13413_ = ~new_n13412_ | ~new_n13411_;
  assign new_n13414_ = ~new_n13413_ | ~new_n13397_;
  assign new_n13415_ = ~new_n1482_ | ~new_n13312_;
  assign new_n13416_ = ~new_n1481_ | ~new_n13309_;
  assign new_n13417_ = ~new_n13414_ | ~new_n13356_;
  assign new_n13418_ = ~new_n13351_ | ~new_n13390_;
  assign new_n13419_ = ~new_n13352_ | ~new_n13280_;
  assign new_n13420_ = ~new_n13359_ | ~new_n13417_;
  assign new_n13421_ = ~new_n1478_ | ~new_n13305_;
  assign new_n13422_ = ~new_n1477_ | ~new_n13324_;
  assign new_n13423_ = ~new_n13420_ | ~new_n13360_;
  assign new_n13424_ = ~new_n13363_ | ~new_n13281_;
  assign new_n13425_ = ~new_n1443_ | ~new_n13304_;
  assign new_n13426_ = ~new_n1475_ | ~new_n13325_;
  assign new_n13427_ = ~new_n13364_ | ~new_n13426_;
  assign new_n13428_ = ~new_n1442_ | ~new_n13328_;
  assign new_n13429_ = ~new_n13423_ | ~new_n13365_;
  assign new_n13430_ = ~new_n1474_ | ~new_n13327_;
  assign new_n13431_ = ~new_n13430_ | ~new_n13429_;
  assign new_n13432_ = ~new_n13431_ | ~new_n13389_;
  assign new_n13433_ = ~new_n1473_ | ~new_n13302_;
  assign new_n13434_ = ~new_n13433_ | ~new_n13432_;
  assign new_n13435_ = ~new_n13434_ | ~new_n13386_;
  assign new_n13436_ = ~new_n1472_ | ~new_n13301_;
  assign new_n13437_ = ~new_n1471_ | ~new_n13332_;
  assign new_n13438_ = ~new_n13435_ | ~new_n13367_;
  assign new_n13439_ = ~new_n13369_ | ~new_n13279_;
  assign new_n13440_ = ~new_n1469_ | ~new_n13334_;
  assign new_n13441_ = ~new_n13370_ | ~new_n13440_;
  assign new_n13442_ = ~new_n1437_ | ~new_n13300_;
  assign new_n13443_ = ~new_n1436_ | ~new_n13336_;
  assign new_n13444_ = ~new_n13438_ | ~new_n13371_;
  assign new_n13445_ = ~new_n1468_ | ~new_n13335_;
  assign new_n13446_ = ~new_n13445_ | ~new_n13444_;
  assign new_n13447_ = ~new_n13446_ | ~new_n13385_;
  assign new_n13448_ = ~new_n1467_ | ~new_n13298_;
  assign new_n13449_ = ~new_n13448_ | ~new_n13447_;
  assign new_n13450_ = ~new_n13449_ | ~new_n13382_;
  assign new_n13451_ = ~new_n1466_ | ~new_n13297_;
  assign new_n13452_ = ~new_n1465_ | ~new_n13343_;
  assign new_n13453_ = ~new_n13278_ | ~new_n13373_ | ~new_n13450_;
  assign new_n13454_ = ~new_n1425_ | ~new_n13294_;
  assign new_n13455_ = ~new_n1426_ | ~new_n13289_;
  assign new_n13456_ = ~new_n1427_ | ~new_n13293_;
  assign new_n13457_ = ~new_n1429_ | ~new_n13346_;
  assign new_n13458_ = ~new_n1428_ | ~new_n13292_;
  assign new_n13459_ = ~new_n13374_ | ~new_n13383_;
  assign new_n13460_ = ~new_n13375_ | ~new_n13278_;
  assign new_n13461_ = ~new_n1430_ | ~new_n13347_;
  assign new_n13462_ = ~new_n1431_ | ~new_n13296_;
  assign new_n13463_ = ~new_n1460_ | ~new_n13341_;
  assign new_n13464_ = ~new_n1459_ | ~new_n13291_;
  assign new_n13465_ = ~new_n13464_ | ~new_n13463_;
  assign new_n13466_ = ~new_n13454_ | ~new_n13349_ | ~new_n13284_;
  assign new_n13467_ = ~new_n13454_ | ~new_n13350_ | ~new_n13284_ | ~new_n13465_;
  assign new_n13468_ = ~new_n1457_ | ~new_n13284_ | ~new_n13287_;
  assign new_n13469_ = ~new_n1461_ | ~new_n13340_;
  assign new_n13470_ = ~new_n1462_ | ~new_n13344_;
  assign new_n13471_ = ~new_n13470_ | ~new_n13469_;
  assign new_n13472_ = ~new_n13454_ | ~new_n13284_ | ~new_n13283_;
  assign new_n13473_ = ~new_n13454_ | ~new_n13284_ | ~new_n13282_;
  assign new_n13474_ = ~new_n1424_ | ~new_n13381_;
  assign new_n13475_ = ~new_n1456_ | ~new_n13288_;
  assign new_n13476_ = ~new_n13381_ | ~new_n1489_ | ~new_n1424_;
  assign new_n13477_ = ~new_n1456_ | ~new_n13348_ | ~new_n13288_;
  assign new_n13478_ = new_n13650_ & new_n13649_;
  assign new_n13479_ = new_n13651_ & new_n13652_;
  assign new_n13480_ = new_n13668_ & new_n13667_;
  assign new_n13481_ = new_n13708_ & new_n13707_;
  assign new_n13482_ = new_n13717_ & new_n13716_;
  assign new_n13483_ = new_n13735_ & new_n13734_;
  assign new_n13484_ = new_n13743_ & new_n13742_;
  assign new_n13485_ = new_n13822_ & new_n13819_;
  assign new_n13486_ = new_n13815_ & new_n13812_;
  assign new_n13487_ = new_n13806_ & new_n13803_;
  assign new_n13488_ = new_n13797_ & new_n13794_;
  assign new_n13489_ = new_n13791_ & new_n13789_;
  assign new_n13490_ = new_n13784_ & new_n13781_;
  assign new_n13491_ = new_n13706_ & new_n13703_;
  assign new_n13492_ = new_n13698_ & new_n13695_;
  assign new_n13493_ = new_n13684_ & new_n13681_;
  assign new_n13494_ = ~new_n1810_;
  assign new_n13495_ = ~new_n1408_;
  assign new_n13496_ = ~new_n1407_;
  assign new_n13497_ = ~new_n1408_ | ~new_n1810_;
  assign new_n13498_ = ~new_n1813_;
  assign new_n13499_ = ~new_n1804_;
  assign new_n13500_ = ~new_n1397_;
  assign new_n13501_ = ~new_n1404_;
  assign new_n13502_ = ~new_n1798_;
  assign new_n13503_ = ~new_n1405_;
  assign new_n13504_ = ~new_n1790_;
  assign new_n13505_ = ~new_n1414_;
  assign new_n13506_ = ~new_n1414_ | ~new_n1790_;
  assign new_n13507_ = ~new_n1801_;
  assign new_n13508_ = ~new_n1401_;
  assign new_n13509_ = ~new_n1397_ | ~new_n1804_;
  assign new_n13510_ = ~new_n1807_;
  assign new_n13511_ = ~new_n1816_;
  assign new_n13512_ = ~new_n1421_;
  assign new_n13513_ = ~new_n1420_;
  assign new_n13514_ = ~new_n1819_;
  assign new_n13515_ = ~new_n13536_ | ~new_n13676_;
  assign new_n13516_ = ~new_n13592_ | ~new_n13664_;
  assign new_n13517_ = ~new_n13653_ | ~new_n13654_;
  assign new_n13518_ = ~new_n1795_ | ~new_n1415_;
  assign new_n13519_ = ~new_n13596_ | ~new_n13690_;
  assign new_n13520_ = ~new_n13687_ | ~new_n13686_;
  assign new_n13521_ = ~new_n2347_;
  assign new_n13522_ = ~new_n1390_;
  assign new_n13523_ = ~new_n1394_;
  assign new_n13524_ = ~new_n2348_;
  assign new_n13525_ = ~new_n2349_;
  assign new_n13526_ = ~new_n1395_;
  assign new_n13527_ = ~new_n2350_;
  assign new_n13528_ = ~new_n1402_;
  assign new_n13529_ = ~new_n2353_;
  assign new_n13530_ = ~new_n1412_;
  assign new_n13531_ = ~new_n1840_;
  assign new_n13532_ = ~new_n1410_;
  assign new_n13533_ = ~new_n1406_;
  assign new_n13534_ = ~new_n1410_ | ~new_n1840_;
  assign new_n13535_ = ~new_n1843_;
  assign new_n13536_ = ~new_n1421_ | ~new_n1816_;
  assign new_n13537_ = ~new_n1822_;
  assign new_n13538_ = ~new_n1399_;
  assign new_n13539_ = ~new_n1828_;
  assign new_n13540_ = ~new_n1409_;
  assign new_n13541_ = ~new_n1825_;
  assign new_n13542_ = ~new_n1400_;
  assign new_n13543_ = ~new_n1400_ | ~new_n1825_;
  assign new_n13544_ = ~new_n1831_;
  assign new_n13545_ = ~new_n1417_;
  assign new_n13546_ = ~new_n1834_;
  assign new_n13547_ = ~new_n1416_;
  assign new_n13548_ = ~new_n1837_;
  assign new_n13549_ = ~new_n1411_;
  assign new_n13550_ = ~new_n1846_;
  assign new_n13551_ = ~new_n1419_;
  assign new_n13552_ = ~new_n1419_ | ~new_n1846_;
  assign new_n13553_ = ~new_n1848_;
  assign new_n13554_ = ~new_n1418_;
  assign new_n13555_ = ~new_n1418_ | ~new_n1848_;
  assign new_n13556_ = ~new_n2354_;
  assign new_n13557_ = ~new_n2352_;
  assign new_n13558_ = ~new_n1398_;
  assign new_n13559_ = ~new_n2351_;
  assign new_n13560_ = ~new_n1403_;
  assign new_n13561_ = ~new_n2348_ | ~new_n1394_;
  assign new_n13562_ = ~new_n1391_;
  assign new_n13563_ = ~new_n2346_;
  assign new_n13564_ = ~new_n13777_ | ~new_n13647_;
  assign new_n13565_ = ~new_n1413_;
  assign new_n13566_ = ~new_n13552_ | ~new_n13786_;
  assign new_n13567_ = ~new_n13732_ | ~new_n13731_;
  assign new_n13568_ = ~new_n13543_ | ~new_n13808_;
  assign new_n13569_ = ~new_n13928_ | ~new_n13927_;
  assign new_n13570_ = ~new_n13975_ | ~new_n13974_;
  assign new_n13571_ = ~new_n13846_ | ~new_n13845_;
  assign new_n13572_ = ~new_n13851_ | ~new_n13850_;
  assign new_n13573_ = ~new_n13858_ | ~new_n13857_;
  assign new_n13574_ = ~new_n13865_ | ~new_n13864_;
  assign new_n13575_ = ~new_n13870_ | ~new_n13869_;
  assign new_n13576_ = ~new_n13879_ | ~new_n13878_;
  assign new_n13577_ = ~new_n13886_ | ~new_n13885_;
  assign new_n13578_ = ~new_n13893_ | ~new_n13892_;
  assign new_n13579_ = ~new_n13900_ | ~new_n13899_;
  assign new_n13580_ = ~new_n13905_ | ~new_n13904_;
  assign new_n13581_ = ~new_n13912_ | ~new_n13911_;
  assign new_n13582_ = ~new_n13919_ | ~new_n13918_;
  assign new_n13583_ = ~new_n13933_ | ~new_n13932_;
  assign new_n13584_ = ~new_n13938_ | ~new_n13937_;
  assign new_n13585_ = ~new_n13945_ | ~new_n13944_;
  assign new_n13586_ = ~new_n13952_ | ~new_n13951_;
  assign new_n13587_ = ~new_n13959_ | ~new_n13958_;
  assign new_n13588_ = ~new_n13966_ | ~new_n13965_;
  assign new_n13589_ = ~new_n13971_ | ~new_n13970_;
  assign new_n13590_ = new_n1798_ & new_n1405_;
  assign new_n13591_ = new_n13660_ & new_n13658_;
  assign new_n13592_ = new_n13665_ & new_n13663_;
  assign new_n13593_ = new_n13672_ & new_n13671_;
  assign new_n13594_ = new_n13497_ & new_n13853_ & new_n13852_;
  assign new_n13595_ = new_n13683_ & new_n13480_;
  assign new_n13596_ = new_n13691_ & new_n13689_;
  assign new_n13597_ = new_n13509_ & new_n13860_ & new_n13859_;
  assign new_n13598_ = new_n13697_ & new_n13478_;
  assign new_n13599_ = new_n13705_ & new_n13652_;
  assign new_n13600_ = new_n13675_ & new_n13481_;
  assign new_n13601_ = new_n13710_ & new_n13642_;
  assign new_n13602_ = new_n13719_ & new_n13643_;
  assign new_n13603_ = new_n13739_ & new_n13738_;
  assign new_n13604_ = new_n13484_ & new_n13753_;
  assign new_n13605_ = new_n13756_ & new_n13751_;
  assign new_n13606_ = new_n13772_ & new_n13769_;
  assign new_n13607_ = new_n13839_ & new_n13773_;
  assign new_n13608_ = new_n13630_ & new_n13749_;
  assign new_n13609_ = new_n13534_ & new_n13940_ & new_n13939_;
  assign new_n13610_ = new_n13643_ & new_n13961_ & new_n13960_;
  assign new_n13611_ = new_n13814_ & new_n13482_;
  assign new_n13612_ = new_n13642_ & new_n13973_ & new_n13972_;
  assign new_n13613_ = new_n13821_ & new_n13481_;
  assign new_n13614_ = ~new_n13593_ | ~new_n13673_;
  assign new_n13615_ = ~new_n13688_ | ~new_n13700_;
  assign new_n13616_ = ~new_n1392_;
  assign new_n13617_ = ~new_n2357_;
  assign new_n13618_ = new_n13874_ & new_n13873_;
  assign new_n13619_ = ~new_n13835_ | ~new_n13775_ | ~new_n13640_;
  assign new_n13620_ = new_n13881_ & new_n13880_;
  assign new_n13621_ = ~new_n13607_ | ~new_n13841_ | ~new_n13840_;
  assign new_n13622_ = new_n13888_ & new_n13887_;
  assign new_n13623_ = ~new_n13561_ | ~new_n13836_ | ~new_n13770_;
  assign new_n13624_ = new_n13895_ & new_n13894_;
  assign new_n13625_ = ~new_n13764_ | ~new_n13763_;
  assign new_n13626_ = new_n13907_ & new_n13906_;
  assign new_n13627_ = ~new_n13760_ | ~new_n13759_;
  assign new_n13628_ = new_n13914_ & new_n13913_;
  assign new_n13629_ = ~new_n13605_ | ~new_n13755_;
  assign new_n13630_ = new_n13921_ & new_n13920_;
  assign new_n13631_ = new_n13926_ & new_n13925_;
  assign new_n13632_ = ~new_n13518_ | ~new_n13798_;
  assign new_n13633_ = ~new_n13603_ | ~new_n13740_;
  assign new_n13634_ = new_n13947_ & new_n13946_;
  assign new_n13635_ = ~new_n13728_ | ~new_n13727_;
  assign new_n13636_ = new_n13954_ & new_n13953_;
  assign new_n13637_ = ~new_n13724_ | ~new_n13723_;
  assign new_n13638_ = ~new_n13714_ | ~new_n13713_;
  assign new_n13639_ = ~new_n13838_ | ~new_n13837_;
  assign new_n13640_ = ~new_n1391_ | ~new_n13621_;
  assign new_n13641_ = ~new_n13509_;
  assign new_n13642_ = ~new_n1819_ | ~new_n1420_;
  assign new_n13643_ = ~new_n1409_ | ~new_n1828_;
  assign new_n13644_ = ~new_n1395_ | ~new_n2349_;
  assign new_n13645_ = ~new_n13543_;
  assign new_n13646_ = ~new_n13552_;
  assign new_n13647_ = ~new_n1402_ | ~new_n2350_;
  assign new_n13648_ = ~new_n13536_;
  assign new_n13649_ = new_n1404_ | new_n1807_;
  assign new_n13650_ = new_n1397_ | new_n1804_;
  assign new_n13651_ = new_n1801_ | new_n1401_;
  assign new_n13652_ = new_n1798_ | new_n1405_;
  assign new_n13653_ = ~new_n13506_;
  assign new_n13654_ = new_n1795_ | new_n1415_;
  assign new_n13655_ = ~new_n13517_;
  assign new_n13656_ = ~new_n13518_;
  assign new_n13657_ = ~new_n13517_ | ~new_n13518_;
  assign new_n13658_ = ~new_n13590_ | ~new_n13651_;
  assign new_n13659_ = ~new_n13479_ | ~new_n13657_;
  assign new_n13660_ = ~new_n1401_ | ~new_n1801_;
  assign new_n13661_ = ~new_n13591_ | ~new_n13659_;
  assign new_n13662_ = ~new_n13510_ | ~new_n13509_;
  assign new_n13663_ = ~new_n1404_ | ~new_n13662_;
  assign new_n13664_ = ~new_n13478_ | ~new_n13661_;
  assign new_n13665_ = ~new_n1807_ | ~new_n13641_;
  assign new_n13666_ = ~new_n13516_;
  assign new_n13667_ = new_n1407_ | new_n1813_;
  assign new_n13668_ = new_n1408_ | new_n1810_;
  assign new_n13669_ = ~new_n13497_;
  assign new_n13670_ = ~new_n13498_ | ~new_n13497_;
  assign new_n13671_ = ~new_n1407_ | ~new_n13670_;
  assign new_n13672_ = ~new_n1813_ | ~new_n13669_;
  assign new_n13673_ = ~new_n13480_ | ~new_n13516_;
  assign new_n13674_ = ~new_n13614_;
  assign new_n13675_ = new_n1816_ | new_n1421_;
  assign new_n13676_ = ~new_n13675_ | ~new_n13614_;
  assign new_n13677_ = ~new_n13515_;
  assign new_n13678_ = new_n1420_ | new_n1819_;
  assign new_n13679_ = new_n1810_ | new_n1408_;
  assign new_n13680_ = ~new_n13679_ | ~new_n13516_;
  assign new_n13681_ = ~new_n13594_ | ~new_n13680_;
  assign new_n13682_ = ~new_n13666_ | ~new_n13497_;
  assign new_n13683_ = ~new_n1813_ | ~new_n1407_;
  assign new_n13684_ = ~new_n13595_ | ~new_n13682_;
  assign new_n13685_ = new_n1408_ | new_n1810_;
  assign new_n13686_ = ~new_n13656_ | ~new_n13652_;
  assign new_n13687_ = ~new_n1405_ | ~new_n1798_;
  assign new_n13688_ = ~new_n13520_;
  assign new_n13689_ = ~new_n13655_ | ~new_n13479_;
  assign new_n13690_ = ~new_n13520_ | ~new_n13651_;
  assign new_n13691_ = ~new_n1401_ | ~new_n1801_;
  assign new_n13692_ = ~new_n13519_;
  assign new_n13693_ = new_n1804_ | new_n1397_;
  assign new_n13694_ = ~new_n13693_ | ~new_n13519_;
  assign new_n13695_ = ~new_n13597_ | ~new_n13694_;
  assign new_n13696_ = ~new_n13692_ | ~new_n13509_;
  assign new_n13697_ = ~new_n1807_ | ~new_n1404_;
  assign new_n13698_ = ~new_n13598_ | ~new_n13696_;
  assign new_n13699_ = new_n1397_ | new_n1804_;
  assign new_n13700_ = ~new_n13655_ | ~new_n13652_;
  assign new_n13701_ = ~new_n13615_;
  assign new_n13702_ = ~new_n1401_ | ~new_n1801_;
  assign new_n13703_ = ~new_n13517_ | ~new_n13518_ | ~new_n13872_ | ~new_n13871_;
  assign new_n13704_ = ~new_n13518_ | ~new_n13517_;
  assign new_n13705_ = ~new_n1405_ | ~new_n1798_;
  assign new_n13706_ = ~new_n13599_ | ~new_n13704_;
  assign new_n13707_ = new_n1420_ | new_n1819_;
  assign new_n13708_ = new_n1399_ | new_n1822_;
  assign new_n13709_ = ~new_n13648_ | ~new_n13481_;
  assign new_n13710_ = ~new_n1399_ | ~new_n1822_;
  assign new_n13711_ = ~new_n13601_ | ~new_n13709_;
  assign new_n13712_ = new_n1822_ | new_n1399_;
  assign new_n13713_ = ~new_n13600_ | ~new_n13614_;
  assign new_n13714_ = ~new_n13712_ | ~new_n13711_;
  assign new_n13715_ = ~new_n13638_;
  assign new_n13716_ = new_n1417_ | new_n1831_;
  assign new_n13717_ = new_n1409_ | new_n1828_;
  assign new_n13718_ = ~new_n13645_ | ~new_n13482_;
  assign new_n13719_ = ~new_n1417_ | ~new_n1831_;
  assign new_n13720_ = ~new_n13602_ | ~new_n13718_;
  assign new_n13721_ = new_n1825_ | new_n1400_;
  assign new_n13722_ = new_n1831_ | new_n1417_;
  assign new_n13723_ = ~new_n13482_ | ~new_n13721_ | ~new_n13638_;
  assign new_n13724_ = ~new_n13722_ | ~new_n13720_;
  assign new_n13725_ = ~new_n13637_;
  assign new_n13726_ = new_n1834_ | new_n1416_;
  assign new_n13727_ = ~new_n13726_ | ~new_n13637_;
  assign new_n13728_ = ~new_n1416_ | ~new_n1834_;
  assign new_n13729_ = ~new_n13635_;
  assign new_n13730_ = new_n1837_ | new_n1411_;
  assign new_n13731_ = ~new_n13730_ | ~new_n13635_;
  assign new_n13732_ = ~new_n1411_ | ~new_n1837_;
  assign new_n13733_ = ~new_n13567_;
  assign new_n13734_ = new_n1406_ | new_n1843_;
  assign new_n13735_ = new_n1410_ | new_n1840_;
  assign new_n13736_ = ~new_n13534_;
  assign new_n13737_ = ~new_n13535_ | ~new_n13534_;
  assign new_n13738_ = ~new_n1406_ | ~new_n13737_;
  assign new_n13739_ = ~new_n1843_ | ~new_n13736_;
  assign new_n13740_ = ~new_n13483_ | ~new_n13567_;
  assign new_n13741_ = ~new_n13633_;
  assign new_n13742_ = new_n1413_ | new_n2354_;
  assign new_n13743_ = new_n1418_ | new_n1848_;
  assign new_n13744_ = new_n1412_ | new_n2353_;
  assign new_n13745_ = ~new_n13555_;
  assign new_n13746_ = ~new_n2354_ | ~new_n13745_;
  assign new_n13747_ = ~new_n13746_ | ~new_n13565_;
  assign new_n13748_ = ~new_n13555_ | ~new_n13556_;
  assign new_n13749_ = ~new_n13748_ | ~new_n13747_;
  assign new_n13750_ = ~new_n13646_ | ~new_n13484_;
  assign new_n13751_ = ~new_n1412_ | ~new_n2353_;
  assign new_n13752_ = ~new_n13749_ | ~new_n13750_;
  assign new_n13753_ = new_n1846_ | new_n1419_;
  assign new_n13754_ = new_n2353_ | new_n1412_;
  assign new_n13755_ = ~new_n13604_ | ~new_n13744_ | ~new_n13633_;
  assign new_n13756_ = ~new_n13754_ | ~new_n13752_;
  assign new_n13757_ = ~new_n13629_;
  assign new_n13758_ = new_n2352_ | new_n1398_;
  assign new_n13759_ = ~new_n13758_ | ~new_n13629_;
  assign new_n13760_ = ~new_n1398_ | ~new_n2352_;
  assign new_n13761_ = ~new_n13627_;
  assign new_n13762_ = new_n2351_ | new_n1403_;
  assign new_n13763_ = ~new_n13762_ | ~new_n13627_;
  assign new_n13764_ = ~new_n1403_ | ~new_n2351_;
  assign new_n13765_ = ~new_n13625_;
  assign new_n13766_ = new_n1395_ | new_n2349_;
  assign new_n13767_ = ~new_n13647_ | ~new_n13644_;
  assign new_n13768_ = ~new_n13561_;
  assign new_n13769_ = new_n2350_ | new_n1402_;
  assign new_n13770_ = ~new_n13639_ | ~new_n13625_ | ~new_n13769_;
  assign new_n13771_ = ~new_n13623_;
  assign new_n13772_ = new_n2347_ | new_n1390_;
  assign new_n13773_ = ~new_n1390_ | ~new_n2347_;
  assign new_n13774_ = ~new_n13621_;
  assign new_n13775_ = ~new_n2346_ | ~new_n13621_;
  assign new_n13776_ = ~new_n13619_;
  assign new_n13777_ = ~new_n13769_ | ~new_n13625_;
  assign new_n13778_ = ~new_n13564_;
  assign new_n13779_ = new_n2349_ | new_n1395_;
  assign new_n13780_ = ~new_n13779_ | ~new_n13564_;
  assign new_n13781_ = ~new_n13624_ | ~new_n13780_ | ~new_n13644_;
  assign new_n13782_ = ~new_n13778_ | ~new_n13644_;
  assign new_n13783_ = ~new_n2348_ | ~new_n1394_;
  assign new_n13784_ = ~new_n13639_ | ~new_n13782_ | ~new_n13783_;
  assign new_n13785_ = new_n1395_ | new_n2349_;
  assign new_n13786_ = ~new_n13753_ | ~new_n13633_;
  assign new_n13787_ = ~new_n13566_;
  assign new_n13788_ = ~new_n13484_ | ~new_n13566_;
  assign new_n13789_ = ~new_n13608_ | ~new_n13788_;
  assign new_n13790_ = ~new_n13788_ | ~new_n13749_;
  assign new_n13791_ = ~new_n13924_ | ~new_n13790_;
  assign new_n13792_ = new_n1848_ | new_n1418_;
  assign new_n13793_ = ~new_n13792_ | ~new_n13566_;
  assign new_n13794_ = ~new_n13631_ | ~new_n13793_ | ~new_n13555_;
  assign new_n13795_ = ~new_n13787_ | ~new_n13555_;
  assign new_n13796_ = ~new_n1413_ | ~new_n2354_;
  assign new_n13797_ = ~new_n13484_ | ~new_n13796_ | ~new_n13795_;
  assign new_n13798_ = new_n1795_ | new_n1415_;
  assign new_n13799_ = ~new_n13632_;
  assign new_n13800_ = new_n1418_ | new_n1848_;
  assign new_n13801_ = new_n1840_ | new_n1410_;
  assign new_n13802_ = ~new_n13801_ | ~new_n13567_;
  assign new_n13803_ = ~new_n13609_ | ~new_n13802_;
  assign new_n13804_ = ~new_n13733_ | ~new_n13534_;
  assign new_n13805_ = ~new_n1843_ | ~new_n1406_;
  assign new_n13806_ = ~new_n13483_ | ~new_n13805_ | ~new_n13804_;
  assign new_n13807_ = new_n1410_ | new_n1840_;
  assign new_n13808_ = ~new_n13721_ | ~new_n13638_;
  assign new_n13809_ = ~new_n13568_;
  assign new_n13810_ = new_n1828_ | new_n1409_;
  assign new_n13811_ = ~new_n13810_ | ~new_n13568_;
  assign new_n13812_ = ~new_n13610_ | ~new_n13811_;
  assign new_n13813_ = ~new_n13809_ | ~new_n13643_;
  assign new_n13814_ = ~new_n1417_ | ~new_n1831_;
  assign new_n13815_ = ~new_n13611_ | ~new_n13813_;
  assign new_n13816_ = new_n1409_ | new_n1828_;
  assign new_n13817_ = new_n1819_ | new_n1420_;
  assign new_n13818_ = ~new_n13817_ | ~new_n13515_;
  assign new_n13819_ = ~new_n13612_ | ~new_n13818_;
  assign new_n13820_ = ~new_n13677_ | ~new_n13642_;
  assign new_n13821_ = ~new_n1399_ | ~new_n1822_;
  assign new_n13822_ = ~new_n13613_ | ~new_n13820_;
  assign new_n13823_ = ~new_n13678_ | ~new_n13642_;
  assign new_n13824_ = ~new_n13675_ | ~new_n13536_;
  assign new_n13825_ = ~new_n13685_ | ~new_n13497_;
  assign new_n13826_ = ~new_n13699_ | ~new_n13509_;
  assign new_n13827_ = ~new_n13702_ | ~new_n13651_;
  assign new_n13828_ = ~new_n13785_ | ~new_n13644_;
  assign new_n13829_ = ~new_n13769_ | ~new_n13647_;
  assign new_n13830_ = ~new_n13800_ | ~new_n13555_;
  assign new_n13831_ = ~new_n13753_ | ~new_n13552_;
  assign new_n13832_ = ~new_n13807_ | ~new_n13534_;
  assign new_n13833_ = ~new_n13816_ | ~new_n13643_;
  assign new_n13834_ = ~new_n13721_ | ~new_n13543_;
  assign new_n13835_ = ~new_n2346_ | ~new_n1391_;
  assign new_n13836_ = ~new_n13767_ | ~new_n13639_;
  assign new_n13837_ = ~new_n1394_ | ~new_n13766_;
  assign new_n13838_ = ~new_n2348_ | ~new_n13766_;
  assign new_n13839_ = ~new_n13772_ | ~new_n13767_ | ~new_n13639_;
  assign new_n13840_ = ~new_n13606_ | ~new_n13625_ | ~new_n13639_;
  assign new_n13841_ = ~new_n13768_ | ~new_n13772_;
  assign new_n13842_ = ~new_n1420_ | ~new_n13514_;
  assign new_n13843_ = ~new_n1819_ | ~new_n13513_;
  assign new_n13844_ = ~new_n13843_ | ~new_n13842_;
  assign new_n13845_ = ~new_n13823_ | ~new_n13515_;
  assign new_n13846_ = ~new_n13844_ | ~new_n13677_;
  assign new_n13847_ = ~new_n1421_ | ~new_n13511_;
  assign new_n13848_ = ~new_n1816_ | ~new_n13512_;
  assign new_n13849_ = ~new_n13848_ | ~new_n13847_;
  assign new_n13850_ = ~new_n13824_ | ~new_n13614_;
  assign new_n13851_ = ~new_n13674_ | ~new_n13849_;
  assign new_n13852_ = ~new_n1407_ | ~new_n13498_;
  assign new_n13853_ = ~new_n1813_ | ~new_n13496_;
  assign new_n13854_ = ~new_n1408_ | ~new_n13494_;
  assign new_n13855_ = ~new_n1810_ | ~new_n13495_;
  assign new_n13856_ = ~new_n13855_ | ~new_n13854_;
  assign new_n13857_ = ~new_n13825_ | ~new_n13516_;
  assign new_n13858_ = ~new_n13856_ | ~new_n13666_;
  assign new_n13859_ = ~new_n1404_ | ~new_n13510_;
  assign new_n13860_ = ~new_n1807_ | ~new_n13501_;
  assign new_n13861_ = ~new_n1397_ | ~new_n13499_;
  assign new_n13862_ = ~new_n1804_ | ~new_n13500_;
  assign new_n13863_ = ~new_n13862_ | ~new_n13861_;
  assign new_n13864_ = ~new_n13826_ | ~new_n13519_;
  assign new_n13865_ = ~new_n13863_ | ~new_n13692_;
  assign new_n13866_ = ~new_n1401_ | ~new_n13507_;
  assign new_n13867_ = ~new_n1801_ | ~new_n13508_;
  assign new_n13868_ = ~new_n13867_ | ~new_n13866_;
  assign new_n13869_ = ~new_n13827_ | ~new_n13615_;
  assign new_n13870_ = ~new_n13701_ | ~new_n13868_;
  assign new_n13871_ = ~new_n1405_ | ~new_n13502_;
  assign new_n13872_ = ~new_n1798_ | ~new_n13503_;
  assign new_n13873_ = ~new_n1392_ | ~new_n13617_;
  assign new_n13874_ = ~new_n2357_ | ~new_n13616_;
  assign new_n13875_ = ~new_n1392_ | ~new_n13617_;
  assign new_n13876_ = ~new_n2357_ | ~new_n13616_;
  assign new_n13877_ = ~new_n13876_ | ~new_n13875_;
  assign new_n13878_ = ~new_n13618_ | ~new_n13619_;
  assign new_n13879_ = ~new_n13776_ | ~new_n13877_;
  assign new_n13880_ = ~new_n1391_ | ~new_n13563_;
  assign new_n13881_ = ~new_n2346_ | ~new_n13562_;
  assign new_n13882_ = ~new_n1391_ | ~new_n13563_;
  assign new_n13883_ = ~new_n2346_ | ~new_n13562_;
  assign new_n13884_ = ~new_n13883_ | ~new_n13882_;
  assign new_n13885_ = ~new_n13620_ | ~new_n13621_;
  assign new_n13886_ = ~new_n13774_ | ~new_n13884_;
  assign new_n13887_ = ~new_n1390_ | ~new_n13521_;
  assign new_n13888_ = ~new_n2347_ | ~new_n13522_;
  assign new_n13889_ = ~new_n1390_ | ~new_n13521_;
  assign new_n13890_ = ~new_n2347_ | ~new_n13522_;
  assign new_n13891_ = ~new_n13890_ | ~new_n13889_;
  assign new_n13892_ = ~new_n13622_ | ~new_n13623_;
  assign new_n13893_ = ~new_n13771_ | ~new_n13891_;
  assign new_n13894_ = ~new_n1394_ | ~new_n13524_;
  assign new_n13895_ = ~new_n2348_ | ~new_n13523_;
  assign new_n13896_ = ~new_n1395_ | ~new_n13525_;
  assign new_n13897_ = ~new_n2349_ | ~new_n13526_;
  assign new_n13898_ = ~new_n13897_ | ~new_n13896_;
  assign new_n13899_ = ~new_n13828_ | ~new_n13564_;
  assign new_n13900_ = ~new_n13898_ | ~new_n13778_;
  assign new_n13901_ = ~new_n1402_ | ~new_n13527_;
  assign new_n13902_ = ~new_n2350_ | ~new_n13528_;
  assign new_n13903_ = ~new_n13902_ | ~new_n13901_;
  assign new_n13904_ = ~new_n13829_ | ~new_n13625_;
  assign new_n13905_ = ~new_n13765_ | ~new_n13903_;
  assign new_n13906_ = ~new_n1403_ | ~new_n13559_;
  assign new_n13907_ = ~new_n2351_ | ~new_n13560_;
  assign new_n13908_ = ~new_n1403_ | ~new_n13559_;
  assign new_n13909_ = ~new_n2351_ | ~new_n13560_;
  assign new_n13910_ = ~new_n13909_ | ~new_n13908_;
  assign new_n13911_ = ~new_n13626_ | ~new_n13627_;
  assign new_n13912_ = ~new_n13761_ | ~new_n13910_;
  assign new_n13913_ = ~new_n1398_ | ~new_n13557_;
  assign new_n13914_ = ~new_n2352_ | ~new_n13558_;
  assign new_n13915_ = ~new_n1398_ | ~new_n13557_;
  assign new_n13916_ = ~new_n2352_ | ~new_n13558_;
  assign new_n13917_ = ~new_n13916_ | ~new_n13915_;
  assign new_n13918_ = ~new_n13628_ | ~new_n13629_;
  assign new_n13919_ = ~new_n13757_ | ~new_n13917_;
  assign new_n13920_ = ~new_n1412_ | ~new_n13529_;
  assign new_n13921_ = ~new_n2353_ | ~new_n13530_;
  assign new_n13922_ = ~new_n1412_ | ~new_n13529_;
  assign new_n13923_ = ~new_n2353_ | ~new_n13530_;
  assign new_n13924_ = ~new_n13923_ | ~new_n13922_;
  assign new_n13925_ = ~new_n1413_ | ~new_n13556_;
  assign new_n13926_ = ~new_n2354_ | ~new_n13565_;
  assign new_n13927_ = ~new_n13653_ | ~new_n13632_;
  assign new_n13928_ = ~new_n13799_ | ~new_n13506_;
  assign new_n13929_ = ~new_n1418_ | ~new_n13553_;
  assign new_n13930_ = ~new_n1848_ | ~new_n13554_;
  assign new_n13931_ = ~new_n13930_ | ~new_n13929_;
  assign new_n13932_ = ~new_n13830_ | ~new_n13566_;
  assign new_n13933_ = ~new_n13931_ | ~new_n13787_;
  assign new_n13934_ = ~new_n1419_ | ~new_n13550_;
  assign new_n13935_ = ~new_n1846_ | ~new_n13551_;
  assign new_n13936_ = ~new_n13935_ | ~new_n13934_;
  assign new_n13937_ = ~new_n13831_ | ~new_n13633_;
  assign new_n13938_ = ~new_n13741_ | ~new_n13936_;
  assign new_n13939_ = ~new_n1406_ | ~new_n13535_;
  assign new_n13940_ = ~new_n1843_ | ~new_n13533_;
  assign new_n13941_ = ~new_n1410_ | ~new_n13531_;
  assign new_n13942_ = ~new_n1840_ | ~new_n13532_;
  assign new_n13943_ = ~new_n13942_ | ~new_n13941_;
  assign new_n13944_ = ~new_n13832_ | ~new_n13567_;
  assign new_n13945_ = ~new_n13943_ | ~new_n13733_;
  assign new_n13946_ = ~new_n1411_ | ~new_n13548_;
  assign new_n13947_ = ~new_n1837_ | ~new_n13549_;
  assign new_n13948_ = ~new_n1411_ | ~new_n13548_;
  assign new_n13949_ = ~new_n1837_ | ~new_n13549_;
  assign new_n13950_ = ~new_n13949_ | ~new_n13948_;
  assign new_n13951_ = ~new_n13634_ | ~new_n13635_;
  assign new_n13952_ = ~new_n13729_ | ~new_n13950_;
  assign new_n13953_ = ~new_n1416_ | ~new_n13546_;
  assign new_n13954_ = ~new_n1834_ | ~new_n13547_;
  assign new_n13955_ = ~new_n1416_ | ~new_n13546_;
  assign new_n13956_ = ~new_n1834_ | ~new_n13547_;
  assign new_n13957_ = ~new_n13956_ | ~new_n13955_;
  assign new_n13958_ = ~new_n13636_ | ~new_n13637_;
  assign new_n13959_ = ~new_n13725_ | ~new_n13957_;
  assign new_n13960_ = ~new_n1417_ | ~new_n13544_;
  assign new_n13961_ = ~new_n1831_ | ~new_n13545_;
  assign new_n13962_ = ~new_n1409_ | ~new_n13539_;
  assign new_n13963_ = ~new_n1828_ | ~new_n13540_;
  assign new_n13964_ = ~new_n13963_ | ~new_n13962_;
  assign new_n13965_ = ~new_n13833_ | ~new_n13568_;
  assign new_n13966_ = ~new_n13964_ | ~new_n13809_;
  assign new_n13967_ = ~new_n1400_ | ~new_n13541_;
  assign new_n13968_ = ~new_n1825_ | ~new_n13542_;
  assign new_n13969_ = ~new_n13968_ | ~new_n13967_;
  assign new_n13970_ = ~new_n13834_ | ~new_n13638_;
  assign new_n13971_ = ~new_n13715_ | ~new_n13969_;
  assign new_n13972_ = ~new_n1399_ | ~new_n13537_;
  assign new_n13973_ = ~new_n1822_ | ~new_n13538_;
  assign new_n13974_ = ~new_n1414_ | ~new_n13504_;
  assign new_n13975_ = ~new_n1790_ | ~new_n13505_;
  assign new_n13976_ = new_n14148_ & new_n14147_;
  assign new_n13977_ = new_n14149_ & new_n14150_;
  assign new_n13978_ = new_n14166_ & new_n14165_;
  assign new_n13979_ = new_n14206_ & new_n14205_;
  assign new_n13980_ = new_n14215_ & new_n14214_;
  assign new_n13981_ = new_n14233_ & new_n14232_;
  assign new_n13982_ = new_n14241_ & new_n14240_;
  assign new_n13983_ = new_n14320_ & new_n14317_;
  assign new_n13984_ = new_n14313_ & new_n14310_;
  assign new_n13985_ = new_n14304_ & new_n14301_;
  assign new_n13986_ = new_n14295_ & new_n14292_;
  assign new_n13987_ = new_n14289_ & new_n14287_;
  assign new_n13988_ = new_n14282_ & new_n14279_;
  assign new_n13989_ = new_n14204_ & new_n14201_;
  assign new_n13990_ = new_n14196_ & new_n14193_;
  assign new_n13991_ = new_n14182_ & new_n14179_;
  assign new_n13992_ = ~new_n1810_;
  assign new_n13993_ = ~new_n1408_;
  assign new_n13994_ = ~new_n1407_;
  assign new_n13995_ = ~new_n1408_ | ~new_n1810_;
  assign new_n13996_ = ~new_n1813_;
  assign new_n13997_ = ~new_n1804_;
  assign new_n13998_ = ~new_n1397_;
  assign new_n13999_ = ~new_n1404_;
  assign new_n14000_ = ~new_n1798_;
  assign new_n14001_ = ~new_n1405_;
  assign new_n14002_ = ~new_n1790_;
  assign new_n14003_ = ~new_n1414_;
  assign new_n14004_ = ~new_n1414_ | ~new_n1790_;
  assign new_n14005_ = ~new_n1801_;
  assign new_n14006_ = ~new_n1401_;
  assign new_n14007_ = ~new_n1397_ | ~new_n1804_;
  assign new_n14008_ = ~new_n1807_;
  assign new_n14009_ = ~new_n1816_;
  assign new_n14010_ = ~new_n1421_;
  assign new_n14011_ = ~new_n1420_;
  assign new_n14012_ = ~new_n1819_;
  assign new_n14013_ = ~new_n14034_ | ~new_n14174_;
  assign new_n14014_ = ~new_n14090_ | ~new_n14162_;
  assign new_n14015_ = ~new_n14151_ | ~new_n14152_;
  assign new_n14016_ = ~new_n1795_ | ~new_n1415_;
  assign new_n14017_ = ~new_n14094_ | ~new_n14188_;
  assign new_n14018_ = ~new_n14185_ | ~new_n14184_;
  assign new_n14019_ = ~new_n2347_;
  assign new_n14020_ = ~new_n1390_;
  assign new_n14021_ = ~new_n1394_;
  assign new_n14022_ = ~new_n2348_;
  assign new_n14023_ = ~new_n2349_;
  assign new_n14024_ = ~new_n1395_;
  assign new_n14025_ = ~new_n2350_;
  assign new_n14026_ = ~new_n1402_;
  assign new_n14027_ = ~new_n2353_;
  assign new_n14028_ = ~new_n1412_;
  assign new_n14029_ = ~new_n1840_;
  assign new_n14030_ = ~new_n1410_;
  assign new_n14031_ = ~new_n1406_;
  assign new_n14032_ = ~new_n1410_ | ~new_n1840_;
  assign new_n14033_ = ~new_n1843_;
  assign new_n14034_ = ~new_n1421_ | ~new_n1816_;
  assign new_n14035_ = ~new_n1822_;
  assign new_n14036_ = ~new_n1399_;
  assign new_n14037_ = ~new_n1828_;
  assign new_n14038_ = ~new_n1409_;
  assign new_n14039_ = ~new_n1825_;
  assign new_n14040_ = ~new_n1400_;
  assign new_n14041_ = ~new_n1400_ | ~new_n1825_;
  assign new_n14042_ = ~new_n1831_;
  assign new_n14043_ = ~new_n1417_;
  assign new_n14044_ = ~new_n1834_;
  assign new_n14045_ = ~new_n1416_;
  assign new_n14046_ = ~new_n1837_;
  assign new_n14047_ = ~new_n1411_;
  assign new_n14048_ = ~new_n1846_;
  assign new_n14049_ = ~new_n1419_;
  assign new_n14050_ = ~new_n1419_ | ~new_n1846_;
  assign new_n14051_ = ~new_n1848_;
  assign new_n14052_ = ~new_n1418_;
  assign new_n14053_ = ~new_n1418_ | ~new_n1848_;
  assign new_n14054_ = ~new_n2354_;
  assign new_n14055_ = ~new_n2352_;
  assign new_n14056_ = ~new_n1398_;
  assign new_n14057_ = ~new_n2351_;
  assign new_n14058_ = ~new_n1403_;
  assign new_n14059_ = ~new_n2348_ | ~new_n1394_;
  assign new_n14060_ = ~new_n1391_;
  assign new_n14061_ = ~new_n2346_;
  assign new_n14062_ = ~new_n14275_ | ~new_n14145_;
  assign new_n14063_ = ~new_n1413_;
  assign new_n14064_ = ~new_n14050_ | ~new_n14284_;
  assign new_n14065_ = ~new_n14230_ | ~new_n14229_;
  assign new_n14066_ = ~new_n14041_ | ~new_n14306_;
  assign new_n14067_ = ~new_n14426_ | ~new_n14425_;
  assign new_n14068_ = ~new_n14473_ | ~new_n14472_;
  assign new_n14069_ = ~new_n14344_ | ~new_n14343_;
  assign new_n14070_ = ~new_n14349_ | ~new_n14348_;
  assign new_n14071_ = ~new_n14356_ | ~new_n14355_;
  assign new_n14072_ = ~new_n14363_ | ~new_n14362_;
  assign new_n14073_ = ~new_n14368_ | ~new_n14367_;
  assign new_n14074_ = ~new_n14377_ | ~new_n14376_;
  assign new_n14075_ = ~new_n14384_ | ~new_n14383_;
  assign new_n14076_ = ~new_n14391_ | ~new_n14390_;
  assign new_n14077_ = ~new_n14398_ | ~new_n14397_;
  assign new_n14078_ = ~new_n14403_ | ~new_n14402_;
  assign new_n14079_ = ~new_n14410_ | ~new_n14409_;
  assign new_n14080_ = ~new_n14417_ | ~new_n14416_;
  assign new_n14081_ = ~new_n14431_ | ~new_n14430_;
  assign new_n14082_ = ~new_n14436_ | ~new_n14435_;
  assign new_n14083_ = ~new_n14443_ | ~new_n14442_;
  assign new_n14084_ = ~new_n14450_ | ~new_n14449_;
  assign new_n14085_ = ~new_n14457_ | ~new_n14456_;
  assign new_n14086_ = ~new_n14464_ | ~new_n14463_;
  assign new_n14087_ = ~new_n14469_ | ~new_n14468_;
  assign new_n14088_ = new_n1798_ & new_n1405_;
  assign new_n14089_ = new_n14158_ & new_n14156_;
  assign new_n14090_ = new_n14163_ & new_n14161_;
  assign new_n14091_ = new_n14170_ & new_n14169_;
  assign new_n14092_ = new_n13995_ & new_n14351_ & new_n14350_;
  assign new_n14093_ = new_n14181_ & new_n13978_;
  assign new_n14094_ = new_n14189_ & new_n14187_;
  assign new_n14095_ = new_n14007_ & new_n14358_ & new_n14357_;
  assign new_n14096_ = new_n14195_ & new_n13976_;
  assign new_n14097_ = new_n14203_ & new_n14150_;
  assign new_n14098_ = new_n14173_ & new_n13979_;
  assign new_n14099_ = new_n14208_ & new_n14140_;
  assign new_n14100_ = new_n14217_ & new_n14141_;
  assign new_n14101_ = new_n14237_ & new_n14236_;
  assign new_n14102_ = new_n13982_ & new_n14251_;
  assign new_n14103_ = new_n14254_ & new_n14249_;
  assign new_n14104_ = new_n14270_ & new_n14267_;
  assign new_n14105_ = new_n14337_ & new_n14271_;
  assign new_n14106_ = new_n14128_ & new_n14247_;
  assign new_n14107_ = new_n14032_ & new_n14438_ & new_n14437_;
  assign new_n14108_ = new_n14141_ & new_n14459_ & new_n14458_;
  assign new_n14109_ = new_n14312_ & new_n13980_;
  assign new_n14110_ = new_n14140_ & new_n14471_ & new_n14470_;
  assign new_n14111_ = new_n14319_ & new_n13979_;
  assign new_n14112_ = ~new_n14091_ | ~new_n14171_;
  assign new_n14113_ = ~new_n14186_ | ~new_n14198_;
  assign new_n14114_ = ~new_n1392_;
  assign new_n14115_ = ~new_n2357_;
  assign new_n14116_ = new_n14372_ & new_n14371_;
  assign new_n14117_ = ~new_n14333_ | ~new_n14273_ | ~new_n14138_;
  assign new_n14118_ = new_n14379_ & new_n14378_;
  assign new_n14119_ = ~new_n14105_ | ~new_n14339_ | ~new_n14338_;
  assign new_n14120_ = new_n14386_ & new_n14385_;
  assign new_n14121_ = ~new_n14059_ | ~new_n14334_ | ~new_n14268_;
  assign new_n14122_ = new_n14393_ & new_n14392_;
  assign new_n14123_ = ~new_n14262_ | ~new_n14261_;
  assign new_n14124_ = new_n14405_ & new_n14404_;
  assign new_n14125_ = ~new_n14258_ | ~new_n14257_;
  assign new_n14126_ = new_n14412_ & new_n14411_;
  assign new_n14127_ = ~new_n14103_ | ~new_n14253_;
  assign new_n14128_ = new_n14419_ & new_n14418_;
  assign new_n14129_ = new_n14424_ & new_n14423_;
  assign new_n14130_ = ~new_n14016_ | ~new_n14296_;
  assign new_n14131_ = ~new_n14101_ | ~new_n14238_;
  assign new_n14132_ = new_n14445_ & new_n14444_;
  assign new_n14133_ = ~new_n14226_ | ~new_n14225_;
  assign new_n14134_ = new_n14452_ & new_n14451_;
  assign new_n14135_ = ~new_n14222_ | ~new_n14221_;
  assign new_n14136_ = ~new_n14212_ | ~new_n14211_;
  assign new_n14137_ = ~new_n14336_ | ~new_n14335_;
  assign new_n14138_ = ~new_n1391_ | ~new_n14119_;
  assign new_n14139_ = ~new_n14007_;
  assign new_n14140_ = ~new_n1819_ | ~new_n1420_;
  assign new_n14141_ = ~new_n1409_ | ~new_n1828_;
  assign new_n14142_ = ~new_n1395_ | ~new_n2349_;
  assign new_n14143_ = ~new_n14041_;
  assign new_n14144_ = ~new_n14050_;
  assign new_n14145_ = ~new_n1402_ | ~new_n2350_;
  assign new_n14146_ = ~new_n14034_;
  assign new_n14147_ = new_n1404_ | new_n1807_;
  assign new_n14148_ = new_n1397_ | new_n1804_;
  assign new_n14149_ = new_n1801_ | new_n1401_;
  assign new_n14150_ = new_n1798_ | new_n1405_;
  assign new_n14151_ = ~new_n14004_;
  assign new_n14152_ = new_n1795_ | new_n1415_;
  assign new_n14153_ = ~new_n14015_;
  assign new_n14154_ = ~new_n14016_;
  assign new_n14155_ = ~new_n14015_ | ~new_n14016_;
  assign new_n14156_ = ~new_n14088_ | ~new_n14149_;
  assign new_n14157_ = ~new_n13977_ | ~new_n14155_;
  assign new_n14158_ = ~new_n1401_ | ~new_n1801_;
  assign new_n14159_ = ~new_n14089_ | ~new_n14157_;
  assign new_n14160_ = ~new_n14008_ | ~new_n14007_;
  assign new_n14161_ = ~new_n1404_ | ~new_n14160_;
  assign new_n14162_ = ~new_n13976_ | ~new_n14159_;
  assign new_n14163_ = ~new_n1807_ | ~new_n14139_;
  assign new_n14164_ = ~new_n14014_;
  assign new_n14165_ = new_n1407_ | new_n1813_;
  assign new_n14166_ = new_n1408_ | new_n1810_;
  assign new_n14167_ = ~new_n13995_;
  assign new_n14168_ = ~new_n13996_ | ~new_n13995_;
  assign new_n14169_ = ~new_n1407_ | ~new_n14168_;
  assign new_n14170_ = ~new_n1813_ | ~new_n14167_;
  assign new_n14171_ = ~new_n13978_ | ~new_n14014_;
  assign new_n14172_ = ~new_n14112_;
  assign new_n14173_ = new_n1816_ | new_n1421_;
  assign new_n14174_ = ~new_n14173_ | ~new_n14112_;
  assign new_n14175_ = ~new_n14013_;
  assign new_n14176_ = new_n1420_ | new_n1819_;
  assign new_n14177_ = new_n1810_ | new_n1408_;
  assign new_n14178_ = ~new_n14177_ | ~new_n14014_;
  assign new_n14179_ = ~new_n14092_ | ~new_n14178_;
  assign new_n14180_ = ~new_n14164_ | ~new_n13995_;
  assign new_n14181_ = ~new_n1813_ | ~new_n1407_;
  assign new_n14182_ = ~new_n14093_ | ~new_n14180_;
  assign new_n14183_ = new_n1408_ | new_n1810_;
  assign new_n14184_ = ~new_n14154_ | ~new_n14150_;
  assign new_n14185_ = ~new_n1405_ | ~new_n1798_;
  assign new_n14186_ = ~new_n14018_;
  assign new_n14187_ = ~new_n14153_ | ~new_n13977_;
  assign new_n14188_ = ~new_n14018_ | ~new_n14149_;
  assign new_n14189_ = ~new_n1401_ | ~new_n1801_;
  assign new_n14190_ = ~new_n14017_;
  assign new_n14191_ = new_n1804_ | new_n1397_;
  assign new_n14192_ = ~new_n14191_ | ~new_n14017_;
  assign new_n14193_ = ~new_n14095_ | ~new_n14192_;
  assign new_n14194_ = ~new_n14190_ | ~new_n14007_;
  assign new_n14195_ = ~new_n1807_ | ~new_n1404_;
  assign new_n14196_ = ~new_n14096_ | ~new_n14194_;
  assign new_n14197_ = new_n1397_ | new_n1804_;
  assign new_n14198_ = ~new_n14153_ | ~new_n14150_;
  assign new_n14199_ = ~new_n14113_;
  assign new_n14200_ = ~new_n1401_ | ~new_n1801_;
  assign new_n14201_ = ~new_n14015_ | ~new_n14016_ | ~new_n14370_ | ~new_n14369_;
  assign new_n14202_ = ~new_n14016_ | ~new_n14015_;
  assign new_n14203_ = ~new_n1405_ | ~new_n1798_;
  assign new_n14204_ = ~new_n14097_ | ~new_n14202_;
  assign new_n14205_ = new_n1420_ | new_n1819_;
  assign new_n14206_ = new_n1399_ | new_n1822_;
  assign new_n14207_ = ~new_n14146_ | ~new_n13979_;
  assign new_n14208_ = ~new_n1399_ | ~new_n1822_;
  assign new_n14209_ = ~new_n14099_ | ~new_n14207_;
  assign new_n14210_ = new_n1822_ | new_n1399_;
  assign new_n14211_ = ~new_n14098_ | ~new_n14112_;
  assign new_n14212_ = ~new_n14210_ | ~new_n14209_;
  assign new_n14213_ = ~new_n14136_;
  assign new_n14214_ = new_n1417_ | new_n1831_;
  assign new_n14215_ = new_n1409_ | new_n1828_;
  assign new_n14216_ = ~new_n14143_ | ~new_n13980_;
  assign new_n14217_ = ~new_n1417_ | ~new_n1831_;
  assign new_n14218_ = ~new_n14100_ | ~new_n14216_;
  assign new_n14219_ = new_n1825_ | new_n1400_;
  assign new_n14220_ = new_n1831_ | new_n1417_;
  assign new_n14221_ = ~new_n13980_ | ~new_n14219_ | ~new_n14136_;
  assign new_n14222_ = ~new_n14220_ | ~new_n14218_;
  assign new_n14223_ = ~new_n14135_;
  assign new_n14224_ = new_n1834_ | new_n1416_;
  assign new_n14225_ = ~new_n14224_ | ~new_n14135_;
  assign new_n14226_ = ~new_n1416_ | ~new_n1834_;
  assign new_n14227_ = ~new_n14133_;
  assign new_n14228_ = new_n1837_ | new_n1411_;
  assign new_n14229_ = ~new_n14228_ | ~new_n14133_;
  assign new_n14230_ = ~new_n1411_ | ~new_n1837_;
  assign new_n14231_ = ~new_n14065_;
  assign new_n14232_ = new_n1406_ | new_n1843_;
  assign new_n14233_ = new_n1410_ | new_n1840_;
  assign new_n14234_ = ~new_n14032_;
  assign new_n14235_ = ~new_n14033_ | ~new_n14032_;
  assign new_n14236_ = ~new_n1406_ | ~new_n14235_;
  assign new_n14237_ = ~new_n1843_ | ~new_n14234_;
  assign new_n14238_ = ~new_n13981_ | ~new_n14065_;
  assign new_n14239_ = ~new_n14131_;
  assign new_n14240_ = new_n1413_ | new_n2354_;
  assign new_n14241_ = new_n1418_ | new_n1848_;
  assign new_n14242_ = new_n1412_ | new_n2353_;
  assign new_n14243_ = ~new_n14053_;
  assign new_n14244_ = ~new_n2354_ | ~new_n14243_;
  assign new_n14245_ = ~new_n14244_ | ~new_n14063_;
  assign new_n14246_ = ~new_n14053_ | ~new_n14054_;
  assign new_n14247_ = ~new_n14246_ | ~new_n14245_;
  assign new_n14248_ = ~new_n14144_ | ~new_n13982_;
  assign new_n14249_ = ~new_n1412_ | ~new_n2353_;
  assign new_n14250_ = ~new_n14247_ | ~new_n14248_;
  assign new_n14251_ = new_n1846_ | new_n1419_;
  assign new_n14252_ = new_n2353_ | new_n1412_;
  assign new_n14253_ = ~new_n14102_ | ~new_n14242_ | ~new_n14131_;
  assign new_n14254_ = ~new_n14252_ | ~new_n14250_;
  assign new_n14255_ = ~new_n14127_;
  assign new_n14256_ = new_n2352_ | new_n1398_;
  assign new_n14257_ = ~new_n14256_ | ~new_n14127_;
  assign new_n14258_ = ~new_n1398_ | ~new_n2352_;
  assign new_n14259_ = ~new_n14125_;
  assign new_n14260_ = new_n2351_ | new_n1403_;
  assign new_n14261_ = ~new_n14260_ | ~new_n14125_;
  assign new_n14262_ = ~new_n1403_ | ~new_n2351_;
  assign new_n14263_ = ~new_n14123_;
  assign new_n14264_ = new_n1395_ | new_n2349_;
  assign new_n14265_ = ~new_n14145_ | ~new_n14142_;
  assign new_n14266_ = ~new_n14059_;
  assign new_n14267_ = new_n2350_ | new_n1402_;
  assign new_n14268_ = ~new_n14137_ | ~new_n14123_ | ~new_n14267_;
  assign new_n14269_ = ~new_n14121_;
  assign new_n14270_ = new_n2347_ | new_n1390_;
  assign new_n14271_ = ~new_n1390_ | ~new_n2347_;
  assign new_n14272_ = ~new_n14119_;
  assign new_n14273_ = ~new_n2346_ | ~new_n14119_;
  assign new_n14274_ = ~new_n14117_;
  assign new_n14275_ = ~new_n14267_ | ~new_n14123_;
  assign new_n14276_ = ~new_n14062_;
  assign new_n14277_ = new_n2349_ | new_n1395_;
  assign new_n14278_ = ~new_n14277_ | ~new_n14062_;
  assign new_n14279_ = ~new_n14122_ | ~new_n14278_ | ~new_n14142_;
  assign new_n14280_ = ~new_n14276_ | ~new_n14142_;
  assign new_n14281_ = ~new_n2348_ | ~new_n1394_;
  assign new_n14282_ = ~new_n14137_ | ~new_n14280_ | ~new_n14281_;
  assign new_n14283_ = new_n1395_ | new_n2349_;
  assign new_n14284_ = ~new_n14251_ | ~new_n14131_;
  assign new_n14285_ = ~new_n14064_;
  assign new_n14286_ = ~new_n13982_ | ~new_n14064_;
  assign new_n14287_ = ~new_n14106_ | ~new_n14286_;
  assign new_n14288_ = ~new_n14286_ | ~new_n14247_;
  assign new_n14289_ = ~new_n14422_ | ~new_n14288_;
  assign new_n14290_ = new_n1848_ | new_n1418_;
  assign new_n14291_ = ~new_n14290_ | ~new_n14064_;
  assign new_n14292_ = ~new_n14129_ | ~new_n14291_ | ~new_n14053_;
  assign new_n14293_ = ~new_n14285_ | ~new_n14053_;
  assign new_n14294_ = ~new_n1413_ | ~new_n2354_;
  assign new_n14295_ = ~new_n13982_ | ~new_n14294_ | ~new_n14293_;
  assign new_n14296_ = new_n1795_ | new_n1415_;
  assign new_n14297_ = ~new_n14130_;
  assign new_n14298_ = new_n1418_ | new_n1848_;
  assign new_n14299_ = new_n1840_ | new_n1410_;
  assign new_n14300_ = ~new_n14299_ | ~new_n14065_;
  assign new_n14301_ = ~new_n14107_ | ~new_n14300_;
  assign new_n14302_ = ~new_n14231_ | ~new_n14032_;
  assign new_n14303_ = ~new_n1843_ | ~new_n1406_;
  assign new_n14304_ = ~new_n13981_ | ~new_n14303_ | ~new_n14302_;
  assign new_n14305_ = new_n1410_ | new_n1840_;
  assign new_n14306_ = ~new_n14219_ | ~new_n14136_;
  assign new_n14307_ = ~new_n14066_;
  assign new_n14308_ = new_n1828_ | new_n1409_;
  assign new_n14309_ = ~new_n14308_ | ~new_n14066_;
  assign new_n14310_ = ~new_n14108_ | ~new_n14309_;
  assign new_n14311_ = ~new_n14307_ | ~new_n14141_;
  assign new_n14312_ = ~new_n1417_ | ~new_n1831_;
  assign new_n14313_ = ~new_n14109_ | ~new_n14311_;
  assign new_n14314_ = new_n1409_ | new_n1828_;
  assign new_n14315_ = new_n1819_ | new_n1420_;
  assign new_n14316_ = ~new_n14315_ | ~new_n14013_;
  assign new_n14317_ = ~new_n14110_ | ~new_n14316_;
  assign new_n14318_ = ~new_n14175_ | ~new_n14140_;
  assign new_n14319_ = ~new_n1399_ | ~new_n1822_;
  assign new_n14320_ = ~new_n14111_ | ~new_n14318_;
  assign new_n14321_ = ~new_n14176_ | ~new_n14140_;
  assign new_n14322_ = ~new_n14173_ | ~new_n14034_;
  assign new_n14323_ = ~new_n14183_ | ~new_n13995_;
  assign new_n14324_ = ~new_n14197_ | ~new_n14007_;
  assign new_n14325_ = ~new_n14200_ | ~new_n14149_;
  assign new_n14326_ = ~new_n14283_ | ~new_n14142_;
  assign new_n14327_ = ~new_n14267_ | ~new_n14145_;
  assign new_n14328_ = ~new_n14298_ | ~new_n14053_;
  assign new_n14329_ = ~new_n14251_ | ~new_n14050_;
  assign new_n14330_ = ~new_n14305_ | ~new_n14032_;
  assign new_n14331_ = ~new_n14314_ | ~new_n14141_;
  assign new_n14332_ = ~new_n14219_ | ~new_n14041_;
  assign new_n14333_ = ~new_n2346_ | ~new_n1391_;
  assign new_n14334_ = ~new_n14265_ | ~new_n14137_;
  assign new_n14335_ = ~new_n1394_ | ~new_n14264_;
  assign new_n14336_ = ~new_n2348_ | ~new_n14264_;
  assign new_n14337_ = ~new_n14270_ | ~new_n14265_ | ~new_n14137_;
  assign new_n14338_ = ~new_n14104_ | ~new_n14123_ | ~new_n14137_;
  assign new_n14339_ = ~new_n14266_ | ~new_n14270_;
  assign new_n14340_ = ~new_n1420_ | ~new_n14012_;
  assign new_n14341_ = ~new_n1819_ | ~new_n14011_;
  assign new_n14342_ = ~new_n14341_ | ~new_n14340_;
  assign new_n14343_ = ~new_n14321_ | ~new_n14013_;
  assign new_n14344_ = ~new_n14342_ | ~new_n14175_;
  assign new_n14345_ = ~new_n1421_ | ~new_n14009_;
  assign new_n14346_ = ~new_n1816_ | ~new_n14010_;
  assign new_n14347_ = ~new_n14346_ | ~new_n14345_;
  assign new_n14348_ = ~new_n14322_ | ~new_n14112_;
  assign new_n14349_ = ~new_n14172_ | ~new_n14347_;
  assign new_n14350_ = ~new_n1407_ | ~new_n13996_;
  assign new_n14351_ = ~new_n1813_ | ~new_n13994_;
  assign new_n14352_ = ~new_n1408_ | ~new_n13992_;
  assign new_n14353_ = ~new_n1810_ | ~new_n13993_;
  assign new_n14354_ = ~new_n14353_ | ~new_n14352_;
  assign new_n14355_ = ~new_n14323_ | ~new_n14014_;
  assign new_n14356_ = ~new_n14354_ | ~new_n14164_;
  assign new_n14357_ = ~new_n1404_ | ~new_n14008_;
  assign new_n14358_ = ~new_n1807_ | ~new_n13999_;
  assign new_n14359_ = ~new_n1397_ | ~new_n13997_;
  assign new_n14360_ = ~new_n1804_ | ~new_n13998_;
  assign new_n14361_ = ~new_n14360_ | ~new_n14359_;
  assign new_n14362_ = ~new_n14324_ | ~new_n14017_;
  assign new_n14363_ = ~new_n14361_ | ~new_n14190_;
  assign new_n14364_ = ~new_n1401_ | ~new_n14005_;
  assign new_n14365_ = ~new_n1801_ | ~new_n14006_;
  assign new_n14366_ = ~new_n14365_ | ~new_n14364_;
  assign new_n14367_ = ~new_n14325_ | ~new_n14113_;
  assign new_n14368_ = ~new_n14199_ | ~new_n14366_;
  assign new_n14369_ = ~new_n1405_ | ~new_n14000_;
  assign new_n14370_ = ~new_n1798_ | ~new_n14001_;
  assign new_n14371_ = ~new_n1392_ | ~new_n14115_;
  assign new_n14372_ = ~new_n2357_ | ~new_n14114_;
  assign new_n14373_ = ~new_n1392_ | ~new_n14115_;
  assign new_n14374_ = ~new_n2357_ | ~new_n14114_;
  assign new_n14375_ = ~new_n14374_ | ~new_n14373_;
  assign new_n14376_ = ~new_n14116_ | ~new_n14117_;
  assign new_n14377_ = ~new_n14274_ | ~new_n14375_;
  assign new_n14378_ = ~new_n1391_ | ~new_n14061_;
  assign new_n14379_ = ~new_n2346_ | ~new_n14060_;
  assign new_n14380_ = ~new_n1391_ | ~new_n14061_;
  assign new_n14381_ = ~new_n2346_ | ~new_n14060_;
  assign new_n14382_ = ~new_n14381_ | ~new_n14380_;
  assign new_n14383_ = ~new_n14118_ | ~new_n14119_;
  assign new_n14384_ = ~new_n14272_ | ~new_n14382_;
  assign new_n14385_ = ~new_n1390_ | ~new_n14019_;
  assign new_n14386_ = ~new_n2347_ | ~new_n14020_;
  assign new_n14387_ = ~new_n1390_ | ~new_n14019_;
  assign new_n14388_ = ~new_n2347_ | ~new_n14020_;
  assign new_n14389_ = ~new_n14388_ | ~new_n14387_;
  assign new_n14390_ = ~new_n14120_ | ~new_n14121_;
  assign new_n14391_ = ~new_n14269_ | ~new_n14389_;
  assign new_n14392_ = ~new_n1394_ | ~new_n14022_;
  assign new_n14393_ = ~new_n2348_ | ~new_n14021_;
  assign new_n14394_ = ~new_n1395_ | ~new_n14023_;
  assign new_n14395_ = ~new_n2349_ | ~new_n14024_;
  assign new_n14396_ = ~new_n14395_ | ~new_n14394_;
  assign new_n14397_ = ~new_n14326_ | ~new_n14062_;
  assign new_n14398_ = ~new_n14396_ | ~new_n14276_;
  assign new_n14399_ = ~new_n1402_ | ~new_n14025_;
  assign new_n14400_ = ~new_n2350_ | ~new_n14026_;
  assign new_n14401_ = ~new_n14400_ | ~new_n14399_;
  assign new_n14402_ = ~new_n14327_ | ~new_n14123_;
  assign new_n14403_ = ~new_n14263_ | ~new_n14401_;
  assign new_n14404_ = ~new_n1403_ | ~new_n14057_;
  assign new_n14405_ = ~new_n2351_ | ~new_n14058_;
  assign new_n14406_ = ~new_n1403_ | ~new_n14057_;
  assign new_n14407_ = ~new_n2351_ | ~new_n14058_;
  assign new_n14408_ = ~new_n14407_ | ~new_n14406_;
  assign new_n14409_ = ~new_n14124_ | ~new_n14125_;
  assign new_n14410_ = ~new_n14259_ | ~new_n14408_;
  assign new_n14411_ = ~new_n1398_ | ~new_n14055_;
  assign new_n14412_ = ~new_n2352_ | ~new_n14056_;
  assign new_n14413_ = ~new_n1398_ | ~new_n14055_;
  assign new_n14414_ = ~new_n2352_ | ~new_n14056_;
  assign new_n14415_ = ~new_n14414_ | ~new_n14413_;
  assign new_n14416_ = ~new_n14126_ | ~new_n14127_;
  assign new_n14417_ = ~new_n14255_ | ~new_n14415_;
  assign new_n14418_ = ~new_n1412_ | ~new_n14027_;
  assign new_n14419_ = ~new_n2353_ | ~new_n14028_;
  assign new_n14420_ = ~new_n1412_ | ~new_n14027_;
  assign new_n14421_ = ~new_n2353_ | ~new_n14028_;
  assign new_n14422_ = ~new_n14421_ | ~new_n14420_;
  assign new_n14423_ = ~new_n1413_ | ~new_n14054_;
  assign new_n14424_ = ~new_n2354_ | ~new_n14063_;
  assign new_n14425_ = ~new_n14151_ | ~new_n14130_;
  assign new_n14426_ = ~new_n14297_ | ~new_n14004_;
  assign new_n14427_ = ~new_n1418_ | ~new_n14051_;
  assign new_n14428_ = ~new_n1848_ | ~new_n14052_;
  assign new_n14429_ = ~new_n14428_ | ~new_n14427_;
  assign new_n14430_ = ~new_n14328_ | ~new_n14064_;
  assign new_n14431_ = ~new_n14429_ | ~new_n14285_;
  assign new_n14432_ = ~new_n1419_ | ~new_n14048_;
  assign new_n14433_ = ~new_n1846_ | ~new_n14049_;
  assign new_n14434_ = ~new_n14433_ | ~new_n14432_;
  assign new_n14435_ = ~new_n14329_ | ~new_n14131_;
  assign new_n14436_ = ~new_n14239_ | ~new_n14434_;
  assign new_n14437_ = ~new_n1406_ | ~new_n14033_;
  assign new_n14438_ = ~new_n1843_ | ~new_n14031_;
  assign new_n14439_ = ~new_n1410_ | ~new_n14029_;
  assign new_n14440_ = ~new_n1840_ | ~new_n14030_;
  assign new_n14441_ = ~new_n14440_ | ~new_n14439_;
  assign new_n14442_ = ~new_n14330_ | ~new_n14065_;
  assign new_n14443_ = ~new_n14441_ | ~new_n14231_;
  assign new_n14444_ = ~new_n1411_ | ~new_n14046_;
  assign new_n14445_ = ~new_n1837_ | ~new_n14047_;
  assign new_n14446_ = ~new_n1411_ | ~new_n14046_;
  assign new_n14447_ = ~new_n1837_ | ~new_n14047_;
  assign new_n14448_ = ~new_n14447_ | ~new_n14446_;
  assign new_n14449_ = ~new_n14132_ | ~new_n14133_;
  assign new_n14450_ = ~new_n14227_ | ~new_n14448_;
  assign new_n14451_ = ~new_n1416_ | ~new_n14044_;
  assign new_n14452_ = ~new_n1834_ | ~new_n14045_;
  assign new_n14453_ = ~new_n1416_ | ~new_n14044_;
  assign new_n14454_ = ~new_n1834_ | ~new_n14045_;
  assign new_n14455_ = ~new_n14454_ | ~new_n14453_;
  assign new_n14456_ = ~new_n14134_ | ~new_n14135_;
  assign new_n14457_ = ~new_n14223_ | ~new_n14455_;
  assign new_n14458_ = ~new_n1417_ | ~new_n14042_;
  assign new_n14459_ = ~new_n1831_ | ~new_n14043_;
  assign new_n14460_ = ~new_n1409_ | ~new_n14037_;
  assign new_n14461_ = ~new_n1828_ | ~new_n14038_;
  assign new_n14462_ = ~new_n14461_ | ~new_n14460_;
  assign new_n14463_ = ~new_n14331_ | ~new_n14066_;
  assign new_n14464_ = ~new_n14462_ | ~new_n14307_;
  assign new_n14465_ = ~new_n1400_ | ~new_n14039_;
  assign new_n14466_ = ~new_n1825_ | ~new_n14040_;
  assign new_n14467_ = ~new_n14466_ | ~new_n14465_;
  assign new_n14468_ = ~new_n14332_ | ~new_n14136_;
  assign new_n14469_ = ~new_n14213_ | ~new_n14467_;
  assign new_n14470_ = ~new_n1399_ | ~new_n14035_;
  assign new_n14471_ = ~new_n1822_ | ~new_n14036_;
  assign new_n14472_ = ~new_n1414_ | ~new_n14002_;
  assign new_n14473_ = ~new_n1790_ | ~new_n14003_;
  assign new_n14474_ = new_n14646_ & new_n14645_;
  assign new_n14475_ = new_n14647_ & new_n14648_;
  assign new_n14476_ = new_n14664_ & new_n14663_;
  assign new_n14477_ = new_n14704_ & new_n14703_;
  assign new_n14478_ = new_n14713_ & new_n14712_;
  assign new_n14479_ = new_n14731_ & new_n14730_;
  assign new_n14480_ = new_n14739_ & new_n14738_;
  assign new_n14481_ = new_n14818_ & new_n14815_;
  assign new_n14482_ = new_n14811_ & new_n14808_;
  assign new_n14483_ = new_n14802_ & new_n14799_;
  assign new_n14484_ = new_n14793_ & new_n14790_;
  assign new_n14485_ = new_n14787_ & new_n14785_;
  assign new_n14486_ = new_n14780_ & new_n14777_;
  assign new_n14487_ = new_n14702_ & new_n14699_;
  assign new_n14488_ = new_n14694_ & new_n14691_;
  assign new_n14489_ = new_n14680_ & new_n14677_;
  assign new_n14490_ = ~new_n1810_;
  assign new_n14491_ = ~new_n1408_;
  assign new_n14492_ = ~new_n1407_;
  assign new_n14493_ = ~new_n1408_ | ~new_n1810_;
  assign new_n14494_ = ~new_n1813_;
  assign new_n14495_ = ~new_n1804_;
  assign new_n14496_ = ~new_n1397_;
  assign new_n14497_ = ~new_n1404_;
  assign new_n14498_ = ~new_n1798_;
  assign new_n14499_ = ~new_n1405_;
  assign new_n14500_ = ~new_n1790_;
  assign new_n14501_ = ~new_n1414_;
  assign new_n14502_ = ~new_n1414_ | ~new_n1790_;
  assign new_n14503_ = ~new_n1801_;
  assign new_n14504_ = ~new_n1401_;
  assign new_n14505_ = ~new_n1397_ | ~new_n1804_;
  assign new_n14506_ = ~new_n1807_;
  assign new_n14507_ = ~new_n1816_;
  assign new_n14508_ = ~new_n1421_;
  assign new_n14509_ = ~new_n1420_;
  assign new_n14510_ = ~new_n1819_;
  assign new_n14511_ = ~new_n14532_ | ~new_n14672_;
  assign new_n14512_ = ~new_n14588_ | ~new_n14660_;
  assign new_n14513_ = ~new_n14649_ | ~new_n14650_;
  assign new_n14514_ = ~new_n1795_ | ~new_n1415_;
  assign new_n14515_ = ~new_n14592_ | ~new_n14686_;
  assign new_n14516_ = ~new_n14683_ | ~new_n14682_;
  assign new_n14517_ = ~new_n2347_;
  assign new_n14518_ = ~new_n1390_;
  assign new_n14519_ = ~new_n1394_;
  assign new_n14520_ = ~new_n2348_;
  assign new_n14521_ = ~new_n2349_;
  assign new_n14522_ = ~new_n1395_;
  assign new_n14523_ = ~new_n2350_;
  assign new_n14524_ = ~new_n1402_;
  assign new_n14525_ = ~new_n2353_;
  assign new_n14526_ = ~new_n1412_;
  assign new_n14527_ = ~new_n1840_;
  assign new_n14528_ = ~new_n1410_;
  assign new_n14529_ = ~new_n1406_;
  assign new_n14530_ = ~new_n1410_ | ~new_n1840_;
  assign new_n14531_ = ~new_n1843_;
  assign new_n14532_ = ~new_n1421_ | ~new_n1816_;
  assign new_n14533_ = ~new_n1822_;
  assign new_n14534_ = ~new_n1399_;
  assign new_n14535_ = ~new_n1828_;
  assign new_n14536_ = ~new_n1409_;
  assign new_n14537_ = ~new_n1825_;
  assign new_n14538_ = ~new_n1400_;
  assign new_n14539_ = ~new_n1400_ | ~new_n1825_;
  assign new_n14540_ = ~new_n1831_;
  assign new_n14541_ = ~new_n1417_;
  assign new_n14542_ = ~new_n1834_;
  assign new_n14543_ = ~new_n1416_;
  assign new_n14544_ = ~new_n1837_;
  assign new_n14545_ = ~new_n1411_;
  assign new_n14546_ = ~new_n1846_;
  assign new_n14547_ = ~new_n1419_;
  assign new_n14548_ = ~new_n1419_ | ~new_n1846_;
  assign new_n14549_ = ~new_n1848_;
  assign new_n14550_ = ~new_n1418_;
  assign new_n14551_ = ~new_n1418_ | ~new_n1848_;
  assign new_n14552_ = ~new_n2354_;
  assign new_n14553_ = ~new_n2352_;
  assign new_n14554_ = ~new_n1398_;
  assign new_n14555_ = ~new_n2351_;
  assign new_n14556_ = ~new_n1403_;
  assign new_n14557_ = ~new_n2348_ | ~new_n1394_;
  assign new_n14558_ = ~new_n1391_;
  assign new_n14559_ = ~new_n2346_;
  assign new_n14560_ = ~new_n14773_ | ~new_n14643_;
  assign new_n14561_ = ~new_n1413_;
  assign new_n14562_ = ~new_n14548_ | ~new_n14782_;
  assign new_n14563_ = ~new_n14728_ | ~new_n14727_;
  assign new_n14564_ = ~new_n14539_ | ~new_n14804_;
  assign new_n14565_ = ~new_n14924_ | ~new_n14923_;
  assign new_n14566_ = ~new_n14971_ | ~new_n14970_;
  assign new_n14567_ = ~new_n14842_ | ~new_n14841_;
  assign new_n14568_ = ~new_n14847_ | ~new_n14846_;
  assign new_n14569_ = ~new_n14854_ | ~new_n14853_;
  assign new_n14570_ = ~new_n14861_ | ~new_n14860_;
  assign new_n14571_ = ~new_n14866_ | ~new_n14865_;
  assign new_n14572_ = ~new_n14875_ | ~new_n14874_;
  assign new_n14573_ = ~new_n14882_ | ~new_n14881_;
  assign new_n14574_ = ~new_n14889_ | ~new_n14888_;
  assign new_n14575_ = ~new_n14896_ | ~new_n14895_;
  assign new_n14576_ = ~new_n14901_ | ~new_n14900_;
  assign new_n14577_ = ~new_n14908_ | ~new_n14907_;
  assign new_n14578_ = ~new_n14915_ | ~new_n14914_;
  assign new_n14579_ = ~new_n14929_ | ~new_n14928_;
  assign new_n14580_ = ~new_n14934_ | ~new_n14933_;
  assign new_n14581_ = ~new_n14941_ | ~new_n14940_;
  assign new_n14582_ = ~new_n14948_ | ~new_n14947_;
  assign new_n14583_ = ~new_n14955_ | ~new_n14954_;
  assign new_n14584_ = ~new_n14962_ | ~new_n14961_;
  assign new_n14585_ = ~new_n14967_ | ~new_n14966_;
  assign new_n14586_ = new_n1798_ & new_n1405_;
  assign new_n14587_ = new_n14656_ & new_n14654_;
  assign new_n14588_ = new_n14661_ & new_n14659_;
  assign new_n14589_ = new_n14668_ & new_n14667_;
  assign new_n14590_ = new_n14493_ & new_n14849_ & new_n14848_;
  assign new_n14591_ = new_n14679_ & new_n14476_;
  assign new_n14592_ = new_n14687_ & new_n14685_;
  assign new_n14593_ = new_n14505_ & new_n14856_ & new_n14855_;
  assign new_n14594_ = new_n14693_ & new_n14474_;
  assign new_n14595_ = new_n14701_ & new_n14648_;
  assign new_n14596_ = new_n14671_ & new_n14477_;
  assign new_n14597_ = new_n14706_ & new_n14638_;
  assign new_n14598_ = new_n14715_ & new_n14639_;
  assign new_n14599_ = new_n14735_ & new_n14734_;
  assign new_n14600_ = new_n14480_ & new_n14749_;
  assign new_n14601_ = new_n14752_ & new_n14747_;
  assign new_n14602_ = new_n14768_ & new_n14765_;
  assign new_n14603_ = new_n14835_ & new_n14769_;
  assign new_n14604_ = new_n14626_ & new_n14745_;
  assign new_n14605_ = new_n14530_ & new_n14936_ & new_n14935_;
  assign new_n14606_ = new_n14639_ & new_n14957_ & new_n14956_;
  assign new_n14607_ = new_n14810_ & new_n14478_;
  assign new_n14608_ = new_n14638_ & new_n14969_ & new_n14968_;
  assign new_n14609_ = new_n14817_ & new_n14477_;
  assign new_n14610_ = ~new_n14589_ | ~new_n14669_;
  assign new_n14611_ = ~new_n14684_ | ~new_n14696_;
  assign new_n14612_ = ~new_n1392_;
  assign new_n14613_ = ~new_n2357_;
  assign new_n14614_ = new_n14870_ & new_n14869_;
  assign new_n14615_ = ~new_n14831_ | ~new_n14771_ | ~new_n14636_;
  assign new_n14616_ = new_n14877_ & new_n14876_;
  assign new_n14617_ = ~new_n14603_ | ~new_n14837_ | ~new_n14836_;
  assign new_n14618_ = new_n14884_ & new_n14883_;
  assign new_n14619_ = ~new_n14557_ | ~new_n14832_ | ~new_n14766_;
  assign new_n14620_ = new_n14891_ & new_n14890_;
  assign new_n14621_ = ~new_n14760_ | ~new_n14759_;
  assign new_n14622_ = new_n14903_ & new_n14902_;
  assign new_n14623_ = ~new_n14756_ | ~new_n14755_;
  assign new_n14624_ = new_n14910_ & new_n14909_;
  assign new_n14625_ = ~new_n14601_ | ~new_n14751_;
  assign new_n14626_ = new_n14917_ & new_n14916_;
  assign new_n14627_ = new_n14922_ & new_n14921_;
  assign new_n14628_ = ~new_n14514_ | ~new_n14794_;
  assign new_n14629_ = ~new_n14599_ | ~new_n14736_;
  assign new_n14630_ = new_n14943_ & new_n14942_;
  assign new_n14631_ = ~new_n14724_ | ~new_n14723_;
  assign new_n14632_ = new_n14950_ & new_n14949_;
  assign new_n14633_ = ~new_n14720_ | ~new_n14719_;
  assign new_n14634_ = ~new_n14710_ | ~new_n14709_;
  assign new_n14635_ = ~new_n14834_ | ~new_n14833_;
  assign new_n14636_ = ~new_n1391_ | ~new_n14617_;
  assign new_n14637_ = ~new_n14505_;
  assign new_n14638_ = ~new_n1819_ | ~new_n1420_;
  assign new_n14639_ = ~new_n1409_ | ~new_n1828_;
  assign new_n14640_ = ~new_n1395_ | ~new_n2349_;
  assign new_n14641_ = ~new_n14539_;
  assign new_n14642_ = ~new_n14548_;
  assign new_n14643_ = ~new_n1402_ | ~new_n2350_;
  assign new_n14644_ = ~new_n14532_;
  assign new_n14645_ = new_n1404_ | new_n1807_;
  assign new_n14646_ = new_n1397_ | new_n1804_;
  assign new_n14647_ = new_n1801_ | new_n1401_;
  assign new_n14648_ = new_n1798_ | new_n1405_;
  assign new_n14649_ = ~new_n14502_;
  assign new_n14650_ = new_n1795_ | new_n1415_;
  assign new_n14651_ = ~new_n14513_;
  assign new_n14652_ = ~new_n14514_;
  assign new_n14653_ = ~new_n14513_ | ~new_n14514_;
  assign new_n14654_ = ~new_n14586_ | ~new_n14647_;
  assign new_n14655_ = ~new_n14475_ | ~new_n14653_;
  assign new_n14656_ = ~new_n1401_ | ~new_n1801_;
  assign new_n14657_ = ~new_n14587_ | ~new_n14655_;
  assign new_n14658_ = ~new_n14506_ | ~new_n14505_;
  assign new_n14659_ = ~new_n1404_ | ~new_n14658_;
  assign new_n14660_ = ~new_n14474_ | ~new_n14657_;
  assign new_n14661_ = ~new_n1807_ | ~new_n14637_;
  assign new_n14662_ = ~new_n14512_;
  assign new_n14663_ = new_n1407_ | new_n1813_;
  assign new_n14664_ = new_n1408_ | new_n1810_;
  assign new_n14665_ = ~new_n14493_;
  assign new_n14666_ = ~new_n14494_ | ~new_n14493_;
  assign new_n14667_ = ~new_n1407_ | ~new_n14666_;
  assign new_n14668_ = ~new_n1813_ | ~new_n14665_;
  assign new_n14669_ = ~new_n14476_ | ~new_n14512_;
  assign new_n14670_ = ~new_n14610_;
  assign new_n14671_ = new_n1816_ | new_n1421_;
  assign new_n14672_ = ~new_n14671_ | ~new_n14610_;
  assign new_n14673_ = ~new_n14511_;
  assign new_n14674_ = new_n1420_ | new_n1819_;
  assign new_n14675_ = new_n1810_ | new_n1408_;
  assign new_n14676_ = ~new_n14675_ | ~new_n14512_;
  assign new_n14677_ = ~new_n14590_ | ~new_n14676_;
  assign new_n14678_ = ~new_n14662_ | ~new_n14493_;
  assign new_n14679_ = ~new_n1813_ | ~new_n1407_;
  assign new_n14680_ = ~new_n14591_ | ~new_n14678_;
  assign new_n14681_ = new_n1408_ | new_n1810_;
  assign new_n14682_ = ~new_n14652_ | ~new_n14648_;
  assign new_n14683_ = ~new_n1405_ | ~new_n1798_;
  assign new_n14684_ = ~new_n14516_;
  assign new_n14685_ = ~new_n14651_ | ~new_n14475_;
  assign new_n14686_ = ~new_n14516_ | ~new_n14647_;
  assign new_n14687_ = ~new_n1401_ | ~new_n1801_;
  assign new_n14688_ = ~new_n14515_;
  assign new_n14689_ = new_n1804_ | new_n1397_;
  assign new_n14690_ = ~new_n14689_ | ~new_n14515_;
  assign new_n14691_ = ~new_n14593_ | ~new_n14690_;
  assign new_n14692_ = ~new_n14688_ | ~new_n14505_;
  assign new_n14693_ = ~new_n1807_ | ~new_n1404_;
  assign new_n14694_ = ~new_n14594_ | ~new_n14692_;
  assign new_n14695_ = new_n1397_ | new_n1804_;
  assign new_n14696_ = ~new_n14651_ | ~new_n14648_;
  assign new_n14697_ = ~new_n14611_;
  assign new_n14698_ = ~new_n1401_ | ~new_n1801_;
  assign new_n14699_ = ~new_n14513_ | ~new_n14514_ | ~new_n14868_ | ~new_n14867_;
  assign new_n14700_ = ~new_n14514_ | ~new_n14513_;
  assign new_n14701_ = ~new_n1405_ | ~new_n1798_;
  assign new_n14702_ = ~new_n14595_ | ~new_n14700_;
  assign new_n14703_ = new_n1420_ | new_n1819_;
  assign new_n14704_ = new_n1399_ | new_n1822_;
  assign new_n14705_ = ~new_n14644_ | ~new_n14477_;
  assign new_n14706_ = ~new_n1399_ | ~new_n1822_;
  assign new_n14707_ = ~new_n14597_ | ~new_n14705_;
  assign new_n14708_ = new_n1822_ | new_n1399_;
  assign new_n14709_ = ~new_n14596_ | ~new_n14610_;
  assign new_n14710_ = ~new_n14708_ | ~new_n14707_;
  assign new_n14711_ = ~new_n14634_;
  assign new_n14712_ = new_n1417_ | new_n1831_;
  assign new_n14713_ = new_n1409_ | new_n1828_;
  assign new_n14714_ = ~new_n14641_ | ~new_n14478_;
  assign new_n14715_ = ~new_n1417_ | ~new_n1831_;
  assign new_n14716_ = ~new_n14598_ | ~new_n14714_;
  assign new_n14717_ = new_n1825_ | new_n1400_;
  assign new_n14718_ = new_n1831_ | new_n1417_;
  assign new_n14719_ = ~new_n14478_ | ~new_n14717_ | ~new_n14634_;
  assign new_n14720_ = ~new_n14718_ | ~new_n14716_;
  assign new_n14721_ = ~new_n14633_;
  assign new_n14722_ = new_n1834_ | new_n1416_;
  assign new_n14723_ = ~new_n14722_ | ~new_n14633_;
  assign new_n14724_ = ~new_n1416_ | ~new_n1834_;
  assign new_n14725_ = ~new_n14631_;
  assign new_n14726_ = new_n1837_ | new_n1411_;
  assign new_n14727_ = ~new_n14726_ | ~new_n14631_;
  assign new_n14728_ = ~new_n1411_ | ~new_n1837_;
  assign new_n14729_ = ~new_n14563_;
  assign new_n14730_ = new_n1406_ | new_n1843_;
  assign new_n14731_ = new_n1410_ | new_n1840_;
  assign new_n14732_ = ~new_n14530_;
  assign new_n14733_ = ~new_n14531_ | ~new_n14530_;
  assign new_n14734_ = ~new_n1406_ | ~new_n14733_;
  assign new_n14735_ = ~new_n1843_ | ~new_n14732_;
  assign new_n14736_ = ~new_n14479_ | ~new_n14563_;
  assign new_n14737_ = ~new_n14629_;
  assign new_n14738_ = new_n1413_ | new_n2354_;
  assign new_n14739_ = new_n1418_ | new_n1848_;
  assign new_n14740_ = new_n1412_ | new_n2353_;
  assign new_n14741_ = ~new_n14551_;
  assign new_n14742_ = ~new_n2354_ | ~new_n14741_;
  assign new_n14743_ = ~new_n14742_ | ~new_n14561_;
  assign new_n14744_ = ~new_n14551_ | ~new_n14552_;
  assign new_n14745_ = ~new_n14744_ | ~new_n14743_;
  assign new_n14746_ = ~new_n14642_ | ~new_n14480_;
  assign new_n14747_ = ~new_n1412_ | ~new_n2353_;
  assign new_n14748_ = ~new_n14745_ | ~new_n14746_;
  assign new_n14749_ = new_n1846_ | new_n1419_;
  assign new_n14750_ = new_n2353_ | new_n1412_;
  assign new_n14751_ = ~new_n14600_ | ~new_n14740_ | ~new_n14629_;
  assign new_n14752_ = ~new_n14750_ | ~new_n14748_;
  assign new_n14753_ = ~new_n14625_;
  assign new_n14754_ = new_n2352_ | new_n1398_;
  assign new_n14755_ = ~new_n14754_ | ~new_n14625_;
  assign new_n14756_ = ~new_n1398_ | ~new_n2352_;
  assign new_n14757_ = ~new_n14623_;
  assign new_n14758_ = new_n2351_ | new_n1403_;
  assign new_n14759_ = ~new_n14758_ | ~new_n14623_;
  assign new_n14760_ = ~new_n1403_ | ~new_n2351_;
  assign new_n14761_ = ~new_n14621_;
  assign new_n14762_ = new_n1395_ | new_n2349_;
  assign new_n14763_ = ~new_n14643_ | ~new_n14640_;
  assign new_n14764_ = ~new_n14557_;
  assign new_n14765_ = new_n2350_ | new_n1402_;
  assign new_n14766_ = ~new_n14635_ | ~new_n14621_ | ~new_n14765_;
  assign new_n14767_ = ~new_n14619_;
  assign new_n14768_ = new_n2347_ | new_n1390_;
  assign new_n14769_ = ~new_n1390_ | ~new_n2347_;
  assign new_n14770_ = ~new_n14617_;
  assign new_n14771_ = ~new_n2346_ | ~new_n14617_;
  assign new_n14772_ = ~new_n14615_;
  assign new_n14773_ = ~new_n14765_ | ~new_n14621_;
  assign new_n14774_ = ~new_n14560_;
  assign new_n14775_ = new_n2349_ | new_n1395_;
  assign new_n14776_ = ~new_n14775_ | ~new_n14560_;
  assign new_n14777_ = ~new_n14620_ | ~new_n14776_ | ~new_n14640_;
  assign new_n14778_ = ~new_n14774_ | ~new_n14640_;
  assign new_n14779_ = ~new_n2348_ | ~new_n1394_;
  assign new_n14780_ = ~new_n14635_ | ~new_n14778_ | ~new_n14779_;
  assign new_n14781_ = new_n1395_ | new_n2349_;
  assign new_n14782_ = ~new_n14749_ | ~new_n14629_;
  assign new_n14783_ = ~new_n14562_;
  assign new_n14784_ = ~new_n14480_ | ~new_n14562_;
  assign new_n14785_ = ~new_n14604_ | ~new_n14784_;
  assign new_n14786_ = ~new_n14784_ | ~new_n14745_;
  assign new_n14787_ = ~new_n14920_ | ~new_n14786_;
  assign new_n14788_ = new_n1848_ | new_n1418_;
  assign new_n14789_ = ~new_n14788_ | ~new_n14562_;
  assign new_n14790_ = ~new_n14627_ | ~new_n14789_ | ~new_n14551_;
  assign new_n14791_ = ~new_n14783_ | ~new_n14551_;
  assign new_n14792_ = ~new_n1413_ | ~new_n2354_;
  assign new_n14793_ = ~new_n14480_ | ~new_n14792_ | ~new_n14791_;
  assign new_n14794_ = new_n1795_ | new_n1415_;
  assign new_n14795_ = ~new_n14628_;
  assign new_n14796_ = new_n1418_ | new_n1848_;
  assign new_n14797_ = new_n1840_ | new_n1410_;
  assign new_n14798_ = ~new_n14797_ | ~new_n14563_;
  assign new_n14799_ = ~new_n14605_ | ~new_n14798_;
  assign new_n14800_ = ~new_n14729_ | ~new_n14530_;
  assign new_n14801_ = ~new_n1843_ | ~new_n1406_;
  assign new_n14802_ = ~new_n14479_ | ~new_n14801_ | ~new_n14800_;
  assign new_n14803_ = new_n1410_ | new_n1840_;
  assign new_n14804_ = ~new_n14717_ | ~new_n14634_;
  assign new_n14805_ = ~new_n14564_;
  assign new_n14806_ = new_n1828_ | new_n1409_;
  assign new_n14807_ = ~new_n14806_ | ~new_n14564_;
  assign new_n14808_ = ~new_n14606_ | ~new_n14807_;
  assign new_n14809_ = ~new_n14805_ | ~new_n14639_;
  assign new_n14810_ = ~new_n1417_ | ~new_n1831_;
  assign new_n14811_ = ~new_n14607_ | ~new_n14809_;
  assign new_n14812_ = new_n1409_ | new_n1828_;
  assign new_n14813_ = new_n1819_ | new_n1420_;
  assign new_n14814_ = ~new_n14813_ | ~new_n14511_;
  assign new_n14815_ = ~new_n14608_ | ~new_n14814_;
  assign new_n14816_ = ~new_n14673_ | ~new_n14638_;
  assign new_n14817_ = ~new_n1399_ | ~new_n1822_;
  assign new_n14818_ = ~new_n14609_ | ~new_n14816_;
  assign new_n14819_ = ~new_n14674_ | ~new_n14638_;
  assign new_n14820_ = ~new_n14671_ | ~new_n14532_;
  assign new_n14821_ = ~new_n14681_ | ~new_n14493_;
  assign new_n14822_ = ~new_n14695_ | ~new_n14505_;
  assign new_n14823_ = ~new_n14698_ | ~new_n14647_;
  assign new_n14824_ = ~new_n14781_ | ~new_n14640_;
  assign new_n14825_ = ~new_n14765_ | ~new_n14643_;
  assign new_n14826_ = ~new_n14796_ | ~new_n14551_;
  assign new_n14827_ = ~new_n14749_ | ~new_n14548_;
  assign new_n14828_ = ~new_n14803_ | ~new_n14530_;
  assign new_n14829_ = ~new_n14812_ | ~new_n14639_;
  assign new_n14830_ = ~new_n14717_ | ~new_n14539_;
  assign new_n14831_ = ~new_n2346_ | ~new_n1391_;
  assign new_n14832_ = ~new_n14763_ | ~new_n14635_;
  assign new_n14833_ = ~new_n1394_ | ~new_n14762_;
  assign new_n14834_ = ~new_n2348_ | ~new_n14762_;
  assign new_n14835_ = ~new_n14768_ | ~new_n14763_ | ~new_n14635_;
  assign new_n14836_ = ~new_n14602_ | ~new_n14621_ | ~new_n14635_;
  assign new_n14837_ = ~new_n14764_ | ~new_n14768_;
  assign new_n14838_ = ~new_n1420_ | ~new_n14510_;
  assign new_n14839_ = ~new_n1819_ | ~new_n14509_;
  assign new_n14840_ = ~new_n14839_ | ~new_n14838_;
  assign new_n14841_ = ~new_n14819_ | ~new_n14511_;
  assign new_n14842_ = ~new_n14840_ | ~new_n14673_;
  assign new_n14843_ = ~new_n1421_ | ~new_n14507_;
  assign new_n14844_ = ~new_n1816_ | ~new_n14508_;
  assign new_n14845_ = ~new_n14844_ | ~new_n14843_;
  assign new_n14846_ = ~new_n14820_ | ~new_n14610_;
  assign new_n14847_ = ~new_n14670_ | ~new_n14845_;
  assign new_n14848_ = ~new_n1407_ | ~new_n14494_;
  assign new_n14849_ = ~new_n1813_ | ~new_n14492_;
  assign new_n14850_ = ~new_n1408_ | ~new_n14490_;
  assign new_n14851_ = ~new_n1810_ | ~new_n14491_;
  assign new_n14852_ = ~new_n14851_ | ~new_n14850_;
  assign new_n14853_ = ~new_n14821_ | ~new_n14512_;
  assign new_n14854_ = ~new_n14852_ | ~new_n14662_;
  assign new_n14855_ = ~new_n1404_ | ~new_n14506_;
  assign new_n14856_ = ~new_n1807_ | ~new_n14497_;
  assign new_n14857_ = ~new_n1397_ | ~new_n14495_;
  assign new_n14858_ = ~new_n1804_ | ~new_n14496_;
  assign new_n14859_ = ~new_n14858_ | ~new_n14857_;
  assign new_n14860_ = ~new_n14822_ | ~new_n14515_;
  assign new_n14861_ = ~new_n14859_ | ~new_n14688_;
  assign new_n14862_ = ~new_n1401_ | ~new_n14503_;
  assign new_n14863_ = ~new_n1801_ | ~new_n14504_;
  assign new_n14864_ = ~new_n14863_ | ~new_n14862_;
  assign new_n14865_ = ~new_n14823_ | ~new_n14611_;
  assign new_n14866_ = ~new_n14697_ | ~new_n14864_;
  assign new_n14867_ = ~new_n1405_ | ~new_n14498_;
  assign new_n14868_ = ~new_n1798_ | ~new_n14499_;
  assign new_n14869_ = ~new_n1392_ | ~new_n14613_;
  assign new_n14870_ = ~new_n2357_ | ~new_n14612_;
  assign new_n14871_ = ~new_n1392_ | ~new_n14613_;
  assign new_n14872_ = ~new_n2357_ | ~new_n14612_;
  assign new_n14873_ = ~new_n14872_ | ~new_n14871_;
  assign new_n14874_ = ~new_n14614_ | ~new_n14615_;
  assign new_n14875_ = ~new_n14772_ | ~new_n14873_;
  assign new_n14876_ = ~new_n1391_ | ~new_n14559_;
  assign new_n14877_ = ~new_n2346_ | ~new_n14558_;
  assign new_n14878_ = ~new_n1391_ | ~new_n14559_;
  assign new_n14879_ = ~new_n2346_ | ~new_n14558_;
  assign new_n14880_ = ~new_n14879_ | ~new_n14878_;
  assign new_n14881_ = ~new_n14616_ | ~new_n14617_;
  assign new_n14882_ = ~new_n14770_ | ~new_n14880_;
  assign new_n14883_ = ~new_n1390_ | ~new_n14517_;
  assign new_n14884_ = ~new_n2347_ | ~new_n14518_;
  assign new_n14885_ = ~new_n1390_ | ~new_n14517_;
  assign new_n14886_ = ~new_n2347_ | ~new_n14518_;
  assign new_n14887_ = ~new_n14886_ | ~new_n14885_;
  assign new_n14888_ = ~new_n14618_ | ~new_n14619_;
  assign new_n14889_ = ~new_n14767_ | ~new_n14887_;
  assign new_n14890_ = ~new_n1394_ | ~new_n14520_;
  assign new_n14891_ = ~new_n2348_ | ~new_n14519_;
  assign new_n14892_ = ~new_n1395_ | ~new_n14521_;
  assign new_n14893_ = ~new_n2349_ | ~new_n14522_;
  assign new_n14894_ = ~new_n14893_ | ~new_n14892_;
  assign new_n14895_ = ~new_n14824_ | ~new_n14560_;
  assign new_n14896_ = ~new_n14894_ | ~new_n14774_;
  assign new_n14897_ = ~new_n1402_ | ~new_n14523_;
  assign new_n14898_ = ~new_n2350_ | ~new_n14524_;
  assign new_n14899_ = ~new_n14898_ | ~new_n14897_;
  assign new_n14900_ = ~new_n14825_ | ~new_n14621_;
  assign new_n14901_ = ~new_n14761_ | ~new_n14899_;
  assign new_n14902_ = ~new_n1403_ | ~new_n14555_;
  assign new_n14903_ = ~new_n2351_ | ~new_n14556_;
  assign new_n14904_ = ~new_n1403_ | ~new_n14555_;
  assign new_n14905_ = ~new_n2351_ | ~new_n14556_;
  assign new_n14906_ = ~new_n14905_ | ~new_n14904_;
  assign new_n14907_ = ~new_n14622_ | ~new_n14623_;
  assign new_n14908_ = ~new_n14757_ | ~new_n14906_;
  assign new_n14909_ = ~new_n1398_ | ~new_n14553_;
  assign new_n14910_ = ~new_n2352_ | ~new_n14554_;
  assign new_n14911_ = ~new_n1398_ | ~new_n14553_;
  assign new_n14912_ = ~new_n2352_ | ~new_n14554_;
  assign new_n14913_ = ~new_n14912_ | ~new_n14911_;
  assign new_n14914_ = ~new_n14624_ | ~new_n14625_;
  assign new_n14915_ = ~new_n14753_ | ~new_n14913_;
  assign new_n14916_ = ~new_n1412_ | ~new_n14525_;
  assign new_n14917_ = ~new_n2353_ | ~new_n14526_;
  assign new_n14918_ = ~new_n1412_ | ~new_n14525_;
  assign new_n14919_ = ~new_n2353_ | ~new_n14526_;
  assign new_n14920_ = ~new_n14919_ | ~new_n14918_;
  assign new_n14921_ = ~new_n1413_ | ~new_n14552_;
  assign new_n14922_ = ~new_n2354_ | ~new_n14561_;
  assign new_n14923_ = ~new_n14649_ | ~new_n14628_;
  assign new_n14924_ = ~new_n14795_ | ~new_n14502_;
  assign new_n14925_ = ~new_n1418_ | ~new_n14549_;
  assign new_n14926_ = ~new_n1848_ | ~new_n14550_;
  assign new_n14927_ = ~new_n14926_ | ~new_n14925_;
  assign new_n14928_ = ~new_n14826_ | ~new_n14562_;
  assign new_n14929_ = ~new_n14927_ | ~new_n14783_;
  assign new_n14930_ = ~new_n1419_ | ~new_n14546_;
  assign new_n14931_ = ~new_n1846_ | ~new_n14547_;
  assign new_n14932_ = ~new_n14931_ | ~new_n14930_;
  assign new_n14933_ = ~new_n14827_ | ~new_n14629_;
  assign new_n14934_ = ~new_n14737_ | ~new_n14932_;
  assign new_n14935_ = ~new_n1406_ | ~new_n14531_;
  assign new_n14936_ = ~new_n1843_ | ~new_n14529_;
  assign new_n14937_ = ~new_n1410_ | ~new_n14527_;
  assign new_n14938_ = ~new_n1840_ | ~new_n14528_;
  assign new_n14939_ = ~new_n14938_ | ~new_n14937_;
  assign new_n14940_ = ~new_n14828_ | ~new_n14563_;
  assign new_n14941_ = ~new_n14939_ | ~new_n14729_;
  assign new_n14942_ = ~new_n1411_ | ~new_n14544_;
  assign new_n14943_ = ~new_n1837_ | ~new_n14545_;
  assign new_n14944_ = ~new_n1411_ | ~new_n14544_;
  assign new_n14945_ = ~new_n1837_ | ~new_n14545_;
  assign new_n14946_ = ~new_n14945_ | ~new_n14944_;
  assign new_n14947_ = ~new_n14630_ | ~new_n14631_;
  assign new_n14948_ = ~new_n14725_ | ~new_n14946_;
  assign new_n14949_ = ~new_n1416_ | ~new_n14542_;
  assign new_n14950_ = ~new_n1834_ | ~new_n14543_;
  assign new_n14951_ = ~new_n1416_ | ~new_n14542_;
  assign new_n14952_ = ~new_n1834_ | ~new_n14543_;
  assign new_n14953_ = ~new_n14952_ | ~new_n14951_;
  assign new_n14954_ = ~new_n14632_ | ~new_n14633_;
  assign new_n14955_ = ~new_n14721_ | ~new_n14953_;
  assign new_n14956_ = ~new_n1417_ | ~new_n14540_;
  assign new_n14957_ = ~new_n1831_ | ~new_n14541_;
  assign new_n14958_ = ~new_n1409_ | ~new_n14535_;
  assign new_n14959_ = ~new_n1828_ | ~new_n14536_;
  assign new_n14960_ = ~new_n14959_ | ~new_n14958_;
  assign new_n14961_ = ~new_n14829_ | ~new_n14564_;
  assign new_n14962_ = ~new_n14960_ | ~new_n14805_;
  assign new_n14963_ = ~new_n1400_ | ~new_n14537_;
  assign new_n14964_ = ~new_n1825_ | ~new_n14538_;
  assign new_n14965_ = ~new_n14964_ | ~new_n14963_;
  assign new_n14966_ = ~new_n14830_ | ~new_n14634_;
  assign new_n14967_ = ~new_n14711_ | ~new_n14965_;
  assign new_n14968_ = ~new_n1399_ | ~new_n14533_;
  assign new_n14969_ = ~new_n1822_ | ~new_n14534_;
  assign new_n14970_ = ~new_n1414_ | ~new_n14500_;
  assign new_n14971_ = ~new_n1790_ | ~new_n14501_;
  assign new_n14972_ = ~pi514;
  assign new_n14973_ = new_n15044_ & new_n15072_;
  assign new_n14974_ = ~pi519;
  assign new_n14975_ = ~pi493;
  assign new_n14976_ = ~pi505;
  assign new_n14977_ = ~pi502;
  assign new_n14978_ = ~pi505 | ~pi502 | ~pi493 | ~pi519 | ~pi514;
  assign new_n14979_ = ~pi511;
  assign new_n14980_ = ~pi501;
  assign new_n14981_ = ~new_n15042_ | ~new_n15053_;
  assign new_n14982_ = ~pi496;
  assign new_n14983_ = ~pi515;
  assign new_n14984_ = ~new_n15043_ | ~new_n15055_;
  assign new_n14985_ = ~pi508;
  assign new_n14986_ = ~pi508 | ~new_n15057_;
  assign new_n14987_ = ~pi498;
  assign new_n14988_ = ~pi498 | ~new_n15058_;
  assign new_n14989_ = ~pi517;
  assign new_n14990_ = ~pi517 | ~new_n15059_;
  assign new_n14991_ = ~pi491;
  assign new_n14992_ = ~pi491 | ~new_n15060_;
  assign new_n14993_ = ~pi506;
  assign new_n14994_ = ~pi506 | ~new_n15061_;
  assign new_n14995_ = ~pi504;
  assign new_n14996_ = ~pi504 | ~new_n15062_;
  assign new_n14997_ = ~pi494;
  assign new_n14998_ = ~pi494 | ~new_n15063_;
  assign new_n14999_ = ~pi513;
  assign new_n15000_ = ~pi513 | ~new_n15064_;
  assign new_n15001_ = ~pi499;
  assign new_n15002_ = ~pi499 | ~new_n15065_;
  assign new_n15003_ = ~pi509;
  assign new_n15004_ = ~pi509 | ~new_n15066_;
  assign new_n15005_ = ~pi497;
  assign new_n15006_ = ~pi497 | ~new_n15067_;
  assign new_n15007_ = ~pi516;
  assign new_n15008_ = ~pi516 | ~new_n15068_;
  assign new_n15009_ = ~pi503;
  assign new_n15010_ = ~pi503 | ~new_n15069_;
  assign new_n15011_ = ~pi507;
  assign new_n15012_ = ~pi507 | ~new_n15070_;
  assign new_n15013_ = ~pi492;
  assign new_n15014_ = ~pi492 | ~new_n15071_;
  assign new_n15015_ = ~pi512;
  assign new_n15016_ = ~pi518;
  assign new_n15017_ = ~new_n15076_ | ~new_n15075_;
  assign new_n15018_ = ~new_n15078_ | ~new_n15077_;
  assign new_n15019_ = ~new_n15080_ | ~new_n15079_;
  assign new_n15020_ = ~new_n15082_ | ~new_n15081_;
  assign new_n15021_ = ~new_n15084_ | ~new_n15083_;
  assign new_n15022_ = ~new_n15086_ | ~new_n15085_;
  assign new_n15023_ = ~new_n15088_ | ~new_n15087_;
  assign new_n15024_ = ~new_n15090_ | ~new_n15089_;
  assign new_n15025_ = ~new_n15092_ | ~new_n15091_;
  assign new_n15026_ = ~new_n15094_ | ~new_n15093_;
  assign new_n15027_ = ~new_n15096_ | ~new_n15095_;
  assign new_n15028_ = ~new_n15098_ | ~new_n15097_;
  assign new_n15029_ = ~new_n15100_ | ~new_n15099_;
  assign new_n15030_ = ~new_n15102_ | ~new_n15101_;
  assign new_n15031_ = ~new_n15104_ | ~new_n15103_;
  assign new_n15032_ = ~new_n15106_ | ~new_n15105_;
  assign new_n15033_ = ~new_n15108_ | ~new_n15107_;
  assign new_n15034_ = ~new_n15110_ | ~new_n15109_;
  assign new_n15035_ = ~new_n15112_ | ~new_n15111_;
  assign new_n15036_ = ~new_n15114_ | ~new_n15113_;
  assign new_n15037_ = ~new_n15116_ | ~new_n15115_;
  assign new_n15038_ = ~new_n15118_ | ~new_n15117_;
  assign new_n15039_ = ~new_n15120_ | ~new_n15119_;
  assign new_n15040_ = ~new_n15122_ | ~new_n15121_;
  assign new_n15041_ = ~new_n15124_ | ~new_n15123_;
  assign new_n15042_ = pi511 & pi501;
  assign new_n15043_ = pi496 & pi515;
  assign new_n15044_ = pi512 & pi518;
  assign new_n15045_ = ~pi511 | ~new_n15053_;
  assign new_n15046_ = ~pi514 | ~pi493 | ~pi502 | ~pi505;
  assign new_n15047_ = ~pi502 | ~pi505 | ~pi514;
  assign new_n15048_ = ~pi502 | ~pi514;
  assign new_n15049_ = ~pi518 | ~new_n15072_;
  assign new_n15050_ = ~pi515 | ~new_n15055_;
  assign new_n15051_ = ~new_n15048_;
  assign new_n15052_ = ~new_n15046_;
  assign new_n15053_ = ~new_n14978_;
  assign new_n15054_ = ~new_n15045_;
  assign new_n15055_ = ~new_n14981_;
  assign new_n15056_ = ~new_n15050_;
  assign new_n15057_ = ~new_n14984_;
  assign new_n15058_ = ~new_n14986_;
  assign new_n15059_ = ~new_n14988_;
  assign new_n15060_ = ~new_n14990_;
  assign new_n15061_ = ~new_n14992_;
  assign new_n15062_ = ~new_n14994_;
  assign new_n15063_ = ~new_n14996_;
  assign new_n15064_ = ~new_n14998_;
  assign new_n15065_ = ~new_n15000_;
  assign new_n15066_ = ~new_n15002_;
  assign new_n15067_ = ~new_n15004_;
  assign new_n15068_ = ~new_n15006_;
  assign new_n15069_ = ~new_n15008_;
  assign new_n15070_ = ~new_n15010_;
  assign new_n15071_ = ~new_n15012_;
  assign new_n15072_ = ~new_n15014_;
  assign new_n15073_ = ~new_n15049_;
  assign new_n15074_ = ~new_n15047_;
  assign new_n15075_ = ~pi501 | ~new_n15045_;
  assign new_n15076_ = ~new_n15054_ | ~new_n14980_;
  assign new_n15077_ = ~pi511 | ~new_n14978_;
  assign new_n15078_ = ~new_n15053_ | ~new_n14979_;
  assign new_n15079_ = ~pi519 | ~new_n15046_;
  assign new_n15080_ = ~new_n15052_ | ~new_n14974_;
  assign new_n15081_ = ~pi493 | ~new_n15047_;
  assign new_n15082_ = ~new_n15074_ | ~new_n14975_;
  assign new_n15083_ = ~pi505 | ~new_n15048_;
  assign new_n15084_ = ~new_n15051_ | ~new_n14976_;
  assign new_n15085_ = ~pi502 | ~new_n14972_;
  assign new_n15086_ = ~pi514 | ~new_n14977_;
  assign new_n15087_ = ~pi512 | ~new_n15049_;
  assign new_n15088_ = ~new_n15073_ | ~new_n15015_;
  assign new_n15089_ = ~pi518 | ~new_n15014_;
  assign new_n15090_ = ~new_n15072_ | ~new_n15016_;
  assign new_n15091_ = ~pi492 | ~new_n15012_;
  assign new_n15092_ = ~new_n15071_ | ~new_n15013_;
  assign new_n15093_ = ~pi507 | ~new_n15010_;
  assign new_n15094_ = ~new_n15070_ | ~new_n15011_;
  assign new_n15095_ = ~pi503 | ~new_n15008_;
  assign new_n15096_ = ~new_n15069_ | ~new_n15009_;
  assign new_n15097_ = ~pi516 | ~new_n15006_;
  assign new_n15098_ = ~new_n15068_ | ~new_n15007_;
  assign new_n15099_ = ~pi497 | ~new_n15004_;
  assign new_n15100_ = ~new_n15067_ | ~new_n15005_;
  assign new_n15101_ = ~pi509 | ~new_n15002_;
  assign new_n15102_ = ~new_n15066_ | ~new_n15003_;
  assign new_n15103_ = ~pi499 | ~new_n15000_;
  assign new_n15104_ = ~new_n15065_ | ~new_n15001_;
  assign new_n15105_ = ~pi513 | ~new_n14998_;
  assign new_n15106_ = ~new_n15064_ | ~new_n14999_;
  assign new_n15107_ = ~pi494 | ~new_n14996_;
  assign new_n15108_ = ~new_n15063_ | ~new_n14997_;
  assign new_n15109_ = ~pi504 | ~new_n14994_;
  assign new_n15110_ = ~new_n15062_ | ~new_n14995_;
  assign new_n15111_ = ~pi506 | ~new_n14992_;
  assign new_n15112_ = ~new_n15061_ | ~new_n14993_;
  assign new_n15113_ = ~pi491 | ~new_n14990_;
  assign new_n15114_ = ~new_n15060_ | ~new_n14991_;
  assign new_n15115_ = ~pi517 | ~new_n14988_;
  assign new_n15116_ = ~new_n15059_ | ~new_n14989_;
  assign new_n15117_ = ~pi498 | ~new_n14986_;
  assign new_n15118_ = ~new_n15058_ | ~new_n14987_;
  assign new_n15119_ = ~pi508 | ~new_n14984_;
  assign new_n15120_ = ~new_n15057_ | ~new_n14985_;
  assign new_n15121_ = ~pi496 | ~new_n15050_;
  assign new_n15122_ = ~new_n15056_ | ~new_n14982_;
  assign new_n15123_ = ~pi515 | ~new_n14981_;
  assign new_n15124_ = ~new_n15055_ | ~new_n14983_;
  assign new_n15125_ = new_n15292_ & new_n15294_ & new_n15298_ & new_n15295_;
  assign new_n15126_ = ~new_n5072_;
  assign new_n15127_ = ~new_n5075_;
  assign new_n15128_ = ~new_n5078_;
  assign new_n15129_ = ~new_n4798_;
  assign new_n15130_ = ~new_n4797_;
  assign new_n15131_ = ~new_n4796_;
  assign new_n15132_ = ~new_n4795_;
  assign new_n15133_ = ~new_n4794_;
  assign new_n15134_ = ~new_n4793_;
  assign new_n15135_ = ~new_n5081_;
  assign new_n15136_ = ~new_n5084_;
  assign new_n15137_ = ~new_n5087_;
  assign new_n15138_ = ~new_n5090_;
  assign new_n15139_ = ~new_n5093_;
  assign new_n15140_ = ~new_n5096_;
  assign new_n15141_ = ~new_n4792_;
  assign new_n15142_ = ~new_n4791_;
  assign new_n15143_ = ~new_n4790_;
  assign new_n15144_ = ~new_n4789_;
  assign new_n15145_ = ~new_n4788_;
  assign new_n15146_ = ~new_n4787_;
  assign new_n15147_ = ~new_n5099_;
  assign new_n15148_ = ~new_n5102_;
  assign new_n15149_ = ~new_n5105_;
  assign new_n15150_ = ~new_n5108_;
  assign new_n15151_ = ~new_n5111_;
  assign new_n15152_ = ~new_n5114_;
  assign new_n15153_ = ~new_n4786_;
  assign new_n15154_ = ~new_n4785_;
  assign new_n15155_ = ~new_n4784_;
  assign new_n15156_ = ~new_n4783_;
  assign new_n15157_ = ~new_n5117_;
  assign new_n15158_ = ~new_n5120_;
  assign new_n15159_ = ~new_n4782_;
  assign new_n15160_ = ~new_n4781_;
  assign new_n15161_ = ~new_n5122_;
  assign new_n15162_ = ~new_n5592_;
  assign new_n15163_ = ~new_n4780_;
  assign new_n15164_ = ~new_n4779_;
  assign new_n15165_ = ~new_n5591_;
  assign new_n15166_ = ~new_n5590_;
  assign new_n15167_ = ~new_n4778_;
  assign new_n15168_ = ~new_n4777_;
  assign new_n15169_ = ~new_n5589_;
  assign new_n15170_ = ~new_n5588_;
  assign new_n15171_ = ~new_n4776_;
  assign new_n15172_ = ~new_n4775_;
  assign new_n15173_ = ~new_n5587_;
  assign new_n15174_ = ~new_n5586_;
  assign new_n15175_ = ~new_n4774_;
  assign new_n15176_ = ~new_n4773_;
  assign new_n15177_ = ~new_n5585_;
  assign new_n15178_ = ~new_n5584_;
  assign new_n15179_ = ~new_n4772_;
  assign new_n15180_ = ~new_n4771_;
  assign new_n15181_ = ~new_n5595_;
  assign new_n15182_ = ~new_n4769_;
  assign new_n15183_ = ~new_n5593_;
  assign new_n15184_ = new_n15217_ & new_n15218_ & new_n15219_;
  assign new_n15185_ = new_n15297_ & new_n15224_ & new_n15223_;
  assign new_n15186_ = new_n4797_ & new_n15127_;
  assign new_n15187_ = new_n15188_ & new_n15221_ & new_n15225_ & new_n15222_;
  assign new_n15188_ = new_n15231_ & new_n15230_ & new_n15226_;
  assign new_n15189_ = new_n5084_ & new_n15133_;
  assign new_n15190_ = new_n15191_ & new_n15228_ & new_n15232_ & new_n15229_;
  assign new_n15191_ = new_n15238_ & new_n15237_ & new_n15233_;
  assign new_n15192_ = new_n4791_ & new_n15139_;
  assign new_n15193_ = new_n15194_ & new_n15235_ & new_n15239_ & new_n15236_;
  assign new_n15194_ = new_n15245_ & new_n15244_ & new_n15240_;
  assign new_n15195_ = new_n5102_ & new_n15145_;
  assign new_n15196_ = new_n15197_ & new_n15242_ & new_n15246_ & new_n15243_;
  assign new_n15197_ = new_n15252_ & new_n15251_ & new_n15247_;
  assign new_n15198_ = new_n4785_ & new_n15151_;
  assign new_n15199_ = new_n15249_ & new_n15200_ & new_n15250_;
  assign new_n15200_ = new_n15254_ & new_n15253_;
  assign new_n15201_ = new_n15256_ & new_n15257_;
  assign new_n15202_ = new_n15259_ & new_n15260_;
  assign new_n15203_ = new_n15262_ & new_n15263_;
  assign new_n15204_ = new_n15265_ & new_n15266_;
  assign new_n15205_ = new_n15268_ & new_n15269_;
  assign new_n15206_ = new_n15271_ & new_n15272_;
  assign new_n15207_ = new_n15274_ & new_n15275_;
  assign new_n15208_ = new_n15277_ & new_n15278_;
  assign new_n15209_ = new_n15280_ & new_n15281_;
  assign new_n15210_ = new_n15283_ & new_n15284_;
  assign new_n15211_ = new_n15289_ & new_n15290_;
  assign new_n15212_ = new_n15296_ & new_n15293_;
  assign new_n15213_ = new_n4770_ & new_n15296_;
  assign new_n15214_ = ~new_n5594_;
  assign new_n15215_ = ~new_n4799_;
  assign new_n15216_ = ~new_n4800_;
  assign new_n15217_ = ~new_n5064_ | ~new_n15216_ | ~new_n15215_;
  assign new_n15218_ = ~new_n5069_ | ~new_n15215_;
  assign new_n15219_ = ~new_n5072_ | ~new_n15129_;
  assign new_n15220_ = ~new_n15185_ | ~new_n15184_;
  assign new_n15221_ = ~new_n15126_ | ~new_n15223_ | ~new_n4798_ | ~new_n15224_;
  assign new_n15222_ = ~new_n15186_ | ~new_n15224_;
  assign new_n15223_ = ~new_n5075_ | ~new_n15130_;
  assign new_n15224_ = ~new_n5078_ | ~new_n15131_;
  assign new_n15225_ = ~new_n4796_ | ~new_n15128_;
  assign new_n15226_ = ~new_n4795_ | ~new_n15135_;
  assign new_n15227_ = ~new_n15220_ | ~new_n15187_;
  assign new_n15228_ = ~new_n15132_ | ~new_n15230_ | ~new_n5081_ | ~new_n15231_;
  assign new_n15229_ = ~new_n15189_ | ~new_n15231_;
  assign new_n15230_ = ~new_n4794_ | ~new_n15136_;
  assign new_n15231_ = ~new_n4793_ | ~new_n15137_;
  assign new_n15232_ = ~new_n5087_ | ~new_n15134_;
  assign new_n15233_ = ~new_n5090_ | ~new_n15141_;
  assign new_n15234_ = ~new_n15227_ | ~new_n15190_;
  assign new_n15235_ = ~new_n15138_ | ~new_n15237_ | ~new_n4792_ | ~new_n15238_;
  assign new_n15236_ = ~new_n15192_ | ~new_n15238_;
  assign new_n15237_ = ~new_n5093_ | ~new_n15142_;
  assign new_n15238_ = ~new_n5096_ | ~new_n15143_;
  assign new_n15239_ = ~new_n4790_ | ~new_n15140_;
  assign new_n15240_ = ~new_n4789_ | ~new_n15147_;
  assign new_n15241_ = ~new_n15234_ | ~new_n15193_;
  assign new_n15242_ = ~new_n15144_ | ~new_n15244_ | ~new_n5099_ | ~new_n15245_;
  assign new_n15243_ = ~new_n15195_ | ~new_n15245_;
  assign new_n15244_ = ~new_n4788_ | ~new_n15148_;
  assign new_n15245_ = ~new_n4787_ | ~new_n15149_;
  assign new_n15246_ = ~new_n5105_ | ~new_n15146_;
  assign new_n15247_ = ~new_n5108_ | ~new_n15153_;
  assign new_n15248_ = ~new_n15241_ | ~new_n15196_;
  assign new_n15249_ = ~new_n15150_ | ~new_n15251_ | ~new_n4786_ | ~new_n15252_;
  assign new_n15250_ = ~new_n15198_ | ~new_n15252_;
  assign new_n15251_ = ~new_n5111_ | ~new_n15154_;
  assign new_n15252_ = ~new_n5114_ | ~new_n15155_;
  assign new_n15253_ = ~new_n4784_ | ~new_n15152_;
  assign new_n15254_ = ~new_n4783_ | ~new_n15157_;
  assign new_n15255_ = ~new_n15248_ | ~new_n15199_;
  assign new_n15256_ = ~new_n5117_ | ~new_n15156_;
  assign new_n15257_ = ~new_n5120_ | ~new_n15159_;
  assign new_n15258_ = ~new_n15201_ | ~new_n15255_;
  assign new_n15259_ = ~new_n4782_ | ~new_n15158_;
  assign new_n15260_ = ~new_n4781_ | ~new_n15161_;
  assign new_n15261_ = ~new_n15202_ | ~new_n15258_;
  assign new_n15262_ = ~new_n5122_ | ~new_n15160_;
  assign new_n15263_ = ~new_n5592_ | ~new_n15163_;
  assign new_n15264_ = ~new_n15203_ | ~new_n15261_;
  assign new_n15265_ = ~new_n4780_ | ~new_n15162_;
  assign new_n15266_ = ~new_n4779_ | ~new_n15165_;
  assign new_n15267_ = ~new_n15204_ | ~new_n15264_;
  assign new_n15268_ = ~new_n5591_ | ~new_n15164_;
  assign new_n15269_ = ~new_n5590_ | ~new_n15167_;
  assign new_n15270_ = ~new_n15205_ | ~new_n15267_;
  assign new_n15271_ = ~new_n4778_ | ~new_n15166_;
  assign new_n15272_ = ~new_n4777_ | ~new_n15169_;
  assign new_n15273_ = ~new_n15206_ | ~new_n15270_;
  assign new_n15274_ = ~new_n5589_ | ~new_n15168_;
  assign new_n15275_ = ~new_n5588_ | ~new_n15171_;
  assign new_n15276_ = ~new_n15207_ | ~new_n15273_;
  assign new_n15277_ = ~new_n4776_ | ~new_n15170_;
  assign new_n15278_ = ~new_n4775_ | ~new_n15173_;
  assign new_n15279_ = ~new_n15208_ | ~new_n15276_;
  assign new_n15280_ = ~new_n5587_ | ~new_n15172_;
  assign new_n15281_ = ~new_n5586_ | ~new_n15175_;
  assign new_n15282_ = ~new_n15209_ | ~new_n15279_;
  assign new_n15283_ = ~new_n4774_ | ~new_n15174_;
  assign new_n15284_ = ~new_n4773_ | ~new_n15177_;
  assign new_n15285_ = ~new_n15210_ | ~new_n15282_;
  assign new_n15286_ = ~new_n5585_ | ~new_n15176_;
  assign new_n15287_ = ~new_n5584_ | ~new_n15179_;
  assign new_n15288_ = ~new_n15287_ | ~new_n15286_ | ~new_n15285_;
  assign new_n15289_ = ~new_n4772_ | ~new_n15178_;
  assign new_n15290_ = ~new_n4771_ | ~new_n15181_;
  assign new_n15291_ = ~new_n15211_ | ~new_n15288_;
  assign new_n15292_ = ~new_n15212_ | ~new_n15291_ | ~new_n15214_;
  assign new_n15293_ = ~new_n5595_ | ~new_n15180_;
  assign new_n15294_ = ~new_n5593_ | ~new_n15182_;
  assign new_n15295_ = ~new_n15214_ | ~new_n15296_ | ~new_n4770_;
  assign new_n15296_ = ~new_n4769_ | ~new_n15183_;
  assign new_n15297_ = ~new_n15216_ | ~new_n5064_ | ~new_n5069_;
  assign new_n15298_ = ~new_n15213_ | ~new_n15293_ | ~new_n15291_;
  assign new_n15299_ = new_n15350_ & new_n15349_;
  assign new_n15300_ = ~pi304 & ~pi305 & ~pi303;
  assign new_n15301_ = ~pi303 & ~pi304;
  assign new_n15302_ = new_n15345_ & new_n15346_ & new_n15348_ & new_n15347_;
  assign new_n15303_ = ~pi287 & ~pi290 & ~pi289 & ~pi288;
  assign new_n15304_ = new_n15435_ & new_n15340_;
  assign new_n15305_ = new_n15433_ & new_n15404_;
  assign new_n15306_ = new_n15432_ & new_n15336_;
  assign new_n15307_ = new_n15431_ & new_n15337_;
  assign new_n15308_ = new_n15429_ & new_n15407_;
  assign new_n15309_ = new_n15428_ & new_n15389_;
  assign new_n15310_ = new_n15427_ & new_n15418_;
  assign new_n15311_ = new_n15425_ & new_n15419_;
  assign new_n15312_ = new_n15424_ & new_n15384_;
  assign new_n15313_ = new_n15357_ & new_n15437_;
  assign new_n15314_ = new_n15423_ & new_n15382_;
  assign new_n15315_ = new_n15417_ & new_n15409_;
  assign new_n15316_ = new_n15416_ & new_n15410_;
  assign new_n15317_ = new_n15415_ & new_n15327_;
  assign new_n15318_ = new_n15402_ & new_n15394_;
  assign new_n15319_ = new_n15401_ & new_n15323_;
  assign new_n15320_ = new_n15400_ & new_n15325_;
  assign new_n15321_ = new_n15398_ & new_n15396_;
  assign new_n15322_ = new_n15397_ & new_n15324_;
  assign new_n15323_ = pi278 | pi279 | pi280 | pi282 | pi281;
  assign new_n15324_ = ~new_n15343_ | ~new_n15441_;
  assign new_n15325_ = ~new_n15344_ | ~new_n15441_;
  assign new_n15326_ = ~pi285;
  assign new_n15327_ = pi278 | pi280 | pi279;
  assign new_n15328_ = ~pi281;
  assign new_n15329_ = ~new_n15299_ | ~new_n15302_;
  assign new_n15330_ = ~new_n15351_ | ~new_n15440_;
  assign new_n15331_ = ~new_n15411_ | ~new_n15373_;
  assign new_n15332_ = ~pi303;
  assign new_n15333_ = ~new_n15355_ | ~new_n15302_;
  assign new_n15334_ = ~pi301;
  assign new_n15335_ = ~pi299;
  assign new_n15336_ = ~new_n15303_ | ~new_n15442_;
  assign new_n15337_ = ~new_n15362_ | ~new_n15405_;
  assign new_n15338_ = ~pi294;
  assign new_n15339_ = ~pi293;
  assign new_n15340_ = ~new_n15363_ | ~new_n15442_;
  assign new_n15341_ = ~pi289;
  assign new_n15342_ = ~new_n15462_ | ~new_n15461_;
  assign new_n15343_ = ~pi284 & ~pi283 & ~pi286 & ~pi285;
  assign new_n15344_ = ~pi283 & ~pi284;
  assign new_n15345_ = ~pi292 & ~pi291 & ~pi290 & ~pi289 & ~pi288;
  assign new_n15346_ = ~pi294 & ~pi293 & ~pi278 & ~pi279;
  assign new_n15347_ = ~pi281 & ~pi280 & ~pi283 & ~pi282;
  assign new_n15348_ = ~pi285 & ~pi284 & ~pi287 & ~pi286;
  assign new_n15349_ = ~pi296 & ~pi295 & ~pi298 & ~pi297;
  assign new_n15350_ = ~pi300 & ~pi299 & ~pi302 & ~pi301;
  assign new_n15351_ = new_n15300_ & new_n15375_;
  assign new_n15352_ = ~pi295 & ~pi296;
  assign new_n15353_ = ~pi297 & ~pi298;
  assign new_n15354_ = ~pi299 & ~pi300;
  assign new_n15355_ = new_n15354_ & new_n15353_ & new_n15352_;
  assign new_n15356_ = ~pi296 & ~pi295 & ~pi298 & ~pi297;
  assign new_n15357_ = new_n15436_ & new_n15333_;
  assign new_n15358_ = ~pi295 & ~pi296 & ~pi297;
  assign new_n15359_ = ~pi295 & ~pi296;
  assign new_n15360_ = ~pi291 & ~pi292 & ~pi293;
  assign new_n15361_ = new_n15360_ & new_n15303_ & new_n15338_;
  assign new_n15362_ = ~pi291 & ~pi292;
  assign new_n15363_ = ~pi288 & ~pi287;
  assign new_n15364_ = ~pi287;
  assign new_n15365_ = new_n15444_ & new_n15443_;
  assign new_n15366_ = ~pi283;
  assign new_n15367_ = new_n15446_ & new_n15445_;
  assign new_n15368_ = ~pi309;
  assign new_n15369_ = ~new_n15412_ | ~new_n15371_;
  assign new_n15370_ = new_n15448_ & new_n15447_;
  assign new_n15371_ = ~pi308;
  assign new_n15372_ = new_n15450_ & new_n15449_;
  assign new_n15373_ = ~pi307;
  assign new_n15374_ = new_n15452_ & new_n15451_;
  assign new_n15375_ = ~pi306;
  assign new_n15376_ = ~new_n15302_ | ~new_n15299_ | ~new_n15300_;
  assign new_n15377_ = new_n15454_ & new_n15453_;
  assign new_n15378_ = ~pi305;
  assign new_n15379_ = ~new_n15302_ | ~new_n15299_ | ~new_n15301_;
  assign new_n15380_ = new_n15456_ & new_n15455_;
  assign new_n15381_ = ~pi302;
  assign new_n15382_ = ~new_n15421_ | ~new_n15334_;
  assign new_n15383_ = new_n15458_ & new_n15457_;
  assign new_n15384_ = ~new_n15356_ | ~new_n15302_;
  assign new_n15385_ = new_n15460_ & new_n15459_;
  assign new_n15386_ = ~pi279;
  assign new_n15387_ = ~pi278;
  assign new_n15388_ = ~pi295;
  assign new_n15389_ = ~new_n15361_ | ~new_n15442_;
  assign new_n15390_ = new_n15464_ & new_n15463_;
  assign new_n15391_ = ~pi291;
  assign new_n15392_ = new_n15466_ & new_n15465_;
  assign new_n15393_ = ~new_n15327_;
  assign new_n15394_ = ~new_n15393_ | ~new_n15328_;
  assign new_n15395_ = ~new_n15325_;
  assign new_n15396_ = ~new_n15395_ | ~new_n15326_;
  assign new_n15397_ = ~pi286 | ~new_n15396_;
  assign new_n15398_ = ~pi285 | ~new_n15325_;
  assign new_n15399_ = ~new_n15441_ | ~new_n15366_;
  assign new_n15400_ = ~pi284 | ~new_n15399_;
  assign new_n15401_ = ~pi282 | ~new_n15394_;
  assign new_n15402_ = ~pi281 | ~new_n15327_;
  assign new_n15403_ = ~new_n15340_;
  assign new_n15404_ = ~new_n15403_ | ~new_n15341_;
  assign new_n15405_ = ~new_n15336_;
  assign new_n15406_ = ~new_n15337_;
  assign new_n15407_ = ~new_n15406_ | ~new_n15339_;
  assign new_n15408_ = ~new_n15389_;
  assign new_n15409_ = ~new_n15440_ | ~new_n15332_;
  assign new_n15410_ = ~new_n15301_ | ~new_n15440_;
  assign new_n15411_ = ~new_n15330_;
  assign new_n15412_ = ~new_n15331_;
  assign new_n15413_ = ~new_n15369_;
  assign new_n15414_ = pi279 | pi278;
  assign new_n15415_ = ~pi280 | ~new_n15414_;
  assign new_n15416_ = ~pi304 | ~new_n15409_;
  assign new_n15417_ = ~pi303 | ~new_n15329_;
  assign new_n15418_ = ~new_n15359_ | ~new_n15302_;
  assign new_n15419_ = ~new_n15358_ | ~new_n15302_;
  assign new_n15420_ = ~new_n15384_;
  assign new_n15421_ = ~new_n15333_;
  assign new_n15422_ = ~new_n15382_;
  assign new_n15423_ = ~pi301 | ~new_n15333_;
  assign new_n15424_ = ~pi298 | ~new_n15419_;
  assign new_n15425_ = ~pi297 | ~new_n15418_;
  assign new_n15426_ = ~new_n15302_ | ~new_n15388_;
  assign new_n15427_ = ~pi296 | ~new_n15426_;
  assign new_n15428_ = ~pi294 | ~new_n15407_;
  assign new_n15429_ = ~pi293 | ~new_n15337_;
  assign new_n15430_ = ~new_n15405_ | ~new_n15391_;
  assign new_n15431_ = ~pi292 | ~new_n15430_;
  assign new_n15432_ = ~pi290 | ~new_n15404_;
  assign new_n15433_ = ~pi289 | ~new_n15340_;
  assign new_n15434_ = ~new_n15442_ | ~new_n15364_;
  assign new_n15435_ = ~pi288 | ~new_n15434_;
  assign new_n15436_ = ~pi299 | ~pi300;
  assign new_n15437_ = ~pi300 | ~new_n15384_;
  assign new_n15438_ = ~new_n15379_;
  assign new_n15439_ = ~new_n15376_;
  assign new_n15440_ = ~new_n15329_;
  assign new_n15441_ = ~new_n15323_;
  assign new_n15442_ = ~new_n15324_;
  assign new_n15443_ = ~pi287 | ~new_n15324_;
  assign new_n15444_ = ~new_n15442_ | ~new_n15364_;
  assign new_n15445_ = ~pi283 | ~new_n15323_;
  assign new_n15446_ = ~new_n15441_ | ~new_n15366_;
  assign new_n15447_ = ~pi309 | ~new_n15369_;
  assign new_n15448_ = ~new_n15413_ | ~new_n15368_;
  assign new_n15449_ = ~pi308 | ~new_n15331_;
  assign new_n15450_ = ~new_n15412_ | ~new_n15371_;
  assign new_n15451_ = ~pi307 | ~new_n15330_;
  assign new_n15452_ = ~new_n15411_ | ~new_n15373_;
  assign new_n15453_ = ~pi306 | ~new_n15376_;
  assign new_n15454_ = ~new_n15439_ | ~new_n15375_;
  assign new_n15455_ = ~pi305 | ~new_n15379_;
  assign new_n15456_ = ~new_n15438_ | ~new_n15378_;
  assign new_n15457_ = ~pi302 | ~new_n15382_;
  assign new_n15458_ = ~new_n15422_ | ~new_n15381_;
  assign new_n15459_ = ~pi299 | ~new_n15384_;
  assign new_n15460_ = ~new_n15420_ | ~new_n15335_;
  assign new_n15461_ = ~pi279 | ~new_n15387_;
  assign new_n15462_ = ~pi278 | ~new_n15386_;
  assign new_n15463_ = ~pi295 | ~new_n15389_;
  assign new_n15464_ = ~new_n15408_ | ~new_n15388_;
  assign new_n15465_ = ~pi291 | ~new_n15336_;
  assign new_n15466_ = ~new_n15405_ | ~new_n15391_;
  assign new_n15467_ = new_n4675_ & new_n15468_;
  assign new_n15468_ = ~new_n4672_;
  assign new_n15469_ = new_n15592_ & new_n15593_;
  assign new_n15470_ = new_n15594_ & new_n15595_;
  assign new_n15471_ = new_n15470_ & new_n15599_ & new_n15559_ & new_n15597_;
  assign new_n15472_ = new_n15606_ & new_n15607_;
  assign new_n15473_ = new_n15609_ & new_n15608_;
  assign new_n15474_ = new_n15563_ & new_n15562_ & new_n15610_;
  assign new_n15475_ = new_n15564_ & new_n15474_;
  assign new_n15476_ = new_n15625_ & new_n15624_;
  assign new_n15477_ = new_n15591_ & new_n15590_;
  assign new_n15478_ = new_n15548_ & new_n15483_;
  assign new_n15479_ = new_n15550_ & new_n15483_;
  assign new_n15480_ = new_n15552_ & new_n15483_;
  assign new_n15481_ = new_n15553_ & new_n15483_;
  assign new_n15482_ = new_n15582_ & new_n15483_;
  assign new_n15483_ = new_n15670_ & new_n15669_;
  assign new_n15484_ = ~new_n15583_ | ~new_n15477_ | ~new_n15667_ | ~new_n15666_;
  assign new_n15485_ = ~new_n4733_;
  assign new_n15486_ = ~new_n4701_;
  assign new_n15487_ = ~new_n4734_;
  assign new_n15488_ = ~new_n4702_;
  assign new_n15489_ = ~new_n4735_;
  assign new_n15490_ = ~new_n4703_;
  assign new_n15491_ = ~new_n4704_;
  assign new_n15492_ = ~new_n4706_;
  assign new_n15493_ = ~new_n4705_;
  assign new_n15494_ = ~new_n4739_;
  assign new_n15495_ = ~new_n4738_;
  assign new_n15496_ = ~new_n4737_;
  assign new_n15497_ = ~new_n4736_;
  assign new_n15498_ = ~new_n4741_;
  assign new_n15499_ = ~new_n4740_;
  assign new_n15500_ = ~new_n4711_;
  assign new_n15501_ = ~new_n4744_;
  assign new_n15502_ = ~new_n4712_;
  assign new_n15503_ = ~new_n4745_;
  assign new_n15504_ = ~new_n4746_;
  assign new_n15505_ = ~new_n4715_;
  assign new_n15506_ = ~new_n4747_;
  assign new_n15507_ = ~new_n4716_;
  assign new_n15508_ = ~new_n4714_;
  assign new_n15509_ = ~new_n4713_;
  assign new_n15510_ = ~new_n4748_;
  assign new_n15511_ = ~new_n4749_;
  assign new_n15512_ = ~new_n4717_;
  assign new_n15513_ = ~new_n4718_;
  assign new_n15514_ = ~new_n4758_;
  assign new_n15515_ = ~new_n4727_;
  assign new_n15516_ = ~new_n4724_;
  assign new_n15517_ = ~new_n4723_;
  assign new_n15518_ = ~new_n4759_;
  assign new_n15519_ = ~new_n4728_;
  assign new_n15520_ = ~new_n4726_;
  assign new_n15521_ = ~new_n4725_;
  assign new_n15522_ = ~new_n4729_;
  assign new_n15523_ = ~new_n4730_;
  assign new_n15524_ = ~new_n4731_;
  assign new_n15525_ = ~new_n4753_;
  assign new_n15526_ = ~new_n4752_;
  assign new_n15527_ = ~new_n4756_;
  assign new_n15528_ = ~new_n4757_;
  assign new_n15529_ = ~new_n4763_;
  assign new_n15530_ = ~new_n4762_;
  assign new_n15531_ = ~new_n4760_;
  assign new_n15532_ = ~new_n4761_;
  assign new_n15533_ = ~new_n4755_;
  assign new_n15534_ = ~new_n4754_;
  assign new_n15535_ = ~new_n4721_;
  assign new_n15536_ = ~new_n4722_;
  assign new_n15537_ = ~new_n4719_;
  assign new_n15538_ = ~new_n4720_;
  assign new_n15539_ = ~new_n4751_;
  assign new_n15540_ = ~new_n4750_;
  assign new_n15541_ = ~new_n4743_;
  assign new_n15542_ = ~new_n4742_;
  assign new_n15543_ = ~new_n4710_;
  assign new_n15544_ = ~new_n4709_;
  assign new_n15545_ = ~new_n4707_;
  assign new_n15546_ = ~new_n4708_;
  assign new_n15547_ = new_n15490_ & new_n4735_;
  assign new_n15548_ = new_n15586_ & new_n15588_ & new_n4739_ & new_n15587_ & new_n15545_;
  assign new_n15549_ = new_n4738_ & new_n15492_;
  assign new_n15550_ = new_n15586_ & new_n15549_ & new_n15588_;
  assign new_n15551_ = new_n4737_ & new_n15493_;
  assign new_n15552_ = new_n15551_ & new_n15586_;
  assign new_n15553_ = new_n4736_ & new_n15491_;
  assign new_n15554_ = new_n4744_ & new_n15502_;
  assign new_n15555_ = new_n4745_ & new_n15509_;
  assign new_n15556_ = new_n15645_ & new_n15644_;
  assign new_n15557_ = new_n4715_ & new_n15506_;
  assign new_n15558_ = new_n4716_ & new_n15510_;
  assign new_n15559_ = new_n15598_ & new_n15596_;
  assign new_n15560_ = new_n4727_ & new_n15518_;
  assign new_n15561_ = new_n4728_ & new_n15531_;
  assign new_n15562_ = new_n15611_ & new_n15605_;
  assign new_n15563_ = new_n15472_ & new_n15612_;
  assign new_n15564_ = new_n15614_ & new_n15613_;
  assign new_n15565_ = new_n15616_ & new_n15617_ & new_n15618_;
  assign new_n15566_ = new_n4756_ & new_n15516_;
  assign new_n15567_ = new_n4757_ & new_n15521_;
  assign new_n15568_ = new_n4763_ & new_n15524_;
  assign new_n15569_ = new_n4762_ & new_n15523_;
  assign new_n15570_ = new_n15476_ & new_n15571_;
  assign new_n15571_ = new_n15630_ & new_n15631_;
  assign new_n15572_ = new_n15629_ & new_n15570_;
  assign new_n15573_ = new_n4721_ & new_n15525_;
  assign new_n15574_ = new_n4722_ & new_n15534_;
  assign new_n15575_ = new_n15634_ & new_n15577_;
  assign new_n15576_ = new_n15575_ & new_n15635_;
  assign new_n15577_ = new_n15637_ & new_n15636_;
  assign new_n15578_ = new_n15601_ & new_n15648_ & new_n15647_;
  assign new_n15579_ = new_n15580_ & new_n15649_;
  assign new_n15580_ = new_n15652_ & new_n15651_;
  assign new_n15581_ = new_n15658_ & new_n15659_ & new_n15657_;
  assign new_n15582_ = new_n15586_ & new_n15588_ & new_n15581_ & new_n15653_ & new_n15587_;
  assign new_n15583_ = new_n15662_ & new_n15663_ & new_n15665_ & new_n15664_;
  assign new_n15584_ = ~new_n15661_ | ~new_n15660_;
  assign new_n15585_ = ~new_n4703_ | ~new_n15489_;
  assign new_n15586_ = ~new_n4704_ | ~new_n15497_;
  assign new_n15587_ = ~new_n4706_ | ~new_n15495_;
  assign new_n15588_ = ~new_n4705_ | ~new_n15496_;
  assign new_n15589_ = ~new_n4702_ | ~new_n15487_;
  assign new_n15590_ = ~new_n15668_ | ~new_n15672_ | ~new_n15671_;
  assign new_n15591_ = ~new_n15488_ | ~new_n15483_ | ~new_n4734_;
  assign new_n15592_ = ~new_n4746_ | ~new_n15508_;
  assign new_n15593_ = ~new_n4747_ | ~new_n15505_;
  assign new_n15594_ = ~new_n4711_ | ~new_n15541_;
  assign new_n15595_ = ~new_n4712_ | ~new_n15501_;
  assign new_n15596_ = ~new_n15557_ | ~new_n15592_;
  assign new_n15597_ = ~new_n15558_ | ~new_n15469_;
  assign new_n15598_ = ~new_n4714_ | ~new_n15504_;
  assign new_n15599_ = ~new_n4713_ | ~new_n15503_;
  assign new_n15600_ = ~new_n4717_ | ~new_n15511_;
  assign new_n15601_ = ~new_n4741_ | ~new_n15544_;
  assign new_n15602_ = ~new_n4740_ | ~new_n15546_;
  assign new_n15603_ = ~new_n4718_ | ~new_n15540_;
  assign new_n15604_ = ~new_n4758_ | ~new_n15520_;
  assign new_n15605_ = ~new_n15560_ | ~new_n15604_;
  assign new_n15606_ = ~new_n4723_ | ~new_n15533_;
  assign new_n15607_ = ~new_n4724_ | ~new_n15527_;
  assign new_n15608_ = ~new_n4759_ | ~new_n15515_;
  assign new_n15609_ = ~new_n4758_ | ~new_n15520_;
  assign new_n15610_ = ~new_n15561_ | ~new_n15473_;
  assign new_n15611_ = ~new_n4726_ | ~new_n15514_;
  assign new_n15612_ = ~new_n4725_ | ~new_n15528_;
  assign new_n15613_ = ~new_n4729_ | ~new_n15532_;
  assign new_n15614_ = ~new_n4730_ | ~new_n15530_;
  assign new_n15615_ = ~new_n4764_ | ~new_n4765_;
  assign new_n15616_ = ~new_n4732_ | ~new_n15615_;
  assign new_n15617_ = new_n4764_ | new_n4765_;
  assign new_n15618_ = ~new_n4731_ | ~new_n15529_;
  assign new_n15619_ = ~new_n15565_ | ~new_n15475_;
  assign new_n15620_ = ~new_n15569_ | ~new_n15613_;
  assign new_n15621_ = ~new_n4760_ | ~new_n15519_;
  assign new_n15622_ = ~new_n4761_ | ~new_n15522_;
  assign new_n15623_ = ~new_n15620_ | ~new_n15621_ | ~new_n15473_ | ~new_n15622_;
  assign new_n15624_ = ~new_n4753_ | ~new_n15535_;
  assign new_n15625_ = ~new_n4752_ | ~new_n15538_;
  assign new_n15626_ = ~new_n15566_ | ~new_n15606_;
  assign new_n15627_ = ~new_n15567_ | ~new_n15472_;
  assign new_n15628_ = ~new_n15568_ | ~new_n15475_;
  assign new_n15629_ = ~new_n15474_ | ~new_n15623_;
  assign new_n15630_ = ~new_n4755_ | ~new_n15517_;
  assign new_n15631_ = ~new_n4754_ | ~new_n15536_;
  assign new_n15632_ = ~new_n15572_ | ~new_n15619_ | ~new_n15626_ | ~new_n15628_ | ~new_n15627_;
  assign new_n15633_ = ~new_n4752_ | ~new_n15538_;
  assign new_n15634_ = ~new_n15573_ | ~new_n15633_;
  assign new_n15635_ = ~new_n15574_ | ~new_n15476_;
  assign new_n15636_ = ~new_n4719_ | ~new_n15539_;
  assign new_n15637_ = ~new_n4720_ | ~new_n15526_;
  assign new_n15638_ = ~new_n15632_ | ~new_n15576_;
  assign new_n15639_ = ~new_n4751_ | ~new_n15537_;
  assign new_n15640_ = ~new_n15639_ | ~new_n15638_;
  assign new_n15641_ = ~new_n15640_ | ~new_n15603_;
  assign new_n15642_ = ~new_n4750_ | ~new_n15513_;
  assign new_n15643_ = ~new_n15642_ | ~new_n15641_;
  assign new_n15644_ = ~new_n4748_ | ~new_n15507_;
  assign new_n15645_ = ~new_n4749_ | ~new_n15512_;
  assign new_n15646_ = ~new_n15556_ | ~new_n15469_;
  assign new_n15647_ = ~new_n15554_ | ~new_n15594_;
  assign new_n15648_ = ~new_n15555_ | ~new_n15470_;
  assign new_n15649_ = ~new_n15471_ | ~new_n15646_;
  assign new_n15650_ = ~new_n15471_ | ~new_n15643_ | ~new_n15600_;
  assign new_n15651_ = ~new_n4743_ | ~new_n15500_;
  assign new_n15652_ = ~new_n4742_ | ~new_n15543_;
  assign new_n15653_ = ~new_n15602_ | ~new_n15578_ | ~new_n15650_ | ~new_n15579_;
  assign new_n15654_ = ~new_n4710_ | ~new_n15542_;
  assign new_n15655_ = ~new_n4709_ | ~new_n15498_;
  assign new_n15656_ = ~new_n15655_ | ~new_n15654_;
  assign new_n15657_ = ~new_n15602_ | ~new_n15656_ | ~new_n15601_;
  assign new_n15658_ = ~new_n4707_ | ~new_n15494_;
  assign new_n15659_ = ~new_n4708_ | ~new_n15499_;
  assign new_n15660_ = ~new_n4734_ | ~new_n15585_;
  assign new_n15661_ = ~new_n15585_ | ~new_n15488_;
  assign new_n15662_ = ~new_n15589_ | ~new_n15547_ | ~new_n15483_;
  assign new_n15663_ = ~new_n15478_ | ~new_n15584_;
  assign new_n15664_ = ~new_n15479_ | ~new_n15584_;
  assign new_n15665_ = ~new_n15480_ | ~new_n15584_;
  assign new_n15666_ = ~new_n15481_ | ~new_n15584_;
  assign new_n15667_ = ~new_n15482_ | ~new_n15584_;
  assign new_n15668_ = ~new_n4701_ | ~new_n4733_;
  assign new_n15669_ = ~new_n4701_ | ~new_n15485_;
  assign new_n15670_ = ~new_n4733_ | ~new_n15486_;
  assign new_n15671_ = new_n4766_ | new_n4733_;
  assign new_n15672_ = ~new_n4766_ | ~new_n15486_;
  assign new_n15673_ = ~new_n4675_;
  assign new_n15674_ = ~new_n4672_;
  assign new_n15675_ = new_n15677_ & new_n15676_;
  assign new_n15676_ = ~new_n4672_ | ~new_n15673_;
  assign new_n15677_ = ~new_n4675_ | ~new_n15674_;
  assign new_n15678_ = new_n15769_ & new_n15768_;
  assign new_n15679_ = new_n15770_ & new_n15771_;
  assign new_n15680_ = new_n15787_ & new_n15786_;
  assign new_n15681_ = new_n15829_ & new_n15828_;
  assign new_n15682_ = new_n15838_ & new_n15837_;
  assign new_n15683_ = new_n15856_ & new_n15855_;
  assign new_n15684_ = new_n15892_ & new_n15889_;
  assign new_n15685_ = new_n15885_ & new_n15882_;
  assign new_n15686_ = new_n15876_ & new_n15873_;
  assign new_n15687_ = new_n15870_ & new_n15866_;
  assign new_n15688_ = new_n15825_ & new_n15822_;
  assign new_n15689_ = new_n15817_ & new_n15814_;
  assign new_n15690_ = new_n15803_ & new_n15800_;
  assign new_n15691_ = ~pi380;
  assign new_n15692_ = ~new_n5083_;
  assign new_n15693_ = ~new_n5086_;
  assign new_n15694_ = ~new_n5083_ | ~pi380;
  assign new_n15695_ = ~pi381;
  assign new_n15696_ = ~pi378;
  assign new_n15697_ = ~new_n5077_;
  assign new_n15698_ = ~new_n5080_;
  assign new_n15699_ = ~pi376;
  assign new_n15700_ = ~new_n5071_;
  assign new_n15701_ = ~pi374;
  assign new_n15702_ = ~new_n5062_;
  assign new_n15703_ = ~new_n5062_ | ~pi374;
  assign new_n15704_ = ~pi377;
  assign new_n15705_ = ~new_n5074_;
  assign new_n15706_ = ~new_n5077_ | ~pi378;
  assign new_n15707_ = ~pi379;
  assign new_n15708_ = ~pi382;
  assign new_n15709_ = ~new_n5089_;
  assign new_n15710_ = ~new_n5092_;
  assign new_n15711_ = ~pi383;
  assign new_n15712_ = ~new_n15723_ | ~new_n15795_;
  assign new_n15713_ = ~new_n15783_ | ~new_n15784_ | ~new_n15782_;
  assign new_n15714_ = ~new_n15772_ | ~new_n15773_;
  assign new_n15715_ = ~pi375 | ~new_n5068_;
  assign new_n15716_ = ~new_n15809_ | ~new_n15810_ | ~new_n15808_;
  assign new_n15717_ = ~new_n15806_ | ~new_n15805_;
  assign new_n15718_ = ~pi390;
  assign new_n15719_ = ~new_n5113_;
  assign new_n15720_ = ~new_n5116_;
  assign new_n15721_ = ~new_n5113_ | ~pi390;
  assign new_n15722_ = ~pi391;
  assign new_n15723_ = ~new_n5089_ | ~pi382;
  assign new_n15724_ = ~pi384;
  assign new_n15725_ = ~new_n5095_;
  assign new_n15726_ = ~pi386;
  assign new_n15727_ = ~new_n5101_;
  assign new_n15728_ = ~pi385;
  assign new_n15729_ = ~new_n5098_;
  assign new_n15730_ = ~new_n5098_ | ~pi385;
  assign new_n15731_ = ~pi387;
  assign new_n15732_ = ~new_n5104_;
  assign new_n15733_ = ~pi388;
  assign new_n15734_ = ~new_n5107_;
  assign new_n15735_ = ~pi389;
  assign new_n15736_ = ~new_n5110_;
  assign new_n15737_ = ~pi392;
  assign new_n15738_ = ~new_n5119_;
  assign new_n15739_ = ~new_n15861_ | ~new_n15860_ | ~new_n15859_;
  assign new_n15740_ = ~new_n15853_ | ~new_n15852_;
  assign new_n15741_ = ~new_n15730_ | ~new_n15878_;
  assign new_n15742_ = ~new_n15933_ | ~new_n15932_;
  assign new_n15743_ = ~new_n15982_ | ~new_n15981_;
  assign new_n15744_ = ~new_n15905_ | ~new_n15904_;
  assign new_n15745_ = ~new_n15910_ | ~new_n15909_;
  assign new_n15746_ = ~new_n15917_ | ~new_n15916_;
  assign new_n15747_ = ~new_n15924_ | ~new_n15923_;
  assign new_n15748_ = ~new_n15929_ | ~new_n15928_;
  assign new_n15749_ = ~new_n15945_ | ~new_n15944_;
  assign new_n15750_ = ~new_n15952_ | ~new_n15951_;
  assign new_n15751_ = ~new_n15959_ | ~new_n15958_;
  assign new_n15752_ = ~new_n15966_ | ~new_n15965_;
  assign new_n15753_ = ~new_n15973_ | ~new_n15972_;
  assign new_n15754_ = ~new_n15978_ | ~new_n15977_;
  assign new_n15755_ = ~new_n15792_ | ~new_n15791_ | ~new_n15790_;
  assign new_n15756_ = ~new_n15807_ | ~new_n15819_;
  assign new_n15757_ = ~new_n15715_ | ~new_n15826_;
  assign new_n15758_ = ~new_n5061_;
  assign new_n15759_ = ~pi393;
  assign new_n15760_ = ~new_n15849_ | ~new_n15848_;
  assign new_n15761_ = ~new_n15845_ | ~new_n15844_;
  assign new_n15762_ = ~new_n15835_ | ~new_n15834_;
  assign new_n15763_ = ~new_n15706_;
  assign new_n15764_ = ~pi383 | ~new_n5092_;
  assign new_n15765_ = ~new_n5101_ | ~pi386;
  assign new_n15766_ = ~new_n15730_;
  assign new_n15767_ = ~new_n15723_;
  assign new_n15768_ = new_n5080_ | pi379;
  assign new_n15769_ = new_n5077_ | pi378;
  assign new_n15770_ = pi377 | new_n5074_;
  assign new_n15771_ = pi376 | new_n5071_;
  assign new_n15772_ = ~new_n15703_;
  assign new_n15773_ = pi375 | new_n5068_;
  assign new_n15774_ = ~new_n15714_;
  assign new_n15775_ = ~new_n15715_;
  assign new_n15776_ = ~new_n15714_ | ~new_n15715_;
  assign new_n15777_ = ~new_n15770_ | ~pi376 | ~new_n5071_;
  assign new_n15778_ = ~new_n15679_ | ~new_n15776_;
  assign new_n15779_ = ~new_n5074_ | ~pi377;
  assign new_n15780_ = ~new_n15778_ | ~new_n15779_ | ~new_n15777_;
  assign new_n15781_ = ~new_n15707_ | ~new_n15706_;
  assign new_n15782_ = ~new_n5080_ | ~new_n15781_;
  assign new_n15783_ = ~new_n15678_ | ~new_n15780_;
  assign new_n15784_ = ~pi379 | ~new_n15763_;
  assign new_n15785_ = ~new_n15713_;
  assign new_n15786_ = new_n5086_ | pi381;
  assign new_n15787_ = new_n5083_ | pi380;
  assign new_n15788_ = ~new_n15694_;
  assign new_n15789_ = ~new_n15695_ | ~new_n15694_;
  assign new_n15790_ = ~new_n5086_ | ~new_n15789_;
  assign new_n15791_ = ~pi381 | ~new_n15788_;
  assign new_n15792_ = ~new_n15680_ | ~new_n15713_;
  assign new_n15793_ = ~new_n15755_;
  assign new_n15794_ = pi382 | new_n5089_;
  assign new_n15795_ = ~new_n15794_ | ~new_n15755_;
  assign new_n15796_ = ~new_n15712_;
  assign new_n15797_ = new_n5092_ | pi383;
  assign new_n15798_ = pi380 | new_n5083_;
  assign new_n15799_ = ~new_n15798_ | ~new_n15713_;
  assign new_n15800_ = ~new_n15799_ | ~new_n15694_ | ~new_n15912_ | ~new_n15911_;
  assign new_n15801_ = ~new_n15785_ | ~new_n15694_;
  assign new_n15802_ = ~pi381 | ~new_n5086_;
  assign new_n15803_ = ~new_n15801_ | ~new_n15802_ | ~new_n15680_;
  assign new_n15804_ = new_n5083_ | pi380;
  assign new_n15805_ = ~new_n15775_ | ~new_n15771_;
  assign new_n15806_ = ~new_n5071_ | ~pi376;
  assign new_n15807_ = ~new_n15717_;
  assign new_n15808_ = ~new_n15774_ | ~new_n15679_;
  assign new_n15809_ = ~new_n15717_ | ~new_n15770_;
  assign new_n15810_ = ~new_n5074_ | ~pi377;
  assign new_n15811_ = ~new_n15716_;
  assign new_n15812_ = pi378 | new_n5077_;
  assign new_n15813_ = ~new_n15812_ | ~new_n15716_;
  assign new_n15814_ = ~new_n15813_ | ~new_n15706_ | ~new_n15919_ | ~new_n15918_;
  assign new_n15815_ = ~new_n15811_ | ~new_n15706_;
  assign new_n15816_ = ~pi379 | ~new_n5080_;
  assign new_n15817_ = ~new_n15815_ | ~new_n15816_ | ~new_n15678_;
  assign new_n15818_ = new_n5077_ | pi378;
  assign new_n15819_ = ~new_n15774_ | ~new_n15771_;
  assign new_n15820_ = ~new_n15756_;
  assign new_n15821_ = ~new_n5074_ | ~pi377;
  assign new_n15822_ = ~new_n15714_ | ~new_n15715_ | ~new_n15931_ | ~new_n15930_;
  assign new_n15823_ = ~new_n15715_ | ~new_n15714_;
  assign new_n15824_ = ~new_n5071_ | ~pi376;
  assign new_n15825_ = ~new_n15823_ | ~new_n15824_ | ~new_n15771_;
  assign new_n15826_ = pi375 | new_n5068_;
  assign new_n15827_ = ~new_n15757_;
  assign new_n15828_ = new_n5092_ | pi383;
  assign new_n15829_ = new_n5095_ | pi384;
  assign new_n15830_ = ~new_n15767_ | ~new_n15681_;
  assign new_n15831_ = ~new_n5095_ | ~pi384;
  assign new_n15832_ = ~new_n15830_ | ~new_n15831_ | ~new_n15764_;
  assign new_n15833_ = pi384 | new_n5095_;
  assign new_n15834_ = ~new_n15755_ | ~new_n15794_ | ~new_n15681_;
  assign new_n15835_ = ~new_n15833_ | ~new_n15832_;
  assign new_n15836_ = ~new_n15762_;
  assign new_n15837_ = new_n5104_ | pi387;
  assign new_n15838_ = new_n5101_ | pi386;
  assign new_n15839_ = ~new_n15766_ | ~new_n15682_;
  assign new_n15840_ = ~new_n5104_ | ~pi387;
  assign new_n15841_ = ~new_n15839_ | ~new_n15840_ | ~new_n15765_;
  assign new_n15842_ = pi385 | new_n5098_;
  assign new_n15843_ = pi387 | new_n5104_;
  assign new_n15844_ = ~new_n15762_ | ~new_n15842_ | ~new_n15682_;
  assign new_n15845_ = ~new_n15843_ | ~new_n15841_;
  assign new_n15846_ = ~new_n15761_;
  assign new_n15847_ = pi388 | new_n5107_;
  assign new_n15848_ = ~new_n15847_ | ~new_n15761_;
  assign new_n15849_ = ~new_n5107_ | ~pi388;
  assign new_n15850_ = ~new_n15760_;
  assign new_n15851_ = pi389 | new_n5110_;
  assign new_n15852_ = ~new_n15851_ | ~new_n15760_;
  assign new_n15853_ = ~new_n5110_ | ~pi389;
  assign new_n15854_ = ~new_n15740_;
  assign new_n15855_ = new_n5116_ | pi391;
  assign new_n15856_ = new_n5113_ | pi390;
  assign new_n15857_ = ~new_n15721_;
  assign new_n15858_ = ~new_n15722_ | ~new_n15721_;
  assign new_n15859_ = ~new_n5116_ | ~new_n15858_;
  assign new_n15860_ = ~pi391 | ~new_n15857_;
  assign new_n15861_ = ~new_n15683_ | ~new_n15740_;
  assign new_n15862_ = ~new_n15739_;
  assign new_n15863_ = pi392 | new_n5119_;
  assign new_n15864_ = ~new_n15863_ | ~new_n15739_;
  assign new_n15865_ = ~new_n5119_ | ~pi392;
  assign new_n15866_ = ~new_n15864_ | ~new_n15865_ | ~new_n15935_ | ~new_n15934_;
  assign new_n15867_ = ~new_n5119_ | ~pi392;
  assign new_n15868_ = ~new_n15862_ | ~new_n15867_;
  assign new_n15869_ = new_n5119_ | pi392;
  assign new_n15870_ = ~new_n15868_ | ~new_n15869_ | ~new_n15938_;
  assign new_n15871_ = pi390 | new_n5113_;
  assign new_n15872_ = ~new_n15871_ | ~new_n15740_;
  assign new_n15873_ = ~new_n15872_ | ~new_n15721_ | ~new_n15947_ | ~new_n15946_;
  assign new_n15874_ = ~new_n15854_ | ~new_n15721_;
  assign new_n15875_ = ~pi391 | ~new_n5116_;
  assign new_n15876_ = ~new_n15874_ | ~new_n15875_ | ~new_n15683_;
  assign new_n15877_ = new_n5113_ | pi390;
  assign new_n15878_ = ~new_n15842_ | ~new_n15762_;
  assign new_n15879_ = ~new_n15741_;
  assign new_n15880_ = pi386 | new_n5101_;
  assign new_n15881_ = ~new_n15880_ | ~new_n15741_;
  assign new_n15882_ = ~new_n15881_ | ~new_n15765_ | ~new_n15968_ | ~new_n15967_;
  assign new_n15883_ = ~new_n15879_ | ~new_n15765_;
  assign new_n15884_ = ~new_n5104_ | ~pi387;
  assign new_n15885_ = ~new_n15883_ | ~new_n15884_ | ~new_n15682_;
  assign new_n15886_ = new_n5101_ | pi386;
  assign new_n15887_ = pi383 | new_n5092_;
  assign new_n15888_ = ~new_n15887_ | ~new_n15712_;
  assign new_n15889_ = ~new_n15888_ | ~new_n15764_ | ~new_n15980_ | ~new_n15979_;
  assign new_n15890_ = ~new_n15796_ | ~new_n15764_;
  assign new_n15891_ = ~new_n5095_ | ~pi384;
  assign new_n15892_ = ~new_n15890_ | ~new_n15891_ | ~new_n15681_;
  assign new_n15893_ = ~new_n15797_ | ~new_n15764_;
  assign new_n15894_ = ~new_n15794_ | ~new_n15723_;
  assign new_n15895_ = ~new_n15804_ | ~new_n15694_;
  assign new_n15896_ = ~new_n15818_ | ~new_n15706_;
  assign new_n15897_ = ~new_n15821_ | ~new_n15770_;
  assign new_n15898_ = ~new_n15877_ | ~new_n15721_;
  assign new_n15899_ = ~new_n15886_ | ~new_n15765_;
  assign new_n15900_ = ~new_n15842_ | ~new_n15730_;
  assign new_n15901_ = ~new_n5092_ | ~new_n15711_;
  assign new_n15902_ = ~pi383 | ~new_n15710_;
  assign new_n15903_ = ~new_n15902_ | ~new_n15901_;
  assign new_n15904_ = ~new_n15893_ | ~new_n15712_;
  assign new_n15905_ = ~new_n15903_ | ~new_n15796_;
  assign new_n15906_ = ~new_n5089_ | ~new_n15708_;
  assign new_n15907_ = ~pi382 | ~new_n15709_;
  assign new_n15908_ = ~new_n15907_ | ~new_n15906_;
  assign new_n15909_ = ~new_n15894_ | ~new_n15755_;
  assign new_n15910_ = ~new_n15793_ | ~new_n15908_;
  assign new_n15911_ = ~new_n5086_ | ~new_n15695_;
  assign new_n15912_ = ~pi381 | ~new_n15693_;
  assign new_n15913_ = ~new_n5083_ | ~new_n15691_;
  assign new_n15914_ = ~pi380 | ~new_n15692_;
  assign new_n15915_ = ~new_n15914_ | ~new_n15913_;
  assign new_n15916_ = ~new_n15895_ | ~new_n15713_;
  assign new_n15917_ = ~new_n15915_ | ~new_n15785_;
  assign new_n15918_ = ~new_n5080_ | ~new_n15707_;
  assign new_n15919_ = ~pi379 | ~new_n15698_;
  assign new_n15920_ = ~new_n5077_ | ~new_n15696_;
  assign new_n15921_ = ~pi378 | ~new_n15697_;
  assign new_n15922_ = ~new_n15921_ | ~new_n15920_;
  assign new_n15923_ = ~new_n15896_ | ~new_n15716_;
  assign new_n15924_ = ~new_n15922_ | ~new_n15811_;
  assign new_n15925_ = ~new_n5074_ | ~new_n15704_;
  assign new_n15926_ = ~pi377 | ~new_n15705_;
  assign new_n15927_ = ~new_n15926_ | ~new_n15925_;
  assign new_n15928_ = ~new_n15897_ | ~new_n15756_;
  assign new_n15929_ = ~new_n15820_ | ~new_n15927_;
  assign new_n15930_ = ~new_n5071_ | ~new_n15699_;
  assign new_n15931_ = ~pi376 | ~new_n15700_;
  assign new_n15932_ = ~new_n15772_ | ~new_n15757_;
  assign new_n15933_ = ~new_n15827_ | ~new_n15703_;
  assign new_n15934_ = ~new_n5061_ | ~new_n15759_;
  assign new_n15935_ = ~pi393 | ~new_n15758_;
  assign new_n15936_ = ~new_n5061_ | ~new_n15759_;
  assign new_n15937_ = ~pi393 | ~new_n15758_;
  assign new_n15938_ = ~new_n15937_ | ~new_n15936_;
  assign new_n15939_ = ~new_n5119_ | ~new_n15737_;
  assign new_n15940_ = ~pi392 | ~new_n15738_;
  assign new_n15941_ = ~new_n5119_ | ~new_n15737_;
  assign new_n15942_ = ~pi392 | ~new_n15738_;
  assign new_n15943_ = ~new_n15942_ | ~new_n15941_;
  assign new_n15944_ = ~new_n15739_ | ~new_n15940_ | ~new_n15939_;
  assign new_n15945_ = ~new_n15943_ | ~new_n15862_;
  assign new_n15946_ = ~new_n5116_ | ~new_n15722_;
  assign new_n15947_ = ~pi391 | ~new_n15720_;
  assign new_n15948_ = ~new_n5113_ | ~new_n15718_;
  assign new_n15949_ = ~pi390 | ~new_n15719_;
  assign new_n15950_ = ~new_n15949_ | ~new_n15948_;
  assign new_n15951_ = ~new_n15898_ | ~new_n15740_;
  assign new_n15952_ = ~new_n15950_ | ~new_n15854_;
  assign new_n15953_ = ~new_n5110_ | ~new_n15735_;
  assign new_n15954_ = ~pi389 | ~new_n15736_;
  assign new_n15955_ = ~new_n5110_ | ~new_n15735_;
  assign new_n15956_ = ~pi389 | ~new_n15736_;
  assign new_n15957_ = ~new_n15956_ | ~new_n15955_;
  assign new_n15958_ = ~new_n15760_ | ~new_n15954_ | ~new_n15953_;
  assign new_n15959_ = ~new_n15850_ | ~new_n15957_;
  assign new_n15960_ = ~new_n5107_ | ~new_n15733_;
  assign new_n15961_ = ~pi388 | ~new_n15734_;
  assign new_n15962_ = ~new_n5107_ | ~new_n15733_;
  assign new_n15963_ = ~pi388 | ~new_n15734_;
  assign new_n15964_ = ~new_n15963_ | ~new_n15962_;
  assign new_n15965_ = ~new_n15761_ | ~new_n15961_ | ~new_n15960_;
  assign new_n15966_ = ~new_n15846_ | ~new_n15964_;
  assign new_n15967_ = ~new_n5104_ | ~new_n15731_;
  assign new_n15968_ = ~pi387 | ~new_n15732_;
  assign new_n15969_ = ~new_n5101_ | ~new_n15726_;
  assign new_n15970_ = ~pi386 | ~new_n15727_;
  assign new_n15971_ = ~new_n15970_ | ~new_n15969_;
  assign new_n15972_ = ~new_n15899_ | ~new_n15741_;
  assign new_n15973_ = ~new_n15971_ | ~new_n15879_;
  assign new_n15974_ = ~new_n5098_ | ~new_n15728_;
  assign new_n15975_ = ~pi385 | ~new_n15729_;
  assign new_n15976_ = ~new_n15975_ | ~new_n15974_;
  assign new_n15977_ = ~new_n15900_ | ~new_n15762_;
  assign new_n15978_ = ~new_n15836_ | ~new_n15976_;
  assign new_n15979_ = ~new_n5095_ | ~new_n15724_;
  assign new_n15980_ = ~pi384 | ~new_n15725_;
  assign new_n15981_ = ~new_n5062_ | ~new_n15701_;
  assign new_n15982_ = ~pi374 | ~new_n15702_;
  assign new_n15983_ = new_n16074_ & new_n16073_;
  assign new_n15984_ = new_n16075_ & new_n16076_;
  assign new_n15985_ = new_n16092_ & new_n16091_;
  assign new_n15986_ = new_n16134_ & new_n16133_;
  assign new_n15987_ = new_n16143_ & new_n16142_;
  assign new_n15988_ = new_n16161_ & new_n16160_;
  assign new_n15989_ = new_n16197_ & new_n16194_;
  assign new_n15990_ = new_n16190_ & new_n16187_;
  assign new_n15991_ = new_n16181_ & new_n16178_;
  assign new_n15992_ = new_n16175_ & new_n16171_;
  assign new_n15993_ = new_n16130_ & new_n16127_;
  assign new_n15994_ = new_n16122_ & new_n16119_;
  assign new_n15995_ = new_n16108_ & new_n16105_;
  assign new_n15996_ = ~pi412;
  assign new_n15997_ = ~new_n5083_;
  assign new_n15998_ = ~new_n5086_;
  assign new_n15999_ = ~new_n5083_ | ~pi412;
  assign new_n16000_ = ~pi413;
  assign new_n16001_ = ~pi410;
  assign new_n16002_ = ~new_n5077_;
  assign new_n16003_ = ~new_n5080_;
  assign new_n16004_ = ~pi408;
  assign new_n16005_ = ~new_n5071_;
  assign new_n16006_ = ~pi406;
  assign new_n16007_ = ~new_n5062_;
  assign new_n16008_ = ~new_n5062_ | ~pi406;
  assign new_n16009_ = ~pi409;
  assign new_n16010_ = ~new_n5074_;
  assign new_n16011_ = ~new_n5077_ | ~pi410;
  assign new_n16012_ = ~pi411;
  assign new_n16013_ = ~pi414;
  assign new_n16014_ = ~new_n5089_;
  assign new_n16015_ = ~new_n5092_;
  assign new_n16016_ = ~pi415;
  assign new_n16017_ = ~new_n16028_ | ~new_n16100_;
  assign new_n16018_ = ~new_n16088_ | ~new_n16089_ | ~new_n16087_;
  assign new_n16019_ = ~new_n16077_ | ~new_n16078_;
  assign new_n16020_ = ~pi407 | ~new_n5068_;
  assign new_n16021_ = ~new_n16114_ | ~new_n16115_ | ~new_n16113_;
  assign new_n16022_ = ~new_n16111_ | ~new_n16110_;
  assign new_n16023_ = ~pi422;
  assign new_n16024_ = ~new_n5113_;
  assign new_n16025_ = ~new_n5116_;
  assign new_n16026_ = ~new_n5113_ | ~pi422;
  assign new_n16027_ = ~pi423;
  assign new_n16028_ = ~new_n5089_ | ~pi414;
  assign new_n16029_ = ~pi416;
  assign new_n16030_ = ~new_n5095_;
  assign new_n16031_ = ~pi418;
  assign new_n16032_ = ~new_n5101_;
  assign new_n16033_ = ~pi417;
  assign new_n16034_ = ~new_n5098_;
  assign new_n16035_ = ~new_n5098_ | ~pi417;
  assign new_n16036_ = ~pi419;
  assign new_n16037_ = ~new_n5104_;
  assign new_n16038_ = ~pi420;
  assign new_n16039_ = ~new_n5107_;
  assign new_n16040_ = ~pi421;
  assign new_n16041_ = ~new_n5110_;
  assign new_n16042_ = ~pi424;
  assign new_n16043_ = ~new_n5119_;
  assign new_n16044_ = ~new_n16166_ | ~new_n16165_ | ~new_n16164_;
  assign new_n16045_ = ~new_n16158_ | ~new_n16157_;
  assign new_n16046_ = ~new_n16035_ | ~new_n16183_;
  assign new_n16047_ = ~new_n16238_ | ~new_n16237_;
  assign new_n16048_ = ~new_n16287_ | ~new_n16286_;
  assign new_n16049_ = ~new_n16210_ | ~new_n16209_;
  assign new_n16050_ = ~new_n16215_ | ~new_n16214_;
  assign new_n16051_ = ~new_n16222_ | ~new_n16221_;
  assign new_n16052_ = ~new_n16229_ | ~new_n16228_;
  assign new_n16053_ = ~new_n16234_ | ~new_n16233_;
  assign new_n16054_ = ~new_n16250_ | ~new_n16249_;
  assign new_n16055_ = ~new_n16257_ | ~new_n16256_;
  assign new_n16056_ = ~new_n16264_ | ~new_n16263_;
  assign new_n16057_ = ~new_n16271_ | ~new_n16270_;
  assign new_n16058_ = ~new_n16278_ | ~new_n16277_;
  assign new_n16059_ = ~new_n16283_ | ~new_n16282_;
  assign new_n16060_ = ~new_n16097_ | ~new_n16096_ | ~new_n16095_;
  assign new_n16061_ = ~new_n16112_ | ~new_n16124_;
  assign new_n16062_ = ~new_n16020_ | ~new_n16131_;
  assign new_n16063_ = ~new_n5061_;
  assign new_n16064_ = ~pi425;
  assign new_n16065_ = ~new_n16154_ | ~new_n16153_;
  assign new_n16066_ = ~new_n16150_ | ~new_n16149_;
  assign new_n16067_ = ~new_n16140_ | ~new_n16139_;
  assign new_n16068_ = ~new_n16011_;
  assign new_n16069_ = ~pi415 | ~new_n5092_;
  assign new_n16070_ = ~new_n5101_ | ~pi418;
  assign new_n16071_ = ~new_n16035_;
  assign new_n16072_ = ~new_n16028_;
  assign new_n16073_ = new_n5080_ | pi411;
  assign new_n16074_ = new_n5077_ | pi410;
  assign new_n16075_ = pi409 | new_n5074_;
  assign new_n16076_ = pi408 | new_n5071_;
  assign new_n16077_ = ~new_n16008_;
  assign new_n16078_ = pi407 | new_n5068_;
  assign new_n16079_ = ~new_n16019_;
  assign new_n16080_ = ~new_n16020_;
  assign new_n16081_ = ~new_n16019_ | ~new_n16020_;
  assign new_n16082_ = ~new_n16075_ | ~pi408 | ~new_n5071_;
  assign new_n16083_ = ~new_n15984_ | ~new_n16081_;
  assign new_n16084_ = ~new_n5074_ | ~pi409;
  assign new_n16085_ = ~new_n16083_ | ~new_n16084_ | ~new_n16082_;
  assign new_n16086_ = ~new_n16012_ | ~new_n16011_;
  assign new_n16087_ = ~new_n5080_ | ~new_n16086_;
  assign new_n16088_ = ~new_n15983_ | ~new_n16085_;
  assign new_n16089_ = ~pi411 | ~new_n16068_;
  assign new_n16090_ = ~new_n16018_;
  assign new_n16091_ = new_n5086_ | pi413;
  assign new_n16092_ = new_n5083_ | pi412;
  assign new_n16093_ = ~new_n15999_;
  assign new_n16094_ = ~new_n16000_ | ~new_n15999_;
  assign new_n16095_ = ~new_n5086_ | ~new_n16094_;
  assign new_n16096_ = ~pi413 | ~new_n16093_;
  assign new_n16097_ = ~new_n15985_ | ~new_n16018_;
  assign new_n16098_ = ~new_n16060_;
  assign new_n16099_ = pi414 | new_n5089_;
  assign new_n16100_ = ~new_n16099_ | ~new_n16060_;
  assign new_n16101_ = ~new_n16017_;
  assign new_n16102_ = new_n5092_ | pi415;
  assign new_n16103_ = pi412 | new_n5083_;
  assign new_n16104_ = ~new_n16103_ | ~new_n16018_;
  assign new_n16105_ = ~new_n16104_ | ~new_n15999_ | ~new_n16217_ | ~new_n16216_;
  assign new_n16106_ = ~new_n16090_ | ~new_n15999_;
  assign new_n16107_ = ~pi413 | ~new_n5086_;
  assign new_n16108_ = ~new_n16106_ | ~new_n16107_ | ~new_n15985_;
  assign new_n16109_ = new_n5083_ | pi412;
  assign new_n16110_ = ~new_n16080_ | ~new_n16076_;
  assign new_n16111_ = ~new_n5071_ | ~pi408;
  assign new_n16112_ = ~new_n16022_;
  assign new_n16113_ = ~new_n16079_ | ~new_n15984_;
  assign new_n16114_ = ~new_n16022_ | ~new_n16075_;
  assign new_n16115_ = ~new_n5074_ | ~pi409;
  assign new_n16116_ = ~new_n16021_;
  assign new_n16117_ = pi410 | new_n5077_;
  assign new_n16118_ = ~new_n16117_ | ~new_n16021_;
  assign new_n16119_ = ~new_n16118_ | ~new_n16011_ | ~new_n16224_ | ~new_n16223_;
  assign new_n16120_ = ~new_n16116_ | ~new_n16011_;
  assign new_n16121_ = ~pi411 | ~new_n5080_;
  assign new_n16122_ = ~new_n16120_ | ~new_n16121_ | ~new_n15983_;
  assign new_n16123_ = new_n5077_ | pi410;
  assign new_n16124_ = ~new_n16079_ | ~new_n16076_;
  assign new_n16125_ = ~new_n16061_;
  assign new_n16126_ = ~new_n5074_ | ~pi409;
  assign new_n16127_ = ~new_n16019_ | ~new_n16020_ | ~new_n16236_ | ~new_n16235_;
  assign new_n16128_ = ~new_n16020_ | ~new_n16019_;
  assign new_n16129_ = ~new_n5071_ | ~pi408;
  assign new_n16130_ = ~new_n16128_ | ~new_n16129_ | ~new_n16076_;
  assign new_n16131_ = pi407 | new_n5068_;
  assign new_n16132_ = ~new_n16062_;
  assign new_n16133_ = new_n5092_ | pi415;
  assign new_n16134_ = new_n5095_ | pi416;
  assign new_n16135_ = ~new_n16072_ | ~new_n15986_;
  assign new_n16136_ = ~new_n5095_ | ~pi416;
  assign new_n16137_ = ~new_n16135_ | ~new_n16136_ | ~new_n16069_;
  assign new_n16138_ = pi416 | new_n5095_;
  assign new_n16139_ = ~new_n16060_ | ~new_n16099_ | ~new_n15986_;
  assign new_n16140_ = ~new_n16138_ | ~new_n16137_;
  assign new_n16141_ = ~new_n16067_;
  assign new_n16142_ = new_n5104_ | pi419;
  assign new_n16143_ = new_n5101_ | pi418;
  assign new_n16144_ = ~new_n16071_ | ~new_n15987_;
  assign new_n16145_ = ~new_n5104_ | ~pi419;
  assign new_n16146_ = ~new_n16144_ | ~new_n16145_ | ~new_n16070_;
  assign new_n16147_ = pi417 | new_n5098_;
  assign new_n16148_ = pi419 | new_n5104_;
  assign new_n16149_ = ~new_n16067_ | ~new_n16147_ | ~new_n15987_;
  assign new_n16150_ = ~new_n16148_ | ~new_n16146_;
  assign new_n16151_ = ~new_n16066_;
  assign new_n16152_ = pi420 | new_n5107_;
  assign new_n16153_ = ~new_n16152_ | ~new_n16066_;
  assign new_n16154_ = ~new_n5107_ | ~pi420;
  assign new_n16155_ = ~new_n16065_;
  assign new_n16156_ = pi421 | new_n5110_;
  assign new_n16157_ = ~new_n16156_ | ~new_n16065_;
  assign new_n16158_ = ~new_n5110_ | ~pi421;
  assign new_n16159_ = ~new_n16045_;
  assign new_n16160_ = new_n5116_ | pi423;
  assign new_n16161_ = new_n5113_ | pi422;
  assign new_n16162_ = ~new_n16026_;
  assign new_n16163_ = ~new_n16027_ | ~new_n16026_;
  assign new_n16164_ = ~new_n5116_ | ~new_n16163_;
  assign new_n16165_ = ~pi423 | ~new_n16162_;
  assign new_n16166_ = ~new_n15988_ | ~new_n16045_;
  assign new_n16167_ = ~new_n16044_;
  assign new_n16168_ = pi424 | new_n5119_;
  assign new_n16169_ = ~new_n16168_ | ~new_n16044_;
  assign new_n16170_ = ~new_n5119_ | ~pi424;
  assign new_n16171_ = ~new_n16169_ | ~new_n16170_ | ~new_n16240_ | ~new_n16239_;
  assign new_n16172_ = ~new_n5119_ | ~pi424;
  assign new_n16173_ = ~new_n16167_ | ~new_n16172_;
  assign new_n16174_ = new_n5119_ | pi424;
  assign new_n16175_ = ~new_n16173_ | ~new_n16174_ | ~new_n16243_;
  assign new_n16176_ = pi422 | new_n5113_;
  assign new_n16177_ = ~new_n16176_ | ~new_n16045_;
  assign new_n16178_ = ~new_n16177_ | ~new_n16026_ | ~new_n16252_ | ~new_n16251_;
  assign new_n16179_ = ~new_n16159_ | ~new_n16026_;
  assign new_n16180_ = ~pi423 | ~new_n5116_;
  assign new_n16181_ = ~new_n16179_ | ~new_n16180_ | ~new_n15988_;
  assign new_n16182_ = new_n5113_ | pi422;
  assign new_n16183_ = ~new_n16147_ | ~new_n16067_;
  assign new_n16184_ = ~new_n16046_;
  assign new_n16185_ = pi418 | new_n5101_;
  assign new_n16186_ = ~new_n16185_ | ~new_n16046_;
  assign new_n16187_ = ~new_n16186_ | ~new_n16070_ | ~new_n16273_ | ~new_n16272_;
  assign new_n16188_ = ~new_n16184_ | ~new_n16070_;
  assign new_n16189_ = ~new_n5104_ | ~pi419;
  assign new_n16190_ = ~new_n16188_ | ~new_n16189_ | ~new_n15987_;
  assign new_n16191_ = new_n5101_ | pi418;
  assign new_n16192_ = pi415 | new_n5092_;
  assign new_n16193_ = ~new_n16192_ | ~new_n16017_;
  assign new_n16194_ = ~new_n16193_ | ~new_n16069_ | ~new_n16285_ | ~new_n16284_;
  assign new_n16195_ = ~new_n16101_ | ~new_n16069_;
  assign new_n16196_ = ~new_n5095_ | ~pi416;
  assign new_n16197_ = ~new_n16195_ | ~new_n16196_ | ~new_n15986_;
  assign new_n16198_ = ~new_n16102_ | ~new_n16069_;
  assign new_n16199_ = ~new_n16099_ | ~new_n16028_;
  assign new_n16200_ = ~new_n16109_ | ~new_n15999_;
  assign new_n16201_ = ~new_n16123_ | ~new_n16011_;
  assign new_n16202_ = ~new_n16126_ | ~new_n16075_;
  assign new_n16203_ = ~new_n16182_ | ~new_n16026_;
  assign new_n16204_ = ~new_n16191_ | ~new_n16070_;
  assign new_n16205_ = ~new_n16147_ | ~new_n16035_;
  assign new_n16206_ = ~new_n5092_ | ~new_n16016_;
  assign new_n16207_ = ~pi415 | ~new_n16015_;
  assign new_n16208_ = ~new_n16207_ | ~new_n16206_;
  assign new_n16209_ = ~new_n16198_ | ~new_n16017_;
  assign new_n16210_ = ~new_n16208_ | ~new_n16101_;
  assign new_n16211_ = ~new_n5089_ | ~new_n16013_;
  assign new_n16212_ = ~pi414 | ~new_n16014_;
  assign new_n16213_ = ~new_n16212_ | ~new_n16211_;
  assign new_n16214_ = ~new_n16199_ | ~new_n16060_;
  assign new_n16215_ = ~new_n16098_ | ~new_n16213_;
  assign new_n16216_ = ~new_n5086_ | ~new_n16000_;
  assign new_n16217_ = ~pi413 | ~new_n15998_;
  assign new_n16218_ = ~new_n5083_ | ~new_n15996_;
  assign new_n16219_ = ~pi412 | ~new_n15997_;
  assign new_n16220_ = ~new_n16219_ | ~new_n16218_;
  assign new_n16221_ = ~new_n16200_ | ~new_n16018_;
  assign new_n16222_ = ~new_n16220_ | ~new_n16090_;
  assign new_n16223_ = ~new_n5080_ | ~new_n16012_;
  assign new_n16224_ = ~pi411 | ~new_n16003_;
  assign new_n16225_ = ~new_n5077_ | ~new_n16001_;
  assign new_n16226_ = ~pi410 | ~new_n16002_;
  assign new_n16227_ = ~new_n16226_ | ~new_n16225_;
  assign new_n16228_ = ~new_n16201_ | ~new_n16021_;
  assign new_n16229_ = ~new_n16227_ | ~new_n16116_;
  assign new_n16230_ = ~new_n5074_ | ~new_n16009_;
  assign new_n16231_ = ~pi409 | ~new_n16010_;
  assign new_n16232_ = ~new_n16231_ | ~new_n16230_;
  assign new_n16233_ = ~new_n16202_ | ~new_n16061_;
  assign new_n16234_ = ~new_n16125_ | ~new_n16232_;
  assign new_n16235_ = ~new_n5071_ | ~new_n16004_;
  assign new_n16236_ = ~pi408 | ~new_n16005_;
  assign new_n16237_ = ~new_n16077_ | ~new_n16062_;
  assign new_n16238_ = ~new_n16132_ | ~new_n16008_;
  assign new_n16239_ = ~new_n5061_ | ~new_n16064_;
  assign new_n16240_ = ~pi425 | ~new_n16063_;
  assign new_n16241_ = ~new_n5061_ | ~new_n16064_;
  assign new_n16242_ = ~pi425 | ~new_n16063_;
  assign new_n16243_ = ~new_n16242_ | ~new_n16241_;
  assign new_n16244_ = ~new_n5119_ | ~new_n16042_;
  assign new_n16245_ = ~pi424 | ~new_n16043_;
  assign new_n16246_ = ~new_n5119_ | ~new_n16042_;
  assign new_n16247_ = ~pi424 | ~new_n16043_;
  assign new_n16248_ = ~new_n16247_ | ~new_n16246_;
  assign new_n16249_ = ~new_n16044_ | ~new_n16245_ | ~new_n16244_;
  assign new_n16250_ = ~new_n16248_ | ~new_n16167_;
  assign new_n16251_ = ~new_n5116_ | ~new_n16027_;
  assign new_n16252_ = ~pi423 | ~new_n16025_;
  assign new_n16253_ = ~new_n5113_ | ~new_n16023_;
  assign new_n16254_ = ~pi422 | ~new_n16024_;
  assign new_n16255_ = ~new_n16254_ | ~new_n16253_;
  assign new_n16256_ = ~new_n16203_ | ~new_n16045_;
  assign new_n16257_ = ~new_n16255_ | ~new_n16159_;
  assign new_n16258_ = ~new_n5110_ | ~new_n16040_;
  assign new_n16259_ = ~pi421 | ~new_n16041_;
  assign new_n16260_ = ~new_n5110_ | ~new_n16040_;
  assign new_n16261_ = ~pi421 | ~new_n16041_;
  assign new_n16262_ = ~new_n16261_ | ~new_n16260_;
  assign new_n16263_ = ~new_n16065_ | ~new_n16259_ | ~new_n16258_;
  assign new_n16264_ = ~new_n16155_ | ~new_n16262_;
  assign new_n16265_ = ~new_n5107_ | ~new_n16038_;
  assign new_n16266_ = ~pi420 | ~new_n16039_;
  assign new_n16267_ = ~new_n5107_ | ~new_n16038_;
  assign new_n16268_ = ~pi420 | ~new_n16039_;
  assign new_n16269_ = ~new_n16268_ | ~new_n16267_;
  assign new_n16270_ = ~new_n16066_ | ~new_n16266_ | ~new_n16265_;
  assign new_n16271_ = ~new_n16151_ | ~new_n16269_;
  assign new_n16272_ = ~new_n5104_ | ~new_n16036_;
  assign new_n16273_ = ~pi419 | ~new_n16037_;
  assign new_n16274_ = ~new_n5101_ | ~new_n16031_;
  assign new_n16275_ = ~pi418 | ~new_n16032_;
  assign new_n16276_ = ~new_n16275_ | ~new_n16274_;
  assign new_n16277_ = ~new_n16204_ | ~new_n16046_;
  assign new_n16278_ = ~new_n16276_ | ~new_n16184_;
  assign new_n16279_ = ~new_n5098_ | ~new_n16033_;
  assign new_n16280_ = ~pi417 | ~new_n16034_;
  assign new_n16281_ = ~new_n16280_ | ~new_n16279_;
  assign new_n16282_ = ~new_n16205_ | ~new_n16067_;
  assign new_n16283_ = ~new_n16141_ | ~new_n16281_;
  assign new_n16284_ = ~new_n5095_ | ~new_n16029_;
  assign new_n16285_ = ~pi416 | ~new_n16030_;
  assign new_n16286_ = ~new_n5062_ | ~new_n16006_;
  assign new_n16287_ = ~pi406 | ~new_n16007_;
  assign new_n16288_ = new_n16417_ & new_n16317_;
  assign new_n16289_ = new_n16415_ & new_n16318_;
  assign new_n16290_ = new_n16414_ & new_n16319_;
  assign new_n16291_ = new_n16413_ & new_n16320_;
  assign new_n16292_ = new_n16411_ & new_n16321_;
  assign new_n16293_ = new_n16410_ & new_n16322_;
  assign new_n16294_ = new_n16409_ & new_n16323_;
  assign new_n16295_ = new_n16407_ & new_n16324_;
  assign new_n16296_ = new_n16405_ & new_n16325_;
  assign new_n16297_ = new_n16403_ & new_n16326_;
  assign new_n16298_ = new_n16401_ & new_n16327_;
  assign new_n16299_ = new_n16399_ & new_n16328_;
  assign new_n16300_ = new_n16397_ & new_n16307_;
  assign new_n16301_ = new_n16395_ & new_n16349_;
  assign new_n16302_ = new_n16380_ & new_n16308_;
  assign new_n16303_ = new_n16379_ & new_n16309_;
  assign new_n16304_ = new_n16378_ & new_n16310_;
  assign new_n16305_ = new_n16376_ & new_n16311_;
  assign new_n16306_ = new_n16375_ & new_n16312_;
  assign new_n16307_ = new_n5064_ | new_n5072_ | new_n5069_;
  assign new_n16308_ = ~new_n16369_ | ~new_n16316_;
  assign new_n16309_ = ~new_n16370_ | ~new_n16315_;
  assign new_n16310_ = ~new_n16338_ | ~new_n16371_;
  assign new_n16311_ = ~new_n16372_ | ~new_n16314_;
  assign new_n16312_ = ~new_n16373_ | ~new_n16313_;
  assign new_n16313_ = ~new_n5090_;
  assign new_n16314_ = ~new_n5087_;
  assign new_n16315_ = ~new_n5078_;
  assign new_n16316_ = ~new_n5075_;
  assign new_n16317_ = ~new_n16339_ | ~new_n16374_;
  assign new_n16318_ = ~new_n16381_ | ~new_n16336_;
  assign new_n16319_ = ~new_n16382_ | ~new_n16335_;
  assign new_n16320_ = ~new_n16340_ | ~new_n16383_;
  assign new_n16321_ = ~new_n16384_ | ~new_n16334_;
  assign new_n16322_ = ~new_n16385_ | ~new_n16333_;
  assign new_n16323_ = ~new_n16341_ | ~new_n16386_;
  assign new_n16324_ = ~new_n16342_ | ~new_n16387_;
  assign new_n16325_ = ~new_n16343_ | ~new_n16388_;
  assign new_n16326_ = ~new_n16332_ | ~new_n16389_ | ~new_n16357_;
  assign new_n16327_ = ~new_n16331_ | ~new_n16390_ | ~new_n16355_;
  assign new_n16328_ = ~new_n16330_ | ~new_n16391_ | ~new_n16353_;
  assign new_n16329_ = ~new_n5594_;
  assign new_n16330_ = ~new_n5584_;
  assign new_n16331_ = ~new_n5586_;
  assign new_n16332_ = ~new_n5588_;
  assign new_n16333_ = ~new_n5114_;
  assign new_n16334_ = ~new_n5111_;
  assign new_n16335_ = ~new_n5102_;
  assign new_n16336_ = ~new_n5099_;
  assign new_n16337_ = ~new_n16435_ | ~new_n16434_;
  assign new_n16338_ = ~new_n5081_ & ~new_n5084_;
  assign new_n16339_ = ~new_n5096_ & ~new_n5093_;
  assign new_n16340_ = ~new_n5105_ & ~new_n5108_;
  assign new_n16341_ = ~new_n5117_ & ~new_n5120_;
  assign new_n16342_ = ~new_n5122_ & ~new_n5592_;
  assign new_n16343_ = ~new_n5591_ & ~new_n5590_;
  assign new_n16344_ = ~new_n5093_;
  assign new_n16345_ = new_n16419_ & new_n16418_;
  assign new_n16346_ = ~new_n5081_;
  assign new_n16347_ = new_n16421_ & new_n16420_;
  assign new_n16348_ = ~new_n5593_;
  assign new_n16349_ = ~new_n16329_ | ~new_n16392_ | ~new_n16351_;
  assign new_n16350_ = new_n16423_ & new_n16422_;
  assign new_n16351_ = ~new_n5595_;
  assign new_n16352_ = new_n16425_ & new_n16424_;
  assign new_n16353_ = ~new_n5585_;
  assign new_n16354_ = new_n16427_ & new_n16426_;
  assign new_n16355_ = ~new_n5587_;
  assign new_n16356_ = new_n16429_ & new_n16428_;
  assign new_n16357_ = ~new_n5589_;
  assign new_n16358_ = new_n16431_ & new_n16430_;
  assign new_n16359_ = ~new_n5591_;
  assign new_n16360_ = new_n16433_ & new_n16432_;
  assign new_n16361_ = ~new_n5069_;
  assign new_n16362_ = ~new_n5064_;
  assign new_n16363_ = ~new_n5122_;
  assign new_n16364_ = new_n16437_ & new_n16436_;
  assign new_n16365_ = ~new_n5117_;
  assign new_n16366_ = new_n16439_ & new_n16438_;
  assign new_n16367_ = ~new_n5105_;
  assign new_n16368_ = new_n16441_ & new_n16440_;
  assign new_n16369_ = ~new_n16307_;
  assign new_n16370_ = ~new_n16308_;
  assign new_n16371_ = ~new_n16309_;
  assign new_n16372_ = ~new_n16310_;
  assign new_n16373_ = ~new_n16311_;
  assign new_n16374_ = ~new_n16312_;
  assign new_n16375_ = ~new_n5090_ | ~new_n16311_;
  assign new_n16376_ = ~new_n5087_ | ~new_n16310_;
  assign new_n16377_ = ~new_n16371_ | ~new_n16346_;
  assign new_n16378_ = ~new_n5084_ | ~new_n16377_;
  assign new_n16379_ = ~new_n5078_ | ~new_n16308_;
  assign new_n16380_ = ~new_n5075_ | ~new_n16307_;
  assign new_n16381_ = ~new_n16317_;
  assign new_n16382_ = ~new_n16318_;
  assign new_n16383_ = ~new_n16319_;
  assign new_n16384_ = ~new_n16320_;
  assign new_n16385_ = ~new_n16321_;
  assign new_n16386_ = ~new_n16322_;
  assign new_n16387_ = ~new_n16323_;
  assign new_n16388_ = ~new_n16324_;
  assign new_n16389_ = ~new_n16325_;
  assign new_n16390_ = ~new_n16326_;
  assign new_n16391_ = ~new_n16327_;
  assign new_n16392_ = ~new_n16328_;
  assign new_n16393_ = ~new_n16349_;
  assign new_n16394_ = ~new_n16392_ | ~new_n16351_;
  assign new_n16395_ = ~new_n5594_ | ~new_n16394_;
  assign new_n16396_ = new_n5069_ | new_n5064_;
  assign new_n16397_ = ~new_n5072_ | ~new_n16396_;
  assign new_n16398_ = ~new_n16391_ | ~new_n16353_;
  assign new_n16399_ = ~new_n5584_ | ~new_n16398_;
  assign new_n16400_ = ~new_n16390_ | ~new_n16355_;
  assign new_n16401_ = ~new_n5586_ | ~new_n16400_;
  assign new_n16402_ = ~new_n16389_ | ~new_n16357_;
  assign new_n16403_ = ~new_n5588_ | ~new_n16402_;
  assign new_n16404_ = ~new_n16388_ | ~new_n16359_;
  assign new_n16405_ = ~new_n5590_ | ~new_n16404_;
  assign new_n16406_ = ~new_n16387_ | ~new_n16363_;
  assign new_n16407_ = ~new_n5592_ | ~new_n16406_;
  assign new_n16408_ = ~new_n16386_ | ~new_n16365_;
  assign new_n16409_ = ~new_n5120_ | ~new_n16408_;
  assign new_n16410_ = ~new_n5114_ | ~new_n16321_;
  assign new_n16411_ = ~new_n5111_ | ~new_n16320_;
  assign new_n16412_ = ~new_n16383_ | ~new_n16367_;
  assign new_n16413_ = ~new_n5108_ | ~new_n16412_;
  assign new_n16414_ = ~new_n5102_ | ~new_n16318_;
  assign new_n16415_ = ~new_n5099_ | ~new_n16317_;
  assign new_n16416_ = ~new_n16374_ | ~new_n16344_;
  assign new_n16417_ = ~new_n5096_ | ~new_n16416_;
  assign new_n16418_ = ~new_n5093_ | ~new_n16312_;
  assign new_n16419_ = ~new_n16374_ | ~new_n16344_;
  assign new_n16420_ = ~new_n5081_ | ~new_n16309_;
  assign new_n16421_ = ~new_n16371_ | ~new_n16346_;
  assign new_n16422_ = ~new_n5593_ | ~new_n16349_;
  assign new_n16423_ = ~new_n16393_ | ~new_n16348_;
  assign new_n16424_ = ~new_n5595_ | ~new_n16328_;
  assign new_n16425_ = ~new_n16392_ | ~new_n16351_;
  assign new_n16426_ = ~new_n5585_ | ~new_n16327_;
  assign new_n16427_ = ~new_n16391_ | ~new_n16353_;
  assign new_n16428_ = ~new_n5587_ | ~new_n16326_;
  assign new_n16429_ = ~new_n16390_ | ~new_n16355_;
  assign new_n16430_ = ~new_n5589_ | ~new_n16325_;
  assign new_n16431_ = ~new_n16389_ | ~new_n16357_;
  assign new_n16432_ = ~new_n5591_ | ~new_n16324_;
  assign new_n16433_ = ~new_n16388_ | ~new_n16359_;
  assign new_n16434_ = ~new_n5069_ | ~new_n16362_;
  assign new_n16435_ = ~new_n5064_ | ~new_n16361_;
  assign new_n16436_ = ~new_n5122_ | ~new_n16323_;
  assign new_n16437_ = ~new_n16387_ | ~new_n16363_;
  assign new_n16438_ = ~new_n5117_ | ~new_n16322_;
  assign new_n16439_ = ~new_n16386_ | ~new_n16365_;
  assign new_n16440_ = ~new_n5105_ | ~new_n16319_;
  assign new_n16441_ = ~new_n16383_ | ~new_n16367_;
  assign new_n16442_ = new_n16551_ & new_n16552_;
  assign new_n16443_ = new_n16554_ & new_n16556_ & new_n16558_ & new_n16557_;
  assign new_n16444_ = new_n16511_ & new_n16443_;
  assign new_n16445_ = new_n16444_ & new_n16562_;
  assign new_n16446_ = new_n16545_ & new_n16547_ & new_n16548_;
  assign new_n16447_ = new_n16542_ & new_n16541_ & new_n16622_ & new_n16621_;
  assign new_n16448_ = ~new_n5595_;
  assign new_n16449_ = ~new_n5208_;
  assign new_n16450_ = ~new_n5215_;
  assign new_n16451_ = ~new_n5216_;
  assign new_n16452_ = ~new_n5590_;
  assign new_n16453_ = ~new_n5222_;
  assign new_n16454_ = ~new_n5221_;
  assign new_n16455_ = ~new_n5114_;
  assign new_n16456_ = ~new_n5111_;
  assign new_n16457_ = ~new_n5108_;
  assign new_n16458_ = ~new_n5227_;
  assign new_n16459_ = ~new_n5096_;
  assign new_n16460_ = ~new_n5093_;
  assign new_n16461_ = ~new_n5087_;
  assign new_n16462_ = ~new_n5090_;
  assign new_n16463_ = ~new_n5084_;
  assign new_n16464_ = ~new_n5081_;
  assign new_n16465_ = ~new_n5078_;
  assign new_n16466_ = ~new_n5075_;
  assign new_n16467_ = ~new_n5220_;
  assign new_n16468_ = ~new_n5072_;
  assign new_n16469_ = ~new_n5069_;
  assign new_n16470_ = ~new_n5228_;
  assign new_n16471_ = ~new_n5209_;
  assign new_n16472_ = ~new_n5206_;
  assign new_n16473_ = ~new_n5205_;
  assign new_n16474_ = ~new_n5204_;
  assign new_n16475_ = ~new_n5203_;
  assign new_n16476_ = ~new_n5202_;
  assign new_n16477_ = ~new_n5201_;
  assign new_n16478_ = ~new_n5200_;
  assign new_n16479_ = ~new_n5230_;
  assign new_n16480_ = ~new_n5229_;
  assign new_n16481_ = ~new_n5102_;
  assign new_n16482_ = ~new_n5099_;
  assign new_n16483_ = ~new_n5105_;
  assign new_n16484_ = ~new_n5226_;
  assign new_n16485_ = ~new_n5225_;
  assign new_n16486_ = ~new_n5224_;
  assign new_n16487_ = ~new_n5223_;
  assign new_n16488_ = ~new_n5591_;
  assign new_n16489_ = ~new_n5120_;
  assign new_n16490_ = ~new_n5117_;
  assign new_n16491_ = ~new_n5122_;
  assign new_n16492_ = ~new_n5592_;
  assign new_n16493_ = ~new_n5219_;
  assign new_n16494_ = ~new_n5218_;
  assign new_n16495_ = ~new_n5217_;
  assign new_n16496_ = ~new_n5589_;
  assign new_n16497_ = ~new_n5588_;
  assign new_n16498_ = ~new_n16615_ | ~new_n16614_;
  assign new_n16499_ = ~new_n5214_;
  assign new_n16500_ = ~new_n5586_;
  assign new_n16501_ = ~new_n5207_;
  assign new_n16502_ = ~new_n5585_;
  assign new_n16503_ = ~new_n5584_;
  assign new_n16504_ = ~new_n5594_;
  assign new_n16505_ = ~new_n5210_;
  assign new_n16506_ = ~new_n5212_;
  assign new_n16507_ = ~new_n5213_;
  assign new_n16508_ = ~new_n5593_;
  assign new_n16509_ = ~new_n5211_;
  assign new_n16510_ = new_n5064_ & new_n16543_;
  assign new_n16511_ = new_n16561_ & new_n16560_ & new_n16559_;
  assign new_n16512_ = new_n16564_ & new_n16565_;
  assign new_n16513_ = new_n16512_ & new_n16563_;
  assign new_n16514_ = new_n5209_ & new_n16468_;
  assign new_n16515_ = new_n5206_ & new_n16466_;
  assign new_n16516_ = new_n16560_ & new_n16559_;
  assign new_n16517_ = new_n16576_ & new_n16577_;
  assign new_n16518_ = new_n16556_ & new_n16554_;
  assign new_n16519_ = new_n16582_ & new_n16520_;
  assign new_n16520_ = new_n16584_ & new_n16583_;
  assign new_n16521_ = new_n16581_ & new_n16519_;
  assign new_n16522_ = new_n5099_ & new_n16480_;
  assign new_n16523_ = new_n16587_ & new_n16524_;
  assign new_n16524_ = new_n16588_ & new_n16586_;
  assign new_n16525_ = new_n16591_ & new_n16568_;
  assign new_n16526_ = new_n16589_ & new_n16553_;
  assign new_n16527_ = new_n16442_ & new_n16528_;
  assign new_n16528_ = new_n16597_ & new_n16598_;
  assign new_n16529_ = new_n5120_ & new_n16453_;
  assign new_n16530_ = new_n5117_ & new_n16487_;
  assign new_n16531_ = new_n16600_ & new_n16602_;
  assign new_n16532_ = new_n16531_ & new_n16605_ & new_n16604_ & new_n16603_;
  assign new_n16533_ = new_n5219_ & new_n16492_;
  assign new_n16534_ = new_n16609_ & new_n16607_ & new_n16608_;
  assign new_n16535_ = new_n16612_ & new_n16601_;
  assign new_n16536_ = new_n16610_ & new_n16549_;
  assign new_n16537_ = new_n16446_ & new_n16620_;
  assign new_n16538_ = new_n5210_ & new_n16448_;
  assign new_n16539_ = new_n16540_ & new_n16545_;
  assign new_n16540_ = new_n5211_ & new_n16503_;
  assign new_n16541_ = new_n16625_ & new_n16624_;
  assign new_n16542_ = new_n16626_ & new_n16627_ & new_n16628_;
  assign new_n16543_ = ~new_n5231_;
  assign new_n16544_ = ~new_n16630_ | ~new_n16629_;
  assign new_n16545_ = ~new_n5207_ | ~new_n16508_;
  assign new_n16546_ = ~new_n5595_ | ~new_n16505_;
  assign new_n16547_ = ~new_n5585_ | ~new_n16506_;
  assign new_n16548_ = ~new_n5584_ | ~new_n16509_;
  assign new_n16549_ = ~new_n5215_ | ~new_n16497_;
  assign new_n16550_ = ~new_n5114_ | ~new_n16486_;
  assign new_n16551_ = ~new_n5221_ | ~new_n16491_;
  assign new_n16552_ = ~new_n5222_ | ~new_n16489_;
  assign new_n16553_ = ~new_n5111_ | ~new_n16485_;
  assign new_n16554_ = ~new_n5096_ | ~new_n16479_;
  assign new_n16555_ = ~new_n5220_ | ~new_n16469_;
  assign new_n16556_ = ~new_n5093_ | ~new_n16478_;
  assign new_n16557_ = ~new_n5087_ | ~new_n16476_;
  assign new_n16558_ = ~new_n5090_ | ~new_n16477_;
  assign new_n16559_ = ~new_n5084_ | ~new_n16475_;
  assign new_n16560_ = ~new_n5081_ | ~new_n16474_;
  assign new_n16561_ = ~new_n5078_ | ~new_n16473_;
  assign new_n16562_ = ~new_n5075_ | ~new_n16472_;
  assign new_n16563_ = ~new_n16510_ | ~new_n16555_;
  assign new_n16564_ = ~new_n5072_ | ~new_n16471_;
  assign new_n16565_ = ~new_n5069_ | ~new_n16467_;
  assign new_n16566_ = ~new_n16513_ | ~new_n16445_;
  assign new_n16567_ = ~new_n5228_ | ~new_n16481_;
  assign new_n16568_ = ~new_n5227_ | ~new_n16483_;
  assign new_n16569_ = ~new_n5201_ | ~new_n16462_;
  assign new_n16570_ = ~new_n5200_ | ~new_n16460_;
  assign new_n16571_ = ~new_n16570_ | ~new_n16569_;
  assign new_n16572_ = ~new_n5205_ | ~new_n16465_;
  assign new_n16573_ = ~new_n5204_ | ~new_n16464_;
  assign new_n16574_ = ~new_n16573_ | ~new_n16572_;
  assign new_n16575_ = ~new_n16516_ | ~new_n16574_;
  assign new_n16576_ = ~new_n5203_ | ~new_n16463_;
  assign new_n16577_ = ~new_n5202_ | ~new_n16461_;
  assign new_n16578_ = ~new_n16517_ | ~new_n16575_;
  assign new_n16579_ = ~new_n16514_ | ~new_n16445_;
  assign new_n16580_ = ~new_n16515_ | ~new_n16444_;
  assign new_n16581_ = ~new_n16443_ | ~new_n16578_;
  assign new_n16582_ = ~new_n16518_ | ~new_n16571_;
  assign new_n16583_ = ~new_n5230_ | ~new_n16459_;
  assign new_n16584_ = ~new_n5229_ | ~new_n16482_;
  assign new_n16585_ = ~new_n16521_ | ~new_n16566_ | ~new_n16567_ | ~new_n16580_ | ~new_n16579_;
  assign new_n16586_ = ~new_n5102_ | ~new_n16470_;
  assign new_n16587_ = ~new_n16522_ | ~new_n16567_;
  assign new_n16588_ = ~new_n5105_ | ~new_n16458_;
  assign new_n16589_ = ~new_n5108_ | ~new_n16484_;
  assign new_n16590_ = ~new_n16585_ | ~new_n16523_;
  assign new_n16591_ = ~new_n5226_ | ~new_n16457_;
  assign new_n16592_ = ~new_n16525_ | ~new_n16590_;
  assign new_n16593_ = ~new_n16526_ | ~new_n16592_;
  assign new_n16594_ = ~new_n5225_ | ~new_n16456_;
  assign new_n16595_ = ~new_n16594_ | ~new_n16593_;
  assign new_n16596_ = ~new_n16595_ | ~new_n16550_;
  assign new_n16597_ = ~new_n5224_ | ~new_n16455_;
  assign new_n16598_ = ~new_n5223_ | ~new_n16490_;
  assign new_n16599_ = ~new_n16596_ | ~new_n16527_;
  assign new_n16600_ = ~new_n5591_ | ~new_n16494_;
  assign new_n16601_ = ~new_n5590_ | ~new_n16495_;
  assign new_n16602_ = ~new_n16529_ | ~new_n16551_;
  assign new_n16603_ = ~new_n16530_ | ~new_n16442_;
  assign new_n16604_ = ~new_n5122_ | ~new_n16454_;
  assign new_n16605_ = ~new_n5592_ | ~new_n16493_;
  assign new_n16606_ = ~new_n16599_ | ~new_n16532_;
  assign new_n16607_ = ~new_n16533_ | ~new_n16600_;
  assign new_n16608_ = ~new_n5218_ | ~new_n16488_;
  assign new_n16609_ = ~new_n5217_ | ~new_n16452_;
  assign new_n16610_ = ~new_n5216_ | ~new_n16496_;
  assign new_n16611_ = ~new_n16606_ | ~new_n16534_;
  assign new_n16612_ = ~new_n5589_ | ~new_n16451_;
  assign new_n16613_ = ~new_n16535_ | ~new_n16611_;
  assign new_n16614_ = ~new_n16536_ | ~new_n16613_;
  assign new_n16615_ = ~new_n5588_ | ~new_n16450_;
  assign new_n16616_ = ~new_n16498_;
  assign new_n16617_ = ~new_n5214_ | ~new_n16616_;
  assign new_n16618_ = ~new_n5587_ | ~new_n16617_;
  assign new_n16619_ = ~new_n16498_ | ~new_n16499_;
  assign new_n16620_ = ~new_n5586_ | ~new_n16507_;
  assign new_n16621_ = ~new_n16537_ | ~new_n16544_ | ~new_n16618_ | ~new_n16619_;
  assign new_n16622_ = ~new_n16504_ | ~new_n16545_ | ~new_n5208_;
  assign new_n16623_ = ~new_n5594_ | ~new_n16449_;
  assign new_n16624_ = ~new_n16623_ | ~new_n16545_ | ~new_n16538_;
  assign new_n16625_ = ~new_n16502_ | ~new_n16544_ | ~new_n5212_ | ~new_n16446_;
  assign new_n16626_ = ~new_n16500_ | ~new_n16544_ | ~new_n5213_ | ~new_n16446_;
  assign new_n16627_ = ~new_n5593_ | ~new_n16501_;
  assign new_n16628_ = ~new_n16544_ | ~new_n16539_;
  assign new_n16629_ = ~new_n5208_ | ~new_n16546_;
  assign new_n16630_ = ~new_n16546_ | ~new_n16504_;
  assign new_n16631_ = new_n16830_ & new_n16829_;
  assign new_n16632_ = new_n16869_ & new_n16868_;
  assign new_n16633_ = new_n16886_ & new_n16885_;
  assign new_n16634_ = new_n16910_ & new_n16909_;
  assign new_n16635_ = new_n17009_ & new_n17008_;
  assign new_n16636_ = ~new_n16965_ | ~new_n16968_;
  assign new_n16637_ = ~new_n16954_ | ~new_n16957_;
  assign new_n16638_ = ~new_n16943_ | ~new_n16946_;
  assign new_n16639_ = ~new_n16935_ | ~new_n16937_;
  assign new_n16640_ = ~new_n16781_ | ~new_n16974_ | ~new_n16802_;
  assign new_n16641_ = ~new_n16863_ | ~new_n16865_;
  assign new_n16642_ = ~new_n16855_ | ~new_n16858_;
  assign new_n16643_ = ~new_n16847_ | ~new_n16849_;
  assign new_n16644_ = ~new_n16791_ | ~new_n16971_;
  assign new_n16645_ = ~new_n5087_;
  assign new_n16646_ = ~new_n5081_;
  assign new_n16647_ = ~new_n5072_;
  assign new_n16648_ = ~new_n5064_;
  assign new_n16649_ = ~new_n4694_;
  assign new_n16650_ = ~new_n5075_;
  assign new_n16651_ = ~new_n4684_;
  assign new_n16652_ = ~new_n4684_ | ~new_n16647_;
  assign new_n16653_ = ~new_n4680_;
  assign new_n16654_ = ~new_n5084_;
  assign new_n16655_ = ~new_n5078_;
  assign new_n16656_ = ~new_n4687_;
  assign new_n16657_ = ~new_n4683_;
  assign new_n16658_ = ~new_n4676_;
  assign new_n16659_ = ~new_n4676_ | ~new_n16655_;
  assign new_n16660_ = ~new_n5090_;
  assign new_n16661_ = ~new_n4686_;
  assign new_n16662_ = ~new_n4686_ | ~new_n16645_;
  assign new_n16663_ = ~new_n4700_;
  assign new_n16664_ = ~new_n5093_;
  assign new_n16665_ = ~new_n4699_;
  assign new_n16666_ = ~new_n16836_ | ~new_n16835_;
  assign new_n16667_ = ~new_n16659_ | ~new_n16851_;
  assign new_n16668_ = ~new_n16972_ | ~new_n16820_ | ~new_n16804_;
  assign new_n16669_ = ~new_n5586_;
  assign new_n16670_ = ~new_n5590_;
  assign new_n16671_ = ~new_n5111_;
  assign new_n16672_ = ~new_n5096_;
  assign new_n16673_ = ~new_n5099_;
  assign new_n16674_ = ~new_n4679_;
  assign new_n16675_ = ~new_n4678_;
  assign new_n16676_ = ~new_n4699_ | ~new_n16664_;
  assign new_n16677_ = ~new_n5102_;
  assign new_n16678_ = ~new_n4688_;
  assign new_n16679_ = ~new_n5105_;
  assign new_n16680_ = ~new_n4696_;
  assign new_n16681_ = ~new_n5114_;
  assign new_n16682_ = ~new_n5108_;
  assign new_n16683_ = ~new_n4689_;
  assign new_n16684_ = ~new_n4690_;
  assign new_n16685_ = ~new_n4695_;
  assign new_n16686_ = ~new_n4695_ | ~new_n16682_;
  assign new_n16687_ = ~new_n5117_;
  assign new_n16688_ = ~new_n4685_;
  assign new_n16689_ = ~new_n4698_;
  assign new_n16690_ = ~new_n5122_;
  assign new_n16691_ = ~new_n4697_;
  assign new_n16692_ = ~new_n5592_;
  assign new_n16693_ = ~new_n4692_;
  assign new_n16694_ = ~new_n5589_;
  assign new_n16695_ = ~new_n5591_;
  assign new_n16696_ = ~new_n4682_;
  assign new_n16697_ = ~new_n4677_;
  assign new_n16698_ = ~new_n4691_;
  assign new_n16699_ = ~new_n4691_ | ~new_n16695_;
  assign new_n16700_ = ~new_n5588_;
  assign new_n16701_ = ~new_n4681_;
  assign new_n16702_ = ~new_n5587_;
  assign new_n16703_ = ~new_n4674_;
  assign new_n16704_ = ~new_n5585_;
  assign new_n16705_ = ~new_n4673_;
  assign new_n16706_ = ~new_n4673_ | ~new_n16669_;
  assign new_n16707_ = ~new_n4669_;
  assign new_n16708_ = ~new_n5584_;
  assign new_n16709_ = ~new_n4670_;
  assign new_n16710_ = ~new_n16924_ | ~new_n16923_;
  assign new_n16711_ = ~new_n16699_ | ~new_n16939_;
  assign new_n16712_ = ~new_n16686_ | ~new_n16950_;
  assign new_n16713_ = ~new_n16676_ | ~new_n16961_;
  assign new_n16714_ = ~new_n4693_;
  assign new_n16715_ = ~new_n17019_ | ~new_n17018_;
  assign new_n16716_ = ~new_n17033_ | ~new_n17032_;
  assign new_n16717_ = ~new_n17038_ | ~new_n17037_;
  assign new_n16718_ = ~new_n17054_ | ~new_n17053_;
  assign new_n16719_ = ~new_n17059_ | ~new_n17058_;
  assign new_n16720_ = ~new_n17064_ | ~new_n17063_;
  assign new_n16721_ = ~new_n17069_ | ~new_n17068_;
  assign new_n16722_ = ~new_n17074_ | ~new_n17073_;
  assign new_n16723_ = ~new_n17090_ | ~new_n17089_;
  assign new_n16724_ = ~new_n17095_ | ~new_n17094_;
  assign new_n16725_ = ~new_n16978_ | ~new_n16977_;
  assign new_n16726_ = ~new_n16987_ | ~new_n16986_;
  assign new_n16727_ = ~new_n16994_ | ~new_n16993_;
  assign new_n16728_ = ~new_n16998_ | ~new_n16997_;
  assign new_n16729_ = ~new_n17007_ | ~new_n17006_;
  assign new_n16730_ = ~new_n17028_ | ~new_n17027_;
  assign new_n16731_ = ~new_n17045_ | ~new_n17044_;
  assign new_n16732_ = ~new_n17049_ | ~new_n17048_;
  assign new_n16733_ = ~new_n17081_ | ~new_n17080_;
  assign new_n16734_ = ~new_n17085_ | ~new_n17084_;
  assign new_n16735_ = ~new_n17102_ | ~new_n17101_;
  assign new_n16736_ = new_n16822_ & new_n16812_;
  assign new_n16737_ = new_n16825_ & new_n16826_;
  assign new_n16738_ = new_n16813_ & new_n16833_ & new_n16828_;
  assign new_n16739_ = new_n16838_ & new_n16814_;
  assign new_n16740_ = new_n16841_ & new_n16842_;
  assign new_n16741_ = new_n16662_ & new_n16980_ & new_n16979_;
  assign new_n16742_ = new_n16983_ & new_n16814_;
  assign new_n16743_ = new_n16857_ & new_n16631_;
  assign new_n16744_ = new_n16990_ & new_n16813_;
  assign new_n16745_ = new_n16652_ & new_n17000_ & new_n16999_;
  assign new_n16746_ = new_n17003_ & new_n16812_;
  assign new_n16747_ = new_n16808_ & new_n16867_ & new_n16844_;
  assign new_n16748_ = new_n16884_ & new_n16889_ & new_n16809_;
  assign new_n16749_ = new_n16908_ & new_n16913_ & new_n16810_;
  assign new_n16750_ = new_n16926_ & new_n16811_;
  assign new_n16751_ = new_n16929_ & new_n16930_;
  assign new_n16752_ = new_n16929_ & new_n16930_;
  assign new_n16753_ = new_n16635_ & new_n16933_;
  assign new_n16754_ = ~new_n17016_ | ~new_n17015_;
  assign new_n16755_ = new_n16706_ & new_n17021_ & new_n17020_;
  assign new_n16756_ = new_n17024_ & new_n16811_;
  assign new_n16757_ = ~new_n17030_ | ~new_n17029_;
  assign new_n16758_ = ~new_n17035_ | ~new_n17034_;
  assign new_n16759_ = new_n16945_ & new_n16634_;
  assign new_n16760_ = new_n17041_ & new_n16810_;
  assign new_n16761_ = ~new_n17051_ | ~new_n17050_;
  assign new_n16762_ = ~new_n17056_ | ~new_n17055_;
  assign new_n16763_ = ~new_n17061_ | ~new_n17060_;
  assign new_n16764_ = ~new_n17066_ | ~new_n17065_;
  assign new_n16765_ = ~new_n17071_ | ~new_n17070_;
  assign new_n16766_ = new_n16956_ & new_n16633_;
  assign new_n16767_ = new_n17077_ & new_n16809_;
  assign new_n16768_ = ~new_n17087_ | ~new_n17086_;
  assign new_n16769_ = ~new_n17092_ | ~new_n17091_;
  assign new_n16770_ = new_n16967_ & new_n16632_;
  assign new_n16771_ = new_n17098_ & new_n16808_;
  assign new_n16772_ = new_n16976_ & new_n16975_;
  assign new_n16773_ = ~new_n16740_ | ~new_n16839_;
  assign new_n16774_ = new_n16985_ & new_n16984_;
  assign new_n16775_ = new_n16992_ & new_n16991_;
  assign new_n16776_ = new_n16996_ & new_n16995_;
  assign new_n16777_ = ~new_n16737_ | ~new_n16823_;
  assign new_n16778_ = new_n17005_ & new_n17004_;
  assign new_n16779_ = ~new_n5595_;
  assign new_n16780_ = ~new_n4671_;
  assign new_n16781_ = new_n17014_ & new_n17013_;
  assign new_n16782_ = ~new_n16751_ | ~new_n16927_;
  assign new_n16783_ = new_n17026_ & new_n17025_;
  assign new_n16784_ = ~new_n16920_ | ~new_n16919_;
  assign new_n16785_ = ~new_n16916_ | ~new_n16915_;
  assign new_n16786_ = new_n17043_ & new_n17042_;
  assign new_n16787_ = new_n17047_ & new_n17046_;
  assign new_n16788_ = ~new_n16906_ | ~new_n16905_;
  assign new_n16789_ = ~new_n16902_ | ~new_n16901_;
  assign new_n16790_ = ~new_n5069_;
  assign new_n16791_ = ~new_n5064_ | ~new_n16714_;
  assign new_n16792_ = ~new_n16973_ | ~new_n16898_ | ~new_n16803_;
  assign new_n16793_ = ~new_n5120_;
  assign new_n16794_ = ~new_n16896_ | ~new_n16895_;
  assign new_n16795_ = ~new_n16892_ | ~new_n16891_;
  assign new_n16796_ = new_n17079_ & new_n17078_;
  assign new_n16797_ = new_n17083_ & new_n17082_;
  assign new_n16798_ = ~new_n16882_ | ~new_n16881_;
  assign new_n16799_ = ~new_n16878_ | ~new_n16877_;
  assign new_n16800_ = ~new_n16874_ | ~new_n16873_;
  assign new_n16801_ = new_n17100_ & new_n17099_;
  assign new_n16802_ = ~new_n17012_ | ~new_n16932_ | ~new_n16782_;
  assign new_n16803_ = ~new_n16794_ | ~new_n16793_;
  assign new_n16804_ = ~new_n16791_ | ~new_n16790_;
  assign new_n16805_ = ~new_n16706_;
  assign new_n16806_ = ~new_n16652_;
  assign new_n16807_ = ~new_n16662_;
  assign new_n16808_ = ~new_n5096_ | ~new_n16675_;
  assign new_n16809_ = ~new_n5111_ | ~new_n16684_;
  assign new_n16810_ = ~new_n5590_ | ~new_n16697_;
  assign new_n16811_ = ~new_n5586_ | ~new_n16705_;
  assign new_n16812_ = ~new_n5072_ | ~new_n16651_;
  assign new_n16813_ = ~new_n5081_ | ~new_n16657_;
  assign new_n16814_ = ~new_n5087_ | ~new_n16661_;
  assign new_n16815_ = ~new_n16686_;
  assign new_n16816_ = ~new_n16699_;
  assign new_n16817_ = ~new_n16659_;
  assign new_n16818_ = ~new_n16676_;
  assign new_n16819_ = ~new_n16791_;
  assign new_n16820_ = ~new_n4694_ | ~new_n16791_;
  assign new_n16821_ = ~new_n16668_;
  assign new_n16822_ = ~new_n5075_ | ~new_n16653_;
  assign new_n16823_ = ~new_n16736_ | ~new_n16668_;
  assign new_n16824_ = ~new_n16653_ | ~new_n16652_;
  assign new_n16825_ = ~new_n16824_ | ~new_n16650_;
  assign new_n16826_ = ~new_n4680_ | ~new_n16806_;
  assign new_n16827_ = ~new_n16777_;
  assign new_n16828_ = ~new_n5084_ | ~new_n16656_;
  assign new_n16829_ = ~new_n4687_ | ~new_n16654_;
  assign new_n16830_ = ~new_n4683_ | ~new_n16646_;
  assign new_n16831_ = ~new_n16817_ | ~new_n16813_;
  assign new_n16832_ = ~new_n16631_ | ~new_n16831_;
  assign new_n16833_ = ~new_n5078_ | ~new_n16658_;
  assign new_n16834_ = ~new_n5084_ | ~new_n16656_;
  assign new_n16835_ = ~new_n16777_ | ~new_n16738_;
  assign new_n16836_ = ~new_n16834_ | ~new_n16832_;
  assign new_n16837_ = ~new_n16666_;
  assign new_n16838_ = ~new_n5090_ | ~new_n16663_;
  assign new_n16839_ = ~new_n16739_ | ~new_n16666_;
  assign new_n16840_ = ~new_n16663_ | ~new_n16662_;
  assign new_n16841_ = ~new_n16840_ | ~new_n16660_;
  assign new_n16842_ = ~new_n4700_ | ~new_n16807_;
  assign new_n16843_ = ~new_n16773_;
  assign new_n16844_ = ~new_n5093_ | ~new_n16665_;
  assign new_n16845_ = ~new_n16844_ | ~new_n16676_;
  assign new_n16846_ = ~new_n16837_ | ~new_n16662_;
  assign new_n16847_ = ~new_n16742_ | ~new_n16846_;
  assign new_n16848_ = ~new_n16666_ | ~new_n16814_;
  assign new_n16849_ = ~new_n16741_ | ~new_n16848_;
  assign new_n16850_ = ~new_n16662_ | ~new_n16814_;
  assign new_n16851_ = ~new_n16833_ | ~new_n16777_;
  assign new_n16852_ = ~new_n16667_;
  assign new_n16853_ = ~new_n4683_ | ~new_n16646_;
  assign new_n16854_ = ~new_n16852_ | ~new_n16853_;
  assign new_n16855_ = ~new_n16744_ | ~new_n16854_;
  assign new_n16856_ = ~new_n16667_ | ~new_n16813_;
  assign new_n16857_ = ~new_n5084_ | ~new_n16656_;
  assign new_n16858_ = ~new_n16743_ | ~new_n16856_;
  assign new_n16859_ = ~new_n4683_ | ~new_n16646_;
  assign new_n16860_ = ~new_n16813_ | ~new_n16859_;
  assign new_n16861_ = ~new_n16833_ | ~new_n16659_;
  assign new_n16862_ = ~new_n16821_ | ~new_n16652_;
  assign new_n16863_ = ~new_n16746_ | ~new_n16862_;
  assign new_n16864_ = ~new_n16668_ | ~new_n16812_;
  assign new_n16865_ = ~new_n16745_ | ~new_n16864_;
  assign new_n16866_ = ~new_n16652_ | ~new_n16812_;
  assign new_n16867_ = ~new_n5099_ | ~new_n16674_;
  assign new_n16868_ = ~new_n4679_ | ~new_n16673_;
  assign new_n16869_ = ~new_n4678_ | ~new_n16672_;
  assign new_n16870_ = ~new_n16818_ | ~new_n16808_;
  assign new_n16871_ = ~new_n16632_ | ~new_n16870_;
  assign new_n16872_ = ~new_n5099_ | ~new_n16674_;
  assign new_n16873_ = ~new_n16773_ | ~new_n16747_;
  assign new_n16874_ = ~new_n16872_ | ~new_n16871_;
  assign new_n16875_ = ~new_n16800_;
  assign new_n16876_ = ~new_n5102_ | ~new_n16678_;
  assign new_n16877_ = ~new_n16876_ | ~new_n16800_;
  assign new_n16878_ = ~new_n4688_ | ~new_n16677_;
  assign new_n16879_ = ~new_n16799_;
  assign new_n16880_ = ~new_n5105_ | ~new_n16680_;
  assign new_n16881_ = ~new_n16880_ | ~new_n16799_;
  assign new_n16882_ = ~new_n4696_ | ~new_n16679_;
  assign new_n16883_ = ~new_n16798_;
  assign new_n16884_ = ~new_n5114_ | ~new_n16683_;
  assign new_n16885_ = ~new_n4689_ | ~new_n16681_;
  assign new_n16886_ = ~new_n4690_ | ~new_n16671_;
  assign new_n16887_ = ~new_n16815_ | ~new_n16809_;
  assign new_n16888_ = ~new_n16633_ | ~new_n16887_;
  assign new_n16889_ = ~new_n5108_ | ~new_n16685_;
  assign new_n16890_ = ~new_n5114_ | ~new_n16683_;
  assign new_n16891_ = ~new_n16798_ | ~new_n16748_;
  assign new_n16892_ = ~new_n16890_ | ~new_n16888_;
  assign new_n16893_ = ~new_n16795_;
  assign new_n16894_ = ~new_n5117_ | ~new_n16688_;
  assign new_n16895_ = ~new_n16894_ | ~new_n16795_;
  assign new_n16896_ = ~new_n4685_ | ~new_n16687_;
  assign new_n16897_ = ~new_n16794_;
  assign new_n16898_ = ~new_n4698_ | ~new_n16794_;
  assign new_n16899_ = ~new_n16792_;
  assign new_n16900_ = ~new_n5122_ | ~new_n16691_;
  assign new_n16901_ = ~new_n16900_ | ~new_n16792_;
  assign new_n16902_ = ~new_n4697_ | ~new_n16690_;
  assign new_n16903_ = ~new_n16789_;
  assign new_n16904_ = ~new_n5592_ | ~new_n16693_;
  assign new_n16905_ = ~new_n16904_ | ~new_n16789_;
  assign new_n16906_ = ~new_n4692_ | ~new_n16692_;
  assign new_n16907_ = ~new_n16788_;
  assign new_n16908_ = ~new_n5589_ | ~new_n16696_;
  assign new_n16909_ = ~new_n4682_ | ~new_n16694_;
  assign new_n16910_ = ~new_n4677_ | ~new_n16670_;
  assign new_n16911_ = ~new_n16816_ | ~new_n16810_;
  assign new_n16912_ = ~new_n16634_ | ~new_n16911_;
  assign new_n16913_ = ~new_n5591_ | ~new_n16698_;
  assign new_n16914_ = ~new_n5589_ | ~new_n16696_;
  assign new_n16915_ = ~new_n16788_ | ~new_n16749_;
  assign new_n16916_ = ~new_n16914_ | ~new_n16912_;
  assign new_n16917_ = ~new_n16785_;
  assign new_n16918_ = ~new_n5588_ | ~new_n16701_;
  assign new_n16919_ = ~new_n16918_ | ~new_n16785_;
  assign new_n16920_ = ~new_n4681_ | ~new_n16700_;
  assign new_n16921_ = ~new_n16784_;
  assign new_n16922_ = ~new_n5587_ | ~new_n16703_;
  assign new_n16923_ = ~new_n16922_ | ~new_n16784_;
  assign new_n16924_ = ~new_n4674_ | ~new_n16702_;
  assign new_n16925_ = ~new_n16710_;
  assign new_n16926_ = ~new_n5585_ | ~new_n16707_;
  assign new_n16927_ = ~new_n16750_ | ~new_n16710_;
  assign new_n16928_ = ~new_n16707_ | ~new_n16706_;
  assign new_n16929_ = ~new_n16928_ | ~new_n16704_;
  assign new_n16930_ = ~new_n4669_ | ~new_n16805_;
  assign new_n16931_ = ~new_n16782_;
  assign new_n16932_ = ~new_n5584_ | ~new_n16709_;
  assign new_n16933_ = ~new_n4670_ | ~new_n16708_;
  assign new_n16934_ = ~new_n16925_ | ~new_n16706_;
  assign new_n16935_ = ~new_n16756_ | ~new_n16934_;
  assign new_n16936_ = ~new_n16710_ | ~new_n16811_;
  assign new_n16937_ = ~new_n16755_ | ~new_n16936_;
  assign new_n16938_ = ~new_n16706_ | ~new_n16811_;
  assign new_n16939_ = ~new_n16913_ | ~new_n16788_;
  assign new_n16940_ = ~new_n16711_;
  assign new_n16941_ = ~new_n4677_ | ~new_n16670_;
  assign new_n16942_ = ~new_n16940_ | ~new_n16941_;
  assign new_n16943_ = ~new_n16760_ | ~new_n16942_;
  assign new_n16944_ = ~new_n16711_ | ~new_n16810_;
  assign new_n16945_ = ~new_n5589_ | ~new_n16696_;
  assign new_n16946_ = ~new_n16759_ | ~new_n16944_;
  assign new_n16947_ = ~new_n4677_ | ~new_n16670_;
  assign new_n16948_ = ~new_n16810_ | ~new_n16947_;
  assign new_n16949_ = ~new_n16913_ | ~new_n16699_;
  assign new_n16950_ = ~new_n16889_ | ~new_n16798_;
  assign new_n16951_ = ~new_n16712_;
  assign new_n16952_ = ~new_n4690_ | ~new_n16671_;
  assign new_n16953_ = ~new_n16951_ | ~new_n16952_;
  assign new_n16954_ = ~new_n16767_ | ~new_n16953_;
  assign new_n16955_ = ~new_n16712_ | ~new_n16809_;
  assign new_n16956_ = ~new_n5114_ | ~new_n16683_;
  assign new_n16957_ = ~new_n16766_ | ~new_n16955_;
  assign new_n16958_ = ~new_n4690_ | ~new_n16671_;
  assign new_n16959_ = ~new_n16809_ | ~new_n16958_;
  assign new_n16960_ = ~new_n16889_ | ~new_n16686_;
  assign new_n16961_ = ~new_n16844_ | ~new_n16773_;
  assign new_n16962_ = ~new_n16713_;
  assign new_n16963_ = ~new_n4678_ | ~new_n16672_;
  assign new_n16964_ = ~new_n16962_ | ~new_n16963_;
  assign new_n16965_ = ~new_n16771_ | ~new_n16964_;
  assign new_n16966_ = ~new_n16713_ | ~new_n16808_;
  assign new_n16967_ = ~new_n5099_ | ~new_n16674_;
  assign new_n16968_ = ~new_n16770_ | ~new_n16966_;
  assign new_n16969_ = ~new_n4678_ | ~new_n16672_;
  assign new_n16970_ = ~new_n16808_ | ~new_n16969_;
  assign new_n16971_ = ~new_n4693_ | ~new_n16648_;
  assign new_n16972_ = ~new_n4694_ | ~new_n16790_;
  assign new_n16973_ = ~new_n4698_ | ~new_n16793_;
  assign new_n16974_ = ~new_n16753_ | ~new_n16752_ | ~new_n16927_;
  assign new_n16975_ = ~new_n5093_ | ~new_n16665_;
  assign new_n16976_ = ~new_n4699_ | ~new_n16664_;
  assign new_n16977_ = ~new_n16845_ | ~new_n16773_;
  assign new_n16978_ = ~new_n16843_ | ~new_n16772_;
  assign new_n16979_ = ~new_n5090_ | ~new_n16663_;
  assign new_n16980_ = ~new_n4700_ | ~new_n16660_;
  assign new_n16981_ = ~new_n5090_ | ~new_n16663_;
  assign new_n16982_ = ~new_n4700_ | ~new_n16660_;
  assign new_n16983_ = ~new_n16982_ | ~new_n16981_;
  assign new_n16984_ = ~new_n5087_ | ~new_n16661_;
  assign new_n16985_ = ~new_n4686_ | ~new_n16645_;
  assign new_n16986_ = ~new_n16850_ | ~new_n16666_;
  assign new_n16987_ = ~new_n16774_ | ~new_n16837_;
  assign new_n16988_ = ~new_n5084_ | ~new_n16656_;
  assign new_n16989_ = ~new_n4687_ | ~new_n16654_;
  assign new_n16990_ = ~new_n16989_ | ~new_n16988_;
  assign new_n16991_ = ~new_n5081_ | ~new_n16657_;
  assign new_n16992_ = ~new_n4683_ | ~new_n16646_;
  assign new_n16993_ = ~new_n16860_ | ~new_n16667_;
  assign new_n16994_ = ~new_n16775_ | ~new_n16852_;
  assign new_n16995_ = ~new_n5078_ | ~new_n16658_;
  assign new_n16996_ = ~new_n4676_ | ~new_n16655_;
  assign new_n16997_ = ~new_n16861_ | ~new_n16777_;
  assign new_n16998_ = ~new_n16827_ | ~new_n16776_;
  assign new_n16999_ = ~new_n5075_ | ~new_n16653_;
  assign new_n17000_ = ~new_n4680_ | ~new_n16650_;
  assign new_n17001_ = ~new_n5075_ | ~new_n16653_;
  assign new_n17002_ = ~new_n4680_ | ~new_n16650_;
  assign new_n17003_ = ~new_n17002_ | ~new_n17001_;
  assign new_n17004_ = ~new_n5072_ | ~new_n16651_;
  assign new_n17005_ = ~new_n4684_ | ~new_n16647_;
  assign new_n17006_ = ~new_n16866_ | ~new_n16668_;
  assign new_n17007_ = ~new_n16778_ | ~new_n16821_;
  assign new_n17008_ = ~new_n5595_ | ~new_n16780_;
  assign new_n17009_ = ~new_n4671_ | ~new_n16779_;
  assign new_n17010_ = ~new_n5595_ | ~new_n16780_;
  assign new_n17011_ = ~new_n4671_ | ~new_n16779_;
  assign new_n17012_ = ~new_n17011_ | ~new_n17010_;
  assign new_n17013_ = ~new_n16709_ | ~new_n5584_ | ~new_n16635_;
  assign new_n17014_ = ~new_n4670_ | ~new_n17012_ | ~new_n16708_;
  assign new_n17015_ = ~new_n5584_ | ~new_n16709_;
  assign new_n17016_ = ~new_n4670_ | ~new_n16708_;
  assign new_n17017_ = ~new_n16754_;
  assign new_n17018_ = ~new_n16931_ | ~new_n17017_;
  assign new_n17019_ = ~new_n16754_ | ~new_n16782_;
  assign new_n17020_ = ~new_n5585_ | ~new_n16707_;
  assign new_n17021_ = ~new_n4669_ | ~new_n16704_;
  assign new_n17022_ = ~new_n5585_ | ~new_n16707_;
  assign new_n17023_ = ~new_n4669_ | ~new_n16704_;
  assign new_n17024_ = ~new_n17023_ | ~new_n17022_;
  assign new_n17025_ = ~new_n5586_ | ~new_n16705_;
  assign new_n17026_ = ~new_n4673_ | ~new_n16669_;
  assign new_n17027_ = ~new_n16938_ | ~new_n16710_;
  assign new_n17028_ = ~new_n16783_ | ~new_n16925_;
  assign new_n17029_ = ~new_n5587_ | ~new_n16703_;
  assign new_n17030_ = ~new_n4674_ | ~new_n16702_;
  assign new_n17031_ = ~new_n16757_;
  assign new_n17032_ = ~new_n16921_ | ~new_n17031_;
  assign new_n17033_ = ~new_n16757_ | ~new_n16784_;
  assign new_n17034_ = ~new_n5588_ | ~new_n16701_;
  assign new_n17035_ = ~new_n4681_ | ~new_n16700_;
  assign new_n17036_ = ~new_n16758_;
  assign new_n17037_ = ~new_n16917_ | ~new_n17036_;
  assign new_n17038_ = ~new_n16758_ | ~new_n16785_;
  assign new_n17039_ = ~new_n5589_ | ~new_n16696_;
  assign new_n17040_ = ~new_n4682_ | ~new_n16694_;
  assign new_n17041_ = ~new_n17040_ | ~new_n17039_;
  assign new_n17042_ = ~new_n5590_ | ~new_n16697_;
  assign new_n17043_ = ~new_n4677_ | ~new_n16670_;
  assign new_n17044_ = ~new_n16948_ | ~new_n16711_;
  assign new_n17045_ = ~new_n16786_ | ~new_n16940_;
  assign new_n17046_ = ~new_n5591_ | ~new_n16698_;
  assign new_n17047_ = ~new_n4691_ | ~new_n16695_;
  assign new_n17048_ = ~new_n16949_ | ~new_n16788_;
  assign new_n17049_ = ~new_n16907_ | ~new_n16787_;
  assign new_n17050_ = ~new_n5592_ | ~new_n16693_;
  assign new_n17051_ = ~new_n4692_ | ~new_n16692_;
  assign new_n17052_ = ~new_n16761_;
  assign new_n17053_ = ~new_n16903_ | ~new_n17052_;
  assign new_n17054_ = ~new_n16761_ | ~new_n16789_;
  assign new_n17055_ = ~new_n5069_ | ~new_n16649_;
  assign new_n17056_ = ~new_n4694_ | ~new_n16790_;
  assign new_n17057_ = ~new_n16762_;
  assign new_n17058_ = ~new_n16819_ | ~new_n17057_;
  assign new_n17059_ = ~new_n16762_ | ~new_n16791_;
  assign new_n17060_ = ~new_n5122_ | ~new_n16691_;
  assign new_n17061_ = ~new_n4697_ | ~new_n16690_;
  assign new_n17062_ = ~new_n16763_;
  assign new_n17063_ = ~new_n16899_ | ~new_n17062_;
  assign new_n17064_ = ~new_n16763_ | ~new_n16792_;
  assign new_n17065_ = ~new_n5120_ | ~new_n16689_;
  assign new_n17066_ = ~new_n4698_ | ~new_n16793_;
  assign new_n17067_ = ~new_n16764_;
  assign new_n17068_ = ~new_n16897_ | ~new_n17067_;
  assign new_n17069_ = ~new_n16764_ | ~new_n16794_;
  assign new_n17070_ = ~new_n5117_ | ~new_n16688_;
  assign new_n17071_ = ~new_n4685_ | ~new_n16687_;
  assign new_n17072_ = ~new_n16765_;
  assign new_n17073_ = ~new_n16893_ | ~new_n17072_;
  assign new_n17074_ = ~new_n16765_ | ~new_n16795_;
  assign new_n17075_ = ~new_n5114_ | ~new_n16683_;
  assign new_n17076_ = ~new_n4689_ | ~new_n16681_;
  assign new_n17077_ = ~new_n17076_ | ~new_n17075_;
  assign new_n17078_ = ~new_n5111_ | ~new_n16684_;
  assign new_n17079_ = ~new_n4690_ | ~new_n16671_;
  assign new_n17080_ = ~new_n16959_ | ~new_n16712_;
  assign new_n17081_ = ~new_n16796_ | ~new_n16951_;
  assign new_n17082_ = ~new_n5108_ | ~new_n16685_;
  assign new_n17083_ = ~new_n4695_ | ~new_n16682_;
  assign new_n17084_ = ~new_n16960_ | ~new_n16798_;
  assign new_n17085_ = ~new_n16883_ | ~new_n16797_;
  assign new_n17086_ = ~new_n5105_ | ~new_n16680_;
  assign new_n17087_ = ~new_n4696_ | ~new_n16679_;
  assign new_n17088_ = ~new_n16768_;
  assign new_n17089_ = ~new_n16879_ | ~new_n17088_;
  assign new_n17090_ = ~new_n16768_ | ~new_n16799_;
  assign new_n17091_ = ~new_n5102_ | ~new_n16678_;
  assign new_n17092_ = ~new_n4688_ | ~new_n16677_;
  assign new_n17093_ = ~new_n16769_;
  assign new_n17094_ = ~new_n16875_ | ~new_n17093_;
  assign new_n17095_ = ~new_n16769_ | ~new_n16800_;
  assign new_n17096_ = ~new_n5099_ | ~new_n16674_;
  assign new_n17097_ = ~new_n4679_ | ~new_n16673_;
  assign new_n17098_ = ~new_n17097_ | ~new_n17096_;
  assign new_n17099_ = ~new_n5096_ | ~new_n16675_;
  assign new_n17100_ = ~new_n4678_ | ~new_n16672_;
  assign new_n17101_ = ~new_n16970_ | ~new_n16713_;
  assign new_n17102_ = ~new_n16801_ | ~new_n16962_;
  assign new_n17103_ = new_n17278_ & new_n17277_;
  assign new_n17104_ = new_n17296_ & new_n17295_;
  assign new_n17105_ = new_n17336_ & new_n17335_;
  assign new_n17106_ = new_n17345_ & new_n17344_;
  assign new_n17107_ = new_n17363_ & new_n17362_;
  assign new_n17108_ = new_n17371_ & new_n17370_;
  assign new_n17109_ = new_n17450_ & new_n17447_;
  assign new_n17110_ = new_n17443_ & new_n17440_;
  assign new_n17111_ = new_n17434_ & new_n17431_;
  assign new_n17112_ = new_n17425_ & new_n17422_;
  assign new_n17113_ = new_n17419_ & new_n17417_;
  assign new_n17114_ = new_n17412_ & new_n17409_;
  assign new_n17115_ = new_n17334_ & new_n17331_;
  assign new_n17116_ = new_n17326_ & new_n17323_;
  assign new_n17117_ = new_n17312_ & new_n17309_;
  assign new_n17118_ = ~new_n5084_;
  assign new_n17119_ = ~new_n4687_;
  assign new_n17120_ = ~new_n4686_;
  assign new_n17121_ = ~new_n4687_ | ~new_n5084_;
  assign new_n17122_ = ~new_n5087_;
  assign new_n17123_ = ~new_n5078_;
  assign new_n17124_ = ~new_n4676_;
  assign new_n17125_ = ~new_n4683_;
  assign new_n17126_ = ~new_n5072_;
  assign new_n17127_ = ~new_n4684_;
  assign new_n17128_ = ~new_n5064_;
  assign new_n17129_ = ~new_n4693_;
  assign new_n17130_ = ~new_n4693_ | ~new_n5064_;
  assign new_n17131_ = ~new_n5075_;
  assign new_n17132_ = ~new_n4680_;
  assign new_n17133_ = ~new_n4676_ | ~new_n5078_;
  assign new_n17134_ = ~new_n5081_;
  assign new_n17135_ = ~new_n5090_;
  assign new_n17136_ = ~new_n4700_;
  assign new_n17137_ = ~new_n4699_;
  assign new_n17138_ = ~new_n5093_;
  assign new_n17139_ = ~new_n17160_ | ~new_n17304_;
  assign new_n17140_ = ~new_n17216_ | ~new_n17292_;
  assign new_n17141_ = ~new_n17281_ | ~new_n17282_;
  assign new_n17142_ = ~new_n5069_ | ~new_n4694_;
  assign new_n17143_ = ~new_n17221_ | ~new_n17318_;
  assign new_n17144_ = ~new_n17315_ | ~new_n17314_;
  assign new_n17145_ = ~new_n5585_;
  assign new_n17146_ = ~new_n4669_;
  assign new_n17147_ = ~new_n4673_;
  assign new_n17148_ = ~new_n5586_;
  assign new_n17149_ = ~new_n5587_;
  assign new_n17150_ = ~new_n4674_;
  assign new_n17151_ = ~new_n5588_;
  assign new_n17152_ = ~new_n4681_;
  assign new_n17153_ = ~new_n5591_;
  assign new_n17154_ = ~new_n4691_;
  assign new_n17155_ = ~new_n5114_;
  assign new_n17156_ = ~new_n4689_;
  assign new_n17157_ = ~new_n4685_;
  assign new_n17158_ = ~new_n4689_ | ~new_n5114_;
  assign new_n17159_ = ~new_n5117_;
  assign new_n17160_ = ~new_n4700_ | ~new_n5090_;
  assign new_n17161_ = ~new_n5096_;
  assign new_n17162_ = ~new_n4678_;
  assign new_n17163_ = ~new_n5102_;
  assign new_n17164_ = ~new_n4688_;
  assign new_n17165_ = ~new_n5099_;
  assign new_n17166_ = ~new_n4679_;
  assign new_n17167_ = ~new_n4679_ | ~new_n5099_;
  assign new_n17168_ = ~new_n5105_;
  assign new_n17169_ = ~new_n4696_;
  assign new_n17170_ = ~new_n5108_;
  assign new_n17171_ = ~new_n4695_;
  assign new_n17172_ = ~new_n5111_;
  assign new_n17173_ = ~new_n4690_;
  assign new_n17174_ = ~new_n5120_;
  assign new_n17175_ = ~new_n4698_;
  assign new_n17176_ = ~new_n4698_ | ~new_n5120_;
  assign new_n17177_ = ~new_n5122_;
  assign new_n17178_ = ~new_n4697_;
  assign new_n17179_ = ~new_n4697_ | ~new_n5122_;
  assign new_n17180_ = ~new_n5592_;
  assign new_n17181_ = ~new_n5590_;
  assign new_n17182_ = ~new_n4677_;
  assign new_n17183_ = ~new_n5589_;
  assign new_n17184_ = ~new_n4682_;
  assign new_n17185_ = ~new_n5586_ | ~new_n4673_;
  assign new_n17186_ = ~new_n4670_;
  assign new_n17187_ = ~new_n5584_;
  assign new_n17188_ = ~new_n17405_ | ~new_n17275_;
  assign new_n17189_ = ~new_n4692_;
  assign new_n17190_ = ~new_n17176_ | ~new_n17414_;
  assign new_n17191_ = ~new_n17360_ | ~new_n17359_;
  assign new_n17192_ = ~new_n17167_ | ~new_n17436_;
  assign new_n17193_ = ~new_n17556_ | ~new_n17555_;
  assign new_n17194_ = ~new_n17603_ | ~new_n17602_;
  assign new_n17195_ = ~new_n17474_ | ~new_n17473_;
  assign new_n17196_ = ~new_n17479_ | ~new_n17478_;
  assign new_n17197_ = ~new_n17486_ | ~new_n17485_;
  assign new_n17198_ = ~new_n17493_ | ~new_n17492_;
  assign new_n17199_ = ~new_n17498_ | ~new_n17497_;
  assign new_n17200_ = ~new_n17507_ | ~new_n17506_;
  assign new_n17201_ = ~new_n17514_ | ~new_n17513_;
  assign new_n17202_ = ~new_n17521_ | ~new_n17520_;
  assign new_n17203_ = ~new_n17528_ | ~new_n17527_;
  assign new_n17204_ = ~new_n17533_ | ~new_n17532_;
  assign new_n17205_ = ~new_n17540_ | ~new_n17539_;
  assign new_n17206_ = ~new_n17547_ | ~new_n17546_;
  assign new_n17207_ = ~new_n17561_ | ~new_n17560_;
  assign new_n17208_ = ~new_n17566_ | ~new_n17565_;
  assign new_n17209_ = ~new_n17573_ | ~new_n17572_;
  assign new_n17210_ = ~new_n17580_ | ~new_n17579_;
  assign new_n17211_ = ~new_n17587_ | ~new_n17586_;
  assign new_n17212_ = ~new_n17594_ | ~new_n17593_;
  assign new_n17213_ = ~new_n17599_ | ~new_n17598_;
  assign new_n17214_ = new_n17288_ & new_n17286_;
  assign new_n17215_ = new_n17103_ & new_n17279_;
  assign new_n17216_ = new_n17293_ & new_n17291_;
  assign new_n17217_ = new_n17300_ & new_n17299_;
  assign new_n17218_ = new_n17121_ & new_n17481_ & new_n17480_;
  assign new_n17219_ = new_n17311_ & new_n17104_;
  assign new_n17220_ = new_n17280_ & new_n17279_;
  assign new_n17221_ = new_n17319_ & new_n17317_;
  assign new_n17222_ = new_n17133_ & new_n17488_ & new_n17487_;
  assign new_n17223_ = new_n17325_ & new_n17103_;
  assign new_n17224_ = new_n17333_ & new_n17280_;
  assign new_n17225_ = new_n17303_ & new_n17105_;
  assign new_n17226_ = new_n17338_ & new_n17270_;
  assign new_n17227_ = new_n17349_ & new_n17106_;
  assign new_n17228_ = new_n17347_ & new_n17271_;
  assign new_n17229_ = new_n17367_ & new_n17366_;
  assign new_n17230_ = new_n17372_ & new_n17108_ & new_n17381_;
  assign new_n17231_ = new_n17384_ & new_n17379_;
  assign new_n17232_ = new_n17400_ & new_n17397_;
  assign new_n17233_ = new_n17467_ & new_n17401_;
  assign new_n17234_ = new_n17272_ & new_n17523_ & new_n17522_;
  assign new_n17235_ = new_n17259_ & new_n17377_;
  assign new_n17236_ = new_n17179_ & new_n17554_ & new_n17553_;
  assign new_n17237_ = new_n17424_ & new_n17108_;
  assign new_n17238_ = new_n17158_ & new_n17568_ & new_n17567_;
  assign new_n17239_ = new_n17433_ & new_n17107_;
  assign new_n17240_ = new_n17271_ & new_n17589_ & new_n17588_;
  assign new_n17241_ = new_n17442_ & new_n17106_;
  assign new_n17242_ = new_n17270_ & new_n17601_ & new_n17600_;
  assign new_n17243_ = new_n17449_ & new_n17105_;
  assign new_n17244_ = ~new_n17217_ | ~new_n17301_;
  assign new_n17245_ = ~new_n17316_ | ~new_n17328_;
  assign new_n17246_ = ~new_n4671_;
  assign new_n17247_ = ~new_n5595_;
  assign new_n17248_ = new_n17502_ & new_n17501_;
  assign new_n17249_ = ~new_n17463_ | ~new_n17403_ | ~new_n17268_;
  assign new_n17250_ = new_n17509_ & new_n17508_;
  assign new_n17251_ = ~new_n17233_ | ~new_n17469_ | ~new_n17468_;
  assign new_n17252_ = new_n17516_ & new_n17515_;
  assign new_n17253_ = ~new_n17185_ | ~new_n17464_ | ~new_n17398_;
  assign new_n17254_ = ~new_n17392_ | ~new_n17391_;
  assign new_n17255_ = new_n17535_ & new_n17534_;
  assign new_n17256_ = ~new_n17388_ | ~new_n17387_;
  assign new_n17257_ = new_n17542_ & new_n17541_;
  assign new_n17258_ = ~new_n17231_ | ~new_n17383_;
  assign new_n17259_ = new_n17549_ & new_n17548_;
  assign new_n17260_ = ~new_n17142_ | ~new_n17426_;
  assign new_n17261_ = ~new_n17229_ | ~new_n17368_;
  assign new_n17262_ = new_n17575_ & new_n17574_;
  assign new_n17263_ = ~new_n17356_ | ~new_n17355_;
  assign new_n17264_ = new_n17582_ & new_n17581_;
  assign new_n17265_ = ~new_n17352_ | ~new_n17351_;
  assign new_n17266_ = ~new_n17342_ | ~new_n17341_;
  assign new_n17267_ = ~new_n17466_ | ~new_n17465_;
  assign new_n17268_ = ~new_n4670_ | ~new_n17251_;
  assign new_n17269_ = ~new_n17133_;
  assign new_n17270_ = ~new_n5093_ | ~new_n4699_;
  assign new_n17271_ = ~new_n4688_ | ~new_n5102_;
  assign new_n17272_ = ~new_n4674_ | ~new_n5587_;
  assign new_n17273_ = ~new_n17167_;
  assign new_n17274_ = ~new_n17176_;
  assign new_n17275_ = ~new_n4681_ | ~new_n5588_;
  assign new_n17276_ = ~new_n17160_;
  assign new_n17277_ = new_n4683_ | new_n5081_;
  assign new_n17278_ = new_n4676_ | new_n5078_;
  assign new_n17279_ = new_n5075_ | new_n4680_;
  assign new_n17280_ = new_n5072_ | new_n4684_;
  assign new_n17281_ = ~new_n17130_;
  assign new_n17282_ = new_n5069_ | new_n4694_;
  assign new_n17283_ = ~new_n17141_;
  assign new_n17284_ = ~new_n17142_;
  assign new_n17285_ = ~new_n17141_ | ~new_n17142_;
  assign new_n17286_ = ~new_n4684_ | ~new_n5072_;
  assign new_n17287_ = ~new_n17285_ | ~new_n17280_;
  assign new_n17288_ = ~new_n4680_ | ~new_n5075_;
  assign new_n17289_ = ~new_n17214_ | ~new_n17287_;
  assign new_n17290_ = ~new_n17134_ | ~new_n17133_;
  assign new_n17291_ = ~new_n4683_ | ~new_n17290_;
  assign new_n17292_ = ~new_n17215_ | ~new_n17289_;
  assign new_n17293_ = ~new_n5081_ | ~new_n17269_;
  assign new_n17294_ = ~new_n17140_;
  assign new_n17295_ = new_n4686_ | new_n5087_;
  assign new_n17296_ = new_n4687_ | new_n5084_;
  assign new_n17297_ = ~new_n17121_;
  assign new_n17298_ = ~new_n17122_ | ~new_n17121_;
  assign new_n17299_ = ~new_n4686_ | ~new_n17298_;
  assign new_n17300_ = ~new_n5087_ | ~new_n17297_;
  assign new_n17301_ = ~new_n17104_ | ~new_n17140_;
  assign new_n17302_ = ~new_n17244_;
  assign new_n17303_ = new_n5090_ | new_n4700_;
  assign new_n17304_ = ~new_n17303_ | ~new_n17244_;
  assign new_n17305_ = ~new_n17139_;
  assign new_n17306_ = new_n4699_ | new_n5093_;
  assign new_n17307_ = new_n5084_ | new_n4687_;
  assign new_n17308_ = ~new_n17307_ | ~new_n17140_;
  assign new_n17309_ = ~new_n17218_ | ~new_n17308_;
  assign new_n17310_ = ~new_n17294_ | ~new_n17121_;
  assign new_n17311_ = ~new_n5087_ | ~new_n4686_;
  assign new_n17312_ = ~new_n17219_ | ~new_n17310_;
  assign new_n17313_ = new_n4687_ | new_n5084_;
  assign new_n17314_ = ~new_n17284_ | ~new_n17280_;
  assign new_n17315_ = ~new_n4684_ | ~new_n5072_;
  assign new_n17316_ = ~new_n17144_;
  assign new_n17317_ = ~new_n17220_ | ~new_n17283_;
  assign new_n17318_ = ~new_n17144_ | ~new_n17279_;
  assign new_n17319_ = ~new_n4680_ | ~new_n5075_;
  assign new_n17320_ = ~new_n17143_;
  assign new_n17321_ = new_n5078_ | new_n4676_;
  assign new_n17322_ = ~new_n17321_ | ~new_n17143_;
  assign new_n17323_ = ~new_n17222_ | ~new_n17322_;
  assign new_n17324_ = ~new_n17320_ | ~new_n17133_;
  assign new_n17325_ = ~new_n5081_ | ~new_n4683_;
  assign new_n17326_ = ~new_n17223_ | ~new_n17324_;
  assign new_n17327_ = new_n4676_ | new_n5078_;
  assign new_n17328_ = ~new_n17283_ | ~new_n17280_;
  assign new_n17329_ = ~new_n17245_;
  assign new_n17330_ = ~new_n4680_ | ~new_n5075_;
  assign new_n17331_ = ~new_n17141_ | ~new_n17142_ | ~new_n17500_ | ~new_n17499_;
  assign new_n17332_ = ~new_n17142_ | ~new_n17141_;
  assign new_n17333_ = ~new_n4684_ | ~new_n5072_;
  assign new_n17334_ = ~new_n17224_ | ~new_n17332_;
  assign new_n17335_ = new_n4699_ | new_n5093_;
  assign new_n17336_ = new_n4678_ | new_n5096_;
  assign new_n17337_ = ~new_n17276_ | ~new_n17105_;
  assign new_n17338_ = ~new_n4678_ | ~new_n5096_;
  assign new_n17339_ = ~new_n17226_ | ~new_n17337_;
  assign new_n17340_ = new_n5096_ | new_n4678_;
  assign new_n17341_ = ~new_n17225_ | ~new_n17244_;
  assign new_n17342_ = ~new_n17340_ | ~new_n17339_;
  assign new_n17343_ = ~new_n17266_;
  assign new_n17344_ = new_n4696_ | new_n5105_;
  assign new_n17345_ = new_n4688_ | new_n5102_;
  assign new_n17346_ = ~new_n17273_ | ~new_n17106_;
  assign new_n17347_ = ~new_n4696_ | ~new_n5105_;
  assign new_n17348_ = ~new_n17228_ | ~new_n17346_;
  assign new_n17349_ = new_n5099_ | new_n4679_;
  assign new_n17350_ = new_n5105_ | new_n4696_;
  assign new_n17351_ = ~new_n17227_ | ~new_n17266_;
  assign new_n17352_ = ~new_n17350_ | ~new_n17348_;
  assign new_n17353_ = ~new_n17265_;
  assign new_n17354_ = new_n5108_ | new_n4695_;
  assign new_n17355_ = ~new_n17354_ | ~new_n17265_;
  assign new_n17356_ = ~new_n4695_ | ~new_n5108_;
  assign new_n17357_ = ~new_n17263_;
  assign new_n17358_ = new_n5111_ | new_n4690_;
  assign new_n17359_ = ~new_n17358_ | ~new_n17263_;
  assign new_n17360_ = ~new_n4690_ | ~new_n5111_;
  assign new_n17361_ = ~new_n17191_;
  assign new_n17362_ = new_n4685_ | new_n5117_;
  assign new_n17363_ = new_n4689_ | new_n5114_;
  assign new_n17364_ = ~new_n17158_;
  assign new_n17365_ = ~new_n17159_ | ~new_n17158_;
  assign new_n17366_ = ~new_n4685_ | ~new_n17365_;
  assign new_n17367_ = ~new_n5117_ | ~new_n17364_;
  assign new_n17368_ = ~new_n17107_ | ~new_n17191_;
  assign new_n17369_ = ~new_n17261_;
  assign new_n17370_ = new_n4692_ | new_n5592_;
  assign new_n17371_ = new_n4697_ | new_n5122_;
  assign new_n17372_ = new_n4691_ | new_n5591_;
  assign new_n17373_ = ~new_n17179_;
  assign new_n17374_ = ~new_n5592_ | ~new_n17373_;
  assign new_n17375_ = ~new_n17374_ | ~new_n17189_;
  assign new_n17376_ = ~new_n17179_ | ~new_n17180_;
  assign new_n17377_ = ~new_n17376_ | ~new_n17375_;
  assign new_n17378_ = ~new_n17274_ | ~new_n17108_;
  assign new_n17379_ = ~new_n4691_ | ~new_n5591_;
  assign new_n17380_ = ~new_n17377_ | ~new_n17378_;
  assign new_n17381_ = new_n5120_ | new_n4698_;
  assign new_n17382_ = new_n5591_ | new_n4691_;
  assign new_n17383_ = ~new_n17261_ | ~new_n17230_;
  assign new_n17384_ = ~new_n17382_ | ~new_n17380_;
  assign new_n17385_ = ~new_n17258_;
  assign new_n17386_ = new_n5590_ | new_n4677_;
  assign new_n17387_ = ~new_n17386_ | ~new_n17258_;
  assign new_n17388_ = ~new_n4677_ | ~new_n5590_;
  assign new_n17389_ = ~new_n17256_;
  assign new_n17390_ = new_n5589_ | new_n4682_;
  assign new_n17391_ = ~new_n17390_ | ~new_n17256_;
  assign new_n17392_ = ~new_n4682_ | ~new_n5589_;
  assign new_n17393_ = ~new_n17254_;
  assign new_n17394_ = new_n4674_ | new_n5587_;
  assign new_n17395_ = ~new_n17275_ | ~new_n17272_;
  assign new_n17396_ = ~new_n17185_;
  assign new_n17397_ = new_n5588_ | new_n4681_;
  assign new_n17398_ = ~new_n17267_ | ~new_n17254_ | ~new_n17397_;
  assign new_n17399_ = ~new_n17253_;
  assign new_n17400_ = new_n5585_ | new_n4669_;
  assign new_n17401_ = ~new_n4669_ | ~new_n5585_;
  assign new_n17402_ = ~new_n17251_;
  assign new_n17403_ = ~new_n5584_ | ~new_n17251_;
  assign new_n17404_ = ~new_n17249_;
  assign new_n17405_ = ~new_n17397_ | ~new_n17254_;
  assign new_n17406_ = ~new_n17188_;
  assign new_n17407_ = new_n5587_ | new_n4674_;
  assign new_n17408_ = ~new_n17407_ | ~new_n17188_;
  assign new_n17409_ = ~new_n17234_ | ~new_n17408_;
  assign new_n17410_ = ~new_n17406_ | ~new_n17272_;
  assign new_n17411_ = ~new_n5586_ | ~new_n4673_;
  assign new_n17412_ = ~new_n17267_ | ~new_n17410_ | ~new_n17411_;
  assign new_n17413_ = new_n4674_ | new_n5587_;
  assign new_n17414_ = ~new_n17381_ | ~new_n17261_;
  assign new_n17415_ = ~new_n17190_;
  assign new_n17416_ = ~new_n17108_ | ~new_n17190_;
  assign new_n17417_ = ~new_n17235_ | ~new_n17416_;
  assign new_n17418_ = ~new_n17416_ | ~new_n17377_;
  assign new_n17419_ = ~new_n17552_ | ~new_n17418_;
  assign new_n17420_ = new_n5122_ | new_n4697_;
  assign new_n17421_ = ~new_n17420_ | ~new_n17190_;
  assign new_n17422_ = ~new_n17236_ | ~new_n17421_;
  assign new_n17423_ = ~new_n17415_ | ~new_n17179_;
  assign new_n17424_ = ~new_n4692_ | ~new_n5592_;
  assign new_n17425_ = ~new_n17237_ | ~new_n17423_;
  assign new_n17426_ = new_n5069_ | new_n4694_;
  assign new_n17427_ = ~new_n17260_;
  assign new_n17428_ = new_n4697_ | new_n5122_;
  assign new_n17429_ = new_n5114_ | new_n4689_;
  assign new_n17430_ = ~new_n17429_ | ~new_n17191_;
  assign new_n17431_ = ~new_n17238_ | ~new_n17430_;
  assign new_n17432_ = ~new_n17361_ | ~new_n17158_;
  assign new_n17433_ = ~new_n5117_ | ~new_n4685_;
  assign new_n17434_ = ~new_n17239_ | ~new_n17432_;
  assign new_n17435_ = new_n4689_ | new_n5114_;
  assign new_n17436_ = ~new_n17349_ | ~new_n17266_;
  assign new_n17437_ = ~new_n17192_;
  assign new_n17438_ = new_n5102_ | new_n4688_;
  assign new_n17439_ = ~new_n17438_ | ~new_n17192_;
  assign new_n17440_ = ~new_n17240_ | ~new_n17439_;
  assign new_n17441_ = ~new_n17437_ | ~new_n17271_;
  assign new_n17442_ = ~new_n4696_ | ~new_n5105_;
  assign new_n17443_ = ~new_n17241_ | ~new_n17441_;
  assign new_n17444_ = new_n4688_ | new_n5102_;
  assign new_n17445_ = new_n5093_ | new_n4699_;
  assign new_n17446_ = ~new_n17445_ | ~new_n17139_;
  assign new_n17447_ = ~new_n17242_ | ~new_n17446_;
  assign new_n17448_ = ~new_n17305_ | ~new_n17270_;
  assign new_n17449_ = ~new_n4678_ | ~new_n5096_;
  assign new_n17450_ = ~new_n17243_ | ~new_n17448_;
  assign new_n17451_ = ~new_n17306_ | ~new_n17270_;
  assign new_n17452_ = ~new_n17303_ | ~new_n17160_;
  assign new_n17453_ = ~new_n17313_ | ~new_n17121_;
  assign new_n17454_ = ~new_n17327_ | ~new_n17133_;
  assign new_n17455_ = ~new_n17330_ | ~new_n17279_;
  assign new_n17456_ = ~new_n17413_ | ~new_n17272_;
  assign new_n17457_ = ~new_n17397_ | ~new_n17275_;
  assign new_n17458_ = ~new_n17428_ | ~new_n17179_;
  assign new_n17459_ = ~new_n17381_ | ~new_n17176_;
  assign new_n17460_ = ~new_n17435_ | ~new_n17158_;
  assign new_n17461_ = ~new_n17444_ | ~new_n17271_;
  assign new_n17462_ = ~new_n17349_ | ~new_n17167_;
  assign new_n17463_ = ~new_n5584_ | ~new_n4670_;
  assign new_n17464_ = ~new_n17395_ | ~new_n17267_;
  assign new_n17465_ = ~new_n4673_ | ~new_n17394_;
  assign new_n17466_ = ~new_n5586_ | ~new_n17394_;
  assign new_n17467_ = ~new_n17400_ | ~new_n17395_ | ~new_n17267_;
  assign new_n17468_ = ~new_n17232_ | ~new_n17254_ | ~new_n17267_;
  assign new_n17469_ = ~new_n17396_ | ~new_n17400_;
  assign new_n17470_ = ~new_n4699_ | ~new_n17138_;
  assign new_n17471_ = ~new_n5093_ | ~new_n17137_;
  assign new_n17472_ = ~new_n17471_ | ~new_n17470_;
  assign new_n17473_ = ~new_n17451_ | ~new_n17139_;
  assign new_n17474_ = ~new_n17472_ | ~new_n17305_;
  assign new_n17475_ = ~new_n4700_ | ~new_n17135_;
  assign new_n17476_ = ~new_n5090_ | ~new_n17136_;
  assign new_n17477_ = ~new_n17476_ | ~new_n17475_;
  assign new_n17478_ = ~new_n17452_ | ~new_n17244_;
  assign new_n17479_ = ~new_n17302_ | ~new_n17477_;
  assign new_n17480_ = ~new_n4686_ | ~new_n17122_;
  assign new_n17481_ = ~new_n5087_ | ~new_n17120_;
  assign new_n17482_ = ~new_n4687_ | ~new_n17118_;
  assign new_n17483_ = ~new_n5084_ | ~new_n17119_;
  assign new_n17484_ = ~new_n17483_ | ~new_n17482_;
  assign new_n17485_ = ~new_n17453_ | ~new_n17140_;
  assign new_n17486_ = ~new_n17484_ | ~new_n17294_;
  assign new_n17487_ = ~new_n4683_ | ~new_n17134_;
  assign new_n17488_ = ~new_n5081_ | ~new_n17125_;
  assign new_n17489_ = ~new_n4676_ | ~new_n17123_;
  assign new_n17490_ = ~new_n5078_ | ~new_n17124_;
  assign new_n17491_ = ~new_n17490_ | ~new_n17489_;
  assign new_n17492_ = ~new_n17454_ | ~new_n17143_;
  assign new_n17493_ = ~new_n17491_ | ~new_n17320_;
  assign new_n17494_ = ~new_n4680_ | ~new_n17131_;
  assign new_n17495_ = ~new_n5075_ | ~new_n17132_;
  assign new_n17496_ = ~new_n17495_ | ~new_n17494_;
  assign new_n17497_ = ~new_n17455_ | ~new_n17245_;
  assign new_n17498_ = ~new_n17329_ | ~new_n17496_;
  assign new_n17499_ = ~new_n4684_ | ~new_n17126_;
  assign new_n17500_ = ~new_n5072_ | ~new_n17127_;
  assign new_n17501_ = ~new_n4671_ | ~new_n17247_;
  assign new_n17502_ = ~new_n5595_ | ~new_n17246_;
  assign new_n17503_ = ~new_n4671_ | ~new_n17247_;
  assign new_n17504_ = ~new_n5595_ | ~new_n17246_;
  assign new_n17505_ = ~new_n17504_ | ~new_n17503_;
  assign new_n17506_ = ~new_n17248_ | ~new_n17249_;
  assign new_n17507_ = ~new_n17404_ | ~new_n17505_;
  assign new_n17508_ = ~new_n4670_ | ~new_n17187_;
  assign new_n17509_ = ~new_n5584_ | ~new_n17186_;
  assign new_n17510_ = ~new_n4670_ | ~new_n17187_;
  assign new_n17511_ = ~new_n5584_ | ~new_n17186_;
  assign new_n17512_ = ~new_n17511_ | ~new_n17510_;
  assign new_n17513_ = ~new_n17250_ | ~new_n17251_;
  assign new_n17514_ = ~new_n17402_ | ~new_n17512_;
  assign new_n17515_ = ~new_n4669_ | ~new_n17145_;
  assign new_n17516_ = ~new_n5585_ | ~new_n17146_;
  assign new_n17517_ = ~new_n4669_ | ~new_n17145_;
  assign new_n17518_ = ~new_n5585_ | ~new_n17146_;
  assign new_n17519_ = ~new_n17518_ | ~new_n17517_;
  assign new_n17520_ = ~new_n17252_ | ~new_n17253_;
  assign new_n17521_ = ~new_n17399_ | ~new_n17519_;
  assign new_n17522_ = ~new_n4673_ | ~new_n17148_;
  assign new_n17523_ = ~new_n5586_ | ~new_n17147_;
  assign new_n17524_ = ~new_n4674_ | ~new_n17149_;
  assign new_n17525_ = ~new_n5587_ | ~new_n17150_;
  assign new_n17526_ = ~new_n17525_ | ~new_n17524_;
  assign new_n17527_ = ~new_n17456_ | ~new_n17188_;
  assign new_n17528_ = ~new_n17526_ | ~new_n17406_;
  assign new_n17529_ = ~new_n4681_ | ~new_n17151_;
  assign new_n17530_ = ~new_n5588_ | ~new_n17152_;
  assign new_n17531_ = ~new_n17530_ | ~new_n17529_;
  assign new_n17532_ = ~new_n17457_ | ~new_n17254_;
  assign new_n17533_ = ~new_n17393_ | ~new_n17531_;
  assign new_n17534_ = ~new_n4682_ | ~new_n17183_;
  assign new_n17535_ = ~new_n5589_ | ~new_n17184_;
  assign new_n17536_ = ~new_n4682_ | ~new_n17183_;
  assign new_n17537_ = ~new_n5589_ | ~new_n17184_;
  assign new_n17538_ = ~new_n17537_ | ~new_n17536_;
  assign new_n17539_ = ~new_n17255_ | ~new_n17256_;
  assign new_n17540_ = ~new_n17389_ | ~new_n17538_;
  assign new_n17541_ = ~new_n4677_ | ~new_n17181_;
  assign new_n17542_ = ~new_n5590_ | ~new_n17182_;
  assign new_n17543_ = ~new_n4677_ | ~new_n17181_;
  assign new_n17544_ = ~new_n5590_ | ~new_n17182_;
  assign new_n17545_ = ~new_n17544_ | ~new_n17543_;
  assign new_n17546_ = ~new_n17257_ | ~new_n17258_;
  assign new_n17547_ = ~new_n17385_ | ~new_n17545_;
  assign new_n17548_ = ~new_n4691_ | ~new_n17153_;
  assign new_n17549_ = ~new_n5591_ | ~new_n17154_;
  assign new_n17550_ = ~new_n4691_ | ~new_n17153_;
  assign new_n17551_ = ~new_n5591_ | ~new_n17154_;
  assign new_n17552_ = ~new_n17551_ | ~new_n17550_;
  assign new_n17553_ = ~new_n4692_ | ~new_n17180_;
  assign new_n17554_ = ~new_n5592_ | ~new_n17189_;
  assign new_n17555_ = ~new_n17281_ | ~new_n17260_;
  assign new_n17556_ = ~new_n17427_ | ~new_n17130_;
  assign new_n17557_ = ~new_n4697_ | ~new_n17177_;
  assign new_n17558_ = ~new_n5122_ | ~new_n17178_;
  assign new_n17559_ = ~new_n17558_ | ~new_n17557_;
  assign new_n17560_ = ~new_n17458_ | ~new_n17190_;
  assign new_n17561_ = ~new_n17559_ | ~new_n17415_;
  assign new_n17562_ = ~new_n4698_ | ~new_n17174_;
  assign new_n17563_ = ~new_n5120_ | ~new_n17175_;
  assign new_n17564_ = ~new_n17563_ | ~new_n17562_;
  assign new_n17565_ = ~new_n17459_ | ~new_n17261_;
  assign new_n17566_ = ~new_n17369_ | ~new_n17564_;
  assign new_n17567_ = ~new_n4685_ | ~new_n17159_;
  assign new_n17568_ = ~new_n5117_ | ~new_n17157_;
  assign new_n17569_ = ~new_n4689_ | ~new_n17155_;
  assign new_n17570_ = ~new_n5114_ | ~new_n17156_;
  assign new_n17571_ = ~new_n17570_ | ~new_n17569_;
  assign new_n17572_ = ~new_n17460_ | ~new_n17191_;
  assign new_n17573_ = ~new_n17571_ | ~new_n17361_;
  assign new_n17574_ = ~new_n4690_ | ~new_n17172_;
  assign new_n17575_ = ~new_n5111_ | ~new_n17173_;
  assign new_n17576_ = ~new_n4690_ | ~new_n17172_;
  assign new_n17577_ = ~new_n5111_ | ~new_n17173_;
  assign new_n17578_ = ~new_n17577_ | ~new_n17576_;
  assign new_n17579_ = ~new_n17262_ | ~new_n17263_;
  assign new_n17580_ = ~new_n17357_ | ~new_n17578_;
  assign new_n17581_ = ~new_n4695_ | ~new_n17170_;
  assign new_n17582_ = ~new_n5108_ | ~new_n17171_;
  assign new_n17583_ = ~new_n4695_ | ~new_n17170_;
  assign new_n17584_ = ~new_n5108_ | ~new_n17171_;
  assign new_n17585_ = ~new_n17584_ | ~new_n17583_;
  assign new_n17586_ = ~new_n17264_ | ~new_n17265_;
  assign new_n17587_ = ~new_n17353_ | ~new_n17585_;
  assign new_n17588_ = ~new_n4696_ | ~new_n17168_;
  assign new_n17589_ = ~new_n5105_ | ~new_n17169_;
  assign new_n17590_ = ~new_n4688_ | ~new_n17163_;
  assign new_n17591_ = ~new_n5102_ | ~new_n17164_;
  assign new_n17592_ = ~new_n17591_ | ~new_n17590_;
  assign new_n17593_ = ~new_n17461_ | ~new_n17192_;
  assign new_n17594_ = ~new_n17592_ | ~new_n17437_;
  assign new_n17595_ = ~new_n4679_ | ~new_n17165_;
  assign new_n17596_ = ~new_n5099_ | ~new_n17166_;
  assign new_n17597_ = ~new_n17596_ | ~new_n17595_;
  assign new_n17598_ = ~new_n17462_ | ~new_n17266_;
  assign new_n17599_ = ~new_n17343_ | ~new_n17597_;
  assign new_n17600_ = ~new_n4678_ | ~new_n17161_;
  assign new_n17601_ = ~new_n5096_ | ~new_n17162_;
  assign new_n17602_ = ~new_n4693_ | ~new_n17128_;
  assign new_n17603_ = ~new_n5064_ | ~new_n17129_;
  assign new_n17604_ = new_n17779_ & new_n17778_;
  assign new_n17605_ = new_n17797_ & new_n17796_;
  assign new_n17606_ = new_n17837_ & new_n17836_;
  assign new_n17607_ = new_n17846_ & new_n17845_;
  assign new_n17608_ = new_n17864_ & new_n17863_;
  assign new_n17609_ = new_n17872_ & new_n17871_;
  assign new_n17610_ = new_n17951_ & new_n17948_;
  assign new_n17611_ = new_n17944_ & new_n17941_;
  assign new_n17612_ = new_n17935_ & new_n17932_;
  assign new_n17613_ = new_n17926_ & new_n17923_;
  assign new_n17614_ = new_n17920_ & new_n17918_;
  assign new_n17615_ = new_n17913_ & new_n17910_;
  assign new_n17616_ = new_n17835_ & new_n17832_;
  assign new_n17617_ = new_n17827_ & new_n17824_;
  assign new_n17618_ = new_n17813_ & new_n17810_;
  assign new_n17619_ = ~new_n5084_;
  assign new_n17620_ = ~new_n4687_;
  assign new_n17621_ = ~new_n4686_;
  assign new_n17622_ = ~new_n4687_ | ~new_n5084_;
  assign new_n17623_ = ~new_n5087_;
  assign new_n17624_ = ~new_n5078_;
  assign new_n17625_ = ~new_n4676_;
  assign new_n17626_ = ~new_n4683_;
  assign new_n17627_ = ~new_n5072_;
  assign new_n17628_ = ~new_n4684_;
  assign new_n17629_ = ~new_n5064_;
  assign new_n17630_ = ~new_n4693_;
  assign new_n17631_ = ~new_n4693_ | ~new_n5064_;
  assign new_n17632_ = ~new_n5075_;
  assign new_n17633_ = ~new_n4680_;
  assign new_n17634_ = ~new_n4676_ | ~new_n5078_;
  assign new_n17635_ = ~new_n5081_;
  assign new_n17636_ = ~new_n5090_;
  assign new_n17637_ = ~new_n4700_;
  assign new_n17638_ = ~new_n4699_;
  assign new_n17639_ = ~new_n5093_;
  assign new_n17640_ = ~new_n17663_ | ~new_n17805_;
  assign new_n17641_ = ~new_n17717_ | ~new_n17793_;
  assign new_n17642_ = ~new_n17782_ | ~new_n17783_;
  assign new_n17643_ = ~new_n5069_ | ~new_n4694_;
  assign new_n17644_ = ~new_n17722_ | ~new_n17819_;
  assign new_n17645_ = ~new_n17816_ | ~new_n17815_;
  assign new_n17646_ = ~new_n5585_;
  assign new_n17647_ = ~new_n4669_;
  assign new_n17648_ = ~new_n4673_;
  assign new_n17649_ = ~new_n5586_;
  assign new_n17650_ = ~new_n5587_;
  assign new_n17651_ = ~new_n4674_;
  assign new_n17652_ = ~new_n5588_;
  assign new_n17653_ = ~new_n4681_;
  assign new_n17654_ = ~new_n5591_;
  assign new_n17655_ = ~new_n4691_;
  assign new_n17656_ = ~new_n5114_;
  assign new_n17657_ = ~new_n4689_;
  assign new_n17658_ = ~new_n4685_;
  assign new_n17659_ = ~new_n4689_ | ~new_n5114_;
  assign new_n17660_ = ~new_n5117_;
  assign new_n17661_ = ~new_n5096_;
  assign new_n17662_ = ~new_n4678_;
  assign new_n17663_ = ~new_n4700_ | ~new_n5090_;
  assign new_n17664_ = ~new_n5102_;
  assign new_n17665_ = ~new_n4688_;
  assign new_n17666_ = ~new_n5099_;
  assign new_n17667_ = ~new_n4679_;
  assign new_n17668_ = ~new_n4679_ | ~new_n5099_;
  assign new_n17669_ = ~new_n5105_;
  assign new_n17670_ = ~new_n4696_;
  assign new_n17671_ = ~new_n5108_;
  assign new_n17672_ = ~new_n4695_;
  assign new_n17673_ = ~new_n5111_;
  assign new_n17674_ = ~new_n4690_;
  assign new_n17675_ = ~new_n5120_;
  assign new_n17676_ = ~new_n4698_;
  assign new_n17677_ = ~new_n4698_ | ~new_n5120_;
  assign new_n17678_ = ~new_n5122_;
  assign new_n17679_ = ~new_n4697_;
  assign new_n17680_ = ~new_n4697_ | ~new_n5122_;
  assign new_n17681_ = ~new_n5592_;
  assign new_n17682_ = ~new_n5590_;
  assign new_n17683_ = ~new_n4677_;
  assign new_n17684_ = ~new_n5589_;
  assign new_n17685_ = ~new_n4682_;
  assign new_n17686_ = ~new_n5586_ | ~new_n4673_;
  assign new_n17687_ = ~new_n4670_;
  assign new_n17688_ = ~new_n5584_;
  assign new_n17689_ = ~new_n17906_ | ~new_n17776_;
  assign new_n17690_ = ~new_n4692_;
  assign new_n17691_ = ~new_n17677_ | ~new_n17915_;
  assign new_n17692_ = ~new_n17861_ | ~new_n17860_;
  assign new_n17693_ = ~new_n17668_ | ~new_n17937_;
  assign new_n17694_ = ~new_n18057_ | ~new_n18056_;
  assign new_n17695_ = ~new_n18104_ | ~new_n18103_;
  assign new_n17696_ = ~new_n17975_ | ~new_n17974_;
  assign new_n17697_ = ~new_n17980_ | ~new_n17979_;
  assign new_n17698_ = ~new_n17987_ | ~new_n17986_;
  assign new_n17699_ = ~new_n17994_ | ~new_n17993_;
  assign new_n17700_ = ~new_n17999_ | ~new_n17998_;
  assign new_n17701_ = ~new_n18008_ | ~new_n18007_;
  assign new_n17702_ = ~new_n18015_ | ~new_n18014_;
  assign new_n17703_ = ~new_n18022_ | ~new_n18021_;
  assign new_n17704_ = ~new_n18029_ | ~new_n18028_;
  assign new_n17705_ = ~new_n18034_ | ~new_n18033_;
  assign new_n17706_ = ~new_n18041_ | ~new_n18040_;
  assign new_n17707_ = ~new_n18048_ | ~new_n18047_;
  assign new_n17708_ = ~new_n18062_ | ~new_n18061_;
  assign new_n17709_ = ~new_n18067_ | ~new_n18066_;
  assign new_n17710_ = ~new_n18074_ | ~new_n18073_;
  assign new_n17711_ = ~new_n18081_ | ~new_n18080_;
  assign new_n17712_ = ~new_n18088_ | ~new_n18087_;
  assign new_n17713_ = ~new_n18095_ | ~new_n18094_;
  assign new_n17714_ = ~new_n18100_ | ~new_n18099_;
  assign new_n17715_ = new_n17789_ & new_n17787_;
  assign new_n17716_ = new_n17604_ & new_n17780_;
  assign new_n17717_ = new_n17794_ & new_n17792_;
  assign new_n17718_ = new_n17801_ & new_n17800_;
  assign new_n17719_ = new_n17622_ & new_n17982_ & new_n17981_;
  assign new_n17720_ = new_n17812_ & new_n17605_;
  assign new_n17721_ = new_n17781_ & new_n17780_;
  assign new_n17722_ = new_n17820_ & new_n17818_;
  assign new_n17723_ = new_n17634_ & new_n17989_ & new_n17988_;
  assign new_n17724_ = new_n17826_ & new_n17604_;
  assign new_n17725_ = new_n17834_ & new_n17781_;
  assign new_n17726_ = new_n17804_ & new_n17606_;
  assign new_n17727_ = new_n17843_ & new_n17839_;
  assign new_n17728_ = new_n17850_ & new_n17607_;
  assign new_n17729_ = new_n17848_ & new_n17772_;
  assign new_n17730_ = new_n17868_ & new_n17867_;
  assign new_n17731_ = new_n17873_ & new_n17609_ & new_n17882_;
  assign new_n17732_ = new_n17885_ & new_n17880_;
  assign new_n17733_ = new_n17901_ & new_n17898_;
  assign new_n17734_ = new_n17968_ & new_n17902_;
  assign new_n17735_ = new_n17773_ & new_n18024_ & new_n18023_;
  assign new_n17736_ = new_n17760_ & new_n17878_;
  assign new_n17737_ = new_n17680_ & new_n18055_ & new_n18054_;
  assign new_n17738_ = new_n17925_ & new_n17609_;
  assign new_n17739_ = new_n17659_ & new_n18069_ & new_n18068_;
  assign new_n17740_ = new_n17934_ & new_n17608_;
  assign new_n17741_ = new_n17772_ & new_n18090_ & new_n18089_;
  assign new_n17742_ = new_n17943_ & new_n17607_;
  assign new_n17743_ = new_n17771_ & new_n18102_ & new_n18101_;
  assign new_n17744_ = new_n17950_ & new_n17606_;
  assign new_n17745_ = ~new_n17718_ | ~new_n17802_;
  assign new_n17746_ = ~new_n17817_ | ~new_n17829_;
  assign new_n17747_ = ~new_n4671_;
  assign new_n17748_ = ~new_n5595_;
  assign new_n17749_ = new_n18003_ & new_n18002_;
  assign new_n17750_ = ~new_n17964_ | ~new_n17904_ | ~new_n17769_;
  assign new_n17751_ = new_n18010_ & new_n18009_;
  assign new_n17752_ = ~new_n17734_ | ~new_n17970_ | ~new_n17969_;
  assign new_n17753_ = new_n18017_ & new_n18016_;
  assign new_n17754_ = ~new_n17686_ | ~new_n17965_ | ~new_n17899_;
  assign new_n17755_ = ~new_n17893_ | ~new_n17892_;
  assign new_n17756_ = new_n18036_ & new_n18035_;
  assign new_n17757_ = ~new_n17889_ | ~new_n17888_;
  assign new_n17758_ = new_n18043_ & new_n18042_;
  assign new_n17759_ = ~new_n17732_ | ~new_n17884_;
  assign new_n17760_ = new_n18050_ & new_n18049_;
  assign new_n17761_ = ~new_n17643_ | ~new_n17927_;
  assign new_n17762_ = ~new_n17730_ | ~new_n17869_;
  assign new_n17763_ = new_n18076_ & new_n18075_;
  assign new_n17764_ = ~new_n17857_ | ~new_n17856_;
  assign new_n17765_ = new_n18083_ & new_n18082_;
  assign new_n17766_ = ~new_n17853_ | ~new_n17852_;
  assign new_n17767_ = ~new_n17727_ | ~new_n17842_;
  assign new_n17768_ = ~new_n17967_ | ~new_n17966_;
  assign new_n17769_ = ~new_n4670_ | ~new_n17752_;
  assign new_n17770_ = ~new_n17634_;
  assign new_n17771_ = ~new_n5093_ | ~new_n4699_;
  assign new_n17772_ = ~new_n4688_ | ~new_n5102_;
  assign new_n17773_ = ~new_n4674_ | ~new_n5587_;
  assign new_n17774_ = ~new_n17668_;
  assign new_n17775_ = ~new_n17677_;
  assign new_n17776_ = ~new_n4681_ | ~new_n5588_;
  assign new_n17777_ = ~new_n17663_;
  assign new_n17778_ = new_n4683_ | new_n5081_;
  assign new_n17779_ = new_n4676_ | new_n5078_;
  assign new_n17780_ = new_n5075_ | new_n4680_;
  assign new_n17781_ = new_n5072_ | new_n4684_;
  assign new_n17782_ = ~new_n17631_;
  assign new_n17783_ = new_n5069_ | new_n4694_;
  assign new_n17784_ = ~new_n17642_;
  assign new_n17785_ = ~new_n17643_;
  assign new_n17786_ = ~new_n17642_ | ~new_n17643_;
  assign new_n17787_ = ~new_n4684_ | ~new_n5072_;
  assign new_n17788_ = ~new_n17786_ | ~new_n17781_;
  assign new_n17789_ = ~new_n4680_ | ~new_n5075_;
  assign new_n17790_ = ~new_n17715_ | ~new_n17788_;
  assign new_n17791_ = ~new_n17635_ | ~new_n17634_;
  assign new_n17792_ = ~new_n4683_ | ~new_n17791_;
  assign new_n17793_ = ~new_n17716_ | ~new_n17790_;
  assign new_n17794_ = ~new_n5081_ | ~new_n17770_;
  assign new_n17795_ = ~new_n17641_;
  assign new_n17796_ = new_n4686_ | new_n5087_;
  assign new_n17797_ = new_n4687_ | new_n5084_;
  assign new_n17798_ = ~new_n17622_;
  assign new_n17799_ = ~new_n17623_ | ~new_n17622_;
  assign new_n17800_ = ~new_n4686_ | ~new_n17799_;
  assign new_n17801_ = ~new_n5087_ | ~new_n17798_;
  assign new_n17802_ = ~new_n17605_ | ~new_n17641_;
  assign new_n17803_ = ~new_n17745_;
  assign new_n17804_ = new_n5090_ | new_n4700_;
  assign new_n17805_ = ~new_n17804_ | ~new_n17745_;
  assign new_n17806_ = ~new_n17640_;
  assign new_n17807_ = new_n4699_ | new_n5093_;
  assign new_n17808_ = new_n5084_ | new_n4687_;
  assign new_n17809_ = ~new_n17808_ | ~new_n17641_;
  assign new_n17810_ = ~new_n17719_ | ~new_n17809_;
  assign new_n17811_ = ~new_n17795_ | ~new_n17622_;
  assign new_n17812_ = ~new_n5087_ | ~new_n4686_;
  assign new_n17813_ = ~new_n17720_ | ~new_n17811_;
  assign new_n17814_ = new_n4687_ | new_n5084_;
  assign new_n17815_ = ~new_n17785_ | ~new_n17781_;
  assign new_n17816_ = ~new_n4684_ | ~new_n5072_;
  assign new_n17817_ = ~new_n17645_;
  assign new_n17818_ = ~new_n17721_ | ~new_n17784_;
  assign new_n17819_ = ~new_n17645_ | ~new_n17780_;
  assign new_n17820_ = ~new_n4680_ | ~new_n5075_;
  assign new_n17821_ = ~new_n17644_;
  assign new_n17822_ = new_n5078_ | new_n4676_;
  assign new_n17823_ = ~new_n17822_ | ~new_n17644_;
  assign new_n17824_ = ~new_n17723_ | ~new_n17823_;
  assign new_n17825_ = ~new_n17821_ | ~new_n17634_;
  assign new_n17826_ = ~new_n5081_ | ~new_n4683_;
  assign new_n17827_ = ~new_n17724_ | ~new_n17825_;
  assign new_n17828_ = new_n4676_ | new_n5078_;
  assign new_n17829_ = ~new_n17784_ | ~new_n17781_;
  assign new_n17830_ = ~new_n17746_;
  assign new_n17831_ = ~new_n4680_ | ~new_n5075_;
  assign new_n17832_ = ~new_n17642_ | ~new_n17643_ | ~new_n18001_ | ~new_n18000_;
  assign new_n17833_ = ~new_n17643_ | ~new_n17642_;
  assign new_n17834_ = ~new_n4684_ | ~new_n5072_;
  assign new_n17835_ = ~new_n17725_ | ~new_n17833_;
  assign new_n17836_ = new_n4699_ | new_n5093_;
  assign new_n17837_ = new_n4678_ | new_n5096_;
  assign new_n17838_ = ~new_n17777_ | ~new_n17606_;
  assign new_n17839_ = ~new_n4678_ | ~new_n5096_;
  assign new_n17840_ = ~new_n17771_ | ~new_n17838_;
  assign new_n17841_ = new_n5096_ | new_n4678_;
  assign new_n17842_ = ~new_n17726_ | ~new_n17745_;
  assign new_n17843_ = ~new_n17841_ | ~new_n17840_;
  assign new_n17844_ = ~new_n17767_;
  assign new_n17845_ = new_n4696_ | new_n5105_;
  assign new_n17846_ = new_n4688_ | new_n5102_;
  assign new_n17847_ = ~new_n17774_ | ~new_n17607_;
  assign new_n17848_ = ~new_n4696_ | ~new_n5105_;
  assign new_n17849_ = ~new_n17729_ | ~new_n17847_;
  assign new_n17850_ = new_n5099_ | new_n4679_;
  assign new_n17851_ = new_n5105_ | new_n4696_;
  assign new_n17852_ = ~new_n17728_ | ~new_n17767_;
  assign new_n17853_ = ~new_n17851_ | ~new_n17849_;
  assign new_n17854_ = ~new_n17766_;
  assign new_n17855_ = new_n5108_ | new_n4695_;
  assign new_n17856_ = ~new_n17855_ | ~new_n17766_;
  assign new_n17857_ = ~new_n4695_ | ~new_n5108_;
  assign new_n17858_ = ~new_n17764_;
  assign new_n17859_ = new_n5111_ | new_n4690_;
  assign new_n17860_ = ~new_n17859_ | ~new_n17764_;
  assign new_n17861_ = ~new_n4690_ | ~new_n5111_;
  assign new_n17862_ = ~new_n17692_;
  assign new_n17863_ = new_n4685_ | new_n5117_;
  assign new_n17864_ = new_n4689_ | new_n5114_;
  assign new_n17865_ = ~new_n17659_;
  assign new_n17866_ = ~new_n17660_ | ~new_n17659_;
  assign new_n17867_ = ~new_n4685_ | ~new_n17866_;
  assign new_n17868_ = ~new_n5117_ | ~new_n17865_;
  assign new_n17869_ = ~new_n17608_ | ~new_n17692_;
  assign new_n17870_ = ~new_n17762_;
  assign new_n17871_ = new_n4692_ | new_n5592_;
  assign new_n17872_ = new_n4697_ | new_n5122_;
  assign new_n17873_ = new_n4691_ | new_n5591_;
  assign new_n17874_ = ~new_n17680_;
  assign new_n17875_ = ~new_n5592_ | ~new_n17874_;
  assign new_n17876_ = ~new_n17875_ | ~new_n17690_;
  assign new_n17877_ = ~new_n17680_ | ~new_n17681_;
  assign new_n17878_ = ~new_n17877_ | ~new_n17876_;
  assign new_n17879_ = ~new_n17775_ | ~new_n17609_;
  assign new_n17880_ = ~new_n4691_ | ~new_n5591_;
  assign new_n17881_ = ~new_n17878_ | ~new_n17879_;
  assign new_n17882_ = new_n5120_ | new_n4698_;
  assign new_n17883_ = new_n5591_ | new_n4691_;
  assign new_n17884_ = ~new_n17762_ | ~new_n17731_;
  assign new_n17885_ = ~new_n17883_ | ~new_n17881_;
  assign new_n17886_ = ~new_n17759_;
  assign new_n17887_ = new_n5590_ | new_n4677_;
  assign new_n17888_ = ~new_n17887_ | ~new_n17759_;
  assign new_n17889_ = ~new_n4677_ | ~new_n5590_;
  assign new_n17890_ = ~new_n17757_;
  assign new_n17891_ = new_n5589_ | new_n4682_;
  assign new_n17892_ = ~new_n17891_ | ~new_n17757_;
  assign new_n17893_ = ~new_n4682_ | ~new_n5589_;
  assign new_n17894_ = ~new_n17755_;
  assign new_n17895_ = new_n4674_ | new_n5587_;
  assign new_n17896_ = ~new_n17776_ | ~new_n17773_;
  assign new_n17897_ = ~new_n17686_;
  assign new_n17898_ = new_n5588_ | new_n4681_;
  assign new_n17899_ = ~new_n17768_ | ~new_n17755_ | ~new_n17898_;
  assign new_n17900_ = ~new_n17754_;
  assign new_n17901_ = new_n5585_ | new_n4669_;
  assign new_n17902_ = ~new_n4669_ | ~new_n5585_;
  assign new_n17903_ = ~new_n17752_;
  assign new_n17904_ = ~new_n5584_ | ~new_n17752_;
  assign new_n17905_ = ~new_n17750_;
  assign new_n17906_ = ~new_n17898_ | ~new_n17755_;
  assign new_n17907_ = ~new_n17689_;
  assign new_n17908_ = new_n5587_ | new_n4674_;
  assign new_n17909_ = ~new_n17908_ | ~new_n17689_;
  assign new_n17910_ = ~new_n17735_ | ~new_n17909_;
  assign new_n17911_ = ~new_n17907_ | ~new_n17773_;
  assign new_n17912_ = ~new_n5586_ | ~new_n4673_;
  assign new_n17913_ = ~new_n17768_ | ~new_n17911_ | ~new_n17912_;
  assign new_n17914_ = new_n4674_ | new_n5587_;
  assign new_n17915_ = ~new_n17882_ | ~new_n17762_;
  assign new_n17916_ = ~new_n17691_;
  assign new_n17917_ = ~new_n17609_ | ~new_n17691_;
  assign new_n17918_ = ~new_n17736_ | ~new_n17917_;
  assign new_n17919_ = ~new_n17917_ | ~new_n17878_;
  assign new_n17920_ = ~new_n18053_ | ~new_n17919_;
  assign new_n17921_ = new_n5122_ | new_n4697_;
  assign new_n17922_ = ~new_n17921_ | ~new_n17691_;
  assign new_n17923_ = ~new_n17737_ | ~new_n17922_;
  assign new_n17924_ = ~new_n17916_ | ~new_n17680_;
  assign new_n17925_ = ~new_n4692_ | ~new_n5592_;
  assign new_n17926_ = ~new_n17738_ | ~new_n17924_;
  assign new_n17927_ = new_n5069_ | new_n4694_;
  assign new_n17928_ = ~new_n17761_;
  assign new_n17929_ = new_n4697_ | new_n5122_;
  assign new_n17930_ = new_n5114_ | new_n4689_;
  assign new_n17931_ = ~new_n17930_ | ~new_n17692_;
  assign new_n17932_ = ~new_n17739_ | ~new_n17931_;
  assign new_n17933_ = ~new_n17862_ | ~new_n17659_;
  assign new_n17934_ = ~new_n5117_ | ~new_n4685_;
  assign new_n17935_ = ~new_n17740_ | ~new_n17933_;
  assign new_n17936_ = new_n4689_ | new_n5114_;
  assign new_n17937_ = ~new_n17850_ | ~new_n17767_;
  assign new_n17938_ = ~new_n17693_;
  assign new_n17939_ = new_n5102_ | new_n4688_;
  assign new_n17940_ = ~new_n17939_ | ~new_n17693_;
  assign new_n17941_ = ~new_n17741_ | ~new_n17940_;
  assign new_n17942_ = ~new_n17938_ | ~new_n17772_;
  assign new_n17943_ = ~new_n4696_ | ~new_n5105_;
  assign new_n17944_ = ~new_n17742_ | ~new_n17942_;
  assign new_n17945_ = new_n4688_ | new_n5102_;
  assign new_n17946_ = new_n5093_ | new_n4699_;
  assign new_n17947_ = ~new_n17946_ | ~new_n17640_;
  assign new_n17948_ = ~new_n17743_ | ~new_n17947_;
  assign new_n17949_ = ~new_n17806_ | ~new_n17771_;
  assign new_n17950_ = ~new_n4678_ | ~new_n5096_;
  assign new_n17951_ = ~new_n17744_ | ~new_n17949_;
  assign new_n17952_ = ~new_n17807_ | ~new_n17771_;
  assign new_n17953_ = ~new_n17804_ | ~new_n17663_;
  assign new_n17954_ = ~new_n17814_ | ~new_n17622_;
  assign new_n17955_ = ~new_n17828_ | ~new_n17634_;
  assign new_n17956_ = ~new_n17831_ | ~new_n17780_;
  assign new_n17957_ = ~new_n17914_ | ~new_n17773_;
  assign new_n17958_ = ~new_n17898_ | ~new_n17776_;
  assign new_n17959_ = ~new_n17929_ | ~new_n17680_;
  assign new_n17960_ = ~new_n17882_ | ~new_n17677_;
  assign new_n17961_ = ~new_n17936_ | ~new_n17659_;
  assign new_n17962_ = ~new_n17945_ | ~new_n17772_;
  assign new_n17963_ = ~new_n17850_ | ~new_n17668_;
  assign new_n17964_ = ~new_n5584_ | ~new_n4670_;
  assign new_n17965_ = ~new_n17896_ | ~new_n17768_;
  assign new_n17966_ = ~new_n4673_ | ~new_n17895_;
  assign new_n17967_ = ~new_n5586_ | ~new_n17895_;
  assign new_n17968_ = ~new_n17901_ | ~new_n17896_ | ~new_n17768_;
  assign new_n17969_ = ~new_n17733_ | ~new_n17755_ | ~new_n17768_;
  assign new_n17970_ = ~new_n17897_ | ~new_n17901_;
  assign new_n17971_ = ~new_n4699_ | ~new_n17639_;
  assign new_n17972_ = ~new_n5093_ | ~new_n17638_;
  assign new_n17973_ = ~new_n17972_ | ~new_n17971_;
  assign new_n17974_ = ~new_n17952_ | ~new_n17640_;
  assign new_n17975_ = ~new_n17973_ | ~new_n17806_;
  assign new_n17976_ = ~new_n4700_ | ~new_n17636_;
  assign new_n17977_ = ~new_n5090_ | ~new_n17637_;
  assign new_n17978_ = ~new_n17977_ | ~new_n17976_;
  assign new_n17979_ = ~new_n17953_ | ~new_n17745_;
  assign new_n17980_ = ~new_n17803_ | ~new_n17978_;
  assign new_n17981_ = ~new_n4686_ | ~new_n17623_;
  assign new_n17982_ = ~new_n5087_ | ~new_n17621_;
  assign new_n17983_ = ~new_n4687_ | ~new_n17619_;
  assign new_n17984_ = ~new_n5084_ | ~new_n17620_;
  assign new_n17985_ = ~new_n17984_ | ~new_n17983_;
  assign new_n17986_ = ~new_n17954_ | ~new_n17641_;
  assign new_n17987_ = ~new_n17985_ | ~new_n17795_;
  assign new_n17988_ = ~new_n4683_ | ~new_n17635_;
  assign new_n17989_ = ~new_n5081_ | ~new_n17626_;
  assign new_n17990_ = ~new_n4676_ | ~new_n17624_;
  assign new_n17991_ = ~new_n5078_ | ~new_n17625_;
  assign new_n17992_ = ~new_n17991_ | ~new_n17990_;
  assign new_n17993_ = ~new_n17955_ | ~new_n17644_;
  assign new_n17994_ = ~new_n17992_ | ~new_n17821_;
  assign new_n17995_ = ~new_n4680_ | ~new_n17632_;
  assign new_n17996_ = ~new_n5075_ | ~new_n17633_;
  assign new_n17997_ = ~new_n17996_ | ~new_n17995_;
  assign new_n17998_ = ~new_n17956_ | ~new_n17746_;
  assign new_n17999_ = ~new_n17830_ | ~new_n17997_;
  assign new_n18000_ = ~new_n4684_ | ~new_n17627_;
  assign new_n18001_ = ~new_n5072_ | ~new_n17628_;
  assign new_n18002_ = ~new_n4671_ | ~new_n17748_;
  assign new_n18003_ = ~new_n5595_ | ~new_n17747_;
  assign new_n18004_ = ~new_n4671_ | ~new_n17748_;
  assign new_n18005_ = ~new_n5595_ | ~new_n17747_;
  assign new_n18006_ = ~new_n18005_ | ~new_n18004_;
  assign new_n18007_ = ~new_n17749_ | ~new_n17750_;
  assign new_n18008_ = ~new_n17905_ | ~new_n18006_;
  assign new_n18009_ = ~new_n4670_ | ~new_n17688_;
  assign new_n18010_ = ~new_n5584_ | ~new_n17687_;
  assign new_n18011_ = ~new_n4670_ | ~new_n17688_;
  assign new_n18012_ = ~new_n5584_ | ~new_n17687_;
  assign new_n18013_ = ~new_n18012_ | ~new_n18011_;
  assign new_n18014_ = ~new_n17751_ | ~new_n17752_;
  assign new_n18015_ = ~new_n17903_ | ~new_n18013_;
  assign new_n18016_ = ~new_n4669_ | ~new_n17646_;
  assign new_n18017_ = ~new_n5585_ | ~new_n17647_;
  assign new_n18018_ = ~new_n4669_ | ~new_n17646_;
  assign new_n18019_ = ~new_n5585_ | ~new_n17647_;
  assign new_n18020_ = ~new_n18019_ | ~new_n18018_;
  assign new_n18021_ = ~new_n17753_ | ~new_n17754_;
  assign new_n18022_ = ~new_n17900_ | ~new_n18020_;
  assign new_n18023_ = ~new_n4673_ | ~new_n17649_;
  assign new_n18024_ = ~new_n5586_ | ~new_n17648_;
  assign new_n18025_ = ~new_n4674_ | ~new_n17650_;
  assign new_n18026_ = ~new_n5587_ | ~new_n17651_;
  assign new_n18027_ = ~new_n18026_ | ~new_n18025_;
  assign new_n18028_ = ~new_n17957_ | ~new_n17689_;
  assign new_n18029_ = ~new_n18027_ | ~new_n17907_;
  assign new_n18030_ = ~new_n4681_ | ~new_n17652_;
  assign new_n18031_ = ~new_n5588_ | ~new_n17653_;
  assign new_n18032_ = ~new_n18031_ | ~new_n18030_;
  assign new_n18033_ = ~new_n17958_ | ~new_n17755_;
  assign new_n18034_ = ~new_n17894_ | ~new_n18032_;
  assign new_n18035_ = ~new_n4682_ | ~new_n17684_;
  assign new_n18036_ = ~new_n5589_ | ~new_n17685_;
  assign new_n18037_ = ~new_n4682_ | ~new_n17684_;
  assign new_n18038_ = ~new_n5589_ | ~new_n17685_;
  assign new_n18039_ = ~new_n18038_ | ~new_n18037_;
  assign new_n18040_ = ~new_n17756_ | ~new_n17757_;
  assign new_n18041_ = ~new_n17890_ | ~new_n18039_;
  assign new_n18042_ = ~new_n4677_ | ~new_n17682_;
  assign new_n18043_ = ~new_n5590_ | ~new_n17683_;
  assign new_n18044_ = ~new_n4677_ | ~new_n17682_;
  assign new_n18045_ = ~new_n5590_ | ~new_n17683_;
  assign new_n18046_ = ~new_n18045_ | ~new_n18044_;
  assign new_n18047_ = ~new_n17758_ | ~new_n17759_;
  assign new_n18048_ = ~new_n17886_ | ~new_n18046_;
  assign new_n18049_ = ~new_n4691_ | ~new_n17654_;
  assign new_n18050_ = ~new_n5591_ | ~new_n17655_;
  assign new_n18051_ = ~new_n4691_ | ~new_n17654_;
  assign new_n18052_ = ~new_n5591_ | ~new_n17655_;
  assign new_n18053_ = ~new_n18052_ | ~new_n18051_;
  assign new_n18054_ = ~new_n4692_ | ~new_n17681_;
  assign new_n18055_ = ~new_n5592_ | ~new_n17690_;
  assign new_n18056_ = ~new_n17782_ | ~new_n17761_;
  assign new_n18057_ = ~new_n17928_ | ~new_n17631_;
  assign new_n18058_ = ~new_n4697_ | ~new_n17678_;
  assign new_n18059_ = ~new_n5122_ | ~new_n17679_;
  assign new_n18060_ = ~new_n18059_ | ~new_n18058_;
  assign new_n18061_ = ~new_n17959_ | ~new_n17691_;
  assign new_n18062_ = ~new_n18060_ | ~new_n17916_;
  assign new_n18063_ = ~new_n4698_ | ~new_n17675_;
  assign new_n18064_ = ~new_n5120_ | ~new_n17676_;
  assign new_n18065_ = ~new_n18064_ | ~new_n18063_;
  assign new_n18066_ = ~new_n17960_ | ~new_n17762_;
  assign new_n18067_ = ~new_n17870_ | ~new_n18065_;
  assign new_n18068_ = ~new_n4685_ | ~new_n17660_;
  assign new_n18069_ = ~new_n5117_ | ~new_n17658_;
  assign new_n18070_ = ~new_n4689_ | ~new_n17656_;
  assign new_n18071_ = ~new_n5114_ | ~new_n17657_;
  assign new_n18072_ = ~new_n18071_ | ~new_n18070_;
  assign new_n18073_ = ~new_n17961_ | ~new_n17692_;
  assign new_n18074_ = ~new_n18072_ | ~new_n17862_;
  assign new_n18075_ = ~new_n4690_ | ~new_n17673_;
  assign new_n18076_ = ~new_n5111_ | ~new_n17674_;
  assign new_n18077_ = ~new_n4690_ | ~new_n17673_;
  assign new_n18078_ = ~new_n5111_ | ~new_n17674_;
  assign new_n18079_ = ~new_n18078_ | ~new_n18077_;
  assign new_n18080_ = ~new_n17763_ | ~new_n17764_;
  assign new_n18081_ = ~new_n17858_ | ~new_n18079_;
  assign new_n18082_ = ~new_n4695_ | ~new_n17671_;
  assign new_n18083_ = ~new_n5108_ | ~new_n17672_;
  assign new_n18084_ = ~new_n4695_ | ~new_n17671_;
  assign new_n18085_ = ~new_n5108_ | ~new_n17672_;
  assign new_n18086_ = ~new_n18085_ | ~new_n18084_;
  assign new_n18087_ = ~new_n17765_ | ~new_n17766_;
  assign new_n18088_ = ~new_n17854_ | ~new_n18086_;
  assign new_n18089_ = ~new_n4696_ | ~new_n17669_;
  assign new_n18090_ = ~new_n5105_ | ~new_n17670_;
  assign new_n18091_ = ~new_n4688_ | ~new_n17664_;
  assign new_n18092_ = ~new_n5102_ | ~new_n17665_;
  assign new_n18093_ = ~new_n18092_ | ~new_n18091_;
  assign new_n18094_ = ~new_n17962_ | ~new_n17693_;
  assign new_n18095_ = ~new_n18093_ | ~new_n17938_;
  assign new_n18096_ = ~new_n4679_ | ~new_n17666_;
  assign new_n18097_ = ~new_n5099_ | ~new_n17667_;
  assign new_n18098_ = ~new_n18097_ | ~new_n18096_;
  assign new_n18099_ = ~new_n17963_ | ~new_n17767_;
  assign new_n18100_ = ~new_n17844_ | ~new_n18098_;
  assign new_n18101_ = ~new_n4678_ | ~new_n17661_;
  assign new_n18102_ = ~new_n5096_ | ~new_n17662_;
  assign new_n18103_ = ~new_n4693_ | ~new_n17629_;
  assign new_n18104_ = ~new_n5064_ | ~new_n17630_;
  assign new_n18105_ = new_n18280_ & new_n18279_;
  assign new_n18106_ = new_n18298_ & new_n18297_;
  assign new_n18107_ = new_n18338_ & new_n18337_;
  assign new_n18108_ = new_n18347_ & new_n18346_;
  assign new_n18109_ = new_n18365_ & new_n18364_;
  assign new_n18110_ = new_n18373_ & new_n18372_;
  assign new_n18111_ = new_n18452_ & new_n18449_;
  assign new_n18112_ = new_n18445_ & new_n18442_;
  assign new_n18113_ = new_n18436_ & new_n18433_;
  assign new_n18114_ = new_n18427_ & new_n18424_;
  assign new_n18115_ = new_n18421_ & new_n18419_;
  assign new_n18116_ = new_n18414_ & new_n18411_;
  assign new_n18117_ = new_n18336_ & new_n18333_;
  assign new_n18118_ = new_n18328_ & new_n18325_;
  assign new_n18119_ = new_n18314_ & new_n18311_;
  assign new_n18120_ = ~new_n5084_;
  assign new_n18121_ = ~new_n4687_;
  assign new_n18122_ = ~new_n4686_;
  assign new_n18123_ = ~new_n4687_ | ~new_n5084_;
  assign new_n18124_ = ~new_n5087_;
  assign new_n18125_ = ~new_n5078_;
  assign new_n18126_ = ~new_n4676_;
  assign new_n18127_ = ~new_n4683_;
  assign new_n18128_ = ~new_n5072_;
  assign new_n18129_ = ~new_n4684_;
  assign new_n18130_ = ~new_n5064_;
  assign new_n18131_ = ~new_n4693_;
  assign new_n18132_ = ~new_n4693_ | ~new_n5064_;
  assign new_n18133_ = ~new_n5075_;
  assign new_n18134_ = ~new_n4680_;
  assign new_n18135_ = ~new_n4676_ | ~new_n5078_;
  assign new_n18136_ = ~new_n5081_;
  assign new_n18137_ = ~new_n5090_;
  assign new_n18138_ = ~new_n4700_;
  assign new_n18139_ = ~new_n4699_;
  assign new_n18140_ = ~new_n5093_;
  assign new_n18141_ = ~new_n18164_ | ~new_n18306_;
  assign new_n18142_ = ~new_n18218_ | ~new_n18294_;
  assign new_n18143_ = ~new_n18283_ | ~new_n18284_;
  assign new_n18144_ = ~new_n5069_ | ~new_n4694_;
  assign new_n18145_ = ~new_n18223_ | ~new_n18320_;
  assign new_n18146_ = ~new_n18317_ | ~new_n18316_;
  assign new_n18147_ = ~new_n5585_;
  assign new_n18148_ = ~new_n4669_;
  assign new_n18149_ = ~new_n4673_;
  assign new_n18150_ = ~new_n5586_;
  assign new_n18151_ = ~new_n5587_;
  assign new_n18152_ = ~new_n4674_;
  assign new_n18153_ = ~new_n5588_;
  assign new_n18154_ = ~new_n4681_;
  assign new_n18155_ = ~new_n5591_;
  assign new_n18156_ = ~new_n4691_;
  assign new_n18157_ = ~new_n5114_;
  assign new_n18158_ = ~new_n4689_;
  assign new_n18159_ = ~new_n4685_;
  assign new_n18160_ = ~new_n4689_ | ~new_n5114_;
  assign new_n18161_ = ~new_n5117_;
  assign new_n18162_ = ~new_n5096_;
  assign new_n18163_ = ~new_n4678_;
  assign new_n18164_ = ~new_n4700_ | ~new_n5090_;
  assign new_n18165_ = ~new_n5102_;
  assign new_n18166_ = ~new_n4688_;
  assign new_n18167_ = ~new_n5099_;
  assign new_n18168_ = ~new_n4679_;
  assign new_n18169_ = ~new_n4679_ | ~new_n5099_;
  assign new_n18170_ = ~new_n5105_;
  assign new_n18171_ = ~new_n4696_;
  assign new_n18172_ = ~new_n5108_;
  assign new_n18173_ = ~new_n4695_;
  assign new_n18174_ = ~new_n5111_;
  assign new_n18175_ = ~new_n4690_;
  assign new_n18176_ = ~new_n5120_;
  assign new_n18177_ = ~new_n4698_;
  assign new_n18178_ = ~new_n4698_ | ~new_n5120_;
  assign new_n18179_ = ~new_n5122_;
  assign new_n18180_ = ~new_n4697_;
  assign new_n18181_ = ~new_n4697_ | ~new_n5122_;
  assign new_n18182_ = ~new_n5592_;
  assign new_n18183_ = ~new_n5590_;
  assign new_n18184_ = ~new_n4677_;
  assign new_n18185_ = ~new_n5589_;
  assign new_n18186_ = ~new_n4682_;
  assign new_n18187_ = ~new_n5586_ | ~new_n4673_;
  assign new_n18188_ = ~new_n4670_;
  assign new_n18189_ = ~new_n5584_;
  assign new_n18190_ = ~new_n18407_ | ~new_n18277_;
  assign new_n18191_ = ~new_n4692_;
  assign new_n18192_ = ~new_n18178_ | ~new_n18416_;
  assign new_n18193_ = ~new_n18362_ | ~new_n18361_;
  assign new_n18194_ = ~new_n18169_ | ~new_n18438_;
  assign new_n18195_ = ~new_n18558_ | ~new_n18557_;
  assign new_n18196_ = ~new_n18605_ | ~new_n18604_;
  assign new_n18197_ = ~new_n18476_ | ~new_n18475_;
  assign new_n18198_ = ~new_n18481_ | ~new_n18480_;
  assign new_n18199_ = ~new_n18488_ | ~new_n18487_;
  assign new_n18200_ = ~new_n18495_ | ~new_n18494_;
  assign new_n18201_ = ~new_n18500_ | ~new_n18499_;
  assign new_n18202_ = ~new_n18509_ | ~new_n18508_;
  assign new_n18203_ = ~new_n18516_ | ~new_n18515_;
  assign new_n18204_ = ~new_n18523_ | ~new_n18522_;
  assign new_n18205_ = ~new_n18530_ | ~new_n18529_;
  assign new_n18206_ = ~new_n18535_ | ~new_n18534_;
  assign new_n18207_ = ~new_n18542_ | ~new_n18541_;
  assign new_n18208_ = ~new_n18549_ | ~new_n18548_;
  assign new_n18209_ = ~new_n18563_ | ~new_n18562_;
  assign new_n18210_ = ~new_n18568_ | ~new_n18567_;
  assign new_n18211_ = ~new_n18575_ | ~new_n18574_;
  assign new_n18212_ = ~new_n18582_ | ~new_n18581_;
  assign new_n18213_ = ~new_n18589_ | ~new_n18588_;
  assign new_n18214_ = ~new_n18596_ | ~new_n18595_;
  assign new_n18215_ = ~new_n18601_ | ~new_n18600_;
  assign new_n18216_ = new_n18290_ & new_n18288_;
  assign new_n18217_ = new_n18105_ & new_n18281_;
  assign new_n18218_ = new_n18295_ & new_n18293_;
  assign new_n18219_ = new_n18302_ & new_n18301_;
  assign new_n18220_ = new_n18123_ & new_n18483_ & new_n18482_;
  assign new_n18221_ = new_n18313_ & new_n18106_;
  assign new_n18222_ = new_n18282_ & new_n18281_;
  assign new_n18223_ = new_n18321_ & new_n18319_;
  assign new_n18224_ = new_n18135_ & new_n18490_ & new_n18489_;
  assign new_n18225_ = new_n18327_ & new_n18105_;
  assign new_n18226_ = new_n18335_ & new_n18282_;
  assign new_n18227_ = new_n18305_ & new_n18107_;
  assign new_n18228_ = new_n18344_ & new_n18340_;
  assign new_n18229_ = new_n18351_ & new_n18108_;
  assign new_n18230_ = new_n18349_ & new_n18273_;
  assign new_n18231_ = new_n18369_ & new_n18368_;
  assign new_n18232_ = new_n18374_ & new_n18110_ & new_n18383_;
  assign new_n18233_ = new_n18386_ & new_n18381_;
  assign new_n18234_ = new_n18402_ & new_n18399_;
  assign new_n18235_ = new_n18469_ & new_n18403_;
  assign new_n18236_ = new_n18274_ & new_n18525_ & new_n18524_;
  assign new_n18237_ = new_n18261_ & new_n18379_;
  assign new_n18238_ = new_n18181_ & new_n18556_ & new_n18555_;
  assign new_n18239_ = new_n18426_ & new_n18110_;
  assign new_n18240_ = new_n18160_ & new_n18570_ & new_n18569_;
  assign new_n18241_ = new_n18435_ & new_n18109_;
  assign new_n18242_ = new_n18273_ & new_n18591_ & new_n18590_;
  assign new_n18243_ = new_n18444_ & new_n18108_;
  assign new_n18244_ = new_n18272_ & new_n18603_ & new_n18602_;
  assign new_n18245_ = new_n18451_ & new_n18107_;
  assign new_n18246_ = ~new_n18219_ | ~new_n18303_;
  assign new_n18247_ = ~new_n18318_ | ~new_n18330_;
  assign new_n18248_ = ~new_n4671_;
  assign new_n18249_ = ~new_n5595_;
  assign new_n18250_ = new_n18504_ & new_n18503_;
  assign new_n18251_ = ~new_n18465_ | ~new_n18405_ | ~new_n18270_;
  assign new_n18252_ = new_n18511_ & new_n18510_;
  assign new_n18253_ = ~new_n18235_ | ~new_n18471_ | ~new_n18470_;
  assign new_n18254_ = new_n18518_ & new_n18517_;
  assign new_n18255_ = ~new_n18187_ | ~new_n18466_ | ~new_n18400_;
  assign new_n18256_ = ~new_n18394_ | ~new_n18393_;
  assign new_n18257_ = new_n18537_ & new_n18536_;
  assign new_n18258_ = ~new_n18390_ | ~new_n18389_;
  assign new_n18259_ = new_n18544_ & new_n18543_;
  assign new_n18260_ = ~new_n18233_ | ~new_n18385_;
  assign new_n18261_ = new_n18551_ & new_n18550_;
  assign new_n18262_ = ~new_n18144_ | ~new_n18428_;
  assign new_n18263_ = ~new_n18231_ | ~new_n18370_;
  assign new_n18264_ = new_n18577_ & new_n18576_;
  assign new_n18265_ = ~new_n18358_ | ~new_n18357_;
  assign new_n18266_ = new_n18584_ & new_n18583_;
  assign new_n18267_ = ~new_n18354_ | ~new_n18353_;
  assign new_n18268_ = ~new_n18228_ | ~new_n18343_;
  assign new_n18269_ = ~new_n18468_ | ~new_n18467_;
  assign new_n18270_ = ~new_n4670_ | ~new_n18253_;
  assign new_n18271_ = ~new_n18135_;
  assign new_n18272_ = ~new_n5093_ | ~new_n4699_;
  assign new_n18273_ = ~new_n4688_ | ~new_n5102_;
  assign new_n18274_ = ~new_n4674_ | ~new_n5587_;
  assign new_n18275_ = ~new_n18169_;
  assign new_n18276_ = ~new_n18178_;
  assign new_n18277_ = ~new_n4681_ | ~new_n5588_;
  assign new_n18278_ = ~new_n18164_;
  assign new_n18279_ = new_n4683_ | new_n5081_;
  assign new_n18280_ = new_n4676_ | new_n5078_;
  assign new_n18281_ = new_n5075_ | new_n4680_;
  assign new_n18282_ = new_n5072_ | new_n4684_;
  assign new_n18283_ = ~new_n18132_;
  assign new_n18284_ = new_n5069_ | new_n4694_;
  assign new_n18285_ = ~new_n18143_;
  assign new_n18286_ = ~new_n18144_;
  assign new_n18287_ = ~new_n18143_ | ~new_n18144_;
  assign new_n18288_ = ~new_n4684_ | ~new_n5072_;
  assign new_n18289_ = ~new_n18287_ | ~new_n18282_;
  assign new_n18290_ = ~new_n4680_ | ~new_n5075_;
  assign new_n18291_ = ~new_n18216_ | ~new_n18289_;
  assign new_n18292_ = ~new_n18136_ | ~new_n18135_;
  assign new_n18293_ = ~new_n4683_ | ~new_n18292_;
  assign new_n18294_ = ~new_n18217_ | ~new_n18291_;
  assign new_n18295_ = ~new_n5081_ | ~new_n18271_;
  assign new_n18296_ = ~new_n18142_;
  assign new_n18297_ = new_n4686_ | new_n5087_;
  assign new_n18298_ = new_n4687_ | new_n5084_;
  assign new_n18299_ = ~new_n18123_;
  assign new_n18300_ = ~new_n18124_ | ~new_n18123_;
  assign new_n18301_ = ~new_n4686_ | ~new_n18300_;
  assign new_n18302_ = ~new_n5087_ | ~new_n18299_;
  assign new_n18303_ = ~new_n18106_ | ~new_n18142_;
  assign new_n18304_ = ~new_n18246_;
  assign new_n18305_ = new_n5090_ | new_n4700_;
  assign new_n18306_ = ~new_n18305_ | ~new_n18246_;
  assign new_n18307_ = ~new_n18141_;
  assign new_n18308_ = new_n4699_ | new_n5093_;
  assign new_n18309_ = new_n5084_ | new_n4687_;
  assign new_n18310_ = ~new_n18309_ | ~new_n18142_;
  assign new_n18311_ = ~new_n18220_ | ~new_n18310_;
  assign new_n18312_ = ~new_n18296_ | ~new_n18123_;
  assign new_n18313_ = ~new_n5087_ | ~new_n4686_;
  assign new_n18314_ = ~new_n18221_ | ~new_n18312_;
  assign new_n18315_ = new_n4687_ | new_n5084_;
  assign new_n18316_ = ~new_n18286_ | ~new_n18282_;
  assign new_n18317_ = ~new_n4684_ | ~new_n5072_;
  assign new_n18318_ = ~new_n18146_;
  assign new_n18319_ = ~new_n18222_ | ~new_n18285_;
  assign new_n18320_ = ~new_n18146_ | ~new_n18281_;
  assign new_n18321_ = ~new_n4680_ | ~new_n5075_;
  assign new_n18322_ = ~new_n18145_;
  assign new_n18323_ = new_n5078_ | new_n4676_;
  assign new_n18324_ = ~new_n18323_ | ~new_n18145_;
  assign new_n18325_ = ~new_n18224_ | ~new_n18324_;
  assign new_n18326_ = ~new_n18322_ | ~new_n18135_;
  assign new_n18327_ = ~new_n5081_ | ~new_n4683_;
  assign new_n18328_ = ~new_n18225_ | ~new_n18326_;
  assign new_n18329_ = new_n4676_ | new_n5078_;
  assign new_n18330_ = ~new_n18285_ | ~new_n18282_;
  assign new_n18331_ = ~new_n18247_;
  assign new_n18332_ = ~new_n4680_ | ~new_n5075_;
  assign new_n18333_ = ~new_n18143_ | ~new_n18144_ | ~new_n18502_ | ~new_n18501_;
  assign new_n18334_ = ~new_n18144_ | ~new_n18143_;
  assign new_n18335_ = ~new_n4684_ | ~new_n5072_;
  assign new_n18336_ = ~new_n18226_ | ~new_n18334_;
  assign new_n18337_ = new_n4699_ | new_n5093_;
  assign new_n18338_ = new_n4678_ | new_n5096_;
  assign new_n18339_ = ~new_n18278_ | ~new_n18107_;
  assign new_n18340_ = ~new_n4678_ | ~new_n5096_;
  assign new_n18341_ = ~new_n18272_ | ~new_n18339_;
  assign new_n18342_ = new_n5096_ | new_n4678_;
  assign new_n18343_ = ~new_n18227_ | ~new_n18246_;
  assign new_n18344_ = ~new_n18342_ | ~new_n18341_;
  assign new_n18345_ = ~new_n18268_;
  assign new_n18346_ = new_n4696_ | new_n5105_;
  assign new_n18347_ = new_n4688_ | new_n5102_;
  assign new_n18348_ = ~new_n18275_ | ~new_n18108_;
  assign new_n18349_ = ~new_n4696_ | ~new_n5105_;
  assign new_n18350_ = ~new_n18230_ | ~new_n18348_;
  assign new_n18351_ = new_n5099_ | new_n4679_;
  assign new_n18352_ = new_n5105_ | new_n4696_;
  assign new_n18353_ = ~new_n18229_ | ~new_n18268_;
  assign new_n18354_ = ~new_n18352_ | ~new_n18350_;
  assign new_n18355_ = ~new_n18267_;
  assign new_n18356_ = new_n5108_ | new_n4695_;
  assign new_n18357_ = ~new_n18356_ | ~new_n18267_;
  assign new_n18358_ = ~new_n4695_ | ~new_n5108_;
  assign new_n18359_ = ~new_n18265_;
  assign new_n18360_ = new_n5111_ | new_n4690_;
  assign new_n18361_ = ~new_n18360_ | ~new_n18265_;
  assign new_n18362_ = ~new_n4690_ | ~new_n5111_;
  assign new_n18363_ = ~new_n18193_;
  assign new_n18364_ = new_n4685_ | new_n5117_;
  assign new_n18365_ = new_n4689_ | new_n5114_;
  assign new_n18366_ = ~new_n18160_;
  assign new_n18367_ = ~new_n18161_ | ~new_n18160_;
  assign new_n18368_ = ~new_n4685_ | ~new_n18367_;
  assign new_n18369_ = ~new_n5117_ | ~new_n18366_;
  assign new_n18370_ = ~new_n18109_ | ~new_n18193_;
  assign new_n18371_ = ~new_n18263_;
  assign new_n18372_ = new_n4692_ | new_n5592_;
  assign new_n18373_ = new_n4697_ | new_n5122_;
  assign new_n18374_ = new_n4691_ | new_n5591_;
  assign new_n18375_ = ~new_n18181_;
  assign new_n18376_ = ~new_n5592_ | ~new_n18375_;
  assign new_n18377_ = ~new_n18376_ | ~new_n18191_;
  assign new_n18378_ = ~new_n18181_ | ~new_n18182_;
  assign new_n18379_ = ~new_n18378_ | ~new_n18377_;
  assign new_n18380_ = ~new_n18276_ | ~new_n18110_;
  assign new_n18381_ = ~new_n4691_ | ~new_n5591_;
  assign new_n18382_ = ~new_n18379_ | ~new_n18380_;
  assign new_n18383_ = new_n5120_ | new_n4698_;
  assign new_n18384_ = new_n5591_ | new_n4691_;
  assign new_n18385_ = ~new_n18263_ | ~new_n18232_;
  assign new_n18386_ = ~new_n18384_ | ~new_n18382_;
  assign new_n18387_ = ~new_n18260_;
  assign new_n18388_ = new_n5590_ | new_n4677_;
  assign new_n18389_ = ~new_n18388_ | ~new_n18260_;
  assign new_n18390_ = ~new_n4677_ | ~new_n5590_;
  assign new_n18391_ = ~new_n18258_;
  assign new_n18392_ = new_n5589_ | new_n4682_;
  assign new_n18393_ = ~new_n18392_ | ~new_n18258_;
  assign new_n18394_ = ~new_n4682_ | ~new_n5589_;
  assign new_n18395_ = ~new_n18256_;
  assign new_n18396_ = new_n4674_ | new_n5587_;
  assign new_n18397_ = ~new_n18277_ | ~new_n18274_;
  assign new_n18398_ = ~new_n18187_;
  assign new_n18399_ = new_n5588_ | new_n4681_;
  assign new_n18400_ = ~new_n18269_ | ~new_n18256_ | ~new_n18399_;
  assign new_n18401_ = ~new_n18255_;
  assign new_n18402_ = new_n5585_ | new_n4669_;
  assign new_n18403_ = ~new_n4669_ | ~new_n5585_;
  assign new_n18404_ = ~new_n18253_;
  assign new_n18405_ = ~new_n5584_ | ~new_n18253_;
  assign new_n18406_ = ~new_n18251_;
  assign new_n18407_ = ~new_n18399_ | ~new_n18256_;
  assign new_n18408_ = ~new_n18190_;
  assign new_n18409_ = new_n5587_ | new_n4674_;
  assign new_n18410_ = ~new_n18409_ | ~new_n18190_;
  assign new_n18411_ = ~new_n18236_ | ~new_n18410_;
  assign new_n18412_ = ~new_n18408_ | ~new_n18274_;
  assign new_n18413_ = ~new_n5586_ | ~new_n4673_;
  assign new_n18414_ = ~new_n18269_ | ~new_n18412_ | ~new_n18413_;
  assign new_n18415_ = new_n4674_ | new_n5587_;
  assign new_n18416_ = ~new_n18383_ | ~new_n18263_;
  assign new_n18417_ = ~new_n18192_;
  assign new_n18418_ = ~new_n18110_ | ~new_n18192_;
  assign new_n18419_ = ~new_n18237_ | ~new_n18418_;
  assign new_n18420_ = ~new_n18418_ | ~new_n18379_;
  assign new_n18421_ = ~new_n18554_ | ~new_n18420_;
  assign new_n18422_ = new_n5122_ | new_n4697_;
  assign new_n18423_ = ~new_n18422_ | ~new_n18192_;
  assign new_n18424_ = ~new_n18238_ | ~new_n18423_;
  assign new_n18425_ = ~new_n18417_ | ~new_n18181_;
  assign new_n18426_ = ~new_n4692_ | ~new_n5592_;
  assign new_n18427_ = ~new_n18239_ | ~new_n18425_;
  assign new_n18428_ = new_n5069_ | new_n4694_;
  assign new_n18429_ = ~new_n18262_;
  assign new_n18430_ = new_n4697_ | new_n5122_;
  assign new_n18431_ = new_n5114_ | new_n4689_;
  assign new_n18432_ = ~new_n18431_ | ~new_n18193_;
  assign new_n18433_ = ~new_n18240_ | ~new_n18432_;
  assign new_n18434_ = ~new_n18363_ | ~new_n18160_;
  assign new_n18435_ = ~new_n5117_ | ~new_n4685_;
  assign new_n18436_ = ~new_n18241_ | ~new_n18434_;
  assign new_n18437_ = new_n4689_ | new_n5114_;
  assign new_n18438_ = ~new_n18351_ | ~new_n18268_;
  assign new_n18439_ = ~new_n18194_;
  assign new_n18440_ = new_n5102_ | new_n4688_;
  assign new_n18441_ = ~new_n18440_ | ~new_n18194_;
  assign new_n18442_ = ~new_n18242_ | ~new_n18441_;
  assign new_n18443_ = ~new_n18439_ | ~new_n18273_;
  assign new_n18444_ = ~new_n4696_ | ~new_n5105_;
  assign new_n18445_ = ~new_n18243_ | ~new_n18443_;
  assign new_n18446_ = new_n4688_ | new_n5102_;
  assign new_n18447_ = new_n5093_ | new_n4699_;
  assign new_n18448_ = ~new_n18447_ | ~new_n18141_;
  assign new_n18449_ = ~new_n18244_ | ~new_n18448_;
  assign new_n18450_ = ~new_n18307_ | ~new_n18272_;
  assign new_n18451_ = ~new_n4678_ | ~new_n5096_;
  assign new_n18452_ = ~new_n18245_ | ~new_n18450_;
  assign new_n18453_ = ~new_n18308_ | ~new_n18272_;
  assign new_n18454_ = ~new_n18305_ | ~new_n18164_;
  assign new_n18455_ = ~new_n18315_ | ~new_n18123_;
  assign new_n18456_ = ~new_n18329_ | ~new_n18135_;
  assign new_n18457_ = ~new_n18332_ | ~new_n18281_;
  assign new_n18458_ = ~new_n18415_ | ~new_n18274_;
  assign new_n18459_ = ~new_n18399_ | ~new_n18277_;
  assign new_n18460_ = ~new_n18430_ | ~new_n18181_;
  assign new_n18461_ = ~new_n18383_ | ~new_n18178_;
  assign new_n18462_ = ~new_n18437_ | ~new_n18160_;
  assign new_n18463_ = ~new_n18446_ | ~new_n18273_;
  assign new_n18464_ = ~new_n18351_ | ~new_n18169_;
  assign new_n18465_ = ~new_n5584_ | ~new_n4670_;
  assign new_n18466_ = ~new_n18397_ | ~new_n18269_;
  assign new_n18467_ = ~new_n4673_ | ~new_n18396_;
  assign new_n18468_ = ~new_n5586_ | ~new_n18396_;
  assign new_n18469_ = ~new_n18402_ | ~new_n18397_ | ~new_n18269_;
  assign new_n18470_ = ~new_n18234_ | ~new_n18256_ | ~new_n18269_;
  assign new_n18471_ = ~new_n18398_ | ~new_n18402_;
  assign new_n18472_ = ~new_n4699_ | ~new_n18140_;
  assign new_n18473_ = ~new_n5093_ | ~new_n18139_;
  assign new_n18474_ = ~new_n18473_ | ~new_n18472_;
  assign new_n18475_ = ~new_n18453_ | ~new_n18141_;
  assign new_n18476_ = ~new_n18474_ | ~new_n18307_;
  assign new_n18477_ = ~new_n4700_ | ~new_n18137_;
  assign new_n18478_ = ~new_n5090_ | ~new_n18138_;
  assign new_n18479_ = ~new_n18478_ | ~new_n18477_;
  assign new_n18480_ = ~new_n18454_ | ~new_n18246_;
  assign new_n18481_ = ~new_n18304_ | ~new_n18479_;
  assign new_n18482_ = ~new_n4686_ | ~new_n18124_;
  assign new_n18483_ = ~new_n5087_ | ~new_n18122_;
  assign new_n18484_ = ~new_n4687_ | ~new_n18120_;
  assign new_n18485_ = ~new_n5084_ | ~new_n18121_;
  assign new_n18486_ = ~new_n18485_ | ~new_n18484_;
  assign new_n18487_ = ~new_n18455_ | ~new_n18142_;
  assign new_n18488_ = ~new_n18486_ | ~new_n18296_;
  assign new_n18489_ = ~new_n4683_ | ~new_n18136_;
  assign new_n18490_ = ~new_n5081_ | ~new_n18127_;
  assign new_n18491_ = ~new_n4676_ | ~new_n18125_;
  assign new_n18492_ = ~new_n5078_ | ~new_n18126_;
  assign new_n18493_ = ~new_n18492_ | ~new_n18491_;
  assign new_n18494_ = ~new_n18456_ | ~new_n18145_;
  assign new_n18495_ = ~new_n18493_ | ~new_n18322_;
  assign new_n18496_ = ~new_n4680_ | ~new_n18133_;
  assign new_n18497_ = ~new_n5075_ | ~new_n18134_;
  assign new_n18498_ = ~new_n18497_ | ~new_n18496_;
  assign new_n18499_ = ~new_n18457_ | ~new_n18247_;
  assign new_n18500_ = ~new_n18331_ | ~new_n18498_;
  assign new_n18501_ = ~new_n4684_ | ~new_n18128_;
  assign new_n18502_ = ~new_n5072_ | ~new_n18129_;
  assign new_n18503_ = ~new_n4671_ | ~new_n18249_;
  assign new_n18504_ = ~new_n5595_ | ~new_n18248_;
  assign new_n18505_ = ~new_n4671_ | ~new_n18249_;
  assign new_n18506_ = ~new_n5595_ | ~new_n18248_;
  assign new_n18507_ = ~new_n18506_ | ~new_n18505_;
  assign new_n18508_ = ~new_n18250_ | ~new_n18251_;
  assign new_n18509_ = ~new_n18406_ | ~new_n18507_;
  assign new_n18510_ = ~new_n4670_ | ~new_n18189_;
  assign new_n18511_ = ~new_n5584_ | ~new_n18188_;
  assign new_n18512_ = ~new_n4670_ | ~new_n18189_;
  assign new_n18513_ = ~new_n5584_ | ~new_n18188_;
  assign new_n18514_ = ~new_n18513_ | ~new_n18512_;
  assign new_n18515_ = ~new_n18252_ | ~new_n18253_;
  assign new_n18516_ = ~new_n18404_ | ~new_n18514_;
  assign new_n18517_ = ~new_n4669_ | ~new_n18147_;
  assign new_n18518_ = ~new_n5585_ | ~new_n18148_;
  assign new_n18519_ = ~new_n4669_ | ~new_n18147_;
  assign new_n18520_ = ~new_n5585_ | ~new_n18148_;
  assign new_n18521_ = ~new_n18520_ | ~new_n18519_;
  assign new_n18522_ = ~new_n18254_ | ~new_n18255_;
  assign new_n18523_ = ~new_n18401_ | ~new_n18521_;
  assign new_n18524_ = ~new_n4673_ | ~new_n18150_;
  assign new_n18525_ = ~new_n5586_ | ~new_n18149_;
  assign new_n18526_ = ~new_n4674_ | ~new_n18151_;
  assign new_n18527_ = ~new_n5587_ | ~new_n18152_;
  assign new_n18528_ = ~new_n18527_ | ~new_n18526_;
  assign new_n18529_ = ~new_n18458_ | ~new_n18190_;
  assign new_n18530_ = ~new_n18528_ | ~new_n18408_;
  assign new_n18531_ = ~new_n4681_ | ~new_n18153_;
  assign new_n18532_ = ~new_n5588_ | ~new_n18154_;
  assign new_n18533_ = ~new_n18532_ | ~new_n18531_;
  assign new_n18534_ = ~new_n18459_ | ~new_n18256_;
  assign new_n18535_ = ~new_n18395_ | ~new_n18533_;
  assign new_n18536_ = ~new_n4682_ | ~new_n18185_;
  assign new_n18537_ = ~new_n5589_ | ~new_n18186_;
  assign new_n18538_ = ~new_n4682_ | ~new_n18185_;
  assign new_n18539_ = ~new_n5589_ | ~new_n18186_;
  assign new_n18540_ = ~new_n18539_ | ~new_n18538_;
  assign new_n18541_ = ~new_n18257_ | ~new_n18258_;
  assign new_n18542_ = ~new_n18391_ | ~new_n18540_;
  assign new_n18543_ = ~new_n4677_ | ~new_n18183_;
  assign new_n18544_ = ~new_n5590_ | ~new_n18184_;
  assign new_n18545_ = ~new_n4677_ | ~new_n18183_;
  assign new_n18546_ = ~new_n5590_ | ~new_n18184_;
  assign new_n18547_ = ~new_n18546_ | ~new_n18545_;
  assign new_n18548_ = ~new_n18259_ | ~new_n18260_;
  assign new_n18549_ = ~new_n18387_ | ~new_n18547_;
  assign new_n18550_ = ~new_n4691_ | ~new_n18155_;
  assign new_n18551_ = ~new_n5591_ | ~new_n18156_;
  assign new_n18552_ = ~new_n4691_ | ~new_n18155_;
  assign new_n18553_ = ~new_n5591_ | ~new_n18156_;
  assign new_n18554_ = ~new_n18553_ | ~new_n18552_;
  assign new_n18555_ = ~new_n4692_ | ~new_n18182_;
  assign new_n18556_ = ~new_n5592_ | ~new_n18191_;
  assign new_n18557_ = ~new_n18283_ | ~new_n18262_;
  assign new_n18558_ = ~new_n18429_ | ~new_n18132_;
  assign new_n18559_ = ~new_n4697_ | ~new_n18179_;
  assign new_n18560_ = ~new_n5122_ | ~new_n18180_;
  assign new_n18561_ = ~new_n18560_ | ~new_n18559_;
  assign new_n18562_ = ~new_n18460_ | ~new_n18192_;
  assign new_n18563_ = ~new_n18561_ | ~new_n18417_;
  assign new_n18564_ = ~new_n4698_ | ~new_n18176_;
  assign new_n18565_ = ~new_n5120_ | ~new_n18177_;
  assign new_n18566_ = ~new_n18565_ | ~new_n18564_;
  assign new_n18567_ = ~new_n18461_ | ~new_n18263_;
  assign new_n18568_ = ~new_n18371_ | ~new_n18566_;
  assign new_n18569_ = ~new_n4685_ | ~new_n18161_;
  assign new_n18570_ = ~new_n5117_ | ~new_n18159_;
  assign new_n18571_ = ~new_n4689_ | ~new_n18157_;
  assign new_n18572_ = ~new_n5114_ | ~new_n18158_;
  assign new_n18573_ = ~new_n18572_ | ~new_n18571_;
  assign new_n18574_ = ~new_n18462_ | ~new_n18193_;
  assign new_n18575_ = ~new_n18573_ | ~new_n18363_;
  assign new_n18576_ = ~new_n4690_ | ~new_n18174_;
  assign new_n18577_ = ~new_n5111_ | ~new_n18175_;
  assign new_n18578_ = ~new_n4690_ | ~new_n18174_;
  assign new_n18579_ = ~new_n5111_ | ~new_n18175_;
  assign new_n18580_ = ~new_n18579_ | ~new_n18578_;
  assign new_n18581_ = ~new_n18264_ | ~new_n18265_;
  assign new_n18582_ = ~new_n18359_ | ~new_n18580_;
  assign new_n18583_ = ~new_n4695_ | ~new_n18172_;
  assign new_n18584_ = ~new_n5108_ | ~new_n18173_;
  assign new_n18585_ = ~new_n4695_ | ~new_n18172_;
  assign new_n18586_ = ~new_n5108_ | ~new_n18173_;
  assign new_n18587_ = ~new_n18586_ | ~new_n18585_;
  assign new_n18588_ = ~new_n18266_ | ~new_n18267_;
  assign new_n18589_ = ~new_n18355_ | ~new_n18587_;
  assign new_n18590_ = ~new_n4696_ | ~new_n18170_;
  assign new_n18591_ = ~new_n5105_ | ~new_n18171_;
  assign new_n18592_ = ~new_n4688_ | ~new_n18165_;
  assign new_n18593_ = ~new_n5102_ | ~new_n18166_;
  assign new_n18594_ = ~new_n18593_ | ~new_n18592_;
  assign new_n18595_ = ~new_n18463_ | ~new_n18194_;
  assign new_n18596_ = ~new_n18594_ | ~new_n18439_;
  assign new_n18597_ = ~new_n4679_ | ~new_n18167_;
  assign new_n18598_ = ~new_n5099_ | ~new_n18168_;
  assign new_n18599_ = ~new_n18598_ | ~new_n18597_;
  assign new_n18600_ = ~new_n18464_ | ~new_n18268_;
  assign new_n18601_ = ~new_n18345_ | ~new_n18599_;
  assign new_n18602_ = ~new_n4678_ | ~new_n18162_;
  assign new_n18603_ = ~new_n5096_ | ~new_n18163_;
  assign new_n18604_ = ~new_n4693_ | ~new_n18130_;
  assign new_n18605_ = ~new_n5064_ | ~new_n18131_;
  assign new_n18606_ = new_n18813_ & new_n18812_;
  assign new_n18607_ = new_n18826_ & new_n18825_;
  assign new_n18608_ = new_n18858_ & new_n18857_;
  assign new_n18609_ = new_n18876_ & new_n18875_;
  assign new_n18610_ = new_n18888_ & new_n18887_;
  assign new_n18611_ = new_n18946_ & new_n18943_;
  assign new_n18612_ = new_n18937_ & new_n18934_;
  assign new_n18613_ = new_n18930_ & new_n18927_;
  assign new_n18614_ = new_n18921_ & new_n18918_;
  assign new_n18615_ = new_n18849_ & new_n18846_;
  assign new_n18616_ = new_n18842_ & new_n18839_;
  assign new_n18617_ = ~new_n4830_;
  assign new_n18618_ = ~new_n4823_;
  assign new_n18619_ = ~new_n4823_ | ~new_n18658_;
  assign new_n18620_ = ~new_n4822_;
  assign new_n18621_ = ~new_n4827_;
  assign new_n18622_ = ~new_n4827_ | ~new_n18660_;
  assign new_n18623_ = ~new_n4826_;
  assign new_n18624_ = ~new_n4829_;
  assign new_n18625_ = ~new_n4828_;
  assign new_n18626_ = ~new_n4825_;
  assign new_n18627_ = ~new_n4824_;
  assign new_n18628_ = ~new_n4821_;
  assign new_n18629_ = ~new_n4820_;
  assign new_n18630_ = ~new_n18823_ | ~new_n18822_;
  assign new_n18631_ = ~new_n18810_ | ~new_n18809_;
  assign new_n18632_ = ~new_n4802_;
  assign new_n18633_ = ~new_n4803_;
  assign new_n18634_ = ~new_n4804_;
  assign new_n18635_ = ~new_n4805_;
  assign new_n18636_ = ~new_n4813_;
  assign new_n18637_ = ~new_n4813_ | ~new_n18671_;
  assign new_n18638_ = ~new_n4812_;
  assign new_n18639_ = ~new_n4819_;
  assign new_n18640_ = ~new_n4817_;
  assign new_n18641_ = ~new_n4818_;
  assign new_n18642_ = ~new_n4818_ | ~new_n18674_;
  assign new_n18643_ = ~new_n4816_;
  assign new_n18644_ = ~new_n4815_;
  assign new_n18645_ = ~new_n4814_;
  assign new_n18646_ = ~new_n4811_;
  assign new_n18647_ = ~new_n4809_;
  assign new_n18648_ = ~new_n4810_;
  assign new_n18649_ = ~new_n4810_ | ~new_n18680_;
  assign new_n18650_ = ~new_n4808_;
  assign new_n18651_ = ~new_n4807_;
  assign new_n18652_ = ~new_n4806_;
  assign new_n18653_ = ~new_n4803_ | ~new_n18669_;
  assign new_n18654_ = ~new_n18649_ | ~new_n18923_;
  assign new_n18655_ = ~new_n18873_ | ~new_n18872_;
  assign new_n18656_ = ~new_n18642_ | ~new_n18939_;
  assign new_n18657_ = ~new_n18968_ | ~new_n18967_;
  assign new_n18658_ = ~new_n18997_ | ~new_n18996_;
  assign new_n18659_ = ~new_n18994_ | ~new_n18993_;
  assign new_n18660_ = ~new_n18988_ | ~new_n18987_;
  assign new_n18661_ = ~new_n18985_ | ~new_n18984_;
  assign new_n18662_ = ~new_n18979_ | ~new_n18978_;
  assign new_n18663_ = ~new_n18982_ | ~new_n18981_;
  assign new_n18664_ = ~new_n18976_ | ~new_n18975_;
  assign new_n18665_ = ~new_n18991_ | ~new_n18990_;
  assign new_n18666_ = ~new_n19000_ | ~new_n18999_;
  assign new_n18667_ = ~new_n19040_ | ~new_n19039_;
  assign new_n18668_ = ~new_n19085_ | ~new_n19084_;
  assign new_n18669_ = ~new_n19088_ | ~new_n19087_;
  assign new_n18670_ = ~new_n19091_ | ~new_n19090_;
  assign new_n18671_ = ~new_n19064_ | ~new_n19063_;
  assign new_n18672_ = ~new_n19061_ | ~new_n19060_;
  assign new_n18673_ = ~new_n19043_ | ~new_n19042_;
  assign new_n18674_ = ~new_n19052_ | ~new_n19051_;
  assign new_n18675_ = ~new_n19046_ | ~new_n19045_;
  assign new_n18676_ = ~new_n19049_ | ~new_n19048_;
  assign new_n18677_ = ~new_n19055_ | ~new_n19054_;
  assign new_n18678_ = ~new_n19058_ | ~new_n19057_;
  assign new_n18679_ = ~new_n19067_ | ~new_n19066_;
  assign new_n18680_ = ~new_n19076_ | ~new_n19075_;
  assign new_n18681_ = ~new_n19070_ | ~new_n19069_;
  assign new_n18682_ = ~new_n19073_ | ~new_n19072_;
  assign new_n18683_ = ~new_n19079_ | ~new_n19078_;
  assign new_n18684_ = ~new_n19082_ | ~new_n19081_;
  assign new_n18685_ = ~new_n19097_ | ~new_n19096_;
  assign new_n18686_ = ~new_n19204_ | ~new_n19203_;
  assign new_n18687_ = ~new_n19003_ | ~new_n19002_;
  assign new_n18688_ = ~new_n19010_ | ~new_n19009_;
  assign new_n18689_ = ~new_n19017_ | ~new_n19016_;
  assign new_n18690_ = ~new_n19024_ | ~new_n19023_;
  assign new_n18691_ = ~new_n19031_ | ~new_n19030_;
  assign new_n18692_ = ~new_n19038_ | ~new_n19037_;
  assign new_n18693_ = ~new_n19100_ | ~new_n19099_;
  assign new_n18694_ = ~new_n19107_ | ~new_n19106_;
  assign new_n18695_ = ~new_n19114_ | ~new_n19113_;
  assign new_n18696_ = ~new_n19119_ | ~new_n19118_;
  assign new_n18697_ = ~new_n19126_ | ~new_n19125_;
  assign new_n18698_ = ~new_n19133_ | ~new_n19132_;
  assign new_n18699_ = ~new_n19140_ | ~new_n19139_;
  assign new_n18700_ = ~new_n19147_ | ~new_n19146_;
  assign new_n18701_ = ~new_n19152_ | ~new_n19151_;
  assign new_n18702_ = ~new_n19159_ | ~new_n19158_;
  assign new_n18703_ = ~new_n19166_ | ~new_n19165_;
  assign new_n18704_ = ~new_n19173_ | ~new_n19172_;
  assign new_n18705_ = ~new_n19180_ | ~new_n19179_;
  assign new_n18706_ = ~new_n19187_ | ~new_n19186_;
  assign new_n18707_ = ~new_n19192_ | ~new_n19191_;
  assign new_n18708_ = ~new_n19199_ | ~new_n19198_;
  assign new_n18709_ = new_n18816_ & new_n18815_;
  assign new_n18710_ = new_n18830_ & new_n18829_;
  assign new_n18711_ = new_n18619_ & new_n19012_ & new_n19011_;
  assign new_n18712_ = new_n18841_ & new_n18607_;
  assign new_n18713_ = new_n18622_ & new_n19033_ & new_n19032_;
  assign new_n18714_ = new_n18848_ & new_n18606_;
  assign new_n18715_ = new_n18862_ & new_n18608_;
  assign new_n18716_ = new_n18860_ & new_n18798_;
  assign new_n18717_ = new_n18880_ & new_n18879_;
  assign new_n18718_ = new_n18892_ & new_n18610_;
  assign new_n18719_ = new_n18890_ & new_n18799_;
  assign new_n18720_ = new_n18908_ & new_n18794_;
  assign new_n18721_ = new_n18966_ & new_n18653_;
  assign new_n18722_ = new_n18913_ & new_n18908_;
  assign new_n18723_ = new_n18963_ & new_n18912_;
  assign new_n18724_ = ~new_n19094_ | ~new_n19093_;
  assign new_n18725_ = new_n18959_ & new_n18653_;
  assign new_n18726_ = new_n18800_ & new_n19109_ & new_n19108_;
  assign new_n18727_ = new_n18803_ & new_n18800_;
  assign new_n18728_ = new_n18920_ & new_n18794_;
  assign new_n18729_ = new_n18799_ & new_n19135_ & new_n19134_;
  assign new_n18730_ = new_n18929_ & new_n18610_;
  assign new_n18731_ = new_n18637_ & new_n19161_ & new_n19160_;
  assign new_n18732_ = new_n18936_ & new_n18609_;
  assign new_n18733_ = new_n18798_ & new_n19182_ & new_n19181_;
  assign new_n18734_ = new_n18945_ & new_n18608_;
  assign new_n18735_ = ~new_n19201_ | ~new_n19200_;
  assign new_n18736_ = ~new_n5093_;
  assign new_n18737_ = new_n18971_ & new_n18970_;
  assign new_n18738_ = ~new_n5078_;
  assign new_n18739_ = ~new_n5064_;
  assign new_n18740_ = ~new_n5069_;
  assign new_n18741_ = ~new_n5075_;
  assign new_n18742_ = ~new_n5072_;
  assign new_n18743_ = ~new_n5081_;
  assign new_n18744_ = ~new_n5087_;
  assign new_n18745_ = ~new_n5084_;
  assign new_n18746_ = ~new_n5090_;
  assign new_n18747_ = ~new_n18835_ | ~new_n18834_;
  assign new_n18748_ = new_n19005_ & new_n19004_;
  assign new_n18749_ = ~new_n18710_ | ~new_n18831_;
  assign new_n18750_ = new_n19019_ & new_n19018_;
  assign new_n18751_ = ~new_n18957_ | ~new_n18819_ | ~new_n18796_;
  assign new_n18752_ = new_n19026_ & new_n19025_;
  assign new_n18753_ = ~new_n18709_ | ~new_n18817_;
  assign new_n18754_ = ~new_n5585_;
  assign new_n18755_ = ~new_n5096_;
  assign new_n18756_ = ~new_n5105_;
  assign new_n18757_ = ~new_n5102_;
  assign new_n18758_ = ~new_n5099_;
  assign new_n18759_ = ~new_n5108_;
  assign new_n18760_ = ~new_n5111_;
  assign new_n18761_ = ~new_n5117_;
  assign new_n18762_ = ~new_n5114_;
  assign new_n18763_ = ~new_n5120_;
  assign new_n18764_ = ~new_n5591_;
  assign new_n18765_ = ~new_n5592_;
  assign new_n18766_ = ~new_n5122_;
  assign new_n18767_ = ~new_n5590_;
  assign new_n18768_ = ~new_n5589_;
  assign new_n18769_ = ~new_n5587_;
  assign new_n18770_ = ~new_n5586_;
  assign new_n18771_ = ~new_n5588_;
  assign new_n18772_ = ~new_n4801_;
  assign new_n18773_ = ~new_n5584_;
  assign new_n18774_ = new_n19102_ & new_n19101_;
  assign new_n18775_ = ~new_n18725_ | ~new_n18909_;
  assign new_n18776_ = ~new_n18803_ | ~new_n18914_;
  assign new_n18777_ = ~new_n18903_ | ~new_n18902_;
  assign new_n18778_ = new_n19121_ & new_n19120_;
  assign new_n18779_ = ~new_n18899_ | ~new_n18898_;
  assign new_n18780_ = new_n19128_ & new_n19127_;
  assign new_n18781_ = ~new_n18895_ | ~new_n18894_;
  assign new_n18782_ = new_n19142_ & new_n19141_;
  assign new_n18783_ = ~new_n18806_ | ~new_n18805_;
  assign new_n18784_ = ~new_n18885_ | ~new_n18884_;
  assign new_n18785_ = new_n19154_ & new_n19153_;
  assign new_n18786_ = ~new_n18717_ | ~new_n18881_;
  assign new_n18787_ = new_n19168_ & new_n19167_;
  assign new_n18788_ = ~new_n18869_ | ~new_n18868_;
  assign new_n18789_ = new_n19175_ & new_n19174_;
  assign new_n18790_ = ~new_n18865_ | ~new_n18864_;
  assign new_n18791_ = ~new_n18855_ | ~new_n18854_;
  assign new_n18792_ = new_n19194_ & new_n19193_;
  assign new_n18793_ = ~new_n18962_ | ~new_n18851_ | ~new_n18795_;
  assign new_n18794_ = ~new_n18961_ | ~new_n18960_;
  assign new_n18795_ = ~new_n18657_ | ~new_n18747_;
  assign new_n18796_ = ~new_n18664_ | ~new_n18753_;
  assign new_n18797_ = ~new_n18622_;
  assign new_n18798_ = ~new_n4817_ | ~new_n18676_;
  assign new_n18799_ = ~new_n4809_ | ~new_n18682_;
  assign new_n18800_ = ~new_n4804_ | ~new_n18668_;
  assign new_n18801_ = ~new_n18642_;
  assign new_n18802_ = ~new_n18649_;
  assign new_n18803_ = ~new_n4805_ | ~new_n18670_;
  assign new_n18804_ = ~new_n18980_ | ~new_n18617_;
  assign new_n18805_ = ~new_n4829_ | ~new_n18804_;
  assign new_n18806_ = ~new_n4830_ | ~new_n18662_;
  assign new_n18807_ = ~new_n18783_;
  assign new_n18808_ = ~new_n18983_ | ~new_n18625_;
  assign new_n18809_ = ~new_n18808_ | ~new_n18783_;
  assign new_n18810_ = ~new_n4828_ | ~new_n18663_;
  assign new_n18811_ = ~new_n18631_;
  assign new_n18812_ = ~new_n18986_ | ~new_n18623_;
  assign new_n18813_ = ~new_n18989_ | ~new_n18621_;
  assign new_n18814_ = ~new_n18623_ | ~new_n18622_;
  assign new_n18815_ = ~new_n18661_ | ~new_n18814_;
  assign new_n18816_ = ~new_n4826_ | ~new_n18797_;
  assign new_n18817_ = ~new_n18606_ | ~new_n18631_;
  assign new_n18818_ = ~new_n18753_;
  assign new_n18819_ = ~new_n4825_ | ~new_n18753_;
  assign new_n18820_ = ~new_n18751_;
  assign new_n18821_ = ~new_n18992_ | ~new_n18627_;
  assign new_n18822_ = ~new_n18821_ | ~new_n18751_;
  assign new_n18823_ = ~new_n4824_ | ~new_n18665_;
  assign new_n18824_ = ~new_n18630_;
  assign new_n18825_ = ~new_n18995_ | ~new_n18620_;
  assign new_n18826_ = ~new_n18998_ | ~new_n18618_;
  assign new_n18827_ = ~new_n18619_;
  assign new_n18828_ = ~new_n18620_ | ~new_n18619_;
  assign new_n18829_ = ~new_n18659_ | ~new_n18828_;
  assign new_n18830_ = ~new_n4822_ | ~new_n18827_;
  assign new_n18831_ = ~new_n18607_ | ~new_n18630_;
  assign new_n18832_ = ~new_n18749_;
  assign new_n18833_ = ~new_n19001_ | ~new_n18628_;
  assign new_n18834_ = ~new_n18833_ | ~new_n18749_;
  assign new_n18835_ = ~new_n4821_ | ~new_n18666_;
  assign new_n18836_ = ~new_n18747_;
  assign new_n18837_ = ~new_n18998_ | ~new_n18618_;
  assign new_n18838_ = ~new_n18837_ | ~new_n18630_;
  assign new_n18839_ = ~new_n18711_ | ~new_n18838_;
  assign new_n18840_ = ~new_n18824_ | ~new_n18619_;
  assign new_n18841_ = ~new_n4822_ | ~new_n18659_;
  assign new_n18842_ = ~new_n18712_ | ~new_n18840_;
  assign new_n18843_ = ~new_n18998_ | ~new_n18618_;
  assign new_n18844_ = ~new_n18989_ | ~new_n18621_;
  assign new_n18845_ = ~new_n18844_ | ~new_n18631_;
  assign new_n18846_ = ~new_n18713_ | ~new_n18845_;
  assign new_n18847_ = ~new_n18811_ | ~new_n18622_;
  assign new_n18848_ = ~new_n4826_ | ~new_n18661_;
  assign new_n18849_ = ~new_n18714_ | ~new_n18847_;
  assign new_n18850_ = ~new_n18989_ | ~new_n18621_;
  assign new_n18851_ = ~new_n4820_ | ~new_n18747_;
  assign new_n18852_ = ~new_n18793_;
  assign new_n18853_ = ~new_n19044_ | ~new_n18639_;
  assign new_n18854_ = ~new_n18853_ | ~new_n18793_;
  assign new_n18855_ = ~new_n4819_ | ~new_n18673_;
  assign new_n18856_ = ~new_n18791_;
  assign new_n18857_ = ~new_n19047_ | ~new_n18643_;
  assign new_n18858_ = ~new_n19050_ | ~new_n18640_;
  assign new_n18859_ = ~new_n18801_ | ~new_n18608_;
  assign new_n18860_ = ~new_n4816_ | ~new_n18675_;
  assign new_n18861_ = ~new_n18716_ | ~new_n18859_;
  assign new_n18862_ = ~new_n19053_ | ~new_n18641_;
  assign new_n18863_ = ~new_n19047_ | ~new_n18643_;
  assign new_n18864_ = ~new_n18715_ | ~new_n18791_;
  assign new_n18865_ = ~new_n18863_ | ~new_n18861_;
  assign new_n18866_ = ~new_n18790_;
  assign new_n18867_ = ~new_n19056_ | ~new_n18644_;
  assign new_n18868_ = ~new_n18867_ | ~new_n18790_;
  assign new_n18869_ = ~new_n4815_ | ~new_n18677_;
  assign new_n18870_ = ~new_n18788_;
  assign new_n18871_ = ~new_n19059_ | ~new_n18645_;
  assign new_n18872_ = ~new_n18871_ | ~new_n18788_;
  assign new_n18873_ = ~new_n4814_ | ~new_n18678_;
  assign new_n18874_ = ~new_n18655_;
  assign new_n18875_ = ~new_n19062_ | ~new_n18638_;
  assign new_n18876_ = ~new_n19065_ | ~new_n18636_;
  assign new_n18877_ = ~new_n18637_;
  assign new_n18878_ = ~new_n18638_ | ~new_n18637_;
  assign new_n18879_ = ~new_n18672_ | ~new_n18878_;
  assign new_n18880_ = ~new_n4812_ | ~new_n18877_;
  assign new_n18881_ = ~new_n18609_ | ~new_n18655_;
  assign new_n18882_ = ~new_n18786_;
  assign new_n18883_ = ~new_n19068_ | ~new_n18646_;
  assign new_n18884_ = ~new_n18883_ | ~new_n18786_;
  assign new_n18885_ = ~new_n4811_ | ~new_n18679_;
  assign new_n18886_ = ~new_n18784_;
  assign new_n18887_ = ~new_n19071_ | ~new_n18650_;
  assign new_n18888_ = ~new_n19074_ | ~new_n18647_;
  assign new_n18889_ = ~new_n18802_ | ~new_n18610_;
  assign new_n18890_ = ~new_n4808_ | ~new_n18681_;
  assign new_n18891_ = ~new_n18719_ | ~new_n18889_;
  assign new_n18892_ = ~new_n19077_ | ~new_n18648_;
  assign new_n18893_ = ~new_n19071_ | ~new_n18650_;
  assign new_n18894_ = ~new_n18718_ | ~new_n18784_;
  assign new_n18895_ = ~new_n18893_ | ~new_n18891_;
  assign new_n18896_ = ~new_n18781_;
  assign new_n18897_ = ~new_n19080_ | ~new_n18651_;
  assign new_n18898_ = ~new_n18897_ | ~new_n18781_;
  assign new_n18899_ = ~new_n4807_ | ~new_n18683_;
  assign new_n18900_ = ~new_n18779_;
  assign new_n18901_ = ~new_n19083_ | ~new_n18652_;
  assign new_n18902_ = ~new_n18901_ | ~new_n18779_;
  assign new_n18903_ = ~new_n4806_ | ~new_n18684_;
  assign new_n18904_ = ~new_n18777_;
  assign new_n18905_ = ~new_n19086_ | ~new_n18634_;
  assign new_n18906_ = ~new_n18803_ | ~new_n18800_;
  assign new_n18907_ = ~new_n18653_;
  assign new_n18908_ = ~new_n19092_ | ~new_n18635_;
  assign new_n18909_ = ~new_n18720_ | ~new_n18777_;
  assign new_n18910_ = ~new_n18775_;
  assign new_n18911_ = ~new_n19041_ | ~new_n18632_;
  assign new_n18912_ = ~new_n4802_ | ~new_n18667_;
  assign new_n18913_ = ~new_n19041_ | ~new_n18632_;
  assign new_n18914_ = ~new_n18908_ | ~new_n18777_;
  assign new_n18915_ = ~new_n18776_;
  assign new_n18916_ = ~new_n19086_ | ~new_n18634_;
  assign new_n18917_ = ~new_n18916_ | ~new_n18776_;
  assign new_n18918_ = ~new_n18726_ | ~new_n18917_;
  assign new_n18919_ = ~new_n18727_ | ~new_n18914_;
  assign new_n18920_ = ~new_n4803_ | ~new_n18669_;
  assign new_n18921_ = ~new_n18728_ | ~new_n18919_;
  assign new_n18922_ = ~new_n19086_ | ~new_n18634_;
  assign new_n18923_ = ~new_n18892_ | ~new_n18784_;
  assign new_n18924_ = ~new_n18654_;
  assign new_n18925_ = ~new_n19074_ | ~new_n18647_;
  assign new_n18926_ = ~new_n18925_ | ~new_n18654_;
  assign new_n18927_ = ~new_n18729_ | ~new_n18926_;
  assign new_n18928_ = ~new_n18924_ | ~new_n18799_;
  assign new_n18929_ = ~new_n4808_ | ~new_n18681_;
  assign new_n18930_ = ~new_n18730_ | ~new_n18928_;
  assign new_n18931_ = ~new_n19074_ | ~new_n18647_;
  assign new_n18932_ = ~new_n19065_ | ~new_n18636_;
  assign new_n18933_ = ~new_n18932_ | ~new_n18655_;
  assign new_n18934_ = ~new_n18731_ | ~new_n18933_;
  assign new_n18935_ = ~new_n18874_ | ~new_n18637_;
  assign new_n18936_ = ~new_n4812_ | ~new_n18672_;
  assign new_n18937_ = ~new_n18732_ | ~new_n18935_;
  assign new_n18938_ = ~new_n19065_ | ~new_n18636_;
  assign new_n18939_ = ~new_n18862_ | ~new_n18791_;
  assign new_n18940_ = ~new_n18656_;
  assign new_n18941_ = ~new_n19050_ | ~new_n18640_;
  assign new_n18942_ = ~new_n18941_ | ~new_n18656_;
  assign new_n18943_ = ~new_n18733_ | ~new_n18942_;
  assign new_n18944_ = ~new_n18940_ | ~new_n18798_;
  assign new_n18945_ = ~new_n4816_ | ~new_n18675_;
  assign new_n18946_ = ~new_n18734_ | ~new_n18944_;
  assign new_n18947_ = ~new_n19050_ | ~new_n18640_;
  assign new_n18948_ = ~new_n18843_ | ~new_n18619_;
  assign new_n18949_ = ~new_n18850_ | ~new_n18622_;
  assign new_n18950_ = ~new_n18922_ | ~new_n18800_;
  assign new_n18951_ = ~new_n18908_ | ~new_n18803_;
  assign new_n18952_ = ~new_n18931_ | ~new_n18799_;
  assign new_n18953_ = ~new_n18892_ | ~new_n18649_;
  assign new_n18954_ = ~new_n18938_ | ~new_n18637_;
  assign new_n18955_ = ~new_n18947_ | ~new_n18798_;
  assign new_n18956_ = ~new_n18862_ | ~new_n18642_;
  assign new_n18957_ = ~new_n4825_ | ~new_n18664_;
  assign new_n18958_ = ~new_n18721_ | ~new_n18959_ | ~new_n18909_;
  assign new_n18959_ = ~new_n18906_ | ~new_n18794_;
  assign new_n18960_ = ~new_n18669_ | ~new_n18905_;
  assign new_n18961_ = ~new_n4803_ | ~new_n18905_;
  assign new_n18962_ = ~new_n4820_ | ~new_n18657_;
  assign new_n18963_ = ~new_n18913_ | ~new_n18906_ | ~new_n18794_;
  assign new_n18964_ = ~new_n18722_ | ~new_n18777_ | ~new_n18794_;
  assign new_n18965_ = ~new_n18907_ | ~new_n18913_;
  assign new_n18966_ = ~new_n4802_ | ~new_n18667_;
  assign new_n18967_ = ~new_n4830_ | ~new_n18736_;
  assign new_n18968_ = ~new_n5093_ | ~new_n18617_;
  assign new_n18969_ = ~new_n18657_;
  assign new_n18970_ = ~new_n18969_ | ~new_n4820_;
  assign new_n18971_ = ~new_n18657_ | ~new_n18629_;
  assign new_n18972_ = ~new_n18969_ | ~new_n4820_;
  assign new_n18973_ = ~new_n18657_ | ~new_n18629_;
  assign new_n18974_ = ~new_n18973_ | ~new_n18972_;
  assign new_n18975_ = ~new_n4830_ | ~new_n18738_;
  assign new_n18976_ = ~new_n5078_ | ~new_n18617_;
  assign new_n18977_ = ~new_n18664_;
  assign new_n18978_ = ~new_n4830_ | ~new_n18739_;
  assign new_n18979_ = ~new_n5064_ | ~new_n18617_;
  assign new_n18980_ = ~new_n18662_;
  assign new_n18981_ = ~new_n4830_ | ~new_n18740_;
  assign new_n18982_ = ~new_n5069_ | ~new_n18617_;
  assign new_n18983_ = ~new_n18663_;
  assign new_n18984_ = ~new_n4830_ | ~new_n18741_;
  assign new_n18985_ = ~new_n5075_ | ~new_n18617_;
  assign new_n18986_ = ~new_n18661_;
  assign new_n18987_ = ~new_n4830_ | ~new_n18742_;
  assign new_n18988_ = ~new_n5072_ | ~new_n18617_;
  assign new_n18989_ = ~new_n18660_;
  assign new_n18990_ = ~new_n4830_ | ~new_n18743_;
  assign new_n18991_ = ~new_n5081_ | ~new_n18617_;
  assign new_n18992_ = ~new_n18665_;
  assign new_n18993_ = ~new_n4830_ | ~new_n18744_;
  assign new_n18994_ = ~new_n5087_ | ~new_n18617_;
  assign new_n18995_ = ~new_n18659_;
  assign new_n18996_ = ~new_n4830_ | ~new_n18745_;
  assign new_n18997_ = ~new_n5084_ | ~new_n18617_;
  assign new_n18998_ = ~new_n18658_;
  assign new_n18999_ = ~new_n4830_ | ~new_n18746_;
  assign new_n19000_ = ~new_n5090_ | ~new_n18617_;
  assign new_n19001_ = ~new_n18666_;
  assign new_n19002_ = ~new_n18737_ | ~new_n18747_;
  assign new_n19003_ = ~new_n18836_ | ~new_n18974_;
  assign new_n19004_ = ~new_n19001_ | ~new_n4821_;
  assign new_n19005_ = ~new_n18666_ | ~new_n18628_;
  assign new_n19006_ = ~new_n19001_ | ~new_n4821_;
  assign new_n19007_ = ~new_n18666_ | ~new_n18628_;
  assign new_n19008_ = ~new_n19007_ | ~new_n19006_;
  assign new_n19009_ = ~new_n18748_ | ~new_n18749_;
  assign new_n19010_ = ~new_n18832_ | ~new_n19008_;
  assign new_n19011_ = ~new_n18995_ | ~new_n4822_;
  assign new_n19012_ = ~new_n18659_ | ~new_n18620_;
  assign new_n19013_ = ~new_n18998_ | ~new_n4823_;
  assign new_n19014_ = ~new_n18658_ | ~new_n18618_;
  assign new_n19015_ = ~new_n19014_ | ~new_n19013_;
  assign new_n19016_ = ~new_n18948_ | ~new_n18630_;
  assign new_n19017_ = ~new_n19015_ | ~new_n18824_;
  assign new_n19018_ = ~new_n18992_ | ~new_n4824_;
  assign new_n19019_ = ~new_n18665_ | ~new_n18627_;
  assign new_n19020_ = ~new_n18992_ | ~new_n4824_;
  assign new_n19021_ = ~new_n18665_ | ~new_n18627_;
  assign new_n19022_ = ~new_n19021_ | ~new_n19020_;
  assign new_n19023_ = ~new_n18750_ | ~new_n18751_;
  assign new_n19024_ = ~new_n18820_ | ~new_n19022_;
  assign new_n19025_ = ~new_n18977_ | ~new_n4825_;
  assign new_n19026_ = ~new_n18664_ | ~new_n18626_;
  assign new_n19027_ = ~new_n18977_ | ~new_n4825_;
  assign new_n19028_ = ~new_n18664_ | ~new_n18626_;
  assign new_n19029_ = ~new_n19028_ | ~new_n19027_;
  assign new_n19030_ = ~new_n18752_ | ~new_n18753_;
  assign new_n19031_ = ~new_n18818_ | ~new_n19029_;
  assign new_n19032_ = ~new_n18986_ | ~new_n4826_;
  assign new_n19033_ = ~new_n18661_ | ~new_n18623_;
  assign new_n19034_ = ~new_n18989_ | ~new_n4827_;
  assign new_n19035_ = ~new_n18660_ | ~new_n18621_;
  assign new_n19036_ = ~new_n19035_ | ~new_n19034_;
  assign new_n19037_ = ~new_n18949_ | ~new_n18631_;
  assign new_n19038_ = ~new_n19036_ | ~new_n18811_;
  assign new_n19039_ = ~new_n4830_ | ~new_n18754_;
  assign new_n19040_ = ~new_n5585_ | ~new_n18617_;
  assign new_n19041_ = ~new_n18667_;
  assign new_n19042_ = ~new_n4830_ | ~new_n18755_;
  assign new_n19043_ = ~new_n5096_ | ~new_n18617_;
  assign new_n19044_ = ~new_n18673_;
  assign new_n19045_ = ~new_n4830_ | ~new_n18756_;
  assign new_n19046_ = ~new_n5105_ | ~new_n18617_;
  assign new_n19047_ = ~new_n18675_;
  assign new_n19048_ = ~new_n4830_ | ~new_n18757_;
  assign new_n19049_ = ~new_n5102_ | ~new_n18617_;
  assign new_n19050_ = ~new_n18676_;
  assign new_n19051_ = ~new_n4830_ | ~new_n18758_;
  assign new_n19052_ = ~new_n5099_ | ~new_n18617_;
  assign new_n19053_ = ~new_n18674_;
  assign new_n19054_ = ~new_n4830_ | ~new_n18759_;
  assign new_n19055_ = ~new_n5108_ | ~new_n18617_;
  assign new_n19056_ = ~new_n18677_;
  assign new_n19057_ = ~new_n4830_ | ~new_n18760_;
  assign new_n19058_ = ~new_n5111_ | ~new_n18617_;
  assign new_n19059_ = ~new_n18678_;
  assign new_n19060_ = ~new_n4830_ | ~new_n18761_;
  assign new_n19061_ = ~new_n5117_ | ~new_n18617_;
  assign new_n19062_ = ~new_n18672_;
  assign new_n19063_ = ~new_n4830_ | ~new_n18762_;
  assign new_n19064_ = ~new_n5114_ | ~new_n18617_;
  assign new_n19065_ = ~new_n18671_;
  assign new_n19066_ = ~new_n4830_ | ~new_n18763_;
  assign new_n19067_ = ~new_n5120_ | ~new_n18617_;
  assign new_n19068_ = ~new_n18679_;
  assign new_n19069_ = ~new_n4830_ | ~new_n18764_;
  assign new_n19070_ = ~new_n5591_ | ~new_n18617_;
  assign new_n19071_ = ~new_n18681_;
  assign new_n19072_ = ~new_n4830_ | ~new_n18765_;
  assign new_n19073_ = ~new_n5592_ | ~new_n18617_;
  assign new_n19074_ = ~new_n18682_;
  assign new_n19075_ = ~new_n4830_ | ~new_n18766_;
  assign new_n19076_ = ~new_n5122_ | ~new_n18617_;
  assign new_n19077_ = ~new_n18680_;
  assign new_n19078_ = ~new_n4830_ | ~new_n18767_;
  assign new_n19079_ = ~new_n5590_ | ~new_n18617_;
  assign new_n19080_ = ~new_n18683_;
  assign new_n19081_ = ~new_n4830_ | ~new_n18768_;
  assign new_n19082_ = ~new_n5589_ | ~new_n18617_;
  assign new_n19083_ = ~new_n18684_;
  assign new_n19084_ = ~new_n4830_ | ~new_n18769_;
  assign new_n19085_ = ~new_n5587_ | ~new_n18617_;
  assign new_n19086_ = ~new_n18668_;
  assign new_n19087_ = ~new_n4830_ | ~new_n18770_;
  assign new_n19088_ = ~new_n5586_ | ~new_n18617_;
  assign new_n19089_ = ~new_n18669_;
  assign new_n19090_ = ~new_n4830_ | ~new_n18771_;
  assign new_n19091_ = ~new_n5588_ | ~new_n18617_;
  assign new_n19092_ = ~new_n18670_;
  assign new_n19093_ = ~new_n4830_ | ~new_n18772_;
  assign new_n19094_ = ~new_n4801_ | ~new_n18617_;
  assign new_n19095_ = ~new_n18724_;
  assign new_n19096_ = ~new_n5584_ | ~new_n19095_;
  assign new_n19097_ = ~new_n18724_ | ~new_n18773_;
  assign new_n19098_ = ~new_n18685_;
  assign new_n19099_ = ~new_n19098_ | ~new_n18958_ | ~new_n18911_;
  assign new_n19100_ = ~new_n18685_ | ~new_n18723_ | ~new_n18965_ | ~new_n18964_;
  assign new_n19101_ = ~new_n19041_ | ~new_n4802_;
  assign new_n19102_ = ~new_n18667_ | ~new_n18632_;
  assign new_n19103_ = ~new_n19041_ | ~new_n4802_;
  assign new_n19104_ = ~new_n18667_ | ~new_n18632_;
  assign new_n19105_ = ~new_n19104_ | ~new_n19103_;
  assign new_n19106_ = ~new_n18774_ | ~new_n18775_;
  assign new_n19107_ = ~new_n18910_ | ~new_n19105_;
  assign new_n19108_ = ~new_n19089_ | ~new_n4803_;
  assign new_n19109_ = ~new_n18669_ | ~new_n18633_;
  assign new_n19110_ = ~new_n19086_ | ~new_n4804_;
  assign new_n19111_ = ~new_n18668_ | ~new_n18634_;
  assign new_n19112_ = ~new_n19111_ | ~new_n19110_;
  assign new_n19113_ = ~new_n18950_ | ~new_n18776_;
  assign new_n19114_ = ~new_n18915_ | ~new_n19112_;
  assign new_n19115_ = ~new_n19092_ | ~new_n4805_;
  assign new_n19116_ = ~new_n18670_ | ~new_n18635_;
  assign new_n19117_ = ~new_n19116_ | ~new_n19115_;
  assign new_n19118_ = ~new_n18951_ | ~new_n18777_;
  assign new_n19119_ = ~new_n18904_ | ~new_n19117_;
  assign new_n19120_ = ~new_n19083_ | ~new_n4806_;
  assign new_n19121_ = ~new_n18684_ | ~new_n18652_;
  assign new_n19122_ = ~new_n19083_ | ~new_n4806_;
  assign new_n19123_ = ~new_n18684_ | ~new_n18652_;
  assign new_n19124_ = ~new_n19123_ | ~new_n19122_;
  assign new_n19125_ = ~new_n18778_ | ~new_n18779_;
  assign new_n19126_ = ~new_n18900_ | ~new_n19124_;
  assign new_n19127_ = ~new_n19080_ | ~new_n4807_;
  assign new_n19128_ = ~new_n18683_ | ~new_n18651_;
  assign new_n19129_ = ~new_n19080_ | ~new_n4807_;
  assign new_n19130_ = ~new_n18683_ | ~new_n18651_;
  assign new_n19131_ = ~new_n19130_ | ~new_n19129_;
  assign new_n19132_ = ~new_n18780_ | ~new_n18781_;
  assign new_n19133_ = ~new_n18896_ | ~new_n19131_;
  assign new_n19134_ = ~new_n19071_ | ~new_n4808_;
  assign new_n19135_ = ~new_n18681_ | ~new_n18650_;
  assign new_n19136_ = ~new_n19074_ | ~new_n4809_;
  assign new_n19137_ = ~new_n18682_ | ~new_n18647_;
  assign new_n19138_ = ~new_n19137_ | ~new_n19136_;
  assign new_n19139_ = ~new_n18952_ | ~new_n18654_;
  assign new_n19140_ = ~new_n19138_ | ~new_n18924_;
  assign new_n19141_ = ~new_n18983_ | ~new_n4828_;
  assign new_n19142_ = ~new_n18663_ | ~new_n18625_;
  assign new_n19143_ = ~new_n18983_ | ~new_n4828_;
  assign new_n19144_ = ~new_n18663_ | ~new_n18625_;
  assign new_n19145_ = ~new_n19144_ | ~new_n19143_;
  assign new_n19146_ = ~new_n18782_ | ~new_n18783_;
  assign new_n19147_ = ~new_n18807_ | ~new_n19145_;
  assign new_n19148_ = ~new_n19077_ | ~new_n4810_;
  assign new_n19149_ = ~new_n18680_ | ~new_n18648_;
  assign new_n19150_ = ~new_n19149_ | ~new_n19148_;
  assign new_n19151_ = ~new_n18953_ | ~new_n18784_;
  assign new_n19152_ = ~new_n18886_ | ~new_n19150_;
  assign new_n19153_ = ~new_n19068_ | ~new_n4811_;
  assign new_n19154_ = ~new_n18679_ | ~new_n18646_;
  assign new_n19155_ = ~new_n19068_ | ~new_n4811_;
  assign new_n19156_ = ~new_n18679_ | ~new_n18646_;
  assign new_n19157_ = ~new_n19156_ | ~new_n19155_;
  assign new_n19158_ = ~new_n18785_ | ~new_n18786_;
  assign new_n19159_ = ~new_n18882_ | ~new_n19157_;
  assign new_n19160_ = ~new_n19062_ | ~new_n4812_;
  assign new_n19161_ = ~new_n18672_ | ~new_n18638_;
  assign new_n19162_ = ~new_n19065_ | ~new_n4813_;
  assign new_n19163_ = ~new_n18671_ | ~new_n18636_;
  assign new_n19164_ = ~new_n19163_ | ~new_n19162_;
  assign new_n19165_ = ~new_n18954_ | ~new_n18655_;
  assign new_n19166_ = ~new_n19164_ | ~new_n18874_;
  assign new_n19167_ = ~new_n19059_ | ~new_n4814_;
  assign new_n19168_ = ~new_n18678_ | ~new_n18645_;
  assign new_n19169_ = ~new_n19059_ | ~new_n4814_;
  assign new_n19170_ = ~new_n18678_ | ~new_n18645_;
  assign new_n19171_ = ~new_n19170_ | ~new_n19169_;
  assign new_n19172_ = ~new_n18787_ | ~new_n18788_;
  assign new_n19173_ = ~new_n18870_ | ~new_n19171_;
  assign new_n19174_ = ~new_n19056_ | ~new_n4815_;
  assign new_n19175_ = ~new_n18677_ | ~new_n18644_;
  assign new_n19176_ = ~new_n19056_ | ~new_n4815_;
  assign new_n19177_ = ~new_n18677_ | ~new_n18644_;
  assign new_n19178_ = ~new_n19177_ | ~new_n19176_;
  assign new_n19179_ = ~new_n18789_ | ~new_n18790_;
  assign new_n19180_ = ~new_n18866_ | ~new_n19178_;
  assign new_n19181_ = ~new_n19047_ | ~new_n4816_;
  assign new_n19182_ = ~new_n18675_ | ~new_n18643_;
  assign new_n19183_ = ~new_n19050_ | ~new_n4817_;
  assign new_n19184_ = ~new_n18676_ | ~new_n18640_;
  assign new_n19185_ = ~new_n19184_ | ~new_n19183_;
  assign new_n19186_ = ~new_n18955_ | ~new_n18656_;
  assign new_n19187_ = ~new_n19185_ | ~new_n18940_;
  assign new_n19188_ = ~new_n19053_ | ~new_n4818_;
  assign new_n19189_ = ~new_n18674_ | ~new_n18641_;
  assign new_n19190_ = ~new_n19189_ | ~new_n19188_;
  assign new_n19191_ = ~new_n18956_ | ~new_n18791_;
  assign new_n19192_ = ~new_n18856_ | ~new_n19190_;
  assign new_n19193_ = ~new_n19044_ | ~new_n4819_;
  assign new_n19194_ = ~new_n18673_ | ~new_n18639_;
  assign new_n19195_ = ~new_n19044_ | ~new_n4819_;
  assign new_n19196_ = ~new_n18673_ | ~new_n18639_;
  assign new_n19197_ = ~new_n19196_ | ~new_n19195_;
  assign new_n19198_ = ~new_n18792_ | ~new_n18793_;
  assign new_n19199_ = ~new_n18852_ | ~new_n19197_;
  assign new_n19200_ = ~new_n4829_ | ~new_n18617_;
  assign new_n19201_ = ~new_n4830_ | ~new_n18624_;
  assign new_n19202_ = ~new_n18735_;
  assign new_n19203_ = ~new_n18662_ | ~new_n19202_;
  assign new_n19204_ = ~new_n18735_ | ~new_n18980_;
  assign new_n19205_ = new_n19380_ & new_n19379_;
  assign new_n19206_ = new_n19398_ & new_n19397_;
  assign new_n19207_ = new_n19438_ & new_n19437_;
  assign new_n19208_ = new_n19447_ & new_n19446_;
  assign new_n19209_ = new_n19465_ & new_n19464_;
  assign new_n19210_ = new_n19473_ & new_n19472_;
  assign new_n19211_ = new_n19552_ & new_n19549_;
  assign new_n19212_ = new_n19545_ & new_n19542_;
  assign new_n19213_ = new_n19536_ & new_n19533_;
  assign new_n19214_ = new_n19527_ & new_n19524_;
  assign new_n19215_ = new_n19521_ & new_n19519_;
  assign new_n19216_ = new_n19514_ & new_n19511_;
  assign new_n19217_ = new_n19436_ & new_n19433_;
  assign new_n19218_ = new_n19428_ & new_n19425_;
  assign new_n19219_ = new_n19414_ & new_n19411_;
  assign new_n19220_ = ~new_n5084_;
  assign new_n19221_ = ~new_n4687_;
  assign new_n19222_ = ~new_n4686_;
  assign new_n19223_ = ~new_n4687_ | ~new_n5084_;
  assign new_n19224_ = ~new_n5087_;
  assign new_n19225_ = ~new_n5078_;
  assign new_n19226_ = ~new_n4676_;
  assign new_n19227_ = ~new_n4683_;
  assign new_n19228_ = ~new_n5072_;
  assign new_n19229_ = ~new_n4684_;
  assign new_n19230_ = ~new_n5064_;
  assign new_n19231_ = ~new_n4693_;
  assign new_n19232_ = ~new_n4693_ | ~new_n5064_;
  assign new_n19233_ = ~new_n5075_;
  assign new_n19234_ = ~new_n4680_;
  assign new_n19235_ = ~new_n4676_ | ~new_n5078_;
  assign new_n19236_ = ~new_n5081_;
  assign new_n19237_ = ~new_n5090_;
  assign new_n19238_ = ~new_n4700_;
  assign new_n19239_ = ~new_n4699_;
  assign new_n19240_ = ~new_n5093_;
  assign new_n19241_ = ~new_n19262_ | ~new_n19406_;
  assign new_n19242_ = ~new_n19318_ | ~new_n19394_;
  assign new_n19243_ = ~new_n19383_ | ~new_n19384_;
  assign new_n19244_ = ~new_n5069_ | ~new_n4694_;
  assign new_n19245_ = ~new_n19323_ | ~new_n19420_;
  assign new_n19246_ = ~new_n19417_ | ~new_n19416_;
  assign new_n19247_ = ~new_n5585_;
  assign new_n19248_ = ~new_n4669_;
  assign new_n19249_ = ~new_n4673_;
  assign new_n19250_ = ~new_n5586_;
  assign new_n19251_ = ~new_n5587_;
  assign new_n19252_ = ~new_n4674_;
  assign new_n19253_ = ~new_n5588_;
  assign new_n19254_ = ~new_n4681_;
  assign new_n19255_ = ~new_n5591_;
  assign new_n19256_ = ~new_n4691_;
  assign new_n19257_ = ~new_n5114_;
  assign new_n19258_ = ~new_n4689_;
  assign new_n19259_ = ~new_n4685_;
  assign new_n19260_ = ~new_n4689_ | ~new_n5114_;
  assign new_n19261_ = ~new_n5117_;
  assign new_n19262_ = ~new_n4700_ | ~new_n5090_;
  assign new_n19263_ = ~new_n5096_;
  assign new_n19264_ = ~new_n4678_;
  assign new_n19265_ = ~new_n5102_;
  assign new_n19266_ = ~new_n4688_;
  assign new_n19267_ = ~new_n5099_;
  assign new_n19268_ = ~new_n4679_;
  assign new_n19269_ = ~new_n4679_ | ~new_n5099_;
  assign new_n19270_ = ~new_n5105_;
  assign new_n19271_ = ~new_n4696_;
  assign new_n19272_ = ~new_n5108_;
  assign new_n19273_ = ~new_n4695_;
  assign new_n19274_ = ~new_n5111_;
  assign new_n19275_ = ~new_n4690_;
  assign new_n19276_ = ~new_n5120_;
  assign new_n19277_ = ~new_n4698_;
  assign new_n19278_ = ~new_n4698_ | ~new_n5120_;
  assign new_n19279_ = ~new_n5122_;
  assign new_n19280_ = ~new_n4697_;
  assign new_n19281_ = ~new_n4697_ | ~new_n5122_;
  assign new_n19282_ = ~new_n5592_;
  assign new_n19283_ = ~new_n5590_;
  assign new_n19284_ = ~new_n4677_;
  assign new_n19285_ = ~new_n5589_;
  assign new_n19286_ = ~new_n4682_;
  assign new_n19287_ = ~new_n5586_ | ~new_n4673_;
  assign new_n19288_ = ~new_n4670_;
  assign new_n19289_ = ~new_n5584_;
  assign new_n19290_ = ~new_n19507_ | ~new_n19377_;
  assign new_n19291_ = ~new_n4692_;
  assign new_n19292_ = ~new_n19278_ | ~new_n19516_;
  assign new_n19293_ = ~new_n19462_ | ~new_n19461_;
  assign new_n19294_ = ~new_n19269_ | ~new_n19538_;
  assign new_n19295_ = ~new_n19658_ | ~new_n19657_;
  assign new_n19296_ = ~new_n19705_ | ~new_n19704_;
  assign new_n19297_ = ~new_n19576_ | ~new_n19575_;
  assign new_n19298_ = ~new_n19581_ | ~new_n19580_;
  assign new_n19299_ = ~new_n19588_ | ~new_n19587_;
  assign new_n19300_ = ~new_n19595_ | ~new_n19594_;
  assign new_n19301_ = ~new_n19600_ | ~new_n19599_;
  assign new_n19302_ = ~new_n19609_ | ~new_n19608_;
  assign new_n19303_ = ~new_n19616_ | ~new_n19615_;
  assign new_n19304_ = ~new_n19623_ | ~new_n19622_;
  assign new_n19305_ = ~new_n19630_ | ~new_n19629_;
  assign new_n19306_ = ~new_n19635_ | ~new_n19634_;
  assign new_n19307_ = ~new_n19642_ | ~new_n19641_;
  assign new_n19308_ = ~new_n19649_ | ~new_n19648_;
  assign new_n19309_ = ~new_n19663_ | ~new_n19662_;
  assign new_n19310_ = ~new_n19668_ | ~new_n19667_;
  assign new_n19311_ = ~new_n19675_ | ~new_n19674_;
  assign new_n19312_ = ~new_n19682_ | ~new_n19681_;
  assign new_n19313_ = ~new_n19689_ | ~new_n19688_;
  assign new_n19314_ = ~new_n19696_ | ~new_n19695_;
  assign new_n19315_ = ~new_n19701_ | ~new_n19700_;
  assign new_n19316_ = new_n19390_ & new_n19388_;
  assign new_n19317_ = new_n19205_ & new_n19381_;
  assign new_n19318_ = new_n19395_ & new_n19393_;
  assign new_n19319_ = new_n19402_ & new_n19401_;
  assign new_n19320_ = new_n19223_ & new_n19583_ & new_n19582_;
  assign new_n19321_ = new_n19413_ & new_n19206_;
  assign new_n19322_ = new_n19382_ & new_n19381_;
  assign new_n19323_ = new_n19421_ & new_n19419_;
  assign new_n19324_ = new_n19235_ & new_n19590_ & new_n19589_;
  assign new_n19325_ = new_n19427_ & new_n19205_;
  assign new_n19326_ = new_n19435_ & new_n19382_;
  assign new_n19327_ = new_n19405_ & new_n19207_;
  assign new_n19328_ = new_n19440_ & new_n19372_;
  assign new_n19329_ = new_n19451_ & new_n19208_;
  assign new_n19330_ = new_n19449_ & new_n19373_;
  assign new_n19331_ = new_n19469_ & new_n19468_;
  assign new_n19332_ = new_n19474_ & new_n19210_ & new_n19483_;
  assign new_n19333_ = new_n19486_ & new_n19481_;
  assign new_n19334_ = new_n19502_ & new_n19499_;
  assign new_n19335_ = new_n19569_ & new_n19503_;
  assign new_n19336_ = new_n19374_ & new_n19625_ & new_n19624_;
  assign new_n19337_ = new_n19361_ & new_n19479_;
  assign new_n19338_ = new_n19281_ & new_n19656_ & new_n19655_;
  assign new_n19339_ = new_n19526_ & new_n19210_;
  assign new_n19340_ = new_n19260_ & new_n19670_ & new_n19669_;
  assign new_n19341_ = new_n19535_ & new_n19209_;
  assign new_n19342_ = new_n19373_ & new_n19691_ & new_n19690_;
  assign new_n19343_ = new_n19544_ & new_n19208_;
  assign new_n19344_ = new_n19372_ & new_n19703_ & new_n19702_;
  assign new_n19345_ = new_n19551_ & new_n19207_;
  assign new_n19346_ = ~new_n19319_ | ~new_n19403_;
  assign new_n19347_ = ~new_n19418_ | ~new_n19430_;
  assign new_n19348_ = ~new_n4671_;
  assign new_n19349_ = ~new_n5595_;
  assign new_n19350_ = new_n19604_ & new_n19603_;
  assign new_n19351_ = ~new_n19565_ | ~new_n19505_ | ~new_n19370_;
  assign new_n19352_ = new_n19611_ & new_n19610_;
  assign new_n19353_ = ~new_n19335_ | ~new_n19571_ | ~new_n19570_;
  assign new_n19354_ = new_n19618_ & new_n19617_;
  assign new_n19355_ = ~new_n19287_ | ~new_n19566_ | ~new_n19500_;
  assign new_n19356_ = ~new_n19494_ | ~new_n19493_;
  assign new_n19357_ = new_n19637_ & new_n19636_;
  assign new_n19358_ = ~new_n19490_ | ~new_n19489_;
  assign new_n19359_ = new_n19644_ & new_n19643_;
  assign new_n19360_ = ~new_n19333_ | ~new_n19485_;
  assign new_n19361_ = new_n19651_ & new_n19650_;
  assign new_n19362_ = ~new_n19244_ | ~new_n19528_;
  assign new_n19363_ = ~new_n19331_ | ~new_n19470_;
  assign new_n19364_ = new_n19677_ & new_n19676_;
  assign new_n19365_ = ~new_n19458_ | ~new_n19457_;
  assign new_n19366_ = new_n19684_ & new_n19683_;
  assign new_n19367_ = ~new_n19454_ | ~new_n19453_;
  assign new_n19368_ = ~new_n19444_ | ~new_n19443_;
  assign new_n19369_ = ~new_n19568_ | ~new_n19567_;
  assign new_n19370_ = ~new_n4670_ | ~new_n19353_;
  assign new_n19371_ = ~new_n19235_;
  assign new_n19372_ = ~new_n5093_ | ~new_n4699_;
  assign new_n19373_ = ~new_n4688_ | ~new_n5102_;
  assign new_n19374_ = ~new_n4674_ | ~new_n5587_;
  assign new_n19375_ = ~new_n19269_;
  assign new_n19376_ = ~new_n19278_;
  assign new_n19377_ = ~new_n4681_ | ~new_n5588_;
  assign new_n19378_ = ~new_n19262_;
  assign new_n19379_ = new_n4683_ | new_n5081_;
  assign new_n19380_ = new_n4676_ | new_n5078_;
  assign new_n19381_ = new_n5075_ | new_n4680_;
  assign new_n19382_ = new_n5072_ | new_n4684_;
  assign new_n19383_ = ~new_n19232_;
  assign new_n19384_ = new_n5069_ | new_n4694_;
  assign new_n19385_ = ~new_n19243_;
  assign new_n19386_ = ~new_n19244_;
  assign new_n19387_ = ~new_n19243_ | ~new_n19244_;
  assign new_n19388_ = ~new_n4684_ | ~new_n5072_;
  assign new_n19389_ = ~new_n19387_ | ~new_n19382_;
  assign new_n19390_ = ~new_n4680_ | ~new_n5075_;
  assign new_n19391_ = ~new_n19316_ | ~new_n19389_;
  assign new_n19392_ = ~new_n19236_ | ~new_n19235_;
  assign new_n19393_ = ~new_n4683_ | ~new_n19392_;
  assign new_n19394_ = ~new_n19317_ | ~new_n19391_;
  assign new_n19395_ = ~new_n5081_ | ~new_n19371_;
  assign new_n19396_ = ~new_n19242_;
  assign new_n19397_ = new_n4686_ | new_n5087_;
  assign new_n19398_ = new_n4687_ | new_n5084_;
  assign new_n19399_ = ~new_n19223_;
  assign new_n19400_ = ~new_n19224_ | ~new_n19223_;
  assign new_n19401_ = ~new_n4686_ | ~new_n19400_;
  assign new_n19402_ = ~new_n5087_ | ~new_n19399_;
  assign new_n19403_ = ~new_n19206_ | ~new_n19242_;
  assign new_n19404_ = ~new_n19346_;
  assign new_n19405_ = new_n5090_ | new_n4700_;
  assign new_n19406_ = ~new_n19405_ | ~new_n19346_;
  assign new_n19407_ = ~new_n19241_;
  assign new_n19408_ = new_n4699_ | new_n5093_;
  assign new_n19409_ = new_n5084_ | new_n4687_;
  assign new_n19410_ = ~new_n19409_ | ~new_n19242_;
  assign new_n19411_ = ~new_n19320_ | ~new_n19410_;
  assign new_n19412_ = ~new_n19396_ | ~new_n19223_;
  assign new_n19413_ = ~new_n5087_ | ~new_n4686_;
  assign new_n19414_ = ~new_n19321_ | ~new_n19412_;
  assign new_n19415_ = new_n4687_ | new_n5084_;
  assign new_n19416_ = ~new_n19386_ | ~new_n19382_;
  assign new_n19417_ = ~new_n4684_ | ~new_n5072_;
  assign new_n19418_ = ~new_n19246_;
  assign new_n19419_ = ~new_n19322_ | ~new_n19385_;
  assign new_n19420_ = ~new_n19246_ | ~new_n19381_;
  assign new_n19421_ = ~new_n4680_ | ~new_n5075_;
  assign new_n19422_ = ~new_n19245_;
  assign new_n19423_ = new_n5078_ | new_n4676_;
  assign new_n19424_ = ~new_n19423_ | ~new_n19245_;
  assign new_n19425_ = ~new_n19324_ | ~new_n19424_;
  assign new_n19426_ = ~new_n19422_ | ~new_n19235_;
  assign new_n19427_ = ~new_n5081_ | ~new_n4683_;
  assign new_n19428_ = ~new_n19325_ | ~new_n19426_;
  assign new_n19429_ = new_n4676_ | new_n5078_;
  assign new_n19430_ = ~new_n19385_ | ~new_n19382_;
  assign new_n19431_ = ~new_n19347_;
  assign new_n19432_ = ~new_n4680_ | ~new_n5075_;
  assign new_n19433_ = ~new_n19243_ | ~new_n19244_ | ~new_n19602_ | ~new_n19601_;
  assign new_n19434_ = ~new_n19244_ | ~new_n19243_;
  assign new_n19435_ = ~new_n4684_ | ~new_n5072_;
  assign new_n19436_ = ~new_n19326_ | ~new_n19434_;
  assign new_n19437_ = new_n4699_ | new_n5093_;
  assign new_n19438_ = new_n4678_ | new_n5096_;
  assign new_n19439_ = ~new_n19378_ | ~new_n19207_;
  assign new_n19440_ = ~new_n4678_ | ~new_n5096_;
  assign new_n19441_ = ~new_n19328_ | ~new_n19439_;
  assign new_n19442_ = new_n5096_ | new_n4678_;
  assign new_n19443_ = ~new_n19327_ | ~new_n19346_;
  assign new_n19444_ = ~new_n19442_ | ~new_n19441_;
  assign new_n19445_ = ~new_n19368_;
  assign new_n19446_ = new_n4696_ | new_n5105_;
  assign new_n19447_ = new_n4688_ | new_n5102_;
  assign new_n19448_ = ~new_n19375_ | ~new_n19208_;
  assign new_n19449_ = ~new_n4696_ | ~new_n5105_;
  assign new_n19450_ = ~new_n19330_ | ~new_n19448_;
  assign new_n19451_ = new_n5099_ | new_n4679_;
  assign new_n19452_ = new_n5105_ | new_n4696_;
  assign new_n19453_ = ~new_n19329_ | ~new_n19368_;
  assign new_n19454_ = ~new_n19452_ | ~new_n19450_;
  assign new_n19455_ = ~new_n19367_;
  assign new_n19456_ = new_n5108_ | new_n4695_;
  assign new_n19457_ = ~new_n19456_ | ~new_n19367_;
  assign new_n19458_ = ~new_n4695_ | ~new_n5108_;
  assign new_n19459_ = ~new_n19365_;
  assign new_n19460_ = new_n5111_ | new_n4690_;
  assign new_n19461_ = ~new_n19460_ | ~new_n19365_;
  assign new_n19462_ = ~new_n4690_ | ~new_n5111_;
  assign new_n19463_ = ~new_n19293_;
  assign new_n19464_ = new_n4685_ | new_n5117_;
  assign new_n19465_ = new_n4689_ | new_n5114_;
  assign new_n19466_ = ~new_n19260_;
  assign new_n19467_ = ~new_n19261_ | ~new_n19260_;
  assign new_n19468_ = ~new_n4685_ | ~new_n19467_;
  assign new_n19469_ = ~new_n5117_ | ~new_n19466_;
  assign new_n19470_ = ~new_n19209_ | ~new_n19293_;
  assign new_n19471_ = ~new_n19363_;
  assign new_n19472_ = new_n4692_ | new_n5592_;
  assign new_n19473_ = new_n4697_ | new_n5122_;
  assign new_n19474_ = new_n4691_ | new_n5591_;
  assign new_n19475_ = ~new_n19281_;
  assign new_n19476_ = ~new_n5592_ | ~new_n19475_;
  assign new_n19477_ = ~new_n19476_ | ~new_n19291_;
  assign new_n19478_ = ~new_n19281_ | ~new_n19282_;
  assign new_n19479_ = ~new_n19478_ | ~new_n19477_;
  assign new_n19480_ = ~new_n19376_ | ~new_n19210_;
  assign new_n19481_ = ~new_n4691_ | ~new_n5591_;
  assign new_n19482_ = ~new_n19479_ | ~new_n19480_;
  assign new_n19483_ = new_n5120_ | new_n4698_;
  assign new_n19484_ = new_n5591_ | new_n4691_;
  assign new_n19485_ = ~new_n19363_ | ~new_n19332_;
  assign new_n19486_ = ~new_n19484_ | ~new_n19482_;
  assign new_n19487_ = ~new_n19360_;
  assign new_n19488_ = new_n5590_ | new_n4677_;
  assign new_n19489_ = ~new_n19488_ | ~new_n19360_;
  assign new_n19490_ = ~new_n4677_ | ~new_n5590_;
  assign new_n19491_ = ~new_n19358_;
  assign new_n19492_ = new_n5589_ | new_n4682_;
  assign new_n19493_ = ~new_n19492_ | ~new_n19358_;
  assign new_n19494_ = ~new_n4682_ | ~new_n5589_;
  assign new_n19495_ = ~new_n19356_;
  assign new_n19496_ = new_n4674_ | new_n5587_;
  assign new_n19497_ = ~new_n19377_ | ~new_n19374_;
  assign new_n19498_ = ~new_n19287_;
  assign new_n19499_ = new_n5588_ | new_n4681_;
  assign new_n19500_ = ~new_n19369_ | ~new_n19356_ | ~new_n19499_;
  assign new_n19501_ = ~new_n19355_;
  assign new_n19502_ = new_n5585_ | new_n4669_;
  assign new_n19503_ = ~new_n4669_ | ~new_n5585_;
  assign new_n19504_ = ~new_n19353_;
  assign new_n19505_ = ~new_n5584_ | ~new_n19353_;
  assign new_n19506_ = ~new_n19351_;
  assign new_n19507_ = ~new_n19499_ | ~new_n19356_;
  assign new_n19508_ = ~new_n19290_;
  assign new_n19509_ = new_n5587_ | new_n4674_;
  assign new_n19510_ = ~new_n19509_ | ~new_n19290_;
  assign new_n19511_ = ~new_n19336_ | ~new_n19510_;
  assign new_n19512_ = ~new_n19508_ | ~new_n19374_;
  assign new_n19513_ = ~new_n5586_ | ~new_n4673_;
  assign new_n19514_ = ~new_n19369_ | ~new_n19512_ | ~new_n19513_;
  assign new_n19515_ = new_n4674_ | new_n5587_;
  assign new_n19516_ = ~new_n19483_ | ~new_n19363_;
  assign new_n19517_ = ~new_n19292_;
  assign new_n19518_ = ~new_n19210_ | ~new_n19292_;
  assign new_n19519_ = ~new_n19337_ | ~new_n19518_;
  assign new_n19520_ = ~new_n19518_ | ~new_n19479_;
  assign new_n19521_ = ~new_n19654_ | ~new_n19520_;
  assign new_n19522_ = new_n5122_ | new_n4697_;
  assign new_n19523_ = ~new_n19522_ | ~new_n19292_;
  assign new_n19524_ = ~new_n19338_ | ~new_n19523_;
  assign new_n19525_ = ~new_n19517_ | ~new_n19281_;
  assign new_n19526_ = ~new_n4692_ | ~new_n5592_;
  assign new_n19527_ = ~new_n19339_ | ~new_n19525_;
  assign new_n19528_ = new_n5069_ | new_n4694_;
  assign new_n19529_ = ~new_n19362_;
  assign new_n19530_ = new_n4697_ | new_n5122_;
  assign new_n19531_ = new_n5114_ | new_n4689_;
  assign new_n19532_ = ~new_n19531_ | ~new_n19293_;
  assign new_n19533_ = ~new_n19340_ | ~new_n19532_;
  assign new_n19534_ = ~new_n19463_ | ~new_n19260_;
  assign new_n19535_ = ~new_n5117_ | ~new_n4685_;
  assign new_n19536_ = ~new_n19341_ | ~new_n19534_;
  assign new_n19537_ = new_n4689_ | new_n5114_;
  assign new_n19538_ = ~new_n19451_ | ~new_n19368_;
  assign new_n19539_ = ~new_n19294_;
  assign new_n19540_ = new_n5102_ | new_n4688_;
  assign new_n19541_ = ~new_n19540_ | ~new_n19294_;
  assign new_n19542_ = ~new_n19342_ | ~new_n19541_;
  assign new_n19543_ = ~new_n19539_ | ~new_n19373_;
  assign new_n19544_ = ~new_n4696_ | ~new_n5105_;
  assign new_n19545_ = ~new_n19343_ | ~new_n19543_;
  assign new_n19546_ = new_n4688_ | new_n5102_;
  assign new_n19547_ = new_n5093_ | new_n4699_;
  assign new_n19548_ = ~new_n19547_ | ~new_n19241_;
  assign new_n19549_ = ~new_n19344_ | ~new_n19548_;
  assign new_n19550_ = ~new_n19407_ | ~new_n19372_;
  assign new_n19551_ = ~new_n4678_ | ~new_n5096_;
  assign new_n19552_ = ~new_n19345_ | ~new_n19550_;
  assign new_n19553_ = ~new_n19408_ | ~new_n19372_;
  assign new_n19554_ = ~new_n19405_ | ~new_n19262_;
  assign new_n19555_ = ~new_n19415_ | ~new_n19223_;
  assign new_n19556_ = ~new_n19429_ | ~new_n19235_;
  assign new_n19557_ = ~new_n19432_ | ~new_n19381_;
  assign new_n19558_ = ~new_n19515_ | ~new_n19374_;
  assign new_n19559_ = ~new_n19499_ | ~new_n19377_;
  assign new_n19560_ = ~new_n19530_ | ~new_n19281_;
  assign new_n19561_ = ~new_n19483_ | ~new_n19278_;
  assign new_n19562_ = ~new_n19537_ | ~new_n19260_;
  assign new_n19563_ = ~new_n19546_ | ~new_n19373_;
  assign new_n19564_ = ~new_n19451_ | ~new_n19269_;
  assign new_n19565_ = ~new_n5584_ | ~new_n4670_;
  assign new_n19566_ = ~new_n19497_ | ~new_n19369_;
  assign new_n19567_ = ~new_n4673_ | ~new_n19496_;
  assign new_n19568_ = ~new_n5586_ | ~new_n19496_;
  assign new_n19569_ = ~new_n19502_ | ~new_n19497_ | ~new_n19369_;
  assign new_n19570_ = ~new_n19334_ | ~new_n19356_ | ~new_n19369_;
  assign new_n19571_ = ~new_n19498_ | ~new_n19502_;
  assign new_n19572_ = ~new_n4699_ | ~new_n19240_;
  assign new_n19573_ = ~new_n5093_ | ~new_n19239_;
  assign new_n19574_ = ~new_n19573_ | ~new_n19572_;
  assign new_n19575_ = ~new_n19553_ | ~new_n19241_;
  assign new_n19576_ = ~new_n19574_ | ~new_n19407_;
  assign new_n19577_ = ~new_n4700_ | ~new_n19237_;
  assign new_n19578_ = ~new_n5090_ | ~new_n19238_;
  assign new_n19579_ = ~new_n19578_ | ~new_n19577_;
  assign new_n19580_ = ~new_n19554_ | ~new_n19346_;
  assign new_n19581_ = ~new_n19404_ | ~new_n19579_;
  assign new_n19582_ = ~new_n4686_ | ~new_n19224_;
  assign new_n19583_ = ~new_n5087_ | ~new_n19222_;
  assign new_n19584_ = ~new_n4687_ | ~new_n19220_;
  assign new_n19585_ = ~new_n5084_ | ~new_n19221_;
  assign new_n19586_ = ~new_n19585_ | ~new_n19584_;
  assign new_n19587_ = ~new_n19555_ | ~new_n19242_;
  assign new_n19588_ = ~new_n19586_ | ~new_n19396_;
  assign new_n19589_ = ~new_n4683_ | ~new_n19236_;
  assign new_n19590_ = ~new_n5081_ | ~new_n19227_;
  assign new_n19591_ = ~new_n4676_ | ~new_n19225_;
  assign new_n19592_ = ~new_n5078_ | ~new_n19226_;
  assign new_n19593_ = ~new_n19592_ | ~new_n19591_;
  assign new_n19594_ = ~new_n19556_ | ~new_n19245_;
  assign new_n19595_ = ~new_n19593_ | ~new_n19422_;
  assign new_n19596_ = ~new_n4680_ | ~new_n19233_;
  assign new_n19597_ = ~new_n5075_ | ~new_n19234_;
  assign new_n19598_ = ~new_n19597_ | ~new_n19596_;
  assign new_n19599_ = ~new_n19557_ | ~new_n19347_;
  assign new_n19600_ = ~new_n19431_ | ~new_n19598_;
  assign new_n19601_ = ~new_n4684_ | ~new_n19228_;
  assign new_n19602_ = ~new_n5072_ | ~new_n19229_;
  assign new_n19603_ = ~new_n4671_ | ~new_n19349_;
  assign new_n19604_ = ~new_n5595_ | ~new_n19348_;
  assign new_n19605_ = ~new_n4671_ | ~new_n19349_;
  assign new_n19606_ = ~new_n5595_ | ~new_n19348_;
  assign new_n19607_ = ~new_n19606_ | ~new_n19605_;
  assign new_n19608_ = ~new_n19350_ | ~new_n19351_;
  assign new_n19609_ = ~new_n19506_ | ~new_n19607_;
  assign new_n19610_ = ~new_n4670_ | ~new_n19289_;
  assign new_n19611_ = ~new_n5584_ | ~new_n19288_;
  assign new_n19612_ = ~new_n4670_ | ~new_n19289_;
  assign new_n19613_ = ~new_n5584_ | ~new_n19288_;
  assign new_n19614_ = ~new_n19613_ | ~new_n19612_;
  assign new_n19615_ = ~new_n19352_ | ~new_n19353_;
  assign new_n19616_ = ~new_n19504_ | ~new_n19614_;
  assign new_n19617_ = ~new_n4669_ | ~new_n19247_;
  assign new_n19618_ = ~new_n5585_ | ~new_n19248_;
  assign new_n19619_ = ~new_n4669_ | ~new_n19247_;
  assign new_n19620_ = ~new_n5585_ | ~new_n19248_;
  assign new_n19621_ = ~new_n19620_ | ~new_n19619_;
  assign new_n19622_ = ~new_n19354_ | ~new_n19355_;
  assign new_n19623_ = ~new_n19501_ | ~new_n19621_;
  assign new_n19624_ = ~new_n4673_ | ~new_n19250_;
  assign new_n19625_ = ~new_n5586_ | ~new_n19249_;
  assign new_n19626_ = ~new_n4674_ | ~new_n19251_;
  assign new_n19627_ = ~new_n5587_ | ~new_n19252_;
  assign new_n19628_ = ~new_n19627_ | ~new_n19626_;
  assign new_n19629_ = ~new_n19558_ | ~new_n19290_;
  assign new_n19630_ = ~new_n19628_ | ~new_n19508_;
  assign new_n19631_ = ~new_n4681_ | ~new_n19253_;
  assign new_n19632_ = ~new_n5588_ | ~new_n19254_;
  assign new_n19633_ = ~new_n19632_ | ~new_n19631_;
  assign new_n19634_ = ~new_n19559_ | ~new_n19356_;
  assign new_n19635_ = ~new_n19495_ | ~new_n19633_;
  assign new_n19636_ = ~new_n4682_ | ~new_n19285_;
  assign new_n19637_ = ~new_n5589_ | ~new_n19286_;
  assign new_n19638_ = ~new_n4682_ | ~new_n19285_;
  assign new_n19639_ = ~new_n5589_ | ~new_n19286_;
  assign new_n19640_ = ~new_n19639_ | ~new_n19638_;
  assign new_n19641_ = ~new_n19357_ | ~new_n19358_;
  assign new_n19642_ = ~new_n19491_ | ~new_n19640_;
  assign new_n19643_ = ~new_n4677_ | ~new_n19283_;
  assign new_n19644_ = ~new_n5590_ | ~new_n19284_;
  assign new_n19645_ = ~new_n4677_ | ~new_n19283_;
  assign new_n19646_ = ~new_n5590_ | ~new_n19284_;
  assign new_n19647_ = ~new_n19646_ | ~new_n19645_;
  assign new_n19648_ = ~new_n19359_ | ~new_n19360_;
  assign new_n19649_ = ~new_n19487_ | ~new_n19647_;
  assign new_n19650_ = ~new_n4691_ | ~new_n19255_;
  assign new_n19651_ = ~new_n5591_ | ~new_n19256_;
  assign new_n19652_ = ~new_n4691_ | ~new_n19255_;
  assign new_n19653_ = ~new_n5591_ | ~new_n19256_;
  assign new_n19654_ = ~new_n19653_ | ~new_n19652_;
  assign new_n19655_ = ~new_n4692_ | ~new_n19282_;
  assign new_n19656_ = ~new_n5592_ | ~new_n19291_;
  assign new_n19657_ = ~new_n19383_ | ~new_n19362_;
  assign new_n19658_ = ~new_n19529_ | ~new_n19232_;
  assign new_n19659_ = ~new_n4697_ | ~new_n19279_;
  assign new_n19660_ = ~new_n5122_ | ~new_n19280_;
  assign new_n19661_ = ~new_n19660_ | ~new_n19659_;
  assign new_n19662_ = ~new_n19560_ | ~new_n19292_;
  assign new_n19663_ = ~new_n19661_ | ~new_n19517_;
  assign new_n19664_ = ~new_n4698_ | ~new_n19276_;
  assign new_n19665_ = ~new_n5120_ | ~new_n19277_;
  assign new_n19666_ = ~new_n19665_ | ~new_n19664_;
  assign new_n19667_ = ~new_n19561_ | ~new_n19363_;
  assign new_n19668_ = ~new_n19471_ | ~new_n19666_;
  assign new_n19669_ = ~new_n4685_ | ~new_n19261_;
  assign new_n19670_ = ~new_n5117_ | ~new_n19259_;
  assign new_n19671_ = ~new_n4689_ | ~new_n19257_;
  assign new_n19672_ = ~new_n5114_ | ~new_n19258_;
  assign new_n19673_ = ~new_n19672_ | ~new_n19671_;
  assign new_n19674_ = ~new_n19562_ | ~new_n19293_;
  assign new_n19675_ = ~new_n19673_ | ~new_n19463_;
  assign new_n19676_ = ~new_n4690_ | ~new_n19274_;
  assign new_n19677_ = ~new_n5111_ | ~new_n19275_;
  assign new_n19678_ = ~new_n4690_ | ~new_n19274_;
  assign new_n19679_ = ~new_n5111_ | ~new_n19275_;
  assign new_n19680_ = ~new_n19679_ | ~new_n19678_;
  assign new_n19681_ = ~new_n19364_ | ~new_n19365_;
  assign new_n19682_ = ~new_n19459_ | ~new_n19680_;
  assign new_n19683_ = ~new_n4695_ | ~new_n19272_;
  assign new_n19684_ = ~new_n5108_ | ~new_n19273_;
  assign new_n19685_ = ~new_n4695_ | ~new_n19272_;
  assign new_n19686_ = ~new_n5108_ | ~new_n19273_;
  assign new_n19687_ = ~new_n19686_ | ~new_n19685_;
  assign new_n19688_ = ~new_n19366_ | ~new_n19367_;
  assign new_n19689_ = ~new_n19455_ | ~new_n19687_;
  assign new_n19690_ = ~new_n4696_ | ~new_n19270_;
  assign new_n19691_ = ~new_n5105_ | ~new_n19271_;
  assign new_n19692_ = ~new_n4688_ | ~new_n19265_;
  assign new_n19693_ = ~new_n5102_ | ~new_n19266_;
  assign new_n19694_ = ~new_n19693_ | ~new_n19692_;
  assign new_n19695_ = ~new_n19563_ | ~new_n19294_;
  assign new_n19696_ = ~new_n19694_ | ~new_n19539_;
  assign new_n19697_ = ~new_n4679_ | ~new_n19267_;
  assign new_n19698_ = ~new_n5099_ | ~new_n19268_;
  assign new_n19699_ = ~new_n19698_ | ~new_n19697_;
  assign new_n19700_ = ~new_n19564_ | ~new_n19368_;
  assign new_n19701_ = ~new_n19445_ | ~new_n19699_;
  assign new_n19702_ = ~new_n4678_ | ~new_n19263_;
  assign new_n19703_ = ~new_n5096_ | ~new_n19264_;
  assign new_n19704_ = ~new_n4693_ | ~new_n19230_;
  assign new_n19705_ = ~new_n5064_ | ~new_n19231_;
  assign new_n19706_ = new_n19905_ & new_n19904_;
  assign new_n19707_ = new_n19944_ & new_n19943_;
  assign new_n19708_ = new_n19961_ & new_n19960_;
  assign new_n19709_ = new_n19985_ & new_n19984_;
  assign new_n19710_ = new_n20084_ & new_n20083_;
  assign new_n19711_ = ~new_n20040_ | ~new_n20043_;
  assign new_n19712_ = ~new_n20029_ | ~new_n20032_;
  assign new_n19713_ = ~new_n20018_ | ~new_n20021_;
  assign new_n19714_ = ~new_n20010_ | ~new_n20012_;
  assign new_n19715_ = ~new_n19856_ | ~new_n20049_ | ~new_n19877_;
  assign new_n19716_ = ~new_n19938_ | ~new_n19940_;
  assign new_n19717_ = ~new_n19930_ | ~new_n19933_;
  assign new_n19718_ = ~new_n19922_ | ~new_n19924_;
  assign new_n19719_ = ~new_n19866_ | ~new_n20046_;
  assign new_n19720_ = ~new_n5087_;
  assign new_n19721_ = ~new_n5081_;
  assign new_n19722_ = ~new_n5072_;
  assign new_n19723_ = ~new_n5064_;
  assign new_n19724_ = ~new_n4694_;
  assign new_n19725_ = ~new_n5075_;
  assign new_n19726_ = ~new_n4684_;
  assign new_n19727_ = ~new_n4684_ | ~new_n19722_;
  assign new_n19728_ = ~new_n4680_;
  assign new_n19729_ = ~new_n5084_;
  assign new_n19730_ = ~new_n5078_;
  assign new_n19731_ = ~new_n4687_;
  assign new_n19732_ = ~new_n4683_;
  assign new_n19733_ = ~new_n4676_;
  assign new_n19734_ = ~new_n4676_ | ~new_n19730_;
  assign new_n19735_ = ~new_n5090_;
  assign new_n19736_ = ~new_n4686_;
  assign new_n19737_ = ~new_n4686_ | ~new_n19720_;
  assign new_n19738_ = ~new_n4700_;
  assign new_n19739_ = ~new_n5093_;
  assign new_n19740_ = ~new_n4699_;
  assign new_n19741_ = ~new_n19911_ | ~new_n19910_;
  assign new_n19742_ = ~new_n19734_ | ~new_n19926_;
  assign new_n19743_ = ~new_n20047_ | ~new_n19895_ | ~new_n19879_;
  assign new_n19744_ = ~new_n5586_;
  assign new_n19745_ = ~new_n5590_;
  assign new_n19746_ = ~new_n5111_;
  assign new_n19747_ = ~new_n5096_;
  assign new_n19748_ = ~new_n5099_;
  assign new_n19749_ = ~new_n4679_;
  assign new_n19750_ = ~new_n4678_;
  assign new_n19751_ = ~new_n4699_ | ~new_n19739_;
  assign new_n19752_ = ~new_n5102_;
  assign new_n19753_ = ~new_n4688_;
  assign new_n19754_ = ~new_n5105_;
  assign new_n19755_ = ~new_n4696_;
  assign new_n19756_ = ~new_n5114_;
  assign new_n19757_ = ~new_n5108_;
  assign new_n19758_ = ~new_n4689_;
  assign new_n19759_ = ~new_n4690_;
  assign new_n19760_ = ~new_n4695_;
  assign new_n19761_ = ~new_n4695_ | ~new_n19757_;
  assign new_n19762_ = ~new_n5117_;
  assign new_n19763_ = ~new_n4685_;
  assign new_n19764_ = ~new_n4698_;
  assign new_n19765_ = ~new_n5122_;
  assign new_n19766_ = ~new_n4697_;
  assign new_n19767_ = ~new_n5592_;
  assign new_n19768_ = ~new_n4692_;
  assign new_n19769_ = ~new_n5589_;
  assign new_n19770_ = ~new_n5591_;
  assign new_n19771_ = ~new_n4682_;
  assign new_n19772_ = ~new_n4677_;
  assign new_n19773_ = ~new_n4691_;
  assign new_n19774_ = ~new_n4691_ | ~new_n19770_;
  assign new_n19775_ = ~new_n5588_;
  assign new_n19776_ = ~new_n4681_;
  assign new_n19777_ = ~new_n5587_;
  assign new_n19778_ = ~new_n4674_;
  assign new_n19779_ = ~new_n5585_;
  assign new_n19780_ = ~new_n4673_;
  assign new_n19781_ = ~new_n4673_ | ~new_n19744_;
  assign new_n19782_ = ~new_n4669_;
  assign new_n19783_ = ~new_n5584_;
  assign new_n19784_ = ~new_n4670_;
  assign new_n19785_ = ~new_n19999_ | ~new_n19998_;
  assign new_n19786_ = ~new_n19774_ | ~new_n20014_;
  assign new_n19787_ = ~new_n19761_ | ~new_n20025_;
  assign new_n19788_ = ~new_n19751_ | ~new_n20036_;
  assign new_n19789_ = ~new_n4693_;
  assign new_n19790_ = ~new_n20094_ | ~new_n20093_;
  assign new_n19791_ = ~new_n20108_ | ~new_n20107_;
  assign new_n19792_ = ~new_n20113_ | ~new_n20112_;
  assign new_n19793_ = ~new_n20129_ | ~new_n20128_;
  assign new_n19794_ = ~new_n20134_ | ~new_n20133_;
  assign new_n19795_ = ~new_n20139_ | ~new_n20138_;
  assign new_n19796_ = ~new_n20144_ | ~new_n20143_;
  assign new_n19797_ = ~new_n20149_ | ~new_n20148_;
  assign new_n19798_ = ~new_n20165_ | ~new_n20164_;
  assign new_n19799_ = ~new_n20170_ | ~new_n20169_;
  assign new_n19800_ = ~new_n20053_ | ~new_n20052_;
  assign new_n19801_ = ~new_n20062_ | ~new_n20061_;
  assign new_n19802_ = ~new_n20069_ | ~new_n20068_;
  assign new_n19803_ = ~new_n20073_ | ~new_n20072_;
  assign new_n19804_ = ~new_n20082_ | ~new_n20081_;
  assign new_n19805_ = ~new_n20103_ | ~new_n20102_;
  assign new_n19806_ = ~new_n20120_ | ~new_n20119_;
  assign new_n19807_ = ~new_n20124_ | ~new_n20123_;
  assign new_n19808_ = ~new_n20156_ | ~new_n20155_;
  assign new_n19809_ = ~new_n20160_ | ~new_n20159_;
  assign new_n19810_ = ~new_n20177_ | ~new_n20176_;
  assign new_n19811_ = new_n19897_ & new_n19887_;
  assign new_n19812_ = new_n19900_ & new_n19901_;
  assign new_n19813_ = new_n19888_ & new_n19908_ & new_n19903_;
  assign new_n19814_ = new_n19913_ & new_n19889_;
  assign new_n19815_ = new_n19916_ & new_n19917_;
  assign new_n19816_ = new_n19737_ & new_n20055_ & new_n20054_;
  assign new_n19817_ = new_n20058_ & new_n19889_;
  assign new_n19818_ = new_n19932_ & new_n19706_;
  assign new_n19819_ = new_n20065_ & new_n19888_;
  assign new_n19820_ = new_n19727_ & new_n20075_ & new_n20074_;
  assign new_n19821_ = new_n20078_ & new_n19887_;
  assign new_n19822_ = new_n19883_ & new_n19942_ & new_n19919_;
  assign new_n19823_ = new_n19959_ & new_n19964_ & new_n19884_;
  assign new_n19824_ = new_n19983_ & new_n19988_ & new_n19885_;
  assign new_n19825_ = new_n20001_ & new_n19886_;
  assign new_n19826_ = new_n20004_ & new_n20005_;
  assign new_n19827_ = new_n20004_ & new_n20005_;
  assign new_n19828_ = new_n19710_ & new_n20008_;
  assign new_n19829_ = ~new_n20091_ | ~new_n20090_;
  assign new_n19830_ = new_n19781_ & new_n20096_ & new_n20095_;
  assign new_n19831_ = new_n20099_ & new_n19886_;
  assign new_n19832_ = ~new_n20105_ | ~new_n20104_;
  assign new_n19833_ = ~new_n20110_ | ~new_n20109_;
  assign new_n19834_ = new_n20020_ & new_n19709_;
  assign new_n19835_ = new_n20116_ & new_n19885_;
  assign new_n19836_ = ~new_n20126_ | ~new_n20125_;
  assign new_n19837_ = ~new_n20131_ | ~new_n20130_;
  assign new_n19838_ = ~new_n20136_ | ~new_n20135_;
  assign new_n19839_ = ~new_n20141_ | ~new_n20140_;
  assign new_n19840_ = ~new_n20146_ | ~new_n20145_;
  assign new_n19841_ = new_n20031_ & new_n19708_;
  assign new_n19842_ = new_n20152_ & new_n19884_;
  assign new_n19843_ = ~new_n20162_ | ~new_n20161_;
  assign new_n19844_ = ~new_n20167_ | ~new_n20166_;
  assign new_n19845_ = new_n20042_ & new_n19707_;
  assign new_n19846_ = new_n20173_ & new_n19883_;
  assign new_n19847_ = new_n20051_ & new_n20050_;
  assign new_n19848_ = ~new_n19815_ | ~new_n19914_;
  assign new_n19849_ = new_n20060_ & new_n20059_;
  assign new_n19850_ = new_n20067_ & new_n20066_;
  assign new_n19851_ = new_n20071_ & new_n20070_;
  assign new_n19852_ = ~new_n19812_ | ~new_n19898_;
  assign new_n19853_ = new_n20080_ & new_n20079_;
  assign new_n19854_ = ~new_n5595_;
  assign new_n19855_ = ~new_n4671_;
  assign new_n19856_ = new_n20089_ & new_n20088_;
  assign new_n19857_ = ~new_n19826_ | ~new_n20002_;
  assign new_n19858_ = new_n20101_ & new_n20100_;
  assign new_n19859_ = ~new_n19995_ | ~new_n19994_;
  assign new_n19860_ = ~new_n19991_ | ~new_n19990_;
  assign new_n19861_ = new_n20118_ & new_n20117_;
  assign new_n19862_ = new_n20122_ & new_n20121_;
  assign new_n19863_ = ~new_n19981_ | ~new_n19980_;
  assign new_n19864_ = ~new_n19977_ | ~new_n19976_;
  assign new_n19865_ = ~new_n5069_;
  assign new_n19866_ = ~new_n5064_ | ~new_n19789_;
  assign new_n19867_ = ~new_n20048_ | ~new_n19973_ | ~new_n19878_;
  assign new_n19868_ = ~new_n5120_;
  assign new_n19869_ = ~new_n19971_ | ~new_n19970_;
  assign new_n19870_ = ~new_n19967_ | ~new_n19966_;
  assign new_n19871_ = new_n20154_ & new_n20153_;
  assign new_n19872_ = new_n20158_ & new_n20157_;
  assign new_n19873_ = ~new_n19957_ | ~new_n19956_;
  assign new_n19874_ = ~new_n19953_ | ~new_n19952_;
  assign new_n19875_ = ~new_n19949_ | ~new_n19948_;
  assign new_n19876_ = new_n20175_ & new_n20174_;
  assign new_n19877_ = ~new_n20087_ | ~new_n20007_ | ~new_n19857_;
  assign new_n19878_ = ~new_n19869_ | ~new_n19868_;
  assign new_n19879_ = ~new_n19866_ | ~new_n19865_;
  assign new_n19880_ = ~new_n19781_;
  assign new_n19881_ = ~new_n19727_;
  assign new_n19882_ = ~new_n19737_;
  assign new_n19883_ = ~new_n5096_ | ~new_n19750_;
  assign new_n19884_ = ~new_n5111_ | ~new_n19759_;
  assign new_n19885_ = ~new_n5590_ | ~new_n19772_;
  assign new_n19886_ = ~new_n5586_ | ~new_n19780_;
  assign new_n19887_ = ~new_n5072_ | ~new_n19726_;
  assign new_n19888_ = ~new_n5081_ | ~new_n19732_;
  assign new_n19889_ = ~new_n5087_ | ~new_n19736_;
  assign new_n19890_ = ~new_n19761_;
  assign new_n19891_ = ~new_n19774_;
  assign new_n19892_ = ~new_n19734_;
  assign new_n19893_ = ~new_n19751_;
  assign new_n19894_ = ~new_n19866_;
  assign new_n19895_ = ~new_n4694_ | ~new_n19866_;
  assign new_n19896_ = ~new_n19743_;
  assign new_n19897_ = ~new_n5075_ | ~new_n19728_;
  assign new_n19898_ = ~new_n19811_ | ~new_n19743_;
  assign new_n19899_ = ~new_n19728_ | ~new_n19727_;
  assign new_n19900_ = ~new_n19899_ | ~new_n19725_;
  assign new_n19901_ = ~new_n4680_ | ~new_n19881_;
  assign new_n19902_ = ~new_n19852_;
  assign new_n19903_ = ~new_n5084_ | ~new_n19731_;
  assign new_n19904_ = ~new_n4687_ | ~new_n19729_;
  assign new_n19905_ = ~new_n4683_ | ~new_n19721_;
  assign new_n19906_ = ~new_n19892_ | ~new_n19888_;
  assign new_n19907_ = ~new_n19706_ | ~new_n19906_;
  assign new_n19908_ = ~new_n5078_ | ~new_n19733_;
  assign new_n19909_ = ~new_n5084_ | ~new_n19731_;
  assign new_n19910_ = ~new_n19852_ | ~new_n19813_;
  assign new_n19911_ = ~new_n19909_ | ~new_n19907_;
  assign new_n19912_ = ~new_n19741_;
  assign new_n19913_ = ~new_n5090_ | ~new_n19738_;
  assign new_n19914_ = ~new_n19814_ | ~new_n19741_;
  assign new_n19915_ = ~new_n19738_ | ~new_n19737_;
  assign new_n19916_ = ~new_n19915_ | ~new_n19735_;
  assign new_n19917_ = ~new_n4700_ | ~new_n19882_;
  assign new_n19918_ = ~new_n19848_;
  assign new_n19919_ = ~new_n5093_ | ~new_n19740_;
  assign new_n19920_ = ~new_n19919_ | ~new_n19751_;
  assign new_n19921_ = ~new_n19912_ | ~new_n19737_;
  assign new_n19922_ = ~new_n19817_ | ~new_n19921_;
  assign new_n19923_ = ~new_n19741_ | ~new_n19889_;
  assign new_n19924_ = ~new_n19816_ | ~new_n19923_;
  assign new_n19925_ = ~new_n19737_ | ~new_n19889_;
  assign new_n19926_ = ~new_n19908_ | ~new_n19852_;
  assign new_n19927_ = ~new_n19742_;
  assign new_n19928_ = ~new_n4683_ | ~new_n19721_;
  assign new_n19929_ = ~new_n19927_ | ~new_n19928_;
  assign new_n19930_ = ~new_n19819_ | ~new_n19929_;
  assign new_n19931_ = ~new_n19742_ | ~new_n19888_;
  assign new_n19932_ = ~new_n5084_ | ~new_n19731_;
  assign new_n19933_ = ~new_n19818_ | ~new_n19931_;
  assign new_n19934_ = ~new_n4683_ | ~new_n19721_;
  assign new_n19935_ = ~new_n19888_ | ~new_n19934_;
  assign new_n19936_ = ~new_n19908_ | ~new_n19734_;
  assign new_n19937_ = ~new_n19896_ | ~new_n19727_;
  assign new_n19938_ = ~new_n19821_ | ~new_n19937_;
  assign new_n19939_ = ~new_n19743_ | ~new_n19887_;
  assign new_n19940_ = ~new_n19820_ | ~new_n19939_;
  assign new_n19941_ = ~new_n19727_ | ~new_n19887_;
  assign new_n19942_ = ~new_n5099_ | ~new_n19749_;
  assign new_n19943_ = ~new_n4679_ | ~new_n19748_;
  assign new_n19944_ = ~new_n4678_ | ~new_n19747_;
  assign new_n19945_ = ~new_n19893_ | ~new_n19883_;
  assign new_n19946_ = ~new_n19707_ | ~new_n19945_;
  assign new_n19947_ = ~new_n5099_ | ~new_n19749_;
  assign new_n19948_ = ~new_n19848_ | ~new_n19822_;
  assign new_n19949_ = ~new_n19947_ | ~new_n19946_;
  assign new_n19950_ = ~new_n19875_;
  assign new_n19951_ = ~new_n5102_ | ~new_n19753_;
  assign new_n19952_ = ~new_n19951_ | ~new_n19875_;
  assign new_n19953_ = ~new_n4688_ | ~new_n19752_;
  assign new_n19954_ = ~new_n19874_;
  assign new_n19955_ = ~new_n5105_ | ~new_n19755_;
  assign new_n19956_ = ~new_n19955_ | ~new_n19874_;
  assign new_n19957_ = ~new_n4696_ | ~new_n19754_;
  assign new_n19958_ = ~new_n19873_;
  assign new_n19959_ = ~new_n5114_ | ~new_n19758_;
  assign new_n19960_ = ~new_n4689_ | ~new_n19756_;
  assign new_n19961_ = ~new_n4690_ | ~new_n19746_;
  assign new_n19962_ = ~new_n19890_ | ~new_n19884_;
  assign new_n19963_ = ~new_n19708_ | ~new_n19962_;
  assign new_n19964_ = ~new_n5108_ | ~new_n19760_;
  assign new_n19965_ = ~new_n5114_ | ~new_n19758_;
  assign new_n19966_ = ~new_n19873_ | ~new_n19823_;
  assign new_n19967_ = ~new_n19965_ | ~new_n19963_;
  assign new_n19968_ = ~new_n19870_;
  assign new_n19969_ = ~new_n5117_ | ~new_n19763_;
  assign new_n19970_ = ~new_n19969_ | ~new_n19870_;
  assign new_n19971_ = ~new_n4685_ | ~new_n19762_;
  assign new_n19972_ = ~new_n19869_;
  assign new_n19973_ = ~new_n4698_ | ~new_n19869_;
  assign new_n19974_ = ~new_n19867_;
  assign new_n19975_ = ~new_n5122_ | ~new_n19766_;
  assign new_n19976_ = ~new_n19975_ | ~new_n19867_;
  assign new_n19977_ = ~new_n4697_ | ~new_n19765_;
  assign new_n19978_ = ~new_n19864_;
  assign new_n19979_ = ~new_n5592_ | ~new_n19768_;
  assign new_n19980_ = ~new_n19979_ | ~new_n19864_;
  assign new_n19981_ = ~new_n4692_ | ~new_n19767_;
  assign new_n19982_ = ~new_n19863_;
  assign new_n19983_ = ~new_n5589_ | ~new_n19771_;
  assign new_n19984_ = ~new_n4682_ | ~new_n19769_;
  assign new_n19985_ = ~new_n4677_ | ~new_n19745_;
  assign new_n19986_ = ~new_n19891_ | ~new_n19885_;
  assign new_n19987_ = ~new_n19709_ | ~new_n19986_;
  assign new_n19988_ = ~new_n5591_ | ~new_n19773_;
  assign new_n19989_ = ~new_n5589_ | ~new_n19771_;
  assign new_n19990_ = ~new_n19863_ | ~new_n19824_;
  assign new_n19991_ = ~new_n19989_ | ~new_n19987_;
  assign new_n19992_ = ~new_n19860_;
  assign new_n19993_ = ~new_n5588_ | ~new_n19776_;
  assign new_n19994_ = ~new_n19993_ | ~new_n19860_;
  assign new_n19995_ = ~new_n4681_ | ~new_n19775_;
  assign new_n19996_ = ~new_n19859_;
  assign new_n19997_ = ~new_n5587_ | ~new_n19778_;
  assign new_n19998_ = ~new_n19997_ | ~new_n19859_;
  assign new_n19999_ = ~new_n4674_ | ~new_n19777_;
  assign new_n20000_ = ~new_n19785_;
  assign new_n20001_ = ~new_n5585_ | ~new_n19782_;
  assign new_n20002_ = ~new_n19825_ | ~new_n19785_;
  assign new_n20003_ = ~new_n19782_ | ~new_n19781_;
  assign new_n20004_ = ~new_n20003_ | ~new_n19779_;
  assign new_n20005_ = ~new_n4669_ | ~new_n19880_;
  assign new_n20006_ = ~new_n19857_;
  assign new_n20007_ = ~new_n5584_ | ~new_n19784_;
  assign new_n20008_ = ~new_n4670_ | ~new_n19783_;
  assign new_n20009_ = ~new_n20000_ | ~new_n19781_;
  assign new_n20010_ = ~new_n19831_ | ~new_n20009_;
  assign new_n20011_ = ~new_n19785_ | ~new_n19886_;
  assign new_n20012_ = ~new_n19830_ | ~new_n20011_;
  assign new_n20013_ = ~new_n19781_ | ~new_n19886_;
  assign new_n20014_ = ~new_n19988_ | ~new_n19863_;
  assign new_n20015_ = ~new_n19786_;
  assign new_n20016_ = ~new_n4677_ | ~new_n19745_;
  assign new_n20017_ = ~new_n20015_ | ~new_n20016_;
  assign new_n20018_ = ~new_n19835_ | ~new_n20017_;
  assign new_n20019_ = ~new_n19786_ | ~new_n19885_;
  assign new_n20020_ = ~new_n5589_ | ~new_n19771_;
  assign new_n20021_ = ~new_n19834_ | ~new_n20019_;
  assign new_n20022_ = ~new_n4677_ | ~new_n19745_;
  assign new_n20023_ = ~new_n19885_ | ~new_n20022_;
  assign new_n20024_ = ~new_n19988_ | ~new_n19774_;
  assign new_n20025_ = ~new_n19964_ | ~new_n19873_;
  assign new_n20026_ = ~new_n19787_;
  assign new_n20027_ = ~new_n4690_ | ~new_n19746_;
  assign new_n20028_ = ~new_n20026_ | ~new_n20027_;
  assign new_n20029_ = ~new_n19842_ | ~new_n20028_;
  assign new_n20030_ = ~new_n19787_ | ~new_n19884_;
  assign new_n20031_ = ~new_n5114_ | ~new_n19758_;
  assign new_n20032_ = ~new_n19841_ | ~new_n20030_;
  assign new_n20033_ = ~new_n4690_ | ~new_n19746_;
  assign new_n20034_ = ~new_n19884_ | ~new_n20033_;
  assign new_n20035_ = ~new_n19964_ | ~new_n19761_;
  assign new_n20036_ = ~new_n19919_ | ~new_n19848_;
  assign new_n20037_ = ~new_n19788_;
  assign new_n20038_ = ~new_n4678_ | ~new_n19747_;
  assign new_n20039_ = ~new_n20037_ | ~new_n20038_;
  assign new_n20040_ = ~new_n19846_ | ~new_n20039_;
  assign new_n20041_ = ~new_n19788_ | ~new_n19883_;
  assign new_n20042_ = ~new_n5099_ | ~new_n19749_;
  assign new_n20043_ = ~new_n19845_ | ~new_n20041_;
  assign new_n20044_ = ~new_n4678_ | ~new_n19747_;
  assign new_n20045_ = ~new_n19883_ | ~new_n20044_;
  assign new_n20046_ = ~new_n4693_ | ~new_n19723_;
  assign new_n20047_ = ~new_n4694_ | ~new_n19865_;
  assign new_n20048_ = ~new_n4698_ | ~new_n19868_;
  assign new_n20049_ = ~new_n19828_ | ~new_n19827_ | ~new_n20002_;
  assign new_n20050_ = ~new_n5093_ | ~new_n19740_;
  assign new_n20051_ = ~new_n4699_ | ~new_n19739_;
  assign new_n20052_ = ~new_n19920_ | ~new_n19848_;
  assign new_n20053_ = ~new_n19918_ | ~new_n19847_;
  assign new_n20054_ = ~new_n5090_ | ~new_n19738_;
  assign new_n20055_ = ~new_n4700_ | ~new_n19735_;
  assign new_n20056_ = ~new_n5090_ | ~new_n19738_;
  assign new_n20057_ = ~new_n4700_ | ~new_n19735_;
  assign new_n20058_ = ~new_n20057_ | ~new_n20056_;
  assign new_n20059_ = ~new_n5087_ | ~new_n19736_;
  assign new_n20060_ = ~new_n4686_ | ~new_n19720_;
  assign new_n20061_ = ~new_n19925_ | ~new_n19741_;
  assign new_n20062_ = ~new_n19849_ | ~new_n19912_;
  assign new_n20063_ = ~new_n5084_ | ~new_n19731_;
  assign new_n20064_ = ~new_n4687_ | ~new_n19729_;
  assign new_n20065_ = ~new_n20064_ | ~new_n20063_;
  assign new_n20066_ = ~new_n5081_ | ~new_n19732_;
  assign new_n20067_ = ~new_n4683_ | ~new_n19721_;
  assign new_n20068_ = ~new_n19935_ | ~new_n19742_;
  assign new_n20069_ = ~new_n19850_ | ~new_n19927_;
  assign new_n20070_ = ~new_n5078_ | ~new_n19733_;
  assign new_n20071_ = ~new_n4676_ | ~new_n19730_;
  assign new_n20072_ = ~new_n19936_ | ~new_n19852_;
  assign new_n20073_ = ~new_n19902_ | ~new_n19851_;
  assign new_n20074_ = ~new_n5075_ | ~new_n19728_;
  assign new_n20075_ = ~new_n4680_ | ~new_n19725_;
  assign new_n20076_ = ~new_n5075_ | ~new_n19728_;
  assign new_n20077_ = ~new_n4680_ | ~new_n19725_;
  assign new_n20078_ = ~new_n20077_ | ~new_n20076_;
  assign new_n20079_ = ~new_n5072_ | ~new_n19726_;
  assign new_n20080_ = ~new_n4684_ | ~new_n19722_;
  assign new_n20081_ = ~new_n19941_ | ~new_n19743_;
  assign new_n20082_ = ~new_n19853_ | ~new_n19896_;
  assign new_n20083_ = ~new_n5595_ | ~new_n19855_;
  assign new_n20084_ = ~new_n4671_ | ~new_n19854_;
  assign new_n20085_ = ~new_n5595_ | ~new_n19855_;
  assign new_n20086_ = ~new_n4671_ | ~new_n19854_;
  assign new_n20087_ = ~new_n20086_ | ~new_n20085_;
  assign new_n20088_ = ~new_n19784_ | ~new_n5584_ | ~new_n19710_;
  assign new_n20089_ = ~new_n4670_ | ~new_n20087_ | ~new_n19783_;
  assign new_n20090_ = ~new_n5584_ | ~new_n19784_;
  assign new_n20091_ = ~new_n4670_ | ~new_n19783_;
  assign new_n20092_ = ~new_n19829_;
  assign new_n20093_ = ~new_n20006_ | ~new_n20092_;
  assign new_n20094_ = ~new_n19829_ | ~new_n19857_;
  assign new_n20095_ = ~new_n5585_ | ~new_n19782_;
  assign new_n20096_ = ~new_n4669_ | ~new_n19779_;
  assign new_n20097_ = ~new_n5585_ | ~new_n19782_;
  assign new_n20098_ = ~new_n4669_ | ~new_n19779_;
  assign new_n20099_ = ~new_n20098_ | ~new_n20097_;
  assign new_n20100_ = ~new_n5586_ | ~new_n19780_;
  assign new_n20101_ = ~new_n4673_ | ~new_n19744_;
  assign new_n20102_ = ~new_n20013_ | ~new_n19785_;
  assign new_n20103_ = ~new_n19858_ | ~new_n20000_;
  assign new_n20104_ = ~new_n5587_ | ~new_n19778_;
  assign new_n20105_ = ~new_n4674_ | ~new_n19777_;
  assign new_n20106_ = ~new_n19832_;
  assign new_n20107_ = ~new_n19996_ | ~new_n20106_;
  assign new_n20108_ = ~new_n19832_ | ~new_n19859_;
  assign new_n20109_ = ~new_n5588_ | ~new_n19776_;
  assign new_n20110_ = ~new_n4681_ | ~new_n19775_;
  assign new_n20111_ = ~new_n19833_;
  assign new_n20112_ = ~new_n19992_ | ~new_n20111_;
  assign new_n20113_ = ~new_n19833_ | ~new_n19860_;
  assign new_n20114_ = ~new_n5589_ | ~new_n19771_;
  assign new_n20115_ = ~new_n4682_ | ~new_n19769_;
  assign new_n20116_ = ~new_n20115_ | ~new_n20114_;
  assign new_n20117_ = ~new_n5590_ | ~new_n19772_;
  assign new_n20118_ = ~new_n4677_ | ~new_n19745_;
  assign new_n20119_ = ~new_n20023_ | ~new_n19786_;
  assign new_n20120_ = ~new_n19861_ | ~new_n20015_;
  assign new_n20121_ = ~new_n5591_ | ~new_n19773_;
  assign new_n20122_ = ~new_n4691_ | ~new_n19770_;
  assign new_n20123_ = ~new_n20024_ | ~new_n19863_;
  assign new_n20124_ = ~new_n19982_ | ~new_n19862_;
  assign new_n20125_ = ~new_n5592_ | ~new_n19768_;
  assign new_n20126_ = ~new_n4692_ | ~new_n19767_;
  assign new_n20127_ = ~new_n19836_;
  assign new_n20128_ = ~new_n19978_ | ~new_n20127_;
  assign new_n20129_ = ~new_n19836_ | ~new_n19864_;
  assign new_n20130_ = ~new_n5069_ | ~new_n19724_;
  assign new_n20131_ = ~new_n4694_ | ~new_n19865_;
  assign new_n20132_ = ~new_n19837_;
  assign new_n20133_ = ~new_n19894_ | ~new_n20132_;
  assign new_n20134_ = ~new_n19837_ | ~new_n19866_;
  assign new_n20135_ = ~new_n5122_ | ~new_n19766_;
  assign new_n20136_ = ~new_n4697_ | ~new_n19765_;
  assign new_n20137_ = ~new_n19838_;
  assign new_n20138_ = ~new_n19974_ | ~new_n20137_;
  assign new_n20139_ = ~new_n19838_ | ~new_n19867_;
  assign new_n20140_ = ~new_n5120_ | ~new_n19764_;
  assign new_n20141_ = ~new_n4698_ | ~new_n19868_;
  assign new_n20142_ = ~new_n19839_;
  assign new_n20143_ = ~new_n19972_ | ~new_n20142_;
  assign new_n20144_ = ~new_n19839_ | ~new_n19869_;
  assign new_n20145_ = ~new_n5117_ | ~new_n19763_;
  assign new_n20146_ = ~new_n4685_ | ~new_n19762_;
  assign new_n20147_ = ~new_n19840_;
  assign new_n20148_ = ~new_n19968_ | ~new_n20147_;
  assign new_n20149_ = ~new_n19840_ | ~new_n19870_;
  assign new_n20150_ = ~new_n5114_ | ~new_n19758_;
  assign new_n20151_ = ~new_n4689_ | ~new_n19756_;
  assign new_n20152_ = ~new_n20151_ | ~new_n20150_;
  assign new_n20153_ = ~new_n5111_ | ~new_n19759_;
  assign new_n20154_ = ~new_n4690_ | ~new_n19746_;
  assign new_n20155_ = ~new_n20034_ | ~new_n19787_;
  assign new_n20156_ = ~new_n19871_ | ~new_n20026_;
  assign new_n20157_ = ~new_n5108_ | ~new_n19760_;
  assign new_n20158_ = ~new_n4695_ | ~new_n19757_;
  assign new_n20159_ = ~new_n20035_ | ~new_n19873_;
  assign new_n20160_ = ~new_n19958_ | ~new_n19872_;
  assign new_n20161_ = ~new_n5105_ | ~new_n19755_;
  assign new_n20162_ = ~new_n4696_ | ~new_n19754_;
  assign new_n20163_ = ~new_n19843_;
  assign new_n20164_ = ~new_n19954_ | ~new_n20163_;
  assign new_n20165_ = ~new_n19843_ | ~new_n19874_;
  assign new_n20166_ = ~new_n5102_ | ~new_n19753_;
  assign new_n20167_ = ~new_n4688_ | ~new_n19752_;
  assign new_n20168_ = ~new_n19844_;
  assign new_n20169_ = ~new_n19950_ | ~new_n20168_;
  assign new_n20170_ = ~new_n19844_ | ~new_n19875_;
  assign new_n20171_ = ~new_n5099_ | ~new_n19749_;
  assign new_n20172_ = ~new_n4679_ | ~new_n19748_;
  assign new_n20173_ = ~new_n20172_ | ~new_n20171_;
  assign new_n20174_ = ~new_n5096_ | ~new_n19750_;
  assign new_n20175_ = ~new_n4678_ | ~new_n19747_;
  assign new_n20176_ = ~new_n20045_ | ~new_n19788_;
  assign new_n20177_ = ~new_n19876_ | ~new_n20037_;
  assign new_n20178_ = new_n20377_ & new_n20376_;
  assign new_n20179_ = new_n20416_ & new_n20415_;
  assign new_n20180_ = new_n20433_ & new_n20432_;
  assign new_n20181_ = new_n20457_ & new_n20456_;
  assign new_n20182_ = new_n20556_ & new_n20555_;
  assign new_n20183_ = ~new_n20512_ | ~new_n20515_;
  assign new_n20184_ = ~new_n20501_ | ~new_n20504_;
  assign new_n20185_ = ~new_n20490_ | ~new_n20493_;
  assign new_n20186_ = ~new_n20482_ | ~new_n20484_;
  assign new_n20187_ = ~new_n20328_ | ~new_n20521_ | ~new_n20349_;
  assign new_n20188_ = ~new_n20410_ | ~new_n20412_;
  assign new_n20189_ = ~new_n20402_ | ~new_n20405_;
  assign new_n20190_ = ~new_n20394_ | ~new_n20396_;
  assign new_n20191_ = ~new_n20338_ | ~new_n20518_;
  assign new_n20192_ = ~new_n5087_;
  assign new_n20193_ = ~new_n5081_;
  assign new_n20194_ = ~new_n5072_;
  assign new_n20195_ = ~new_n5064_;
  assign new_n20196_ = ~new_n4694_;
  assign new_n20197_ = ~new_n5075_;
  assign new_n20198_ = ~new_n4684_;
  assign new_n20199_ = ~new_n4684_ | ~new_n20194_;
  assign new_n20200_ = ~new_n4680_;
  assign new_n20201_ = ~new_n5084_;
  assign new_n20202_ = ~new_n5078_;
  assign new_n20203_ = ~new_n4687_;
  assign new_n20204_ = ~new_n4683_;
  assign new_n20205_ = ~new_n4676_;
  assign new_n20206_ = ~new_n4676_ | ~new_n20202_;
  assign new_n20207_ = ~new_n5090_;
  assign new_n20208_ = ~new_n4686_;
  assign new_n20209_ = ~new_n4686_ | ~new_n20192_;
  assign new_n20210_ = ~new_n4700_;
  assign new_n20211_ = ~new_n5093_;
  assign new_n20212_ = ~new_n4699_;
  assign new_n20213_ = ~new_n20383_ | ~new_n20382_;
  assign new_n20214_ = ~new_n20206_ | ~new_n20398_;
  assign new_n20215_ = ~new_n20519_ | ~new_n20367_ | ~new_n20351_;
  assign new_n20216_ = ~new_n5586_;
  assign new_n20217_ = ~new_n5590_;
  assign new_n20218_ = ~new_n5111_;
  assign new_n20219_ = ~new_n5096_;
  assign new_n20220_ = ~new_n5099_;
  assign new_n20221_ = ~new_n4679_;
  assign new_n20222_ = ~new_n4678_;
  assign new_n20223_ = ~new_n4699_ | ~new_n20211_;
  assign new_n20224_ = ~new_n5102_;
  assign new_n20225_ = ~new_n4688_;
  assign new_n20226_ = ~new_n5105_;
  assign new_n20227_ = ~new_n4696_;
  assign new_n20228_ = ~new_n5114_;
  assign new_n20229_ = ~new_n5108_;
  assign new_n20230_ = ~new_n4689_;
  assign new_n20231_ = ~new_n4690_;
  assign new_n20232_ = ~new_n4695_;
  assign new_n20233_ = ~new_n4695_ | ~new_n20229_;
  assign new_n20234_ = ~new_n5117_;
  assign new_n20235_ = ~new_n4685_;
  assign new_n20236_ = ~new_n4698_;
  assign new_n20237_ = ~new_n5122_;
  assign new_n20238_ = ~new_n4697_;
  assign new_n20239_ = ~new_n5592_;
  assign new_n20240_ = ~new_n4692_;
  assign new_n20241_ = ~new_n5589_;
  assign new_n20242_ = ~new_n5591_;
  assign new_n20243_ = ~new_n4682_;
  assign new_n20244_ = ~new_n4677_;
  assign new_n20245_ = ~new_n4691_;
  assign new_n20246_ = ~new_n4691_ | ~new_n20242_;
  assign new_n20247_ = ~new_n5588_;
  assign new_n20248_ = ~new_n4681_;
  assign new_n20249_ = ~new_n5587_;
  assign new_n20250_ = ~new_n4674_;
  assign new_n20251_ = ~new_n5585_;
  assign new_n20252_ = ~new_n4673_;
  assign new_n20253_ = ~new_n4673_ | ~new_n20216_;
  assign new_n20254_ = ~new_n4669_;
  assign new_n20255_ = ~new_n5584_;
  assign new_n20256_ = ~new_n4670_;
  assign new_n20257_ = ~new_n20471_ | ~new_n20470_;
  assign new_n20258_ = ~new_n20246_ | ~new_n20486_;
  assign new_n20259_ = ~new_n20233_ | ~new_n20497_;
  assign new_n20260_ = ~new_n20223_ | ~new_n20508_;
  assign new_n20261_ = ~new_n4693_;
  assign new_n20262_ = ~new_n20566_ | ~new_n20565_;
  assign new_n20263_ = ~new_n20580_ | ~new_n20579_;
  assign new_n20264_ = ~new_n20585_ | ~new_n20584_;
  assign new_n20265_ = ~new_n20601_ | ~new_n20600_;
  assign new_n20266_ = ~new_n20606_ | ~new_n20605_;
  assign new_n20267_ = ~new_n20611_ | ~new_n20610_;
  assign new_n20268_ = ~new_n20616_ | ~new_n20615_;
  assign new_n20269_ = ~new_n20621_ | ~new_n20620_;
  assign new_n20270_ = ~new_n20637_ | ~new_n20636_;
  assign new_n20271_ = ~new_n20642_ | ~new_n20641_;
  assign new_n20272_ = ~new_n20525_ | ~new_n20524_;
  assign new_n20273_ = ~new_n20534_ | ~new_n20533_;
  assign new_n20274_ = ~new_n20541_ | ~new_n20540_;
  assign new_n20275_ = ~new_n20545_ | ~new_n20544_;
  assign new_n20276_ = ~new_n20554_ | ~new_n20553_;
  assign new_n20277_ = ~new_n20575_ | ~new_n20574_;
  assign new_n20278_ = ~new_n20592_ | ~new_n20591_;
  assign new_n20279_ = ~new_n20596_ | ~new_n20595_;
  assign new_n20280_ = ~new_n20628_ | ~new_n20627_;
  assign new_n20281_ = ~new_n20632_ | ~new_n20631_;
  assign new_n20282_ = ~new_n20649_ | ~new_n20648_;
  assign new_n20283_ = new_n20369_ & new_n20359_;
  assign new_n20284_ = new_n20372_ & new_n20373_;
  assign new_n20285_ = new_n20360_ & new_n20380_ & new_n20375_;
  assign new_n20286_ = new_n20385_ & new_n20361_;
  assign new_n20287_ = new_n20388_ & new_n20389_;
  assign new_n20288_ = new_n20209_ & new_n20527_ & new_n20526_;
  assign new_n20289_ = new_n20530_ & new_n20361_;
  assign new_n20290_ = new_n20404_ & new_n20178_;
  assign new_n20291_ = new_n20537_ & new_n20360_;
  assign new_n20292_ = new_n20199_ & new_n20547_ & new_n20546_;
  assign new_n20293_ = new_n20550_ & new_n20359_;
  assign new_n20294_ = new_n20355_ & new_n20414_ & new_n20391_;
  assign new_n20295_ = new_n20431_ & new_n20436_ & new_n20356_;
  assign new_n20296_ = new_n20455_ & new_n20460_ & new_n20357_;
  assign new_n20297_ = new_n20473_ & new_n20358_;
  assign new_n20298_ = new_n20476_ & new_n20477_;
  assign new_n20299_ = new_n20476_ & new_n20477_;
  assign new_n20300_ = new_n20182_ & new_n20480_;
  assign new_n20301_ = ~new_n20563_ | ~new_n20562_;
  assign new_n20302_ = new_n20253_ & new_n20568_ & new_n20567_;
  assign new_n20303_ = new_n20571_ & new_n20358_;
  assign new_n20304_ = ~new_n20577_ | ~new_n20576_;
  assign new_n20305_ = ~new_n20582_ | ~new_n20581_;
  assign new_n20306_ = new_n20492_ & new_n20181_;
  assign new_n20307_ = new_n20588_ & new_n20357_;
  assign new_n20308_ = ~new_n20598_ | ~new_n20597_;
  assign new_n20309_ = ~new_n20603_ | ~new_n20602_;
  assign new_n20310_ = ~new_n20608_ | ~new_n20607_;
  assign new_n20311_ = ~new_n20613_ | ~new_n20612_;
  assign new_n20312_ = ~new_n20618_ | ~new_n20617_;
  assign new_n20313_ = new_n20503_ & new_n20180_;
  assign new_n20314_ = new_n20624_ & new_n20356_;
  assign new_n20315_ = ~new_n20634_ | ~new_n20633_;
  assign new_n20316_ = ~new_n20639_ | ~new_n20638_;
  assign new_n20317_ = new_n20514_ & new_n20179_;
  assign new_n20318_ = new_n20645_ & new_n20355_;
  assign new_n20319_ = new_n20523_ & new_n20522_;
  assign new_n20320_ = ~new_n20287_ | ~new_n20386_;
  assign new_n20321_ = new_n20532_ & new_n20531_;
  assign new_n20322_ = new_n20539_ & new_n20538_;
  assign new_n20323_ = new_n20543_ & new_n20542_;
  assign new_n20324_ = ~new_n20284_ | ~new_n20370_;
  assign new_n20325_ = new_n20552_ & new_n20551_;
  assign new_n20326_ = ~new_n5595_;
  assign new_n20327_ = ~new_n4671_;
  assign new_n20328_ = new_n20561_ & new_n20560_;
  assign new_n20329_ = ~new_n20298_ | ~new_n20474_;
  assign new_n20330_ = new_n20573_ & new_n20572_;
  assign new_n20331_ = ~new_n20467_ | ~new_n20466_;
  assign new_n20332_ = ~new_n20463_ | ~new_n20462_;
  assign new_n20333_ = new_n20590_ & new_n20589_;
  assign new_n20334_ = new_n20594_ & new_n20593_;
  assign new_n20335_ = ~new_n20453_ | ~new_n20452_;
  assign new_n20336_ = ~new_n20449_ | ~new_n20448_;
  assign new_n20337_ = ~new_n5069_;
  assign new_n20338_ = ~new_n5064_ | ~new_n20261_;
  assign new_n20339_ = ~new_n20520_ | ~new_n20445_ | ~new_n20350_;
  assign new_n20340_ = ~new_n5120_;
  assign new_n20341_ = ~new_n20443_ | ~new_n20442_;
  assign new_n20342_ = ~new_n20439_ | ~new_n20438_;
  assign new_n20343_ = new_n20626_ & new_n20625_;
  assign new_n20344_ = new_n20630_ & new_n20629_;
  assign new_n20345_ = ~new_n20429_ | ~new_n20428_;
  assign new_n20346_ = ~new_n20425_ | ~new_n20424_;
  assign new_n20347_ = ~new_n20421_ | ~new_n20420_;
  assign new_n20348_ = new_n20647_ & new_n20646_;
  assign new_n20349_ = ~new_n20559_ | ~new_n20479_ | ~new_n20329_;
  assign new_n20350_ = ~new_n20341_ | ~new_n20340_;
  assign new_n20351_ = ~new_n20338_ | ~new_n20337_;
  assign new_n20352_ = ~new_n20253_;
  assign new_n20353_ = ~new_n20199_;
  assign new_n20354_ = ~new_n20209_;
  assign new_n20355_ = ~new_n5096_ | ~new_n20222_;
  assign new_n20356_ = ~new_n5111_ | ~new_n20231_;
  assign new_n20357_ = ~new_n5590_ | ~new_n20244_;
  assign new_n20358_ = ~new_n5586_ | ~new_n20252_;
  assign new_n20359_ = ~new_n5072_ | ~new_n20198_;
  assign new_n20360_ = ~new_n5081_ | ~new_n20204_;
  assign new_n20361_ = ~new_n5087_ | ~new_n20208_;
  assign new_n20362_ = ~new_n20233_;
  assign new_n20363_ = ~new_n20246_;
  assign new_n20364_ = ~new_n20206_;
  assign new_n20365_ = ~new_n20223_;
  assign new_n20366_ = ~new_n20338_;
  assign new_n20367_ = ~new_n4694_ | ~new_n20338_;
  assign new_n20368_ = ~new_n20215_;
  assign new_n20369_ = ~new_n5075_ | ~new_n20200_;
  assign new_n20370_ = ~new_n20283_ | ~new_n20215_;
  assign new_n20371_ = ~new_n20200_ | ~new_n20199_;
  assign new_n20372_ = ~new_n20371_ | ~new_n20197_;
  assign new_n20373_ = ~new_n4680_ | ~new_n20353_;
  assign new_n20374_ = ~new_n20324_;
  assign new_n20375_ = ~new_n5084_ | ~new_n20203_;
  assign new_n20376_ = ~new_n4687_ | ~new_n20201_;
  assign new_n20377_ = ~new_n4683_ | ~new_n20193_;
  assign new_n20378_ = ~new_n20364_ | ~new_n20360_;
  assign new_n20379_ = ~new_n20178_ | ~new_n20378_;
  assign new_n20380_ = ~new_n5078_ | ~new_n20205_;
  assign new_n20381_ = ~new_n5084_ | ~new_n20203_;
  assign new_n20382_ = ~new_n20324_ | ~new_n20285_;
  assign new_n20383_ = ~new_n20381_ | ~new_n20379_;
  assign new_n20384_ = ~new_n20213_;
  assign new_n20385_ = ~new_n5090_ | ~new_n20210_;
  assign new_n20386_ = ~new_n20286_ | ~new_n20213_;
  assign new_n20387_ = ~new_n20210_ | ~new_n20209_;
  assign new_n20388_ = ~new_n20387_ | ~new_n20207_;
  assign new_n20389_ = ~new_n4700_ | ~new_n20354_;
  assign new_n20390_ = ~new_n20320_;
  assign new_n20391_ = ~new_n5093_ | ~new_n20212_;
  assign new_n20392_ = ~new_n20391_ | ~new_n20223_;
  assign new_n20393_ = ~new_n20384_ | ~new_n20209_;
  assign new_n20394_ = ~new_n20289_ | ~new_n20393_;
  assign new_n20395_ = ~new_n20213_ | ~new_n20361_;
  assign new_n20396_ = ~new_n20288_ | ~new_n20395_;
  assign new_n20397_ = ~new_n20209_ | ~new_n20361_;
  assign new_n20398_ = ~new_n20380_ | ~new_n20324_;
  assign new_n20399_ = ~new_n20214_;
  assign new_n20400_ = ~new_n4683_ | ~new_n20193_;
  assign new_n20401_ = ~new_n20399_ | ~new_n20400_;
  assign new_n20402_ = ~new_n20291_ | ~new_n20401_;
  assign new_n20403_ = ~new_n20214_ | ~new_n20360_;
  assign new_n20404_ = ~new_n5084_ | ~new_n20203_;
  assign new_n20405_ = ~new_n20290_ | ~new_n20403_;
  assign new_n20406_ = ~new_n4683_ | ~new_n20193_;
  assign new_n20407_ = ~new_n20360_ | ~new_n20406_;
  assign new_n20408_ = ~new_n20380_ | ~new_n20206_;
  assign new_n20409_ = ~new_n20368_ | ~new_n20199_;
  assign new_n20410_ = ~new_n20293_ | ~new_n20409_;
  assign new_n20411_ = ~new_n20215_ | ~new_n20359_;
  assign new_n20412_ = ~new_n20292_ | ~new_n20411_;
  assign new_n20413_ = ~new_n20199_ | ~new_n20359_;
  assign new_n20414_ = ~new_n5099_ | ~new_n20221_;
  assign new_n20415_ = ~new_n4679_ | ~new_n20220_;
  assign new_n20416_ = ~new_n4678_ | ~new_n20219_;
  assign new_n20417_ = ~new_n20365_ | ~new_n20355_;
  assign new_n20418_ = ~new_n20179_ | ~new_n20417_;
  assign new_n20419_ = ~new_n5099_ | ~new_n20221_;
  assign new_n20420_ = ~new_n20320_ | ~new_n20294_;
  assign new_n20421_ = ~new_n20419_ | ~new_n20418_;
  assign new_n20422_ = ~new_n20347_;
  assign new_n20423_ = ~new_n5102_ | ~new_n20225_;
  assign new_n20424_ = ~new_n20423_ | ~new_n20347_;
  assign new_n20425_ = ~new_n4688_ | ~new_n20224_;
  assign new_n20426_ = ~new_n20346_;
  assign new_n20427_ = ~new_n5105_ | ~new_n20227_;
  assign new_n20428_ = ~new_n20427_ | ~new_n20346_;
  assign new_n20429_ = ~new_n4696_ | ~new_n20226_;
  assign new_n20430_ = ~new_n20345_;
  assign new_n20431_ = ~new_n5114_ | ~new_n20230_;
  assign new_n20432_ = ~new_n4689_ | ~new_n20228_;
  assign new_n20433_ = ~new_n4690_ | ~new_n20218_;
  assign new_n20434_ = ~new_n20362_ | ~new_n20356_;
  assign new_n20435_ = ~new_n20180_ | ~new_n20434_;
  assign new_n20436_ = ~new_n5108_ | ~new_n20232_;
  assign new_n20437_ = ~new_n5114_ | ~new_n20230_;
  assign new_n20438_ = ~new_n20345_ | ~new_n20295_;
  assign new_n20439_ = ~new_n20437_ | ~new_n20435_;
  assign new_n20440_ = ~new_n20342_;
  assign new_n20441_ = ~new_n5117_ | ~new_n20235_;
  assign new_n20442_ = ~new_n20441_ | ~new_n20342_;
  assign new_n20443_ = ~new_n4685_ | ~new_n20234_;
  assign new_n20444_ = ~new_n20341_;
  assign new_n20445_ = ~new_n4698_ | ~new_n20341_;
  assign new_n20446_ = ~new_n20339_;
  assign new_n20447_ = ~new_n5122_ | ~new_n20238_;
  assign new_n20448_ = ~new_n20447_ | ~new_n20339_;
  assign new_n20449_ = ~new_n4697_ | ~new_n20237_;
  assign new_n20450_ = ~new_n20336_;
  assign new_n20451_ = ~new_n5592_ | ~new_n20240_;
  assign new_n20452_ = ~new_n20451_ | ~new_n20336_;
  assign new_n20453_ = ~new_n4692_ | ~new_n20239_;
  assign new_n20454_ = ~new_n20335_;
  assign new_n20455_ = ~new_n5589_ | ~new_n20243_;
  assign new_n20456_ = ~new_n4682_ | ~new_n20241_;
  assign new_n20457_ = ~new_n4677_ | ~new_n20217_;
  assign new_n20458_ = ~new_n20363_ | ~new_n20357_;
  assign new_n20459_ = ~new_n20181_ | ~new_n20458_;
  assign new_n20460_ = ~new_n5591_ | ~new_n20245_;
  assign new_n20461_ = ~new_n5589_ | ~new_n20243_;
  assign new_n20462_ = ~new_n20335_ | ~new_n20296_;
  assign new_n20463_ = ~new_n20461_ | ~new_n20459_;
  assign new_n20464_ = ~new_n20332_;
  assign new_n20465_ = ~new_n5588_ | ~new_n20248_;
  assign new_n20466_ = ~new_n20465_ | ~new_n20332_;
  assign new_n20467_ = ~new_n4681_ | ~new_n20247_;
  assign new_n20468_ = ~new_n20331_;
  assign new_n20469_ = ~new_n5587_ | ~new_n20250_;
  assign new_n20470_ = ~new_n20469_ | ~new_n20331_;
  assign new_n20471_ = ~new_n4674_ | ~new_n20249_;
  assign new_n20472_ = ~new_n20257_;
  assign new_n20473_ = ~new_n5585_ | ~new_n20254_;
  assign new_n20474_ = ~new_n20297_ | ~new_n20257_;
  assign new_n20475_ = ~new_n20254_ | ~new_n20253_;
  assign new_n20476_ = ~new_n20475_ | ~new_n20251_;
  assign new_n20477_ = ~new_n4669_ | ~new_n20352_;
  assign new_n20478_ = ~new_n20329_;
  assign new_n20479_ = ~new_n5584_ | ~new_n20256_;
  assign new_n20480_ = ~new_n4670_ | ~new_n20255_;
  assign new_n20481_ = ~new_n20472_ | ~new_n20253_;
  assign new_n20482_ = ~new_n20303_ | ~new_n20481_;
  assign new_n20483_ = ~new_n20257_ | ~new_n20358_;
  assign new_n20484_ = ~new_n20302_ | ~new_n20483_;
  assign new_n20485_ = ~new_n20253_ | ~new_n20358_;
  assign new_n20486_ = ~new_n20460_ | ~new_n20335_;
  assign new_n20487_ = ~new_n20258_;
  assign new_n20488_ = ~new_n4677_ | ~new_n20217_;
  assign new_n20489_ = ~new_n20487_ | ~new_n20488_;
  assign new_n20490_ = ~new_n20307_ | ~new_n20489_;
  assign new_n20491_ = ~new_n20258_ | ~new_n20357_;
  assign new_n20492_ = ~new_n5589_ | ~new_n20243_;
  assign new_n20493_ = ~new_n20306_ | ~new_n20491_;
  assign new_n20494_ = ~new_n4677_ | ~new_n20217_;
  assign new_n20495_ = ~new_n20357_ | ~new_n20494_;
  assign new_n20496_ = ~new_n20460_ | ~new_n20246_;
  assign new_n20497_ = ~new_n20436_ | ~new_n20345_;
  assign new_n20498_ = ~new_n20259_;
  assign new_n20499_ = ~new_n4690_ | ~new_n20218_;
  assign new_n20500_ = ~new_n20498_ | ~new_n20499_;
  assign new_n20501_ = ~new_n20314_ | ~new_n20500_;
  assign new_n20502_ = ~new_n20259_ | ~new_n20356_;
  assign new_n20503_ = ~new_n5114_ | ~new_n20230_;
  assign new_n20504_ = ~new_n20313_ | ~new_n20502_;
  assign new_n20505_ = ~new_n4690_ | ~new_n20218_;
  assign new_n20506_ = ~new_n20356_ | ~new_n20505_;
  assign new_n20507_ = ~new_n20436_ | ~new_n20233_;
  assign new_n20508_ = ~new_n20391_ | ~new_n20320_;
  assign new_n20509_ = ~new_n20260_;
  assign new_n20510_ = ~new_n4678_ | ~new_n20219_;
  assign new_n20511_ = ~new_n20509_ | ~new_n20510_;
  assign new_n20512_ = ~new_n20318_ | ~new_n20511_;
  assign new_n20513_ = ~new_n20260_ | ~new_n20355_;
  assign new_n20514_ = ~new_n5099_ | ~new_n20221_;
  assign new_n20515_ = ~new_n20317_ | ~new_n20513_;
  assign new_n20516_ = ~new_n4678_ | ~new_n20219_;
  assign new_n20517_ = ~new_n20355_ | ~new_n20516_;
  assign new_n20518_ = ~new_n4693_ | ~new_n20195_;
  assign new_n20519_ = ~new_n4694_ | ~new_n20337_;
  assign new_n20520_ = ~new_n4698_ | ~new_n20340_;
  assign new_n20521_ = ~new_n20300_ | ~new_n20299_ | ~new_n20474_;
  assign new_n20522_ = ~new_n5093_ | ~new_n20212_;
  assign new_n20523_ = ~new_n4699_ | ~new_n20211_;
  assign new_n20524_ = ~new_n20392_ | ~new_n20320_;
  assign new_n20525_ = ~new_n20390_ | ~new_n20319_;
  assign new_n20526_ = ~new_n5090_ | ~new_n20210_;
  assign new_n20527_ = ~new_n4700_ | ~new_n20207_;
  assign new_n20528_ = ~new_n5090_ | ~new_n20210_;
  assign new_n20529_ = ~new_n4700_ | ~new_n20207_;
  assign new_n20530_ = ~new_n20529_ | ~new_n20528_;
  assign new_n20531_ = ~new_n5087_ | ~new_n20208_;
  assign new_n20532_ = ~new_n4686_ | ~new_n20192_;
  assign new_n20533_ = ~new_n20397_ | ~new_n20213_;
  assign new_n20534_ = ~new_n20321_ | ~new_n20384_;
  assign new_n20535_ = ~new_n5084_ | ~new_n20203_;
  assign new_n20536_ = ~new_n4687_ | ~new_n20201_;
  assign new_n20537_ = ~new_n20536_ | ~new_n20535_;
  assign new_n20538_ = ~new_n5081_ | ~new_n20204_;
  assign new_n20539_ = ~new_n4683_ | ~new_n20193_;
  assign new_n20540_ = ~new_n20407_ | ~new_n20214_;
  assign new_n20541_ = ~new_n20322_ | ~new_n20399_;
  assign new_n20542_ = ~new_n5078_ | ~new_n20205_;
  assign new_n20543_ = ~new_n4676_ | ~new_n20202_;
  assign new_n20544_ = ~new_n20408_ | ~new_n20324_;
  assign new_n20545_ = ~new_n20374_ | ~new_n20323_;
  assign new_n20546_ = ~new_n5075_ | ~new_n20200_;
  assign new_n20547_ = ~new_n4680_ | ~new_n20197_;
  assign new_n20548_ = ~new_n5075_ | ~new_n20200_;
  assign new_n20549_ = ~new_n4680_ | ~new_n20197_;
  assign new_n20550_ = ~new_n20549_ | ~new_n20548_;
  assign new_n20551_ = ~new_n5072_ | ~new_n20198_;
  assign new_n20552_ = ~new_n4684_ | ~new_n20194_;
  assign new_n20553_ = ~new_n20413_ | ~new_n20215_;
  assign new_n20554_ = ~new_n20325_ | ~new_n20368_;
  assign new_n20555_ = ~new_n5595_ | ~new_n20327_;
  assign new_n20556_ = ~new_n4671_ | ~new_n20326_;
  assign new_n20557_ = ~new_n5595_ | ~new_n20327_;
  assign new_n20558_ = ~new_n4671_ | ~new_n20326_;
  assign new_n20559_ = ~new_n20558_ | ~new_n20557_;
  assign new_n20560_ = ~new_n20256_ | ~new_n5584_ | ~new_n20182_;
  assign new_n20561_ = ~new_n4670_ | ~new_n20559_ | ~new_n20255_;
  assign new_n20562_ = ~new_n5584_ | ~new_n20256_;
  assign new_n20563_ = ~new_n4670_ | ~new_n20255_;
  assign new_n20564_ = ~new_n20301_;
  assign new_n20565_ = ~new_n20478_ | ~new_n20564_;
  assign new_n20566_ = ~new_n20301_ | ~new_n20329_;
  assign new_n20567_ = ~new_n5585_ | ~new_n20254_;
  assign new_n20568_ = ~new_n4669_ | ~new_n20251_;
  assign new_n20569_ = ~new_n5585_ | ~new_n20254_;
  assign new_n20570_ = ~new_n4669_ | ~new_n20251_;
  assign new_n20571_ = ~new_n20570_ | ~new_n20569_;
  assign new_n20572_ = ~new_n5586_ | ~new_n20252_;
  assign new_n20573_ = ~new_n4673_ | ~new_n20216_;
  assign new_n20574_ = ~new_n20485_ | ~new_n20257_;
  assign new_n20575_ = ~new_n20330_ | ~new_n20472_;
  assign new_n20576_ = ~new_n5587_ | ~new_n20250_;
  assign new_n20577_ = ~new_n4674_ | ~new_n20249_;
  assign new_n20578_ = ~new_n20304_;
  assign new_n20579_ = ~new_n20468_ | ~new_n20578_;
  assign new_n20580_ = ~new_n20304_ | ~new_n20331_;
  assign new_n20581_ = ~new_n5588_ | ~new_n20248_;
  assign new_n20582_ = ~new_n4681_ | ~new_n20247_;
  assign new_n20583_ = ~new_n20305_;
  assign new_n20584_ = ~new_n20464_ | ~new_n20583_;
  assign new_n20585_ = ~new_n20305_ | ~new_n20332_;
  assign new_n20586_ = ~new_n5589_ | ~new_n20243_;
  assign new_n20587_ = ~new_n4682_ | ~new_n20241_;
  assign new_n20588_ = ~new_n20587_ | ~new_n20586_;
  assign new_n20589_ = ~new_n5590_ | ~new_n20244_;
  assign new_n20590_ = ~new_n4677_ | ~new_n20217_;
  assign new_n20591_ = ~new_n20495_ | ~new_n20258_;
  assign new_n20592_ = ~new_n20333_ | ~new_n20487_;
  assign new_n20593_ = ~new_n5591_ | ~new_n20245_;
  assign new_n20594_ = ~new_n4691_ | ~new_n20242_;
  assign new_n20595_ = ~new_n20496_ | ~new_n20335_;
  assign new_n20596_ = ~new_n20454_ | ~new_n20334_;
  assign new_n20597_ = ~new_n5592_ | ~new_n20240_;
  assign new_n20598_ = ~new_n4692_ | ~new_n20239_;
  assign new_n20599_ = ~new_n20308_;
  assign new_n20600_ = ~new_n20450_ | ~new_n20599_;
  assign new_n20601_ = ~new_n20308_ | ~new_n20336_;
  assign new_n20602_ = ~new_n5069_ | ~new_n20196_;
  assign new_n20603_ = ~new_n4694_ | ~new_n20337_;
  assign new_n20604_ = ~new_n20309_;
  assign new_n20605_ = ~new_n20366_ | ~new_n20604_;
  assign new_n20606_ = ~new_n20309_ | ~new_n20338_;
  assign new_n20607_ = ~new_n5122_ | ~new_n20238_;
  assign new_n20608_ = ~new_n4697_ | ~new_n20237_;
  assign new_n20609_ = ~new_n20310_;
  assign new_n20610_ = ~new_n20446_ | ~new_n20609_;
  assign new_n20611_ = ~new_n20310_ | ~new_n20339_;
  assign new_n20612_ = ~new_n5120_ | ~new_n20236_;
  assign new_n20613_ = ~new_n4698_ | ~new_n20340_;
  assign new_n20614_ = ~new_n20311_;
  assign new_n20615_ = ~new_n20444_ | ~new_n20614_;
  assign new_n20616_ = ~new_n20311_ | ~new_n20341_;
  assign new_n20617_ = ~new_n5117_ | ~new_n20235_;
  assign new_n20618_ = ~new_n4685_ | ~new_n20234_;
  assign new_n20619_ = ~new_n20312_;
  assign new_n20620_ = ~new_n20440_ | ~new_n20619_;
  assign new_n20621_ = ~new_n20312_ | ~new_n20342_;
  assign new_n20622_ = ~new_n5114_ | ~new_n20230_;
  assign new_n20623_ = ~new_n4689_ | ~new_n20228_;
  assign new_n20624_ = ~new_n20623_ | ~new_n20622_;
  assign new_n20625_ = ~new_n5111_ | ~new_n20231_;
  assign new_n20626_ = ~new_n4690_ | ~new_n20218_;
  assign new_n20627_ = ~new_n20506_ | ~new_n20259_;
  assign new_n20628_ = ~new_n20343_ | ~new_n20498_;
  assign new_n20629_ = ~new_n5108_ | ~new_n20232_;
  assign new_n20630_ = ~new_n4695_ | ~new_n20229_;
  assign new_n20631_ = ~new_n20507_ | ~new_n20345_;
  assign new_n20632_ = ~new_n20430_ | ~new_n20344_;
  assign new_n20633_ = ~new_n5105_ | ~new_n20227_;
  assign new_n20634_ = ~new_n4696_ | ~new_n20226_;
  assign new_n20635_ = ~new_n20315_;
  assign new_n20636_ = ~new_n20426_ | ~new_n20635_;
  assign new_n20637_ = ~new_n20315_ | ~new_n20346_;
  assign new_n20638_ = ~new_n5102_ | ~new_n20225_;
  assign new_n20639_ = ~new_n4688_ | ~new_n20224_;
  assign new_n20640_ = ~new_n20316_;
  assign new_n20641_ = ~new_n20422_ | ~new_n20640_;
  assign new_n20642_ = ~new_n20316_ | ~new_n20347_;
  assign new_n20643_ = ~new_n5099_ | ~new_n20221_;
  assign new_n20644_ = ~new_n4679_ | ~new_n20220_;
  assign new_n20645_ = ~new_n20644_ | ~new_n20643_;
  assign new_n20646_ = ~new_n5096_ | ~new_n20222_;
  assign new_n20647_ = ~new_n4678_ | ~new_n20219_;
  assign new_n20648_ = ~new_n20517_ | ~new_n20260_;
  assign new_n20649_ = ~new_n20348_ | ~new_n20509_;
  assign new_n20650_ = new_n20849_ & new_n20848_;
  assign new_n20651_ = new_n20888_ & new_n20887_;
  assign new_n20652_ = new_n20905_ & new_n20904_;
  assign new_n20653_ = new_n20929_ & new_n20928_;
  assign new_n20654_ = new_n21028_ & new_n21027_;
  assign new_n20655_ = ~new_n20984_ | ~new_n20987_;
  assign new_n20656_ = ~new_n20973_ | ~new_n20976_;
  assign new_n20657_ = ~new_n20962_ | ~new_n20965_;
  assign new_n20658_ = ~new_n20954_ | ~new_n20956_;
  assign new_n20659_ = ~new_n20800_ | ~new_n20993_ | ~new_n20821_;
  assign new_n20660_ = ~new_n20882_ | ~new_n20884_;
  assign new_n20661_ = ~new_n20874_ | ~new_n20877_;
  assign new_n20662_ = ~new_n20866_ | ~new_n20868_;
  assign new_n20663_ = ~new_n20810_ | ~new_n20990_;
  assign new_n20664_ = ~new_n5087_;
  assign new_n20665_ = ~new_n5081_;
  assign new_n20666_ = ~new_n5072_;
  assign new_n20667_ = ~new_n5064_;
  assign new_n20668_ = ~new_n4694_;
  assign new_n20669_ = ~new_n5075_;
  assign new_n20670_ = ~new_n4684_;
  assign new_n20671_ = ~new_n4684_ | ~new_n20666_;
  assign new_n20672_ = ~new_n4680_;
  assign new_n20673_ = ~new_n5084_;
  assign new_n20674_ = ~new_n5078_;
  assign new_n20675_ = ~new_n4687_;
  assign new_n20676_ = ~new_n4683_;
  assign new_n20677_ = ~new_n4676_;
  assign new_n20678_ = ~new_n4676_ | ~new_n20674_;
  assign new_n20679_ = ~new_n5090_;
  assign new_n20680_ = ~new_n4686_;
  assign new_n20681_ = ~new_n4686_ | ~new_n20664_;
  assign new_n20682_ = ~new_n4700_;
  assign new_n20683_ = ~new_n5093_;
  assign new_n20684_ = ~new_n4699_;
  assign new_n20685_ = ~new_n20855_ | ~new_n20854_;
  assign new_n20686_ = ~new_n20678_ | ~new_n20870_;
  assign new_n20687_ = ~new_n20991_ | ~new_n20839_ | ~new_n20823_;
  assign new_n20688_ = ~new_n5586_;
  assign new_n20689_ = ~new_n5590_;
  assign new_n20690_ = ~new_n5111_;
  assign new_n20691_ = ~new_n5096_;
  assign new_n20692_ = ~new_n5099_;
  assign new_n20693_ = ~new_n4679_;
  assign new_n20694_ = ~new_n4678_;
  assign new_n20695_ = ~new_n4699_ | ~new_n20683_;
  assign new_n20696_ = ~new_n5102_;
  assign new_n20697_ = ~new_n4688_;
  assign new_n20698_ = ~new_n5105_;
  assign new_n20699_ = ~new_n4696_;
  assign new_n20700_ = ~new_n5114_;
  assign new_n20701_ = ~new_n5108_;
  assign new_n20702_ = ~new_n4689_;
  assign new_n20703_ = ~new_n4690_;
  assign new_n20704_ = ~new_n4695_;
  assign new_n20705_ = ~new_n4695_ | ~new_n20701_;
  assign new_n20706_ = ~new_n5117_;
  assign new_n20707_ = ~new_n4685_;
  assign new_n20708_ = ~new_n4698_;
  assign new_n20709_ = ~new_n5122_;
  assign new_n20710_ = ~new_n4697_;
  assign new_n20711_ = ~new_n5592_;
  assign new_n20712_ = ~new_n4692_;
  assign new_n20713_ = ~new_n5589_;
  assign new_n20714_ = ~new_n5591_;
  assign new_n20715_ = ~new_n4682_;
  assign new_n20716_ = ~new_n4677_;
  assign new_n20717_ = ~new_n4691_;
  assign new_n20718_ = ~new_n4691_ | ~new_n20714_;
  assign new_n20719_ = ~new_n5588_;
  assign new_n20720_ = ~new_n4681_;
  assign new_n20721_ = ~new_n5587_;
  assign new_n20722_ = ~new_n4674_;
  assign new_n20723_ = ~new_n5585_;
  assign new_n20724_ = ~new_n4673_;
  assign new_n20725_ = ~new_n4673_ | ~new_n20688_;
  assign new_n20726_ = ~new_n4669_;
  assign new_n20727_ = ~new_n5584_;
  assign new_n20728_ = ~new_n4670_;
  assign new_n20729_ = ~new_n20943_ | ~new_n20942_;
  assign new_n20730_ = ~new_n20718_ | ~new_n20958_;
  assign new_n20731_ = ~new_n20705_ | ~new_n20969_;
  assign new_n20732_ = ~new_n20695_ | ~new_n20980_;
  assign new_n20733_ = ~new_n4693_;
  assign new_n20734_ = ~new_n21038_ | ~new_n21037_;
  assign new_n20735_ = ~new_n21052_ | ~new_n21051_;
  assign new_n20736_ = ~new_n21057_ | ~new_n21056_;
  assign new_n20737_ = ~new_n7896_ | ~new_n7897_;
  assign new_n20738_ = ~new_n7891_ | ~new_n7892_;
  assign new_n20739_ = ~new_n4629_ | ~new_n7887_;
  assign new_n20740_ = ~new_n4624_ | ~new_n4625_;
  assign new_n20741_ = ~new_n4619_ | ~new_n4620_;
  assign new_n20742_ = ~new_n1350_ | ~new_n1351_;
  assign new_n20743_ = ~new_n1345_ | ~new_n1346_;
  assign new_n20744_ = ~new_n20997_ | ~new_n20996_;
  assign new_n20745_ = ~new_n21006_ | ~new_n21005_;
  assign new_n20746_ = ~new_n21013_ | ~new_n21012_;
  assign new_n20747_ = ~new_n21017_ | ~new_n21016_;
  assign new_n20748_ = ~new_n21026_ | ~new_n21025_;
  assign new_n20749_ = ~new_n21047_ | ~new_n21046_;
  assign new_n20750_ = ~new_n7905_ | ~new_n7906_;
  assign new_n20751_ = ~new_n7901_ | ~new_n7902_;
  assign new_n20752_ = ~new_n4612_ | ~new_n4613_;
  assign new_n20753_ = ~new_n4608_ | ~new_n4609_;
  assign new_n20754_ = ~new_n1036_ | ~new_n1037_;
  assign new_n20755_ = new_n20841_ & new_n20831_;
  assign new_n20756_ = new_n20844_ & new_n20845_;
  assign new_n20757_ = new_n20832_ & new_n20852_ & new_n20847_;
  assign new_n20758_ = new_n20857_ & new_n20833_;
  assign new_n20759_ = new_n20860_ & new_n20861_;
  assign new_n20760_ = new_n20681_ & new_n20999_ & new_n20998_;
  assign new_n20761_ = new_n21002_ & new_n20833_;
  assign new_n20762_ = new_n20876_ & new_n20650_;
  assign new_n20763_ = new_n21009_ & new_n20832_;
  assign new_n20764_ = new_n20671_ & new_n21019_ & new_n21018_;
  assign new_n20765_ = new_n21022_ & new_n20831_;
  assign new_n20766_ = new_n20827_ & new_n20886_ & new_n20863_;
  assign new_n20767_ = new_n20903_ & new_n20908_ & new_n20828_;
  assign new_n20768_ = new_n20927_ & new_n20932_ & new_n20829_;
  assign new_n20769_ = new_n20945_ & new_n20830_;
  assign new_n20770_ = new_n20948_ & new_n20949_;
  assign new_n20771_ = new_n20948_ & new_n20949_;
  assign new_n20772_ = new_n20654_ & new_n20952_;
  assign new_n20773_ = ~new_n21035_ | ~new_n21034_;
  assign new_n20774_ = new_n20725_ & new_n21040_ & new_n21039_;
  assign new_n20775_ = new_n21043_ & new_n20830_;
  assign new_n20776_ = ~new_n21049_ | ~new_n21048_;
  assign new_n20777_ = ~new_n21054_ | ~new_n21053_;
  assign new_n20778_ = new_n20964_ & new_n20653_;
  assign new_n20779_ = new_n21060_ & new_n20829_;
  assign new_n20780_ = ~new_n7899_ | ~new_n7900_;
  assign new_n20781_ = ~new_n7894_ | ~new_n7895_;
  assign new_n20782_ = ~new_n7889_ | ~new_n7890_;
  assign new_n20783_ = ~new_n4627_ | ~new_n4628_;
  assign new_n20784_ = ~new_n4622_ | ~new_n4623_;
  assign new_n20785_ = new_n20975_ & new_n20652_;
  assign new_n20786_ = new_n4616_ & new_n20828_;
  assign new_n20787_ = ~new_n4606_ | ~new_n4607_;
  assign new_n20788_ = ~new_n1348_ | ~new_n1349_;
  assign new_n20789_ = new_n20986_ & new_n20651_;
  assign new_n20790_ = new_n1342_ & new_n20827_;
  assign new_n20791_ = new_n20995_ & new_n20994_;
  assign new_n20792_ = ~new_n20759_ | ~new_n20858_;
  assign new_n20793_ = new_n21004_ & new_n21003_;
  assign new_n20794_ = new_n21011_ & new_n21010_;
  assign new_n20795_ = new_n21015_ & new_n21014_;
  assign new_n20796_ = ~new_n20756_ | ~new_n20842_;
  assign new_n20797_ = new_n21024_ & new_n21023_;
  assign new_n20798_ = ~new_n5595_;
  assign new_n20799_ = ~new_n4671_;
  assign new_n20800_ = new_n21033_ & new_n21032_;
  assign new_n20801_ = ~new_n20770_ | ~new_n20946_;
  assign new_n20802_ = new_n21045_ & new_n21044_;
  assign new_n20803_ = ~new_n20939_ | ~new_n20938_;
  assign new_n20804_ = ~new_n20935_ | ~new_n20934_;
  assign new_n20805_ = new_n21062_ & new_n21061_;
  assign new_n20806_ = new_n7903_ & new_n7904_;
  assign new_n20807_ = ~new_n20925_ | ~new_n20924_;
  assign new_n20808_ = ~new_n20921_ | ~new_n20920_;
  assign new_n20809_ = ~new_n5069_;
  assign new_n20810_ = ~new_n5064_ | ~new_n20733_;
  assign new_n20811_ = ~new_n20992_ | ~new_n20917_ | ~new_n20822_;
  assign new_n20812_ = ~new_n5120_;
  assign new_n20813_ = ~new_n20915_ | ~new_n20914_;
  assign new_n20814_ = ~new_n20911_ | ~new_n20910_;
  assign new_n20815_ = new_n4614_ & new_n4615_;
  assign new_n20816_ = new_n4610_ & new_n4611_;
  assign new_n20817_ = ~new_n20901_ | ~new_n20900_;
  assign new_n20818_ = ~new_n20897_ | ~new_n20896_;
  assign new_n20819_ = ~new_n20893_ | ~new_n20892_;
  assign new_n20820_ = new_n1038_ & new_n1341_;
  assign new_n20821_ = ~new_n21031_ | ~new_n20951_ | ~new_n20801_;
  assign new_n20822_ = ~new_n20813_ | ~new_n20812_;
  assign new_n20823_ = ~new_n20810_ | ~new_n20809_;
  assign new_n20824_ = ~new_n20725_;
  assign new_n20825_ = ~new_n20671_;
  assign new_n20826_ = ~new_n20681_;
  assign new_n20827_ = ~new_n5096_ | ~new_n20694_;
  assign new_n20828_ = ~new_n5111_ | ~new_n20703_;
  assign new_n20829_ = ~new_n5590_ | ~new_n20716_;
  assign new_n20830_ = ~new_n5586_ | ~new_n20724_;
  assign new_n20831_ = ~new_n5072_ | ~new_n20670_;
  assign new_n20832_ = ~new_n5081_ | ~new_n20676_;
  assign new_n20833_ = ~new_n5087_ | ~new_n20680_;
  assign new_n20834_ = ~new_n20705_;
  assign new_n20835_ = ~new_n20718_;
  assign new_n20836_ = ~new_n20678_;
  assign new_n20837_ = ~new_n20695_;
  assign new_n20838_ = ~new_n20810_;
  assign new_n20839_ = ~new_n4694_ | ~new_n20810_;
  assign new_n20840_ = ~new_n20687_;
  assign new_n20841_ = ~new_n5075_ | ~new_n20672_;
  assign new_n20842_ = ~new_n20755_ | ~new_n20687_;
  assign new_n20843_ = ~new_n20672_ | ~new_n20671_;
  assign new_n20844_ = ~new_n20843_ | ~new_n20669_;
  assign new_n20845_ = ~new_n4680_ | ~new_n20825_;
  assign new_n20846_ = ~new_n20796_;
  assign new_n20847_ = ~new_n5084_ | ~new_n20675_;
  assign new_n20848_ = ~new_n4687_ | ~new_n20673_;
  assign new_n20849_ = ~new_n4683_ | ~new_n20665_;
  assign new_n20850_ = ~new_n20836_ | ~new_n20832_;
  assign new_n20851_ = ~new_n20650_ | ~new_n20850_;
  assign new_n20852_ = ~new_n5078_ | ~new_n20677_;
  assign new_n20853_ = ~new_n5084_ | ~new_n20675_;
  assign new_n20854_ = ~new_n20796_ | ~new_n20757_;
  assign new_n20855_ = ~new_n20853_ | ~new_n20851_;
  assign new_n20856_ = ~new_n20685_;
  assign new_n20857_ = ~new_n5090_ | ~new_n20682_;
  assign new_n20858_ = ~new_n20758_ | ~new_n20685_;
  assign new_n20859_ = ~new_n20682_ | ~new_n20681_;
  assign new_n20860_ = ~new_n20859_ | ~new_n20679_;
  assign new_n20861_ = ~new_n4700_ | ~new_n20826_;
  assign new_n20862_ = ~new_n20792_;
  assign new_n20863_ = ~new_n5093_ | ~new_n20684_;
  assign new_n20864_ = ~new_n20863_ | ~new_n20695_;
  assign new_n20865_ = ~new_n20856_ | ~new_n20681_;
  assign new_n20866_ = ~new_n20761_ | ~new_n20865_;
  assign new_n20867_ = ~new_n20685_ | ~new_n20833_;
  assign new_n20868_ = ~new_n20760_ | ~new_n20867_;
  assign new_n20869_ = ~new_n20681_ | ~new_n20833_;
  assign new_n20870_ = ~new_n20852_ | ~new_n20796_;
  assign new_n20871_ = ~new_n20686_;
  assign new_n20872_ = ~new_n4683_ | ~new_n20665_;
  assign new_n20873_ = ~new_n20871_ | ~new_n20872_;
  assign new_n20874_ = ~new_n20763_ | ~new_n20873_;
  assign new_n20875_ = ~new_n20686_ | ~new_n20832_;
  assign new_n20876_ = ~new_n5084_ | ~new_n20675_;
  assign new_n20877_ = ~new_n20762_ | ~new_n20875_;
  assign new_n20878_ = ~new_n4683_ | ~new_n20665_;
  assign new_n20879_ = ~new_n20832_ | ~new_n20878_;
  assign new_n20880_ = ~new_n20852_ | ~new_n20678_;
  assign new_n20881_ = ~new_n20840_ | ~new_n20671_;
  assign new_n20882_ = ~new_n20765_ | ~new_n20881_;
  assign new_n20883_ = ~new_n20687_ | ~new_n20831_;
  assign new_n20884_ = ~new_n20764_ | ~new_n20883_;
  assign new_n20885_ = ~new_n20671_ | ~new_n20831_;
  assign new_n20886_ = ~new_n5099_ | ~new_n20693_;
  assign new_n20887_ = ~new_n4679_ | ~new_n20692_;
  assign new_n20888_ = ~new_n4678_ | ~new_n20691_;
  assign new_n20889_ = ~new_n20837_ | ~new_n20827_;
  assign new_n20890_ = ~new_n20651_ | ~new_n20889_;
  assign new_n20891_ = ~new_n5099_ | ~new_n20693_;
  assign new_n20892_ = ~new_n20792_ | ~new_n20766_;
  assign new_n20893_ = ~new_n20891_ | ~new_n20890_;
  assign new_n20894_ = ~new_n20819_;
  assign new_n20895_ = ~new_n5102_ | ~new_n20697_;
  assign new_n20896_ = ~new_n20895_ | ~new_n20819_;
  assign new_n20897_ = ~new_n4688_ | ~new_n20696_;
  assign new_n20898_ = ~new_n20818_;
  assign new_n20899_ = ~new_n5105_ | ~new_n20699_;
  assign new_n20900_ = ~new_n20899_ | ~new_n20818_;
  assign new_n20901_ = ~new_n4696_ | ~new_n20698_;
  assign new_n20902_ = ~new_n20817_;
  assign new_n20903_ = ~new_n5114_ | ~new_n20702_;
  assign new_n20904_ = ~new_n4689_ | ~new_n20700_;
  assign new_n20905_ = ~new_n4690_ | ~new_n20690_;
  assign new_n20906_ = ~new_n20834_ | ~new_n20828_;
  assign new_n20907_ = ~new_n20652_ | ~new_n20906_;
  assign new_n20908_ = ~new_n5108_ | ~new_n20704_;
  assign new_n20909_ = ~new_n5114_ | ~new_n20702_;
  assign new_n20910_ = ~new_n20817_ | ~new_n20767_;
  assign new_n20911_ = ~new_n20909_ | ~new_n20907_;
  assign new_n20912_ = ~new_n20814_;
  assign new_n20913_ = ~new_n5117_ | ~new_n20707_;
  assign new_n20914_ = ~new_n20913_ | ~new_n20814_;
  assign new_n20915_ = ~new_n4685_ | ~new_n20706_;
  assign new_n20916_ = ~new_n20813_;
  assign new_n20917_ = ~new_n4698_ | ~new_n20813_;
  assign new_n20918_ = ~new_n20811_;
  assign new_n20919_ = ~new_n5122_ | ~new_n20710_;
  assign new_n20920_ = ~new_n20919_ | ~new_n20811_;
  assign new_n20921_ = ~new_n4697_ | ~new_n20709_;
  assign new_n20922_ = ~new_n20808_;
  assign new_n20923_ = ~new_n5592_ | ~new_n20712_;
  assign new_n20924_ = ~new_n20923_ | ~new_n20808_;
  assign new_n20925_ = ~new_n4692_ | ~new_n20711_;
  assign new_n20926_ = ~new_n20807_;
  assign new_n20927_ = ~new_n5589_ | ~new_n20715_;
  assign new_n20928_ = ~new_n4682_ | ~new_n20713_;
  assign new_n20929_ = ~new_n4677_ | ~new_n20689_;
  assign new_n20930_ = ~new_n20835_ | ~new_n20829_;
  assign new_n20931_ = ~new_n20653_ | ~new_n20930_;
  assign new_n20932_ = ~new_n5591_ | ~new_n20717_;
  assign new_n20933_ = ~new_n5589_ | ~new_n20715_;
  assign new_n20934_ = ~new_n20807_ | ~new_n20768_;
  assign new_n20935_ = ~new_n20933_ | ~new_n20931_;
  assign new_n20936_ = ~new_n20804_;
  assign new_n20937_ = ~new_n5588_ | ~new_n20720_;
  assign new_n20938_ = ~new_n20937_ | ~new_n20804_;
  assign new_n20939_ = ~new_n4681_ | ~new_n20719_;
  assign new_n20940_ = ~new_n20803_;
  assign new_n20941_ = ~new_n5587_ | ~new_n20722_;
  assign new_n20942_ = ~new_n20941_ | ~new_n20803_;
  assign new_n20943_ = ~new_n4674_ | ~new_n20721_;
  assign new_n20944_ = ~new_n20729_;
  assign new_n20945_ = ~new_n5585_ | ~new_n20726_;
  assign new_n20946_ = ~new_n20769_ | ~new_n20729_;
  assign new_n20947_ = ~new_n20726_ | ~new_n20725_;
  assign new_n20948_ = ~new_n20947_ | ~new_n20723_;
  assign new_n20949_ = ~new_n4669_ | ~new_n20824_;
  assign new_n20950_ = ~new_n20801_;
  assign new_n20951_ = ~new_n5584_ | ~new_n20728_;
  assign new_n20952_ = ~new_n4670_ | ~new_n20727_;
  assign new_n20953_ = ~new_n20944_ | ~new_n20725_;
  assign new_n20954_ = ~new_n20775_ | ~new_n20953_;
  assign new_n20955_ = ~new_n20729_ | ~new_n20830_;
  assign new_n20956_ = ~new_n20774_ | ~new_n20955_;
  assign new_n20957_ = ~new_n20725_ | ~new_n20830_;
  assign new_n20958_ = ~new_n20932_ | ~new_n20807_;
  assign new_n20959_ = ~new_n20730_;
  assign new_n20960_ = ~new_n4677_ | ~new_n20689_;
  assign new_n20961_ = ~new_n20959_ | ~new_n20960_;
  assign new_n20962_ = ~new_n20779_ | ~new_n20961_;
  assign new_n20963_ = ~new_n20730_ | ~new_n20829_;
  assign new_n20964_ = ~new_n5589_ | ~new_n20715_;
  assign new_n20965_ = ~new_n20778_ | ~new_n20963_;
  assign new_n20966_ = ~new_n4677_ | ~new_n20689_;
  assign new_n20967_ = ~new_n20829_ | ~new_n20966_;
  assign new_n20968_ = ~new_n20932_ | ~new_n20718_;
  assign new_n20969_ = ~new_n20908_ | ~new_n20817_;
  assign new_n20970_ = ~new_n20731_;
  assign new_n20971_ = ~new_n4690_ | ~new_n20690_;
  assign new_n20972_ = ~new_n20970_ | ~new_n20971_;
  assign new_n20973_ = ~new_n20786_ | ~new_n20972_;
  assign new_n20974_ = ~new_n20731_ | ~new_n20828_;
  assign new_n20975_ = ~new_n5114_ | ~new_n20702_;
  assign new_n20976_ = ~new_n20785_ | ~new_n20974_;
  assign new_n20977_ = ~new_n4690_ | ~new_n20690_;
  assign new_n20978_ = ~new_n20828_ | ~new_n20977_;
  assign new_n20979_ = ~new_n20908_ | ~new_n20705_;
  assign new_n20980_ = ~new_n20863_ | ~new_n20792_;
  assign new_n20981_ = ~new_n20732_;
  assign new_n20982_ = ~new_n4678_ | ~new_n20691_;
  assign new_n20983_ = ~new_n20981_ | ~new_n20982_;
  assign new_n20984_ = ~new_n20790_ | ~new_n20983_;
  assign new_n20985_ = ~new_n20732_ | ~new_n20827_;
  assign new_n20986_ = ~new_n5099_ | ~new_n20693_;
  assign new_n20987_ = ~new_n20789_ | ~new_n20985_;
  assign new_n20988_ = ~new_n4678_ | ~new_n20691_;
  assign new_n20989_ = ~new_n20827_ | ~new_n20988_;
  assign new_n20990_ = ~new_n4693_ | ~new_n20667_;
  assign new_n20991_ = ~new_n4694_ | ~new_n20809_;
  assign new_n20992_ = ~new_n4698_ | ~new_n20812_;
  assign new_n20993_ = ~new_n20772_ | ~new_n20771_ | ~new_n20946_;
  assign new_n20994_ = ~new_n5093_ | ~new_n20684_;
  assign new_n20995_ = ~new_n4699_ | ~new_n20683_;
  assign new_n20996_ = ~new_n20864_ | ~new_n20792_;
  assign new_n20997_ = ~new_n20862_ | ~new_n20791_;
  assign new_n20998_ = ~new_n5090_ | ~new_n20682_;
  assign new_n20999_ = ~new_n4700_ | ~new_n20679_;
  assign new_n21000_ = ~new_n5090_ | ~new_n20682_;
  assign new_n21001_ = ~new_n4700_ | ~new_n20679_;
  assign new_n21002_ = ~new_n21001_ | ~new_n21000_;
  assign new_n21003_ = ~new_n5087_ | ~new_n20680_;
  assign new_n21004_ = ~new_n4686_ | ~new_n20664_;
  assign new_n21005_ = ~new_n20869_ | ~new_n20685_;
  assign new_n21006_ = ~new_n20793_ | ~new_n20856_;
  assign new_n21007_ = ~new_n5084_ | ~new_n20675_;
  assign new_n21008_ = ~new_n4687_ | ~new_n20673_;
  assign new_n21009_ = ~new_n21008_ | ~new_n21007_;
  assign new_n21010_ = ~new_n5081_ | ~new_n20676_;
  assign new_n21011_ = ~new_n4683_ | ~new_n20665_;
  assign new_n21012_ = ~new_n20879_ | ~new_n20686_;
  assign new_n21013_ = ~new_n20794_ | ~new_n20871_;
  assign new_n21014_ = ~new_n5078_ | ~new_n20677_;
  assign new_n21015_ = ~new_n4676_ | ~new_n20674_;
  assign new_n21016_ = ~new_n20880_ | ~new_n20796_;
  assign new_n21017_ = ~new_n20846_ | ~new_n20795_;
  assign new_n21018_ = ~new_n5075_ | ~new_n20672_;
  assign new_n21019_ = ~new_n4680_ | ~new_n20669_;
  assign new_n21020_ = ~new_n5075_ | ~new_n20672_;
  assign new_n21021_ = ~new_n4680_ | ~new_n20669_;
  assign new_n21022_ = ~new_n21021_ | ~new_n21020_;
  assign new_n21023_ = ~new_n5072_ | ~new_n20670_;
  assign new_n21024_ = ~new_n4684_ | ~new_n20666_;
  assign new_n21025_ = ~new_n20885_ | ~new_n20687_;
  assign new_n21026_ = ~new_n20797_ | ~new_n20840_;
  assign new_n21027_ = ~new_n5595_ | ~new_n20799_;
  assign new_n21028_ = ~new_n4671_ | ~new_n20798_;
  assign new_n21029_ = ~new_n5595_ | ~new_n20799_;
  assign new_n21030_ = ~new_n4671_ | ~new_n20798_;
  assign new_n21031_ = ~new_n21030_ | ~new_n21029_;
  assign new_n21032_ = ~new_n20728_ | ~new_n5584_ | ~new_n20654_;
  assign new_n21033_ = ~new_n4670_ | ~new_n21031_ | ~new_n20727_;
  assign new_n21034_ = ~new_n5584_ | ~new_n20728_;
  assign new_n21035_ = ~new_n4670_ | ~new_n20727_;
  assign new_n21036_ = ~new_n20773_;
  assign new_n21037_ = ~new_n20950_ | ~new_n21036_;
  assign new_n21038_ = ~new_n20773_ | ~new_n20801_;
  assign new_n21039_ = ~new_n5585_ | ~new_n20726_;
  assign new_n21040_ = ~new_n4669_ | ~new_n20723_;
  assign new_n21041_ = ~new_n5585_ | ~new_n20726_;
  assign new_n21042_ = ~new_n4669_ | ~new_n20723_;
  assign new_n21043_ = ~new_n21042_ | ~new_n21041_;
  assign new_n21044_ = ~new_n5586_ | ~new_n20724_;
  assign new_n21045_ = ~new_n4673_ | ~new_n20688_;
  assign new_n21046_ = ~new_n20957_ | ~new_n20729_;
  assign new_n21047_ = ~new_n20802_ | ~new_n20944_;
  assign new_n21048_ = ~new_n5587_ | ~new_n20722_;
  assign new_n21049_ = ~new_n4674_ | ~new_n20721_;
  assign new_n21050_ = ~new_n20776_;
  assign new_n21051_ = ~new_n20940_ | ~new_n21050_;
  assign new_n21052_ = ~new_n20776_ | ~new_n20803_;
  assign new_n21053_ = ~new_n5588_ | ~new_n20720_;
  assign new_n21054_ = ~new_n4681_ | ~new_n20719_;
  assign new_n21055_ = ~new_n20777_;
  assign new_n21056_ = ~new_n20936_ | ~new_n21055_;
  assign new_n21057_ = ~new_n20777_ | ~new_n20804_;
  assign new_n21058_ = ~new_n5589_ | ~new_n20715_;
  assign new_n21059_ = ~new_n4682_ | ~new_n20713_;
  assign new_n21060_ = ~new_n21059_ | ~new_n21058_;
  assign new_n21061_ = ~new_n5590_ | ~new_n20716_;
  assign new_n21062_ = ~new_n4677_ | ~new_n20689_;
endmodule



// Benchmark "b22" written by ABC on Sun Apr 23 00:37:58 2023

module b22 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519,
    pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549,
    pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559,
    pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569,
    pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579,
    pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589,
    pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599,
    pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609,
    pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639,
    pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649,
    pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659,
    pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669,
    pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679,
    pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689,
    pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699,
    pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729,
    pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739,
    pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749,
    pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759,
    pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518, po519,
    po520, po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548, po549,
    po550, po551, po552, po553, po554, po555, po556, po557, po558, po559,
    po560, po561, po562, po563, po564, po565, po566, po567, po568, po569,
    po570, po571, po572, po573, po574, po575, po576, po577, po578, po579,
    po580, po581, po582, po583, po584, po585, po586, po587, po588, po589,
    po590, po591, po592, po593, po594, po595, po596, po597, po598, po599,
    po600, po601, po602, po603, po604, po605, po606, po607, po608, po609,
    po610, po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638, po639,
    po640, po641, po642, po643, po644, po645, po646, po647, po648, po649,
    po650, po651, po652, po653, po654, po655, po656, po657, po658, po659,
    po660, po661, po662, po663, po664, po665, po666, po667, po668, po669,
    po670, po671, po672, po673, po674, po675, po676, po677, po678, po679,
    po680, po681, po682, po683, po684, po685, po686, po687, po688, po689,
    po690, po691, po692, po693, po694, po695, po696, po697, po698, po699,
    po700, po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728, po729,
    po730, po731, po732, po733, po734, po735, po736, po737, po738, po739,
    po740, po741, po742, po743, po744, po745, po746, po747, po748, po749,
    po750, po751, po752, po753, po754, po755, po756  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518,
    pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528,
    pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558,
    pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568,
    pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578,
    pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588,
    pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598,
    pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608,
    pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618,
    pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648,
    pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658,
    pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668,
    pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678,
    pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688,
    pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698,
    pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708,
    pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738,
    pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748,
    pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758,
    pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518, po519,
    po520, po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548, po549,
    po550, po551, po552, po553, po554, po555, po556, po557, po558, po559,
    po560, po561, po562, po563, po564, po565, po566, po567, po568, po569,
    po570, po571, po572, po573, po574, po575, po576, po577, po578, po579,
    po580, po581, po582, po583, po584, po585, po586, po587, po588, po589,
    po590, po591, po592, po593, po594, po595, po596, po597, po598, po599,
    po600, po601, po602, po603, po604, po605, po606, po607, po608, po609,
    po610, po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638, po639,
    po640, po641, po642, po643, po644, po645, po646, po647, po648, po649,
    po650, po651, po652, po653, po654, po655, po656, po657, po658, po659,
    po660, po661, po662, po663, po664, po665, po666, po667, po668, po669,
    po670, po671, po672, po673, po674, po675, po676, po677, po678, po679,
    po680, po681, po682, po683, po684, po685, po686, po687, po688, po689,
    po690, po691, po692, po693, po694, po695, po696, po697, po698, po699,
    po700, po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728, po729,
    po730, po731, po732, po733, po734, po735, po736, po737, po738, po739,
    po740, po741, po742, po743, po744, po745, po746, po747, po748, po749,
    po750, po751, po752, po753, po754, po755, po756;
  wire new_n1526_, new_n1527_, new_n1528_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_,
    new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_,
    new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2387_, new_n2388_, new_n2390_,
    new_n2391_, new_n2393_, new_n2394_, new_n2396_, new_n2397_, new_n2399_,
    new_n2400_, new_n2402_, new_n2403_, new_n2405_, new_n2406_, new_n2408_,
    new_n2409_, new_n2411_, new_n2412_, new_n2414_, new_n2415_, new_n2417_,
    new_n2418_, new_n2420_, new_n2421_, new_n2423_, new_n2424_, new_n2426_,
    new_n2427_, new_n2429_, new_n2430_, new_n2432_, new_n2433_, new_n2435_,
    new_n2436_, new_n2438_, new_n2439_, new_n2441_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_,
    new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_,
    new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_,
    new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_,
    new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_,
    new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_,
    new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_,
    new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_,
    new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_,
    new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_,
    new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_,
    new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_,
    new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_,
    new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_,
    new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_,
    new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_,
    new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_,
    new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_,
    new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_,
    new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_,
    new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_,
    new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_,
    new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_,
    new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_,
    new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_,
    new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_,
    new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_,
    new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_,
    new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_,
    new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_,
    new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_,
    new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_,
    new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_,
    new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_,
    new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_,
    new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_,
    new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_,
    new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_,
    new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_,
    new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_,
    new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_,
    new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_,
    new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_,
    new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_,
    new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_,
    new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_,
    new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_,
    new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_,
    new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_,
    new_n5404_, new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_,
    new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_,
    new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_,
    new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_,
    new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_,
    new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_,
    new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_,
    new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_,
    new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5651_, new_n5652_,
    new_n5654_, new_n5655_, new_n5657_, new_n5658_, new_n5660_, new_n5661_,
    new_n5663_, new_n5664_, new_n5666_, new_n5667_, new_n5669_, new_n5670_,
    new_n5672_, new_n5673_, new_n5675_, new_n5676_, new_n5678_, new_n5679_,
    new_n5681_, new_n5682_, new_n5684_, new_n5685_, new_n5687_, new_n5688_,
    new_n5690_, new_n5691_, new_n5693_, new_n5694_, new_n5696_, new_n5697_,
    new_n5699_, new_n5700_, new_n5702_, new_n5703_, new_n5705_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_,
    new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_,
    new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_,
    new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_,
    new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_,
    new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_,
    new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_,
    new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_,
    new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_,
    new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_,
    new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_,
    new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_,
    new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_,
    new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_,
    new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_,
    new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_,
    new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_,
    new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_,
    new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_,
    new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_,
    new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_,
    new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_,
    new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_,
    new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_,
    new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_,
    new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_,
    new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_,
    new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_,
    new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_,
    new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_,
    new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_,
    new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_,
    new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_,
    new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_,
    new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_,
    new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_,
    new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_,
    new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_,
    new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_,
    new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_,
    new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_,
    new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_,
    new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_,
    new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_,
    new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_,
    new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_,
    new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_,
    new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_,
    new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_,
    new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_,
    new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_,
    new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_,
    new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_,
    new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_,
    new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_,
    new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_,
    new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_,
    new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_,
    new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_,
    new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_,
    new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_,
    new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_,
    new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_,
    new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_,
    new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_,
    new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_,
    new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_,
    new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_,
    new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_,
    new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_,
    new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_,
    new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_,
    new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_,
    new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_,
    new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_,
    new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_,
    new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_,
    new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_,
    new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_,
    new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_,
    new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_,
    new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_,
    new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_,
    new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_,
    new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_,
    new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_,
    new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_,
    new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_,
    new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_,
    new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_,
    new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_,
    new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_,
    new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_,
    new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_,
    new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_,
    new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_,
    new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_,
    new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_,
    new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_,
    new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_,
    new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_,
    new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_,
    new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_,
    new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_,
    new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_,
    new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_,
    new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_,
    new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_,
    new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_,
    new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_,
    new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_,
    new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_,
    new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_,
    new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_,
    new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_,
    new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_,
    new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_,
    new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_,
    new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_,
    new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_,
    new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_,
    new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_,
    new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_,
    new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_,
    new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_,
    new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_,
    new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_,
    new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_,
    new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_,
    new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_,
    new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_,
    new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_,
    new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_,
    new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_,
    new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_,
    new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_,
    new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_,
    new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_,
    new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_,
    new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_,
    new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_,
    new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_,
    new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_,
    new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_,
    new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_,
    new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_,
    new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_,
    new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_,
    new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_,
    new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_,
    new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_,
    new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_,
    new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_,
    new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_,
    new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_,
    new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_,
    new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_,
    new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_,
    new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_,
    new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_,
    new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_,
    new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_,
    new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_,
    new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_,
    new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_,
    new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_,
    new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_,
    new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_,
    new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_,
    new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_,
    new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_,
    new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_,
    new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_,
    new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_,
    new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_,
    new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_,
    new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_,
    new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_,
    new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_,
    new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_,
    new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_,
    new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_,
    new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_,
    new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_,
    new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_,
    new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_,
    new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_,
    new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_,
    new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_,
    new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_,
    new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_,
    new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_,
    new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_,
    new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_,
    new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_,
    new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_,
    new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_,
    new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_,
    new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_,
    new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_,
    new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_,
    new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_,
    new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_,
    new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_,
    new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_,
    new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8530_, new_n8675_, new_n8676_, new_n8677_, new_n8678_,
    new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_,
    new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_,
    new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_,
    new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_,
    new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_,
    new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_,
    new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_,
    new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_,
    new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_,
    new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_,
    new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_,
    new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_,
    new_n8751_, new_n8752_, new_n8753_, new_n8756_, new_n8757_, new_n8758_,
    new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_,
    new_n8765_, new_n8766_, new_n8767_, new_n8769_, new_n8770_, new_n8772_,
    new_n8773_, new_n8775_, new_n8776_, new_n8778_, new_n8779_, new_n8781_,
    new_n8782_, new_n8784_, new_n8785_, new_n8787_, new_n8788_, new_n8790_,
    new_n8791_, new_n8793_, new_n8794_, new_n8796_, new_n8797_, new_n8799_,
    new_n8800_, new_n8802_, new_n8803_, new_n8805_, new_n8806_, new_n8808_,
    new_n8809_, new_n8811_, new_n8812_, new_n8814_, new_n8815_, new_n8817_,
    new_n8818_, new_n8820_, new_n8821_, new_n8823_, new_n8901_, new_n8902_,
    new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_,
    new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_,
    new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_,
    new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_,
    new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_,
    new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_,
    new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_,
    new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_,
    new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_,
    new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_,
    new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_,
    new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_,
    new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_,
    new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_,
    new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_,
    new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_,
    new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_,
    new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_,
    new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_,
    new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_,
    new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_,
    new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_,
    new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_,
    new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_,
    new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_,
    new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_,
    new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_,
    new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_,
    new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_,
    new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_,
    new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_,
    new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_,
    new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_,
    new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_,
    new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_,
    new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_,
    new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_,
    new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_,
    new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_,
    new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_,
    new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_,
    new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_,
    new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_,
    new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_,
    new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_,
    new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_,
    new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_,
    new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_,
    new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_,
    new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_,
    new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_,
    new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_,
    new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_,
    new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_,
    new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_,
    new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_,
    new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_,
    new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_,
    new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_,
    new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_,
    new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_,
    new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_,
    new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_,
    new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_,
    new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_,
    new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_,
    new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_,
    new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_,
    new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_,
    new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_,
    new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_,
    new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_,
    new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_,
    new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_,
    new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_,
    new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_,
    new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_,
    new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_,
    new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_,
    new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_,
    new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_,
    new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_,
    new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_,
    new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_,
    new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_,
    new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_,
    new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_,
    new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_,
    new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_,
    new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_,
    new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_,
    new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_,
    new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_,
    new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_,
    new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_,
    new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_,
    new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12147_, new_n12148_, new_n12149_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12333_, new_n12334_, new_n12335_,
    new_n12336_, new_n12337_, new_n12338_, new_n12339_, new_n12340_,
    new_n12341_, new_n12342_, new_n12343_, new_n12344_, new_n12345_,
    new_n12346_, new_n12347_, new_n12348_, new_n12349_, new_n12350_,
    new_n12351_, new_n12352_, new_n12353_, new_n12354_, new_n12355_,
    new_n12356_, new_n12357_, new_n12358_, new_n12359_, new_n12360_,
    new_n12361_, new_n12362_, new_n12363_, new_n12364_, new_n12365_,
    new_n12366_, new_n12367_, new_n12368_, new_n12369_, new_n12370_,
    new_n12371_, new_n12372_, new_n12373_, new_n12374_, new_n12375_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12384_, new_n12385_,
    new_n12386_, new_n12387_, new_n12388_, new_n12389_, new_n12390_,
    new_n12391_, new_n12392_, new_n12393_, new_n12394_, new_n12395_,
    new_n12396_, new_n12397_, new_n12398_, new_n12399_, new_n12400_,
    new_n12401_, new_n12402_, new_n12403_, new_n12404_, new_n12405_,
    new_n12406_, new_n12407_, new_n12408_, new_n12409_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12420_,
    new_n12421_, new_n12422_, new_n12423_, new_n12424_, new_n12425_,
    new_n12426_, new_n12427_, new_n12428_, new_n12429_, new_n12430_,
    new_n12431_, new_n12432_, new_n12433_, new_n12434_, new_n12435_,
    new_n12436_, new_n12437_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14075_,
    new_n14076_, new_n14077_, new_n14078_, new_n14079_, new_n14080_,
    new_n14081_, new_n14082_, new_n14083_, new_n14084_, new_n14085_,
    new_n14086_, new_n14087_, new_n14088_, new_n14089_, new_n14090_,
    new_n14091_, new_n14092_, new_n14093_, new_n14094_, new_n14095_,
    new_n14096_, new_n14097_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14103_, new_n14104_, new_n14105_,
    new_n14106_, new_n14107_, new_n14108_, new_n14109_, new_n14110_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14117_, new_n14118_, new_n14119_, new_n14120_,
    new_n14121_, new_n14122_, new_n14123_, new_n14124_, new_n14125_,
    new_n14126_, new_n14127_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14133_, new_n14134_, new_n14135_,
    new_n14136_, new_n14137_, new_n14138_, new_n14139_, new_n14140_,
    new_n14141_, new_n14142_, new_n14143_, new_n14144_, new_n14145_,
    new_n14146_, new_n14147_, new_n14148_, new_n14149_, new_n14150_,
    new_n14151_, new_n14152_, new_n14153_, new_n14154_, new_n14155_,
    new_n14156_, new_n14157_, new_n14158_, new_n14159_, new_n14160_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14205_,
    new_n14206_, new_n14207_, new_n14208_, new_n14209_, new_n14210_,
    new_n14211_, new_n14212_, new_n14213_, new_n14214_, new_n14215_,
    new_n14216_, new_n14217_, new_n14218_, new_n14219_, new_n14220_,
    new_n14221_, new_n14222_, new_n14223_, new_n14224_, new_n14225_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14241_, new_n14242_, new_n14243_, new_n14244_, new_n14245_,
    new_n14246_, new_n14247_, new_n14248_, new_n14249_, new_n14250_,
    new_n14251_, new_n14252_, new_n14253_, new_n14254_, new_n14255_,
    new_n14256_, new_n14257_, new_n14258_, new_n14259_, new_n14260_,
    new_n14261_, new_n14262_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14268_, new_n14269_, new_n14270_,
    new_n14271_, new_n14272_, new_n14273_, new_n14274_, new_n14275_,
    new_n14276_, new_n14277_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14284_, new_n14285_,
    new_n14286_, new_n14287_, new_n14288_, new_n14289_, new_n14290_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14342_, new_n14343_, new_n14344_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14416_, new_n14417_, new_n14418_, new_n14419_, new_n14420_,
    new_n14421_, new_n14422_, new_n14423_, new_n14424_, new_n14425_,
    new_n14426_, new_n14427_, new_n14428_, new_n14429_, new_n14430_,
    new_n14431_, new_n14432_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14465_,
    new_n14466_, new_n14467_, new_n14468_, new_n14469_, new_n14470_,
    new_n14471_, new_n14472_, new_n14473_, new_n14474_, new_n14475_,
    new_n14476_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14481_, new_n14482_, new_n14483_, new_n14484_, new_n14485_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14595_,
    new_n14596_, new_n14597_, new_n14598_, new_n14599_, new_n14600_,
    new_n14601_, new_n14602_, new_n14603_, new_n14604_, new_n14605_,
    new_n14606_, new_n14607_, new_n14608_, new_n14609_, new_n14610_,
    new_n14611_, new_n14612_, new_n14613_, new_n14614_, new_n14615_,
    new_n14616_, new_n14617_, new_n14618_, new_n14619_, new_n14620_,
    new_n14621_, new_n14622_, new_n14623_, new_n14624_, new_n14625_,
    new_n14626_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14840_,
    new_n14841_, new_n14842_, new_n14843_, new_n14844_, new_n14845_,
    new_n14846_, new_n14847_, new_n14848_, new_n14849_, new_n14850_,
    new_n14851_, new_n14852_, new_n14853_, new_n14854_, new_n14855_,
    new_n14856_, new_n14857_, new_n14858_, new_n14859_, new_n14860_,
    new_n14861_, new_n14862_, new_n14863_, new_n14864_, new_n14865_,
    new_n14866_, new_n14867_, new_n14868_, new_n14869_, new_n14870_,
    new_n14871_, new_n14872_, new_n14873_, new_n14874_, new_n14875_,
    new_n14876_, new_n14877_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14887_, new_n14888_, new_n14889_, new_n14890_,
    new_n14891_, new_n14892_, new_n14893_, new_n14894_, new_n14895_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14902_, new_n14903_, new_n14904_, new_n14905_,
    new_n14906_, new_n14907_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15328_, new_n15329_, new_n15330_,
    new_n15331_, new_n15332_, new_n15333_, new_n15334_, new_n15335_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15381_, new_n15382_, new_n15383_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15390_,
    new_n15391_, new_n15392_, new_n15393_, new_n15394_, new_n15395_,
    new_n15396_, new_n15397_, new_n15398_, new_n15399_, new_n15400_,
    new_n15401_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15438_, new_n15439_, new_n15440_,
    new_n15441_, new_n15442_, new_n15443_, new_n15444_, new_n15445_,
    new_n15446_, new_n15447_, new_n15448_, new_n15449_, new_n15450_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15494_, new_n15495_,
    new_n15496_, new_n15497_, new_n15498_, new_n15499_, new_n15500_,
    new_n15501_, new_n15502_, new_n15503_, new_n15504_, new_n15505_,
    new_n15506_, new_n15507_, new_n15508_, new_n15509_, new_n15510_,
    new_n15511_, new_n15512_, new_n15513_, new_n15514_, new_n15515_,
    new_n15516_, new_n15517_, new_n15518_, new_n15519_, new_n15520_,
    new_n15521_, new_n15522_, new_n15523_, new_n15524_, new_n15525_,
    new_n15526_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15531_, new_n15532_, new_n15533_, new_n15534_, new_n15535_,
    new_n15536_, new_n15537_, new_n15538_, new_n15539_, new_n15540_,
    new_n15541_, new_n15542_, new_n15543_, new_n15544_, new_n15545_,
    new_n15546_, new_n15547_, new_n15548_, new_n15549_, new_n15550_,
    new_n15551_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16349_, new_n16350_,
    new_n16351_, new_n16352_, new_n16353_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16361_, new_n16362_, new_n16363_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16489_, new_n16490_,
    new_n16491_, new_n16492_, new_n16493_, new_n16494_, new_n16495_,
    new_n16496_, new_n16497_, new_n16498_, new_n16499_, new_n16500_,
    new_n16501_, new_n16502_, new_n16503_, new_n16504_, new_n16505_,
    new_n16506_, new_n16507_, new_n16508_, new_n16509_, new_n16510_,
    new_n16511_, new_n16512_, new_n16513_, new_n16514_, new_n16515_,
    new_n16516_, new_n16517_, new_n16518_, new_n16519_, new_n16520_,
    new_n16521_, new_n16522_, new_n16523_, new_n16524_, new_n16525_,
    new_n16526_, new_n16527_, new_n16528_, new_n16529_, new_n16530_,
    new_n16531_, new_n16532_, new_n16533_, new_n16534_, new_n16535_,
    new_n16536_, new_n16537_, new_n16538_, new_n16539_, new_n16540_,
    new_n16541_, new_n16542_, new_n16543_, new_n16544_, new_n16545_,
    new_n16546_, new_n16547_, new_n16548_, new_n16549_, new_n16550_,
    new_n16551_, new_n16552_, new_n16553_, new_n16554_, new_n16555_,
    new_n16556_, new_n16557_, new_n16558_, new_n16559_, new_n16560_,
    new_n16561_, new_n16562_, new_n16563_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16618_, new_n16619_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16659_, new_n16660_,
    new_n16661_, new_n16662_, new_n16663_, new_n16664_, new_n16665_,
    new_n16666_, new_n16667_, new_n16668_, new_n16669_, new_n16670_,
    new_n16671_, new_n16672_, new_n16673_, new_n16674_, new_n16675_,
    new_n16676_, new_n16677_, new_n16678_, new_n16679_, new_n16680_,
    new_n16681_, new_n16682_, new_n16683_, new_n16684_, new_n16685_,
    new_n16686_, new_n16687_, new_n16688_, new_n16689_, new_n16690_,
    new_n16691_, new_n16692_, new_n16693_, new_n16694_, new_n16695_,
    new_n16696_, new_n16697_, new_n16698_, new_n16699_, new_n16700_,
    new_n16701_, new_n16702_, new_n16703_, new_n16704_, new_n16705_,
    new_n16706_, new_n16707_, new_n16708_, new_n16709_, new_n16710_,
    new_n16711_, new_n16712_, new_n16713_, new_n16714_, new_n16715_,
    new_n16716_, new_n16717_, new_n16718_, new_n16719_, new_n16720_,
    new_n16721_, new_n16722_, new_n16723_, new_n16724_, new_n16725_,
    new_n16726_, new_n16727_, new_n16728_, new_n16729_, new_n16730_,
    new_n16731_, new_n16732_, new_n16733_, new_n16734_, new_n16735_,
    new_n16736_, new_n16737_, new_n16738_, new_n16739_, new_n16740_,
    new_n16741_, new_n16742_, new_n16743_, new_n16744_, new_n16745_,
    new_n16746_, new_n16747_, new_n16748_, new_n16749_, new_n16750_,
    new_n16751_, new_n16752_, new_n16753_, new_n16754_, new_n16755_,
    new_n16756_, new_n16757_, new_n16758_, new_n16759_, new_n16760_,
    new_n16761_, new_n16762_, new_n16763_, new_n16764_, new_n16765_,
    new_n16766_, new_n16767_, new_n16768_, new_n16769_, new_n16770_,
    new_n16771_, new_n16772_, new_n16773_, new_n16774_, new_n16775_,
    new_n16776_, new_n16777_, new_n16778_, new_n16779_, new_n16780_,
    new_n16781_, new_n16782_, new_n16783_, new_n16784_, new_n16785_,
    new_n16786_, new_n16787_, new_n16788_, new_n16789_, new_n16790_,
    new_n16791_, new_n16792_, new_n16793_, new_n16794_, new_n16795_,
    new_n16796_, new_n16797_, new_n16798_, new_n16799_, new_n16800_,
    new_n16801_, new_n16802_, new_n16803_, new_n16804_, new_n16805_,
    new_n16806_, new_n16807_, new_n16808_, new_n16809_, new_n16810_,
    new_n16811_, new_n16812_, new_n16813_, new_n16814_, new_n16815_,
    new_n16816_, new_n16817_, new_n16818_, new_n16819_, new_n16820_,
    new_n16821_, new_n16822_, new_n16823_, new_n16824_, new_n16825_,
    new_n16826_, new_n16827_, new_n16828_, new_n16829_, new_n16830_,
    new_n16831_, new_n16832_, new_n16833_, new_n16834_, new_n16835_,
    new_n16836_, new_n16837_, new_n16838_, new_n16839_, new_n16840_,
    new_n16841_, new_n16842_, new_n16843_, new_n16844_, new_n16845_,
    new_n16846_, new_n16847_, new_n16848_, new_n16849_, new_n16850_,
    new_n16851_, new_n16852_, new_n16853_, new_n16854_, new_n16855_,
    new_n16856_, new_n16857_, new_n16858_, new_n16859_, new_n16860_,
    new_n16861_, new_n16862_, new_n16863_, new_n16864_, new_n16865_,
    new_n16866_, new_n16867_, new_n16868_, new_n16869_, new_n16870_,
    new_n16871_, new_n16872_, new_n16873_, new_n16874_, new_n16875_,
    new_n16876_, new_n16877_, new_n16878_, new_n16879_, new_n16880_,
    new_n16881_, new_n16882_, new_n16883_, new_n16884_, new_n16885_,
    new_n16886_, new_n16887_, new_n16888_, new_n16889_, new_n16890_,
    new_n16891_, new_n16892_, new_n16893_, new_n16894_, new_n16895_,
    new_n16896_, new_n16897_, new_n16898_, new_n16899_, new_n16900_,
    new_n16901_, new_n16902_, new_n16903_, new_n16904_, new_n16905_,
    new_n16906_, new_n16907_, new_n16908_, new_n16909_, new_n16910_,
    new_n16911_, new_n16912_, new_n16913_, new_n16914_, new_n16915_,
    new_n16916_, new_n16917_, new_n16918_, new_n16919_, new_n16920_,
    new_n16921_, new_n16922_, new_n16923_, new_n16924_, new_n16925_,
    new_n16926_, new_n16927_, new_n16928_, new_n16929_, new_n16930_,
    new_n16931_, new_n16932_, new_n16933_, new_n16934_, new_n16935_,
    new_n16936_, new_n16937_, new_n16938_, new_n16939_, new_n16940_,
    new_n16941_, new_n16942_, new_n16943_, new_n16944_, new_n16945_,
    new_n16946_, new_n16947_, new_n16948_, new_n16949_, new_n16950_,
    new_n16951_, new_n16952_, new_n16953_, new_n16954_, new_n16955_,
    new_n16956_, new_n16957_, new_n16958_, new_n16959_, new_n16960_,
    new_n16961_, new_n16962_, new_n16963_, new_n16964_, new_n16965_,
    new_n16966_, new_n16967_, new_n16968_, new_n16969_, new_n16970_,
    new_n16971_, new_n16972_, new_n16973_, new_n16974_, new_n16975_,
    new_n16976_, new_n16977_, new_n16978_, new_n16979_, new_n16980_,
    new_n16981_, new_n16982_, new_n16983_, new_n16984_, new_n16985_,
    new_n16986_, new_n16987_, new_n16988_, new_n16989_, new_n16990_,
    new_n16991_, new_n16992_, new_n16993_, new_n16994_, new_n16995_,
    new_n16996_, new_n16997_, new_n16998_, new_n16999_, new_n17000_,
    new_n17001_, new_n17002_, new_n17003_, new_n17004_, new_n17005_,
    new_n17006_, new_n17007_, new_n17008_, new_n17009_, new_n17010_,
    new_n17011_, new_n17012_, new_n17013_, new_n17014_, new_n17015_,
    new_n17016_, new_n17017_, new_n17018_, new_n17019_, new_n17020_,
    new_n17021_, new_n17022_, new_n17023_, new_n17024_, new_n17025_,
    new_n17026_, new_n17027_, new_n17028_, new_n17029_, new_n17030_,
    new_n17031_, new_n17032_, new_n17033_, new_n17034_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17039_, new_n17040_,
    new_n17041_, new_n17042_, new_n17043_, new_n17044_, new_n17045_,
    new_n17046_, new_n17047_, new_n17048_, new_n17049_, new_n17050_,
    new_n17051_, new_n17052_, new_n17053_, new_n17054_, new_n17055_,
    new_n17056_, new_n17057_, new_n17058_, new_n17059_, new_n17060_,
    new_n17061_, new_n17062_, new_n17063_, new_n17064_, new_n17065_,
    new_n17066_, new_n17067_, new_n17068_, new_n17069_, new_n17070_,
    new_n17071_, new_n17072_, new_n17073_, new_n17074_, new_n17075_,
    new_n17076_, new_n17077_, new_n17078_, new_n17079_, new_n17080_,
    new_n17081_, new_n17082_, new_n17083_, new_n17084_, new_n17085_,
    new_n17086_, new_n17087_, new_n17088_, new_n17089_, new_n17090_,
    new_n17091_, new_n17092_, new_n17093_, new_n17094_, new_n17095_,
    new_n17096_, new_n17097_, new_n17098_, new_n17099_, new_n17100_,
    new_n17101_, new_n17102_, new_n17103_, new_n17104_, new_n17105_,
    new_n17106_, new_n17107_, new_n17108_, new_n17109_, new_n17110_,
    new_n17111_, new_n17112_, new_n17113_, new_n17114_, new_n17115_,
    new_n17116_, new_n17117_, new_n17118_, new_n17119_, new_n17120_,
    new_n17121_, new_n17122_, new_n17123_, new_n17124_, new_n17125_,
    new_n17126_, new_n17127_, new_n17128_, new_n17129_, new_n17130_,
    new_n17131_, new_n17132_, new_n17133_, new_n17134_, new_n17135_,
    new_n17136_, new_n17137_, new_n17138_, new_n17139_, new_n17140_,
    new_n17141_, new_n17142_, new_n17143_, new_n17144_, new_n17145_,
    new_n17146_, new_n17147_, new_n17148_, new_n17149_, new_n17150_,
    new_n17151_, new_n17152_, new_n17153_, new_n17154_, new_n17155_,
    new_n17156_, new_n17157_, new_n17158_, new_n17159_, new_n17160_,
    new_n17161_, new_n17162_, new_n17163_, new_n17164_, new_n17165_,
    new_n17166_, new_n17167_, new_n17168_, new_n17169_, new_n17170_,
    new_n17171_, new_n17172_, new_n17173_, new_n17174_, new_n17175_,
    new_n17176_, new_n17177_, new_n17178_, new_n17179_, new_n17180_,
    new_n17181_, new_n17182_, new_n17183_, new_n17184_, new_n17185_,
    new_n17186_, new_n17187_, new_n17188_, new_n17189_, new_n17190_,
    new_n17191_, new_n17192_, new_n17193_, new_n17194_, new_n17195_,
    new_n17196_, new_n17197_, new_n17198_, new_n17199_, new_n17200_,
    new_n17201_, new_n17202_, new_n17203_, new_n17204_, new_n17205_,
    new_n17206_, new_n17207_, new_n17208_, new_n17209_, new_n17210_,
    new_n17211_, new_n17212_, new_n17213_, new_n17214_, new_n17215_,
    new_n17216_, new_n17217_, new_n17218_, new_n17219_, new_n17220_,
    new_n17221_, new_n17222_, new_n17223_, new_n17224_, new_n17225_,
    new_n17226_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17233_, new_n17234_, new_n17235_,
    new_n17236_, new_n17237_, new_n17238_, new_n17239_, new_n17240_,
    new_n17241_, new_n17242_, new_n17243_, new_n17244_, new_n17245_,
    new_n17246_, new_n17247_, new_n17248_, new_n17249_, new_n17250_,
    new_n17251_, new_n17252_, new_n17253_, new_n17254_, new_n17255_,
    new_n17256_, new_n17257_, new_n17258_, new_n17259_, new_n17260_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17283_, new_n17284_, new_n17285_,
    new_n17286_, new_n17287_, new_n17288_, new_n17289_, new_n17290_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17345_,
    new_n17346_, new_n17347_, new_n17348_, new_n17349_, new_n17350_,
    new_n17351_, new_n17352_, new_n17353_, new_n17354_, new_n17355_,
    new_n17356_, new_n17357_, new_n17358_, new_n17359_, new_n17360_,
    new_n17361_, new_n17362_, new_n17363_, new_n17364_, new_n17365_,
    new_n17366_, new_n17367_, new_n17368_, new_n17369_, new_n17370_,
    new_n17371_, new_n17372_, new_n17373_, new_n17374_, new_n17375_,
    new_n17376_, new_n17377_, new_n17378_, new_n17379_, new_n17380_,
    new_n17381_, new_n17382_, new_n17383_, new_n17384_, new_n17385_,
    new_n17386_, new_n17387_, new_n17388_, new_n17389_, new_n17390_,
    new_n17391_, new_n17392_, new_n17393_, new_n17394_, new_n17395_,
    new_n17396_, new_n17397_, new_n17398_, new_n17399_, new_n17400_,
    new_n17401_, new_n17402_, new_n17403_, new_n17404_, new_n17405_,
    new_n17406_, new_n17407_, new_n17408_, new_n17409_, new_n17410_,
    new_n17411_, new_n17412_, new_n17413_, new_n17414_, new_n17415_,
    new_n17416_, new_n17417_, new_n17418_, new_n17419_, new_n17420_,
    new_n17421_, new_n17422_, new_n17423_, new_n17424_, new_n17425_,
    new_n17426_, new_n17427_, new_n17428_, new_n17429_, new_n17430_,
    new_n17431_, new_n17432_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17438_, new_n17439_, new_n17440_,
    new_n17441_, new_n17442_, new_n17443_, new_n17444_, new_n17445_,
    new_n17446_, new_n17447_, new_n17448_, new_n17449_, new_n17450_,
    new_n17451_, new_n17452_, new_n17453_, new_n17454_, new_n17455_,
    new_n17456_, new_n17457_, new_n17458_, new_n17459_, new_n17460_,
    new_n17461_, new_n17462_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17468_, new_n17469_, new_n17470_,
    new_n17471_, new_n17472_, new_n17473_, new_n17474_, new_n17475_,
    new_n17476_, new_n17477_, new_n17478_, new_n17479_, new_n17480_,
    new_n17481_, new_n17482_, new_n17483_, new_n17484_, new_n17485_,
    new_n17486_, new_n17487_, new_n17488_, new_n17489_, new_n17490_,
    new_n17491_, new_n17492_, new_n17493_, new_n17494_, new_n17495_,
    new_n17496_, new_n17497_, new_n17498_, new_n17499_, new_n17500_,
    new_n17501_, new_n17502_, new_n17503_, new_n17504_, new_n17505_,
    new_n17506_, new_n17507_, new_n17508_, new_n17509_, new_n17510_,
    new_n17511_, new_n17512_, new_n17513_, new_n17514_, new_n17515_,
    new_n17516_, new_n17517_, new_n17518_, new_n17519_, new_n17520_,
    new_n17521_, new_n17522_, new_n17523_, new_n17524_, new_n17525_,
    new_n17526_, new_n17527_, new_n17528_, new_n17529_, new_n17530_,
    new_n17531_, new_n17532_, new_n17533_, new_n17534_, new_n17535_,
    new_n17536_, new_n17537_, new_n17538_, new_n17539_, new_n17540_,
    new_n17541_, new_n17542_, new_n17543_, new_n17544_, new_n17545_,
    new_n17546_, new_n17547_, new_n17548_, new_n17549_, new_n17550_,
    new_n17551_, new_n17552_, new_n17553_, new_n17554_, new_n17555_,
    new_n17556_, new_n17557_, new_n17558_, new_n17559_, new_n17560_,
    new_n17561_, new_n17562_, new_n17563_, new_n17564_, new_n17565_,
    new_n17566_, new_n17567_, new_n17568_, new_n17569_, new_n17570_,
    new_n17571_, new_n17572_, new_n17573_, new_n17574_, new_n17575_,
    new_n17576_, new_n17577_, new_n17578_, new_n17579_, new_n17580_,
    new_n17581_, new_n17582_, new_n17583_, new_n17584_, new_n17585_,
    new_n17586_, new_n17587_, new_n17588_, new_n17589_, new_n17590_,
    new_n17591_, new_n17592_, new_n17593_, new_n17594_, new_n17595_,
    new_n17596_, new_n17597_, new_n17598_, new_n17599_, new_n17600_,
    new_n17601_, new_n17602_, new_n17603_, new_n17604_, new_n17605_,
    new_n17606_, new_n17607_, new_n17608_, new_n17609_, new_n17610_,
    new_n17611_, new_n17612_, new_n17613_, new_n17614_, new_n17615_,
    new_n17616_, new_n17617_, new_n17618_, new_n17619_, new_n17620_,
    new_n17621_, new_n17622_, new_n17623_, new_n17624_, new_n17625_,
    new_n17626_, new_n17627_, new_n17628_, new_n17629_, new_n17630_,
    new_n17631_, new_n17632_, new_n17633_, new_n17634_, new_n17635_,
    new_n17636_, new_n17637_, new_n17638_, new_n17639_, new_n17640_,
    new_n17641_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17667_, new_n17668_, new_n17669_, new_n17670_,
    new_n17671_, new_n17672_, new_n17673_, new_n17674_, new_n17675_,
    new_n17676_, new_n17677_, new_n17678_, new_n17679_, new_n17680_,
    new_n17681_, new_n17682_, new_n17683_, new_n17684_, new_n17685_,
    new_n17686_, new_n17687_, new_n17688_, new_n17689_, new_n17690_,
    new_n17691_, new_n17692_, new_n17693_, new_n17694_, new_n17695_,
    new_n17696_, new_n17697_, new_n17698_, new_n17699_, new_n17700_,
    new_n17701_, new_n17702_, new_n17703_, new_n17704_, new_n17705_,
    new_n17706_, new_n17707_, new_n17708_, new_n17709_, new_n17710_,
    new_n17711_, new_n17712_, new_n17713_, new_n17714_, new_n17715_,
    new_n17716_, new_n17717_, new_n17718_, new_n17719_, new_n17720_,
    new_n17721_, new_n17722_, new_n17723_, new_n17724_, new_n17725_,
    new_n17726_, new_n17727_, new_n17728_, new_n17729_, new_n17730_,
    new_n17731_, new_n17732_, new_n17733_, new_n17734_, new_n17735_,
    new_n17736_, new_n17737_, new_n17738_, new_n17739_, new_n17740_,
    new_n17741_, new_n17742_, new_n17743_, new_n17744_, new_n17745_,
    new_n17746_, new_n17747_, new_n17748_, new_n17749_, new_n17750_,
    new_n17751_, new_n17752_, new_n17753_, new_n17754_, new_n17755_,
    new_n17756_, new_n17757_, new_n17758_, new_n17759_, new_n17760_,
    new_n17761_, new_n17762_, new_n17763_, new_n17764_, new_n17765_,
    new_n17766_, new_n17767_, new_n17768_, new_n17769_, new_n17770_,
    new_n17771_, new_n17772_, new_n17773_, new_n17774_, new_n17775_,
    new_n17776_, new_n17777_, new_n17778_, new_n17779_, new_n17780_,
    new_n17781_, new_n17782_, new_n17783_, new_n17784_, new_n17785_,
    new_n17786_, new_n17787_, new_n17788_, new_n17789_, new_n17790_,
    new_n17791_, new_n17792_, new_n17793_, new_n17794_, new_n17795_,
    new_n17796_, new_n17797_, new_n17798_, new_n17799_, new_n17800_,
    new_n17801_, new_n17802_, new_n17803_, new_n17804_, new_n17805_,
    new_n17806_, new_n17807_, new_n17808_, new_n17809_, new_n17810_,
    new_n17811_, new_n17812_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17824_, new_n17825_,
    new_n17826_, new_n17827_, new_n17828_, new_n17829_, new_n17830_,
    new_n17831_, new_n17832_, new_n17833_, new_n17834_, new_n17835_,
    new_n17836_, new_n17837_, new_n17838_, new_n17839_, new_n17840_,
    new_n17841_, new_n17842_, new_n17843_, new_n17844_, new_n17845_,
    new_n17846_, new_n17847_, new_n17848_, new_n17849_, new_n17850_,
    new_n17851_, new_n17852_, new_n17853_, new_n17854_, new_n17855_,
    new_n17856_, new_n17857_, new_n17858_, new_n17859_, new_n17860_,
    new_n17861_, new_n17862_, new_n17863_, new_n17864_, new_n17865_,
    new_n17866_, new_n17867_, new_n17868_, new_n17869_, new_n17870_,
    new_n17871_, new_n17872_, new_n17873_, new_n17874_, new_n17875_,
    new_n17876_, new_n17877_, new_n17878_, new_n17879_, new_n17880_,
    new_n17881_, new_n17882_, new_n17883_, new_n17884_, new_n17885_,
    new_n17886_, new_n17887_, new_n17888_, new_n17889_, new_n17890_,
    new_n17891_, new_n17892_, new_n17893_, new_n17894_, new_n17895_,
    new_n17896_, new_n17897_, new_n17898_, new_n17899_, new_n17900_,
    new_n17901_, new_n17902_, new_n17903_, new_n17904_, new_n17905_,
    new_n17906_, new_n17907_, new_n17908_, new_n17909_, new_n17910_,
    new_n17911_, new_n17912_, new_n17913_, new_n17914_, new_n17915_,
    new_n17916_, new_n17917_, new_n17918_, new_n17919_, new_n17920_,
    new_n17921_, new_n17922_, new_n17923_, new_n17924_, new_n17925_,
    new_n17926_, new_n17927_, new_n17928_, new_n17929_, new_n17930_,
    new_n17931_, new_n17932_, new_n17933_, new_n17934_, new_n17935_,
    new_n17936_, new_n17937_, new_n17938_, new_n17939_, new_n17940_,
    new_n17941_, new_n17942_, new_n17943_, new_n17944_, new_n17945_,
    new_n17946_, new_n17947_, new_n17948_, new_n17949_, new_n17950_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17970_,
    new_n17971_, new_n17972_, new_n17973_, new_n17974_, new_n17975_,
    new_n17976_, new_n17977_, new_n17978_, new_n17979_, new_n17980_,
    new_n17981_, new_n17982_, new_n17983_, new_n17984_, new_n17985_,
    new_n17986_, new_n17987_, new_n17988_, new_n17989_, new_n17990_,
    new_n17991_, new_n17992_, new_n17993_, new_n17994_, new_n17995_,
    new_n17996_, new_n17997_, new_n17998_, new_n17999_, new_n18000_,
    new_n18001_, new_n18002_, new_n18003_, new_n18004_, new_n18005_,
    new_n18006_, new_n18007_, new_n18008_, new_n18009_, new_n18010_,
    new_n18011_, new_n18012_, new_n18013_, new_n18014_, new_n18015_,
    new_n18016_, new_n18017_, new_n18018_, new_n18019_, new_n18020_,
    new_n18021_, new_n18022_, new_n18023_, new_n18024_, new_n18025_,
    new_n18026_, new_n18027_, new_n18028_, new_n18029_, new_n18030_,
    new_n18031_, new_n18032_, new_n18033_, new_n18034_, new_n18035_,
    new_n18036_, new_n18037_, new_n18038_, new_n18039_, new_n18040_,
    new_n18041_, new_n18042_, new_n18043_, new_n18044_, new_n18045_,
    new_n18046_, new_n18047_, new_n18048_, new_n18049_, new_n18050_,
    new_n18051_, new_n18052_, new_n18053_, new_n18054_, new_n18055_,
    new_n18056_, new_n18057_, new_n18058_, new_n18059_, new_n18060_,
    new_n18061_, new_n18062_, new_n18063_, new_n18064_, new_n18065_,
    new_n18066_, new_n18067_, new_n18068_, new_n18069_, new_n18070_,
    new_n18071_, new_n18072_, new_n18073_, new_n18074_, new_n18075_,
    new_n18076_, new_n18077_, new_n18078_, new_n18079_, new_n18080_,
    new_n18081_, new_n18082_, new_n18083_, new_n18084_, new_n18085_,
    new_n18086_, new_n18087_, new_n18088_, new_n18089_, new_n18090_,
    new_n18091_, new_n18092_, new_n18093_, new_n18094_, new_n18095_,
    new_n18096_, new_n18097_, new_n18098_, new_n18099_, new_n18100_,
    new_n18101_, new_n18102_, new_n18103_, new_n18104_, new_n18105_,
    new_n18106_, new_n18107_, new_n18108_, new_n18109_, new_n18110_,
    new_n18111_, new_n18112_, new_n18113_, new_n18114_, new_n18115_,
    new_n18116_, new_n18117_, new_n18118_, new_n18119_, new_n18120_,
    new_n18121_, new_n18122_, new_n18123_, new_n18124_, new_n18125_,
    new_n18126_, new_n18127_, new_n18128_, new_n18129_, new_n18130_,
    new_n18131_, new_n18132_, new_n18133_, new_n18134_, new_n18135_,
    new_n18136_, new_n18137_, new_n18138_, new_n18139_, new_n18140_,
    new_n18141_, new_n18142_, new_n18143_, new_n18144_, new_n18145_,
    new_n18146_, new_n18147_, new_n18148_, new_n18149_, new_n18150_,
    new_n18151_, new_n18152_, new_n18153_, new_n18154_, new_n18155_,
    new_n18156_, new_n18157_, new_n18158_, new_n18159_, new_n18160_,
    new_n18161_, new_n18162_, new_n18163_, new_n18164_, new_n18165_,
    new_n18166_, new_n18167_, new_n18168_, new_n18169_, new_n18170_,
    new_n18171_, new_n18172_, new_n18173_, new_n18174_, new_n18175_,
    new_n18176_, new_n18177_, new_n18178_, new_n18179_, new_n18180_,
    new_n18181_, new_n18182_, new_n18183_, new_n18184_, new_n18185_,
    new_n18186_, new_n18187_, new_n18188_, new_n18189_, new_n18190_,
    new_n18191_, new_n18192_, new_n18193_, new_n18194_, new_n18195_,
    new_n18196_, new_n18197_, new_n18198_, new_n18199_, new_n18200_,
    new_n18201_, new_n18202_, new_n18203_, new_n18204_, new_n18205_,
    new_n18206_, new_n18207_, new_n18208_, new_n18209_, new_n18210_,
    new_n18211_, new_n18212_, new_n18213_, new_n18214_, new_n18215_,
    new_n18216_, new_n18217_, new_n18218_, new_n18219_, new_n18220_,
    new_n18221_, new_n18222_, new_n18223_, new_n18224_, new_n18225_,
    new_n18226_, new_n18227_, new_n18228_, new_n18229_, new_n18230_,
    new_n18231_, new_n18232_, new_n18233_, new_n18234_, new_n18235_,
    new_n18236_, new_n18237_, new_n18238_, new_n18239_, new_n18240_,
    new_n18241_, new_n18242_, new_n18243_, new_n18244_, new_n18245_,
    new_n18246_, new_n18247_, new_n18248_, new_n18249_, new_n18250_,
    new_n18251_, new_n18252_, new_n18253_, new_n18254_, new_n18255_,
    new_n18256_, new_n18257_, new_n18258_, new_n18259_, new_n18260_,
    new_n18261_, new_n18262_, new_n18263_, new_n18264_, new_n18265_,
    new_n18266_, new_n18267_, new_n18268_, new_n18269_, new_n18270_,
    new_n18271_, new_n18272_, new_n18273_, new_n18274_, new_n18275_,
    new_n18276_, new_n18277_, new_n18278_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18376_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18381_, new_n18382_, new_n18383_, new_n18384_, new_n18385_,
    new_n18386_, new_n18387_, new_n18388_, new_n18389_, new_n18390_,
    new_n18391_, new_n18392_, new_n18393_, new_n18394_, new_n18395_,
    new_n18396_, new_n18397_, new_n18398_, new_n18399_, new_n18400_,
    new_n18401_, new_n18402_, new_n18403_, new_n18404_, new_n18405_,
    new_n18406_, new_n18407_, new_n18408_, new_n18409_, new_n18410_,
    new_n18411_, new_n18412_, new_n18413_, new_n18414_, new_n18415_,
    new_n18416_, new_n18417_, new_n18418_, new_n18419_, new_n18420_,
    new_n18421_, new_n18422_, new_n18423_, new_n18424_, new_n18425_,
    new_n18426_, new_n18427_, new_n18428_, new_n18429_, new_n18430_,
    new_n18431_, new_n18432_, new_n18433_, new_n18434_, new_n18435_,
    new_n18436_, new_n18437_, new_n18438_, new_n18439_, new_n18440_,
    new_n18441_, new_n18442_, new_n18443_, new_n18444_, new_n18445_,
    new_n18446_, new_n18447_, new_n18448_, new_n18449_, new_n18450_,
    new_n18451_, new_n18452_, new_n18453_, new_n18454_, new_n18455_,
    new_n18456_, new_n18457_, new_n18458_, new_n18459_, new_n18460_,
    new_n18461_, new_n18462_, new_n18463_, new_n18464_, new_n18465_,
    new_n18466_, new_n18467_, new_n18468_, new_n18469_, new_n18470_,
    new_n18471_, new_n18472_, new_n18473_, new_n18474_, new_n18475_,
    new_n18476_, new_n18477_, new_n18478_, new_n18479_, new_n18480_,
    new_n18481_, new_n18482_, new_n18483_, new_n18484_, new_n18485_,
    new_n18486_, new_n18487_, new_n18488_, new_n18489_, new_n18490_,
    new_n18491_, new_n18492_, new_n18493_, new_n18494_, new_n18495_,
    new_n18496_, new_n18497_, new_n18498_, new_n18499_, new_n18500_,
    new_n18501_, new_n18502_, new_n18503_, new_n18504_, new_n18505_,
    new_n18506_, new_n18507_, new_n18508_, new_n18509_, new_n18510_,
    new_n18511_, new_n18512_, new_n18513_, new_n18514_, new_n18515_,
    new_n18516_, new_n18517_, new_n18518_, new_n18519_, new_n18520_,
    new_n18521_, new_n18522_, new_n18523_, new_n18524_, new_n18525_,
    new_n18526_, new_n18527_, new_n18528_, new_n18529_, new_n18530_,
    new_n18531_, new_n18532_, new_n18533_, new_n18534_, new_n18535_,
    new_n18536_, new_n18537_, new_n18538_, new_n18539_, new_n18540_,
    new_n18541_, new_n18542_, new_n18543_, new_n18544_, new_n18545_,
    new_n18546_, new_n18547_, new_n18548_, new_n18549_, new_n18550_,
    new_n18551_, new_n18552_, new_n18553_, new_n18554_, new_n18555_,
    new_n18556_, new_n18557_, new_n18558_, new_n18559_, new_n18560_,
    new_n18561_, new_n18562_, new_n18563_, new_n18564_, new_n18565_,
    new_n18566_, new_n18567_, new_n18568_, new_n18569_, new_n18570_,
    new_n18571_, new_n18572_, new_n18573_, new_n18574_, new_n18575_,
    new_n18576_, new_n18577_, new_n18578_, new_n18579_, new_n18580_,
    new_n18581_, new_n18582_, new_n18583_, new_n18584_, new_n18585_,
    new_n18586_, new_n18587_, new_n18588_, new_n18589_, new_n18590_,
    new_n18591_, new_n18592_, new_n18593_, new_n18594_, new_n18595_,
    new_n18596_, new_n18597_, new_n18598_, new_n18599_, new_n18600_,
    new_n18601_, new_n18602_, new_n18603_, new_n18604_, new_n18605_,
    new_n18606_, new_n18607_, new_n18608_, new_n18609_, new_n18610_,
    new_n18611_, new_n18612_, new_n18613_, new_n18614_, new_n18615_,
    new_n18616_, new_n18617_, new_n18618_, new_n18619_, new_n18620_,
    new_n18621_, new_n18622_, new_n18623_, new_n18624_, new_n18625_,
    new_n18626_, new_n18627_, new_n18628_, new_n18629_, new_n18630_,
    new_n18631_, new_n18632_, new_n18633_, new_n18634_, new_n18635_,
    new_n18636_, new_n18637_, new_n18638_, new_n18639_, new_n18640_,
    new_n18641_, new_n18642_, new_n18643_, new_n18644_, new_n18645_,
    new_n18646_, new_n18647_, new_n18648_, new_n18649_, new_n18650_,
    new_n18651_, new_n18652_, new_n18653_, new_n18654_, new_n18655_,
    new_n18656_, new_n18657_, new_n18658_, new_n18659_, new_n18660_,
    new_n18661_, new_n18662_, new_n18663_, new_n18664_, new_n18665_,
    new_n18666_, new_n18667_, new_n18668_, new_n18669_, new_n18670_,
    new_n18671_, new_n18672_, new_n18673_, new_n18674_, new_n18675_,
    new_n18676_, new_n18677_, new_n18678_, new_n18679_, new_n18680_,
    new_n18681_, new_n18682_, new_n18683_, new_n18684_, new_n18685_,
    new_n18686_, new_n18687_, new_n18688_, new_n18689_, new_n18690_,
    new_n18691_, new_n18692_, new_n18693_, new_n18694_, new_n18695_,
    new_n18696_, new_n18697_, new_n18698_, new_n18699_, new_n18700_,
    new_n18701_, new_n18702_, new_n18703_, new_n18704_, new_n18705_,
    new_n18706_, new_n18707_, new_n18708_, new_n18709_, new_n18710_,
    new_n18711_, new_n18712_, new_n18713_, new_n18714_, new_n18715_,
    new_n18716_, new_n18717_, new_n18718_, new_n18719_, new_n18720_,
    new_n18721_, new_n18722_, new_n18723_, new_n18724_, new_n18725_,
    new_n18726_, new_n18727_, new_n18728_, new_n18729_, new_n18730_,
    new_n18731_, new_n18732_, new_n18733_, new_n18734_, new_n18735_,
    new_n18736_, new_n18737_, new_n18738_, new_n18739_, new_n18740_,
    new_n18741_, new_n18742_, new_n18743_, new_n18744_, new_n18745_,
    new_n18746_, new_n18747_, new_n18748_, new_n18749_, new_n18750_,
    new_n18751_, new_n18752_, new_n18753_, new_n18754_, new_n18755_,
    new_n18756_, new_n18757_, new_n18758_, new_n18759_, new_n18760_,
    new_n18761_, new_n18762_, new_n18763_, new_n18764_, new_n18765_,
    new_n18766_, new_n18767_, new_n18768_, new_n18769_, new_n18770_,
    new_n18771_, new_n18772_, new_n18773_, new_n18774_, new_n18775_,
    new_n18776_, new_n18777_, new_n18778_, new_n18779_, new_n18780_,
    new_n18781_, new_n18782_, new_n18783_, new_n18784_, new_n18785_,
    new_n18786_, new_n18787_, new_n18788_, new_n18789_, new_n18790_,
    new_n18791_, new_n18792_, new_n18793_, new_n18794_, new_n18795_,
    new_n18796_, new_n18797_, new_n18798_, new_n18799_, new_n18800_,
    new_n18801_, new_n18802_, new_n18803_, new_n18804_, new_n18805_,
    new_n18806_, new_n18807_, new_n18808_, new_n18809_, new_n18810_,
    new_n18811_, new_n18812_, new_n18813_, new_n18814_, new_n18815_,
    new_n18816_, new_n18817_, new_n18818_, new_n18819_, new_n18820_,
    new_n18821_, new_n18822_, new_n18823_, new_n18824_, new_n18825_,
    new_n18826_, new_n18827_, new_n18828_, new_n18829_, new_n18830_,
    new_n18831_, new_n18832_, new_n18833_, new_n18834_, new_n18835_,
    new_n18836_, new_n18837_, new_n18838_, new_n18839_, new_n18840_,
    new_n18841_, new_n18842_, new_n18843_, new_n18844_, new_n18845_,
    new_n18846_, new_n18847_, new_n18848_, new_n18849_, new_n18850_,
    new_n18851_, new_n18852_, new_n18853_, new_n18854_, new_n18855_,
    new_n18856_, new_n18857_, new_n18858_, new_n18859_, new_n18860_,
    new_n18861_, new_n18862_, new_n18863_, new_n18864_, new_n18865_,
    new_n18866_, new_n18867_, new_n18868_, new_n18869_, new_n18870_,
    new_n18871_, new_n18872_, new_n18873_, new_n18874_, new_n18875_,
    new_n18876_, new_n18877_, new_n18878_, new_n18879_, new_n18880_,
    new_n18881_, new_n18882_, new_n18883_, new_n18884_, new_n18885_,
    new_n18886_, new_n18887_, new_n18888_, new_n18889_, new_n18890_,
    new_n18891_, new_n18892_, new_n18893_, new_n18894_, new_n18895_,
    new_n18896_, new_n18897_, new_n18898_, new_n18899_, new_n18900_,
    new_n18901_, new_n18902_, new_n18903_, new_n18904_, new_n18905_,
    new_n18906_, new_n18907_, new_n18908_, new_n18909_, new_n18910_,
    new_n18911_, new_n18912_, new_n18913_, new_n18914_, new_n18915_,
    new_n18916_, new_n18917_, new_n18918_, new_n18919_, new_n18920_,
    new_n18921_, new_n18922_, new_n18923_, new_n18924_, new_n18925_,
    new_n18926_, new_n18927_, new_n18928_, new_n18929_, new_n18930_,
    new_n18931_, new_n18932_, new_n18933_, new_n18934_, new_n18935_,
    new_n18936_, new_n18937_, new_n18938_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18944_, new_n18945_,
    new_n18946_, new_n18947_, new_n18948_, new_n18949_, new_n18950_,
    new_n18951_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18992_, new_n18993_, new_n18994_, new_n18995_,
    new_n18996_, new_n18997_, new_n18998_, new_n18999_, new_n19000_,
    new_n19001_, new_n19002_, new_n19003_, new_n19004_, new_n19005_,
    new_n19006_, new_n19007_, new_n19008_, new_n19009_, new_n19010_,
    new_n19011_, new_n19012_, new_n19013_, new_n19014_, new_n19015_,
    new_n19016_, new_n19017_, new_n19018_, new_n19019_, new_n19020_,
    new_n19021_, new_n19022_, new_n19023_, new_n19024_, new_n19025_,
    new_n19026_, new_n19027_, new_n19028_, new_n19029_, new_n19030_,
    new_n19031_, new_n19032_, new_n19033_, new_n19034_, new_n19035_,
    new_n19036_, new_n19037_, new_n19038_, new_n19039_, new_n19040_,
    new_n19041_, new_n19042_, new_n19043_, new_n19044_, new_n19045_,
    new_n19046_, new_n19047_, new_n19048_, new_n19049_, new_n19050_,
    new_n19051_, new_n19052_, new_n19053_, new_n19054_, new_n19055_,
    new_n19056_, new_n19057_, new_n19058_, new_n19059_, new_n19060_,
    new_n19061_, new_n19062_, new_n19063_, new_n19064_, new_n19065_,
    new_n19066_, new_n19067_, new_n19068_, new_n19069_, new_n19070_,
    new_n19071_, new_n19072_, new_n19073_, new_n19074_, new_n19075_,
    new_n19076_, new_n19077_, new_n19078_, new_n19079_, new_n19080_,
    new_n19081_, new_n19082_, new_n19083_, new_n19084_, new_n19085_,
    new_n19086_, new_n19087_, new_n19088_, new_n19089_, new_n19090_,
    new_n19091_, new_n19092_, new_n19093_, new_n19094_, new_n19095_,
    new_n19096_, new_n19097_, new_n19098_, new_n19099_, new_n19100_,
    new_n19101_, new_n19102_, new_n19103_, new_n19104_, new_n19105_,
    new_n19106_, new_n19107_, new_n19108_, new_n19109_, new_n19110_,
    new_n19111_, new_n19112_, new_n19113_, new_n19114_, new_n19115_,
    new_n19116_, new_n19117_, new_n19118_, new_n19119_, new_n19120_,
    new_n19121_, new_n19122_, new_n19123_, new_n19124_, new_n19125_,
    new_n19126_, new_n19127_, new_n19128_, new_n19129_, new_n19130_,
    new_n19131_, new_n19132_, new_n19133_, new_n19134_, new_n19135_,
    new_n19136_, new_n19137_, new_n19138_, new_n19139_, new_n19140_,
    new_n19141_, new_n19142_, new_n19143_, new_n19144_, new_n19145_,
    new_n19146_, new_n19147_, new_n19148_, new_n19149_, new_n19150_,
    new_n19151_, new_n19152_, new_n19153_, new_n19154_, new_n19155_,
    new_n19156_, new_n19157_, new_n19158_, new_n19159_, new_n19160_,
    new_n19161_, new_n19162_, new_n19163_, new_n19164_, new_n19165_,
    new_n19166_, new_n19167_, new_n19168_, new_n19169_, new_n19170_,
    new_n19171_, new_n19172_, new_n19173_, new_n19174_, new_n19175_,
    new_n19176_, new_n19177_, new_n19178_, new_n19179_, new_n19180_,
    new_n19181_, new_n19182_, new_n19183_, new_n19184_, new_n19185_,
    new_n19186_, new_n19187_, new_n19188_, new_n19189_, new_n19190_,
    new_n19191_, new_n19192_, new_n19193_, new_n19194_, new_n19195_,
    new_n19196_, new_n19197_, new_n19198_, new_n19199_, new_n19200_,
    new_n19201_, new_n19202_, new_n19203_, new_n19204_, new_n19205_,
    new_n19206_, new_n19207_, new_n19208_, new_n19209_, new_n19210_,
    new_n19211_, new_n19212_, new_n19213_, new_n19214_, new_n19215_,
    new_n19216_, new_n19217_, new_n19218_, new_n19219_, new_n19220_,
    new_n19221_, new_n19222_, new_n19223_, new_n19224_, new_n19225_,
    new_n19226_, new_n19227_, new_n19228_, new_n19229_, new_n19230_,
    new_n19231_, new_n19232_, new_n19233_, new_n19234_, new_n19235_,
    new_n19236_, new_n19237_, new_n19238_, new_n19239_, new_n19240_,
    new_n19241_, new_n19242_, new_n19243_, new_n19244_, new_n19245_,
    new_n19246_, new_n19247_, new_n19248_, new_n19249_, new_n19250_,
    new_n19251_, new_n19252_, new_n19253_, new_n19254_, new_n19255_,
    new_n19256_, new_n19257_, new_n19258_, new_n19259_, new_n19260_,
    new_n19261_, new_n19262_, new_n19263_, new_n19264_, new_n19265_,
    new_n19266_, new_n19267_, new_n19268_, new_n19269_, new_n19270_,
    new_n19271_, new_n19272_, new_n19273_, new_n19274_, new_n19275_,
    new_n19276_, new_n19277_, new_n19278_, new_n19279_, new_n19280_,
    new_n19281_, new_n19282_, new_n19283_, new_n19284_, new_n19285_,
    new_n19286_, new_n19287_, new_n19288_, new_n19289_, new_n19290_,
    new_n19291_, new_n19292_, new_n19293_, new_n19294_, new_n19295_,
    new_n19296_, new_n19297_, new_n19298_, new_n19299_, new_n19300_,
    new_n19301_, new_n19302_, new_n19303_, new_n19304_, new_n19305_,
    new_n19306_, new_n19307_, new_n19308_, new_n19309_, new_n19310_,
    new_n19311_, new_n19312_, new_n19313_, new_n19314_, new_n19315_,
    new_n19316_, new_n19317_, new_n19318_, new_n19319_, new_n19320_,
    new_n19321_, new_n19322_, new_n19323_, new_n19324_, new_n19325_,
    new_n19326_, new_n19327_, new_n19328_, new_n19329_, new_n19330_,
    new_n19331_, new_n19332_, new_n19333_, new_n19334_, new_n19335_,
    new_n19336_, new_n19337_, new_n19338_, new_n19339_, new_n19340_,
    new_n19341_, new_n19342_, new_n19343_, new_n19344_, new_n19345_,
    new_n19346_, new_n19347_, new_n19348_, new_n19349_, new_n19350_,
    new_n19351_, new_n19352_, new_n19353_, new_n19354_, new_n19355_,
    new_n19356_, new_n19357_, new_n19358_, new_n19359_, new_n19360_,
    new_n19361_, new_n19362_, new_n19363_, new_n19364_, new_n19365_,
    new_n19366_, new_n19367_, new_n19368_, new_n19369_, new_n19370_,
    new_n19371_, new_n19372_, new_n19373_, new_n19374_, new_n19375_,
    new_n19376_, new_n19377_, new_n19378_, new_n19379_, new_n19380_,
    new_n19381_, new_n19382_, new_n19383_, new_n19384_, new_n19385_,
    new_n19386_, new_n19387_, new_n19388_, new_n19389_, new_n19390_,
    new_n19391_, new_n19392_, new_n19393_, new_n19394_, new_n19395_,
    new_n19396_, new_n19397_, new_n19398_, new_n19399_, new_n19400_,
    new_n19401_, new_n19402_, new_n19403_, new_n19404_, new_n19405_,
    new_n19406_, new_n19407_, new_n19408_, new_n19409_, new_n19410_,
    new_n19411_, new_n19412_, new_n19413_, new_n19414_, new_n19415_,
    new_n19416_, new_n19417_, new_n19418_, new_n19419_, new_n19420_,
    new_n19421_, new_n19422_, new_n19423_, new_n19424_, new_n19425_,
    new_n19426_, new_n19427_, new_n19428_, new_n19429_, new_n19430_,
    new_n19431_, new_n19432_, new_n19433_, new_n19434_, new_n19435_,
    new_n19436_, new_n19437_, new_n19438_, new_n19439_, new_n19440_,
    new_n19441_, new_n19442_, new_n19443_, new_n19444_, new_n19445_,
    new_n19446_, new_n19447_, new_n19448_, new_n19449_, new_n19450_,
    new_n19451_, new_n19452_, new_n19453_, new_n19454_, new_n19455_,
    new_n19456_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19513_, new_n19514_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19738_, new_n19739_, new_n19740_,
    new_n19741_, new_n19742_, new_n19743_, new_n19744_, new_n19745_,
    new_n19746_, new_n19747_, new_n19748_, new_n19749_, new_n19750_,
    new_n19751_, new_n19752_, new_n19753_, new_n19754_, new_n19755_,
    new_n19756_, new_n19757_, new_n19758_, new_n19759_, new_n19760_,
    new_n19761_, new_n19762_, new_n19763_, new_n19764_, new_n19765_,
    new_n19766_, new_n19767_, new_n19768_, new_n19769_, new_n19770_,
    new_n19771_, new_n19772_, new_n19773_, new_n19774_, new_n19775_,
    new_n19776_, new_n19777_, new_n19778_, new_n19779_, new_n19780_,
    new_n19781_, new_n19782_, new_n19783_, new_n19784_, new_n19785_,
    new_n19786_, new_n19787_, new_n19788_, new_n19789_, new_n19790_,
    new_n19791_, new_n19792_, new_n19793_, new_n19794_, new_n19795_,
    new_n19796_, new_n19797_, new_n19798_, new_n19799_, new_n19800_,
    new_n19801_, new_n19802_, new_n19803_, new_n19804_, new_n19805_,
    new_n19806_, new_n19807_, new_n19808_, new_n19809_, new_n19810_,
    new_n19811_, new_n19812_, new_n19813_, new_n19814_, new_n19815_,
    new_n19816_, new_n19817_, new_n19818_, new_n19819_, new_n19820_,
    new_n19821_, new_n19822_, new_n19823_, new_n19824_, new_n19825_,
    new_n19826_, new_n19827_, new_n19828_, new_n19829_, new_n19830_,
    new_n19831_, new_n19832_, new_n19833_, new_n19834_, new_n19835_,
    new_n19836_, new_n19837_, new_n19838_, new_n19839_, new_n19840_,
    new_n19841_, new_n19842_, new_n19843_, new_n19844_, new_n19845_,
    new_n19846_, new_n19847_, new_n19848_, new_n19849_, new_n19850_,
    new_n19851_, new_n19852_, new_n19853_, new_n19854_, new_n19855_,
    new_n19856_, new_n19857_, new_n19858_, new_n19859_, new_n19860_,
    new_n19861_, new_n19862_, new_n19863_, new_n19864_, new_n19865_,
    new_n19866_, new_n19867_, new_n19868_, new_n19869_, new_n19870_,
    new_n19871_, new_n19872_, new_n19873_, new_n19874_, new_n19875_,
    new_n19876_, new_n19877_, new_n19878_, new_n19879_, new_n19880_,
    new_n19881_, new_n19882_, new_n19883_, new_n19884_, new_n19885_,
    new_n19886_, new_n19887_, new_n19888_, new_n19889_, new_n19890_,
    new_n19891_, new_n19892_, new_n19893_, new_n19894_, new_n19895_,
    new_n19896_, new_n19897_, new_n19898_, new_n19899_, new_n19900_,
    new_n19901_, new_n19902_, new_n19903_, new_n19904_, new_n19905_,
    new_n19906_, new_n19907_, new_n19908_, new_n19909_, new_n19910_,
    new_n19911_, new_n19912_, new_n19913_, new_n19914_, new_n19915_,
    new_n19916_, new_n19917_, new_n19918_, new_n19919_, new_n19920_,
    new_n19921_, new_n19922_, new_n19923_, new_n19924_, new_n19925_,
    new_n19926_, new_n19927_, new_n19928_, new_n19929_, new_n19930_,
    new_n19931_, new_n19932_, new_n19933_, new_n19934_, new_n19935_,
    new_n19936_, new_n19937_, new_n19938_, new_n19939_, new_n19940_,
    new_n19941_, new_n19942_, new_n19943_, new_n19944_, new_n19945_,
    new_n19946_, new_n19947_, new_n19948_, new_n19949_, new_n19950_,
    new_n19951_, new_n19952_, new_n19953_, new_n19954_, new_n19955_,
    new_n19956_, new_n19957_, new_n19958_, new_n19959_, new_n19960_,
    new_n19961_, new_n19962_, new_n19963_, new_n19964_, new_n19965_,
    new_n19966_, new_n19967_, new_n19968_, new_n19969_, new_n19970_,
    new_n19971_, new_n19972_, new_n19973_, new_n19974_, new_n19975_,
    new_n19976_, new_n19977_, new_n19978_, new_n19979_, new_n19980_,
    new_n19981_, new_n19982_, new_n19983_, new_n19984_, new_n19985_,
    new_n19986_, new_n19987_, new_n19988_, new_n19989_, new_n19990_,
    new_n19991_, new_n19992_, new_n19993_, new_n19994_, new_n19995_,
    new_n19996_, new_n19997_, new_n19998_, new_n19999_, new_n20000_,
    new_n20001_, new_n20002_, new_n20003_, new_n20004_, new_n20005_,
    new_n20006_, new_n20007_, new_n20008_, new_n20009_, new_n20010_,
    new_n20011_, new_n20012_, new_n20013_, new_n20014_, new_n20015_,
    new_n20016_, new_n20017_, new_n20018_, new_n20019_, new_n20020_,
    new_n20021_, new_n20022_, new_n20023_, new_n20024_, new_n20025_,
    new_n20026_, new_n20027_, new_n20028_, new_n20029_, new_n20030_,
    new_n20031_, new_n20032_, new_n20033_, new_n20034_, new_n20035_,
    new_n20036_, new_n20037_, new_n20038_, new_n20039_, new_n20040_,
    new_n20041_, new_n20042_, new_n20043_, new_n20044_, new_n20045_,
    new_n20046_, new_n20047_, new_n20048_, new_n20049_, new_n20050_,
    new_n20051_, new_n20052_, new_n20053_, new_n20054_, new_n20055_,
    new_n20056_, new_n20057_, new_n20058_, new_n20059_, new_n20060_,
    new_n20061_, new_n20062_, new_n20063_, new_n20064_, new_n20065_,
    new_n20066_, new_n20067_, new_n20068_, new_n20069_, new_n20070_,
    new_n20071_, new_n20072_, new_n20073_, new_n20074_, new_n20075_,
    new_n20076_, new_n20077_, new_n20078_, new_n20079_, new_n20080_,
    new_n20081_, new_n20082_, new_n20083_, new_n20084_, new_n20085_,
    new_n20086_, new_n20087_, new_n20088_, new_n20089_, new_n20090_,
    new_n20091_, new_n20092_, new_n20093_, new_n20094_, new_n20095_,
    new_n20096_, new_n20097_, new_n20098_, new_n20099_, new_n20100_,
    new_n20101_, new_n20102_, new_n20103_, new_n20104_, new_n20105_,
    new_n20106_, new_n20107_, new_n20108_, new_n20109_, new_n20110_,
    new_n20111_, new_n20112_, new_n20113_, new_n20114_, new_n20115_,
    new_n20116_, new_n20117_, new_n20118_, new_n20119_, new_n20120_,
    new_n20121_, new_n20122_, new_n20123_, new_n20124_, new_n20125_,
    new_n20126_, new_n20127_, new_n20128_, new_n20129_, new_n20130_,
    new_n20131_, new_n20132_, new_n20133_, new_n20134_, new_n20135_,
    new_n20136_, new_n20137_, new_n20138_, new_n20139_, new_n20140_,
    new_n20141_, new_n20142_, new_n20143_, new_n20144_, new_n20145_,
    new_n20146_, new_n20147_, new_n20148_, new_n20149_, new_n20150_,
    new_n20151_, new_n20152_, new_n20153_, new_n20154_, new_n20155_,
    new_n20156_, new_n20157_, new_n20158_, new_n20159_, new_n20160_,
    new_n20161_, new_n20162_, new_n20163_, new_n20164_, new_n20165_,
    new_n20166_, new_n20167_, new_n20168_, new_n20169_, new_n20170_,
    new_n20171_, new_n20172_, new_n20173_, new_n20174_, new_n20175_,
    new_n20176_, new_n20177_, new_n20178_, new_n20179_, new_n20180_,
    new_n20181_, new_n20182_, new_n20183_, new_n20184_, new_n20185_,
    new_n20186_, new_n20187_, new_n20188_, new_n20189_, new_n20190_,
    new_n20191_, new_n20192_, new_n20193_, new_n20194_, new_n20195_,
    new_n20196_, new_n20197_, new_n20198_, new_n20199_, new_n20200_,
    new_n20201_, new_n20202_, new_n20203_, new_n20204_, new_n20205_,
    new_n20206_, new_n20207_, new_n20208_, new_n20209_, new_n20210_,
    new_n20211_, new_n20212_, new_n20213_, new_n20214_, new_n20215_,
    new_n20216_, new_n20217_, new_n20218_, new_n20219_, new_n20220_,
    new_n20221_, new_n20222_, new_n20223_, new_n20224_, new_n20225_,
    new_n20226_, new_n20227_, new_n20228_, new_n20229_, new_n20230_,
    new_n20231_, new_n20232_, new_n20233_, new_n20234_, new_n20235_,
    new_n20236_, new_n20237_, new_n20238_, new_n20239_, new_n20240_,
    new_n20241_, new_n20242_, new_n20243_, new_n20244_, new_n20245_,
    new_n20246_, new_n20247_, new_n20248_, new_n20249_, new_n20250_,
    new_n20251_, new_n20252_, new_n20253_, new_n20254_, new_n20255_,
    new_n20256_, new_n20257_, new_n20258_, new_n20259_, new_n20260_,
    new_n20261_, new_n20262_, new_n20263_, new_n20264_, new_n20265_,
    new_n20266_, new_n20267_, new_n20268_, new_n20269_, new_n20270_,
    new_n20271_, new_n20272_, new_n20273_, new_n20274_, new_n20275_,
    new_n20276_, new_n20277_, new_n20278_, new_n20279_, new_n20280_,
    new_n20281_, new_n20282_, new_n20283_, new_n20284_, new_n20285_,
    new_n20286_, new_n20287_, new_n20288_, new_n20289_, new_n20290_,
    new_n20291_, new_n20292_, new_n20293_, new_n20294_, new_n20295_,
    new_n20296_, new_n20297_, new_n20298_, new_n20299_, new_n20300_,
    new_n20301_, new_n20302_, new_n20303_, new_n20304_, new_n20305_,
    new_n20306_, new_n20307_, new_n20308_, new_n20309_, new_n20310_,
    new_n20311_, new_n20312_, new_n20313_, new_n20314_, new_n20315_,
    new_n20316_, new_n20317_, new_n20318_, new_n20319_, new_n20320_,
    new_n20321_, new_n20322_, new_n20323_, new_n20324_, new_n20325_,
    new_n20326_, new_n20327_, new_n20328_, new_n20329_, new_n20330_,
    new_n20331_, new_n20332_, new_n20333_, new_n20334_, new_n20335_,
    new_n20336_, new_n20337_, new_n20338_, new_n20339_, new_n20340_,
    new_n20341_, new_n20342_, new_n20343_, new_n20344_, new_n20345_,
    new_n20346_, new_n20347_, new_n20348_, new_n20349_, new_n20350_,
    new_n20351_, new_n20352_, new_n20353_, new_n20354_, new_n20355_,
    new_n20356_, new_n20357_, new_n20358_, new_n20359_, new_n20360_,
    new_n20361_, new_n20362_, new_n20363_, new_n20364_, new_n20365_,
    new_n20366_, new_n20367_, new_n20368_, new_n20369_, new_n20370_,
    new_n20371_, new_n20372_, new_n20373_, new_n20374_, new_n20375_,
    new_n20376_, new_n20377_, new_n20378_, new_n20379_, new_n20380_,
    new_n20381_, new_n20382_, new_n20383_, new_n20384_, new_n20385_,
    new_n20386_, new_n20387_, new_n20388_, new_n20389_, new_n20390_,
    new_n20391_, new_n20392_, new_n20393_, new_n20394_, new_n20395_,
    new_n20396_, new_n20397_, new_n20398_, new_n20399_, new_n20400_,
    new_n20401_, new_n20402_, new_n20403_, new_n20404_, new_n20405_,
    new_n20406_, new_n20407_, new_n20408_, new_n20409_, new_n20410_,
    new_n20411_, new_n20412_, new_n20413_, new_n20414_, new_n20415_,
    new_n20416_, new_n20417_, new_n20418_, new_n20419_, new_n20420_,
    new_n20421_, new_n20422_, new_n20423_, new_n20424_, new_n20425_,
    new_n20426_, new_n20427_, new_n20428_, new_n20429_, new_n20430_,
    new_n20431_, new_n20432_, new_n20433_, new_n20434_, new_n20435_,
    new_n20436_, new_n20437_, new_n20438_, new_n20439_, new_n20440_,
    new_n20441_, new_n20442_, new_n20443_, new_n20444_, new_n20445_,
    new_n20446_, new_n20447_, new_n20448_, new_n20449_, new_n20450_,
    new_n20451_, new_n20452_, new_n20453_, new_n20454_, new_n20455_,
    new_n20456_, new_n20457_, new_n20458_, new_n20459_, new_n20460_,
    new_n20461_, new_n20462_, new_n20463_, new_n20464_, new_n20465_,
    new_n20466_, new_n20467_, new_n20468_, new_n20469_, new_n20470_,
    new_n20471_, new_n20472_, new_n20473_, new_n20474_, new_n20475_,
    new_n20476_, new_n20477_, new_n20478_, new_n20479_, new_n20480_,
    new_n20481_, new_n20482_, new_n20483_, new_n20484_, new_n20485_,
    new_n20486_, new_n20487_, new_n20488_, new_n20489_, new_n20490_,
    new_n20491_, new_n20492_, new_n20493_, new_n20494_, new_n20495_,
    new_n20496_, new_n20497_, new_n20498_, new_n20499_, new_n20500_,
    new_n20501_, new_n20502_, new_n20503_, new_n20504_, new_n20505_,
    new_n20506_, new_n20507_, new_n20508_, new_n20509_, new_n20510_,
    new_n20511_, new_n20512_, new_n20513_, new_n20514_, new_n20515_,
    new_n20516_, new_n20517_, new_n20518_, new_n20519_, new_n20520_,
    new_n20521_, new_n20522_, new_n20523_, new_n20524_, new_n20525_,
    new_n20526_, new_n20527_, new_n20528_, new_n20529_, new_n20530_,
    new_n20531_, new_n20532_, new_n20533_, new_n20534_, new_n20535_,
    new_n20536_, new_n20537_, new_n20538_, new_n20539_, new_n20540_,
    new_n20541_, new_n20542_, new_n20543_, new_n20544_, new_n20545_,
    new_n20546_, new_n20547_, new_n20548_, new_n20549_, new_n20550_,
    new_n20551_, new_n20552_, new_n20553_, new_n20554_, new_n20555_,
    new_n20556_, new_n20557_, new_n20558_, new_n20559_, new_n20560_,
    new_n20561_, new_n20562_, new_n20563_, new_n20564_, new_n20565_,
    new_n20566_, new_n20567_, new_n20568_, new_n20569_, new_n20570_,
    new_n20571_, new_n20572_, new_n20573_, new_n20574_, new_n20575_,
    new_n20576_, new_n20577_, new_n20578_, new_n20579_, new_n20580_,
    new_n20581_, new_n20582_, new_n20583_, new_n20584_, new_n20585_,
    new_n20586_, new_n20587_, new_n20588_, new_n20589_, new_n20590_,
    new_n20591_, new_n20592_, new_n20593_, new_n20594_, new_n20595_,
    new_n20596_, new_n20597_, new_n20598_, new_n20599_, new_n20600_,
    new_n20601_, new_n20602_, new_n20603_, new_n20604_, new_n20605_,
    new_n20606_, new_n20607_, new_n20608_, new_n20609_, new_n20610_,
    new_n20611_, new_n20612_, new_n20613_, new_n20614_, new_n20615_,
    new_n20616_, new_n20617_, new_n20618_, new_n20619_, new_n20620_,
    new_n20621_, new_n20622_, new_n20623_, new_n20624_, new_n20625_,
    new_n20626_, new_n20627_, new_n20628_, new_n20629_, new_n20630_,
    new_n20631_, new_n20632_, new_n20633_, new_n20634_, new_n20635_,
    new_n20636_, new_n20637_, new_n20638_, new_n20639_, new_n20640_,
    new_n20641_, new_n20642_, new_n20643_, new_n20644_, new_n20645_,
    new_n20646_, new_n20647_, new_n20648_, new_n20649_, new_n20650_,
    new_n20651_, new_n20652_, new_n20653_, new_n20654_, new_n20655_,
    new_n20656_, new_n20657_, new_n20658_, new_n20659_, new_n20660_,
    new_n20661_, new_n20662_, new_n20663_, new_n20664_, new_n20665_,
    new_n20666_, new_n20667_, new_n20668_, new_n20669_, new_n20670_,
    new_n20671_, new_n20672_, new_n20673_, new_n20674_, new_n20675_,
    new_n20676_, new_n20677_, new_n20678_, new_n20679_, new_n20680_,
    new_n20681_, new_n20682_, new_n20683_, new_n20684_, new_n20685_,
    new_n20686_, new_n20687_, new_n20688_, new_n20689_, new_n20690_,
    new_n20691_, new_n20692_, new_n20693_, new_n20694_, new_n20695_,
    new_n20696_, new_n20697_, new_n20698_, new_n20699_, new_n20700_,
    new_n20701_, new_n20702_, new_n20703_, new_n20704_, new_n20705_,
    new_n20706_, new_n20707_, new_n20708_, new_n20709_, new_n20710_,
    new_n20711_, new_n20712_, new_n20713_, new_n20714_, new_n20715_,
    new_n20716_, new_n20717_, new_n20718_, new_n20719_, new_n20720_,
    new_n20721_, new_n20722_, new_n20723_, new_n20724_, new_n20725_,
    new_n20726_, new_n20727_, new_n20728_, new_n20729_, new_n20730_,
    new_n20731_, new_n20732_, new_n20733_, new_n20734_, new_n20735_,
    new_n20736_, new_n20737_, new_n20738_, new_n20739_, new_n20740_,
    new_n20741_, new_n20742_, new_n20743_, new_n20744_, new_n20745_,
    new_n20746_, new_n20747_, new_n20748_, new_n20749_, new_n20750_,
    new_n20751_, new_n20752_, new_n20753_, new_n20754_, new_n20755_,
    new_n20756_, new_n20757_, new_n20758_, new_n20759_, new_n20760_,
    new_n20761_, new_n20762_, new_n20763_, new_n20764_, new_n20765_,
    new_n20766_, new_n20767_, new_n20768_, new_n20769_, new_n20770_,
    new_n20771_, new_n20772_, new_n20773_, new_n20774_, new_n20775_,
    new_n20776_, new_n20777_, new_n20778_, new_n20779_, new_n20780_,
    new_n20781_, new_n20782_, new_n20783_, new_n20784_, new_n20785_,
    new_n20786_, new_n20787_, new_n20788_, new_n20789_, new_n20790_,
    new_n20791_, new_n20792_, new_n20793_, new_n20794_, new_n20795_,
    new_n20796_, new_n20797_, new_n20798_, new_n20799_, new_n20800_,
    new_n20801_, new_n20802_, new_n20803_, new_n20804_, new_n20805_,
    new_n20806_, new_n20807_, new_n20808_, new_n20809_, new_n20810_,
    new_n20811_, new_n20812_, new_n20813_, new_n20814_, new_n20815_,
    new_n20816_, new_n20817_, new_n20818_, new_n20819_, new_n20820_,
    new_n20821_, new_n20822_, new_n20823_, new_n20824_, new_n20825_,
    new_n20826_, new_n20827_, new_n20828_, new_n20829_, new_n20830_,
    new_n20831_, new_n20832_, new_n20833_, new_n20834_, new_n20835_,
    new_n20836_, new_n20837_, new_n20838_, new_n20839_, new_n20840_,
    new_n20841_, new_n20842_, new_n20843_, new_n20844_, new_n20845_,
    new_n20846_, new_n20847_, new_n20848_, new_n20849_, new_n20850_,
    new_n20851_, new_n20852_, new_n20853_, new_n20854_, new_n20855_,
    new_n20856_, new_n20857_, new_n20858_, new_n20859_, new_n20860_,
    new_n20861_, new_n20862_, new_n20863_, new_n20864_, new_n20865_,
    new_n20866_, new_n20867_, new_n20868_, new_n20869_, new_n20870_,
    new_n20871_, new_n20872_, new_n20873_, new_n20874_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20888_, new_n20889_, new_n20890_,
    new_n20891_, new_n20892_, new_n20893_, new_n20894_, new_n20895_,
    new_n20896_, new_n20897_, new_n20898_, new_n20899_, new_n20900_,
    new_n20901_, new_n20902_, new_n20903_, new_n20904_, new_n20905_,
    new_n20906_, new_n20907_, new_n20908_, new_n20909_, new_n20910_,
    new_n20911_, new_n20912_, new_n20913_, new_n20914_, new_n20915_,
    new_n20916_, new_n20917_, new_n20918_, new_n20919_, new_n20920_,
    new_n20921_, new_n20922_, new_n20923_, new_n20924_, new_n20925_,
    new_n20926_, new_n20927_, new_n20928_, new_n20929_, new_n20930_,
    new_n20931_, new_n20932_, new_n20933_, new_n20934_, new_n20935_,
    new_n20936_, new_n20937_, new_n20938_, new_n20939_, new_n20940_,
    new_n20941_, new_n20942_, new_n20943_, new_n20944_, new_n20945_,
    new_n20946_, new_n20947_, new_n20948_, new_n20949_, new_n20950_,
    new_n20951_, new_n20952_, new_n20953_, new_n20954_, new_n20955_,
    new_n20956_, new_n20957_, new_n20958_, new_n20959_, new_n20960_,
    new_n20961_, new_n20962_, new_n20963_, new_n20964_, new_n20965_,
    new_n20966_, new_n20967_, new_n20968_, new_n20969_, new_n20970_,
    new_n20971_, new_n20972_, new_n20973_, new_n20974_, new_n20975_,
    new_n20976_, new_n20977_, new_n20978_, new_n20979_, new_n20980_,
    new_n20981_, new_n20982_, new_n20983_, new_n20984_, new_n20985_,
    new_n20986_, new_n20987_, new_n20988_, new_n20989_, new_n20990_,
    new_n20991_, new_n20992_, new_n20993_, new_n20994_, new_n20995_,
    new_n20996_, new_n20997_, new_n20998_, new_n20999_, new_n21000_,
    new_n21001_, new_n21002_, new_n21003_, new_n21004_, new_n21005_,
    new_n21006_, new_n21007_, new_n21008_, new_n21009_, new_n21010_,
    new_n21011_, new_n21012_, new_n21013_, new_n21014_, new_n21015_,
    new_n21016_, new_n21017_, new_n21018_, new_n21019_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21028_, new_n21029_, new_n21030_,
    new_n21031_, new_n21032_, new_n21033_, new_n21034_, new_n21035_,
    new_n21036_, new_n21037_, new_n21038_, new_n21039_, new_n21040_,
    new_n21041_, new_n21042_, new_n21043_, new_n21044_, new_n21045_,
    new_n21046_, new_n21047_, new_n21048_, new_n21049_, new_n21050_,
    new_n21051_, new_n21052_, new_n21053_, new_n21054_, new_n21055_,
    new_n21056_, new_n21057_, new_n21058_, new_n21059_, new_n21060_,
    new_n21061_, new_n21062_, new_n21063_, new_n21064_, new_n21065_,
    new_n21066_, new_n21067_, new_n21068_, new_n21069_, new_n21070_,
    new_n21071_, new_n21072_, new_n21073_, new_n21074_, new_n21075_,
    new_n21076_, new_n21077_, new_n21078_, new_n21079_, new_n21080_,
    new_n21081_, new_n21082_, new_n21083_, new_n21084_, new_n21085_,
    new_n21086_, new_n21087_, new_n21088_, new_n21089_, new_n21090_,
    new_n21091_, new_n21092_, new_n21093_, new_n21094_, new_n21095_,
    new_n21096_, new_n21097_, new_n21098_, new_n21099_, new_n21100_,
    new_n21101_, new_n21102_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21109_, new_n21110_,
    new_n21111_, new_n21112_, new_n21113_, new_n21114_, new_n21115_,
    new_n21116_, new_n21117_, new_n21118_, new_n21119_, new_n21120_,
    new_n21121_, new_n21122_, new_n21123_, new_n21124_, new_n21125_,
    new_n21126_, new_n21127_, new_n21128_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21142_, new_n21143_, new_n21144_, new_n21145_,
    new_n21146_, new_n21147_, new_n21148_, new_n21149_, new_n21150_,
    new_n21151_, new_n21152_, new_n21153_, new_n21154_, new_n21155_,
    new_n21156_, new_n21157_, new_n21158_, new_n21159_, new_n21160_,
    new_n21161_, new_n21162_, new_n21163_, new_n21164_, new_n21165_,
    new_n21166_, new_n21167_, new_n21168_, new_n21169_, new_n21170_,
    new_n21171_, new_n21172_, new_n21173_, new_n21174_, new_n21175_,
    new_n21176_, new_n21177_, new_n21178_, new_n21179_, new_n21180_,
    new_n21181_, new_n21182_, new_n21183_, new_n21184_, new_n21185_,
    new_n21186_, new_n21187_, new_n21188_, new_n21189_, new_n21190_,
    new_n21191_, new_n21192_, new_n21193_, new_n21194_, new_n21195_,
    new_n21196_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21236_, new_n21237_, new_n21238_, new_n21239_, new_n21240_,
    new_n21241_, new_n21242_, new_n21243_, new_n21244_, new_n21245_,
    new_n21246_, new_n21247_, new_n21248_, new_n21249_, new_n21250_,
    new_n21251_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21275_,
    new_n21276_, new_n21277_, new_n21278_, new_n21279_, new_n21280_,
    new_n21281_, new_n21282_, new_n21283_, new_n21284_, new_n21285_,
    new_n21286_, new_n21287_, new_n21288_, new_n21289_, new_n21290_,
    new_n21291_, new_n21292_, new_n21293_, new_n21294_, new_n21295_,
    new_n21296_, new_n21297_, new_n21298_, new_n21299_, new_n21300_,
    new_n21301_, new_n21302_, new_n21303_, new_n21304_, new_n21305_,
    new_n21306_, new_n21307_, new_n21308_, new_n21309_, new_n21310_,
    new_n21311_, new_n21312_, new_n21313_, new_n21314_, new_n21315_,
    new_n21316_, new_n21317_, new_n21318_, new_n21319_, new_n21320_,
    new_n21321_, new_n21322_, new_n21323_, new_n21324_, new_n21325_,
    new_n21326_, new_n21327_, new_n21328_, new_n21329_, new_n21330_,
    new_n21331_, new_n21332_, new_n21333_, new_n21334_, new_n21335_,
    new_n21336_, new_n21337_, new_n21338_, new_n21339_, new_n21340_,
    new_n21341_, new_n21342_, new_n21343_, new_n21344_, new_n21345_,
    new_n21346_, new_n21347_, new_n21348_, new_n21349_, new_n21350_,
    new_n21351_, new_n21352_, new_n21353_, new_n21354_, new_n21355_,
    new_n21356_, new_n21357_, new_n21358_, new_n21359_, new_n21360_,
    new_n21361_, new_n21362_, new_n21363_, new_n21364_, new_n21365_,
    new_n21366_, new_n21367_, new_n21368_, new_n21369_, new_n21370_,
    new_n21371_, new_n21372_, new_n21373_, new_n21374_, new_n21375_,
    new_n21376_, new_n21377_, new_n21378_, new_n21379_, new_n21380_,
    new_n21381_, new_n21382_, new_n21383_, new_n21384_, new_n21385_,
    new_n21386_, new_n21387_, new_n21388_, new_n21389_, new_n21390_,
    new_n21391_, new_n21392_, new_n21393_, new_n21394_, new_n21395_,
    new_n21396_, new_n21397_, new_n21398_, new_n21399_, new_n21400_,
    new_n21401_, new_n21402_, new_n21403_, new_n21404_, new_n21405_,
    new_n21406_, new_n21407_, new_n21408_, new_n21409_, new_n21410_,
    new_n21411_, new_n21412_, new_n21413_, new_n21414_, new_n21415_,
    new_n21416_, new_n21417_, new_n21418_, new_n21419_, new_n21420_,
    new_n21421_, new_n21422_, new_n21423_, new_n21424_, new_n21425_,
    new_n21426_, new_n21427_, new_n21428_, new_n21429_, new_n21430_,
    new_n21431_, new_n21432_, new_n21433_, new_n21434_, new_n21435_,
    new_n21436_, new_n21437_, new_n21438_, new_n21439_, new_n21440_,
    new_n21441_, new_n21442_, new_n21443_, new_n21444_, new_n21445_,
    new_n21446_, new_n21447_, new_n21448_, new_n21449_, new_n21450_,
    new_n21451_, new_n21452_, new_n21453_, new_n21454_, new_n21455_,
    new_n21456_, new_n21457_, new_n21458_, new_n21459_, new_n21460_,
    new_n21461_, new_n21462_, new_n21463_, new_n21464_, new_n21465_,
    new_n21466_, new_n21467_, new_n21468_, new_n21469_, new_n21470_,
    new_n21471_, new_n21472_, new_n21473_, new_n21474_, new_n21475_,
    new_n21476_, new_n21477_, new_n21478_, new_n21479_, new_n21480_,
    new_n21481_, new_n21482_, new_n21483_, new_n21484_, new_n21485_,
    new_n21486_, new_n21487_, new_n21488_, new_n21489_, new_n21490_,
    new_n21491_, new_n21492_, new_n21493_, new_n21494_, new_n21495_,
    new_n21496_, new_n21497_, new_n21498_, new_n21499_, new_n21500_,
    new_n21501_, new_n21502_, new_n21503_, new_n21504_, new_n21505_,
    new_n21506_, new_n21507_, new_n21508_, new_n21509_, new_n21510_,
    new_n21511_, new_n21512_, new_n21513_, new_n21514_, new_n21515_,
    new_n21516_, new_n21517_, new_n21518_, new_n21519_, new_n21520_,
    new_n21521_, new_n21522_, new_n21523_, new_n21524_, new_n21525_,
    new_n21526_, new_n21527_, new_n21528_, new_n21529_, new_n21530_,
    new_n21531_, new_n21532_, new_n21533_, new_n21534_, new_n21535_,
    new_n21536_, new_n21537_, new_n21538_, new_n21539_, new_n21540_,
    new_n21541_, new_n21542_, new_n21543_, new_n21544_, new_n21545_,
    new_n21546_, new_n21547_, new_n21548_, new_n21549_, new_n21550_,
    new_n21551_, new_n21552_, new_n21553_, new_n21554_, new_n21555_,
    new_n21556_, new_n21557_, new_n21558_, new_n21559_, new_n21560_,
    new_n21561_, new_n21562_, new_n21563_, new_n21564_, new_n21565_,
    new_n21566_, new_n21567_, new_n21568_, new_n21569_, new_n21570_,
    new_n21571_, new_n21572_, new_n21573_, new_n21574_, new_n21575_,
    new_n21576_, new_n21577_, new_n21578_, new_n21579_, new_n21580_,
    new_n21581_, new_n21582_, new_n21583_, new_n21584_, new_n21585_,
    new_n21586_, new_n21587_, new_n21588_, new_n21589_, new_n21590_,
    new_n21591_, new_n21592_, new_n21593_, new_n21594_, new_n21595_,
    new_n21596_, new_n21597_, new_n21598_, new_n21599_, new_n21600_,
    new_n21601_, new_n21602_, new_n21603_, new_n21604_, new_n21605_,
    new_n21606_, new_n21607_, new_n21608_, new_n21609_, new_n21610_,
    new_n21611_, new_n21612_, new_n21613_, new_n21614_, new_n21615_,
    new_n21616_, new_n21617_, new_n21618_, new_n21619_, new_n21620_,
    new_n21621_, new_n21622_, new_n21623_, new_n21624_, new_n21625_,
    new_n21626_, new_n21627_, new_n21628_, new_n21629_, new_n21630_,
    new_n21631_, new_n21632_, new_n21633_, new_n21634_, new_n21635_,
    new_n21636_, new_n21637_, new_n21638_, new_n21639_, new_n21640_,
    new_n21641_, new_n21642_, new_n21643_, new_n21644_, new_n21645_,
    new_n21646_, new_n21647_, new_n21648_, new_n21649_, new_n21650_,
    new_n21651_, new_n21652_, new_n21653_, new_n21654_, new_n21655_,
    new_n21656_, new_n21657_, new_n21658_, new_n21659_, new_n21660_,
    new_n21661_, new_n21662_, new_n21663_, new_n21664_, new_n21665_,
    new_n21666_, new_n21667_, new_n21668_, new_n21669_, new_n21670_,
    new_n21671_, new_n21672_, new_n21673_, new_n21674_, new_n21675_,
    new_n21676_, new_n21677_, new_n21678_, new_n21679_, new_n21680_,
    new_n21681_, new_n21682_, new_n21683_, new_n21684_, new_n21685_,
    new_n21686_, new_n21687_, new_n21688_, new_n21689_, new_n21690_,
    new_n21691_, new_n21692_, new_n21693_, new_n21694_, new_n21695_,
    new_n21696_, new_n21697_, new_n21698_, new_n21699_, new_n21700_,
    new_n21701_, new_n21702_, new_n21703_, new_n21704_, new_n21705_,
    new_n21706_, new_n21707_, new_n21708_, new_n21709_, new_n21710_,
    new_n21711_, new_n21712_, new_n21713_, new_n21714_, new_n21715_,
    new_n21716_, new_n21717_, new_n21718_, new_n21719_, new_n21720_,
    new_n21721_, new_n21722_, new_n21723_, new_n21724_, new_n21725_,
    new_n21726_, new_n21727_, new_n21728_, new_n21729_, new_n21730_,
    new_n21731_, new_n21732_, new_n21733_, new_n21734_, new_n21735_,
    new_n21736_, new_n21737_, new_n21738_, new_n21739_, new_n21740_,
    new_n21741_, new_n21742_, new_n21743_, new_n21744_, new_n21745_,
    new_n21746_, new_n21747_, new_n21748_, new_n21749_, new_n21750_,
    new_n21751_, new_n21752_, new_n21753_, new_n21754_, new_n21755_,
    new_n21756_, new_n21757_, new_n21758_, new_n21759_, new_n21760_,
    new_n21761_, new_n21762_, new_n21763_, new_n21764_, new_n21765_,
    new_n21766_, new_n21767_, new_n21768_, new_n21769_, new_n21770_,
    new_n21771_, new_n21772_, new_n21773_, new_n21774_, new_n21775_,
    new_n21776_, new_n21777_, new_n21778_, new_n21779_, new_n21780_,
    new_n21781_, new_n21782_, new_n21783_, new_n21784_, new_n21785_,
    new_n21786_, new_n21787_, new_n21788_, new_n21789_, new_n21790_,
    new_n21791_, new_n21792_, new_n21793_, new_n21794_, new_n21795_,
    new_n21796_, new_n21797_, new_n21798_, new_n21799_, new_n21800_,
    new_n21801_, new_n21802_, new_n21803_, new_n21804_, new_n21805_,
    new_n21806_, new_n21807_, new_n21808_, new_n21809_, new_n21810_,
    new_n21811_, new_n21812_, new_n21813_, new_n21814_, new_n21815_,
    new_n21816_, new_n21817_, new_n21818_, new_n21819_, new_n21820_,
    new_n21821_, new_n21822_, new_n21823_, new_n21824_, new_n21825_,
    new_n21826_, new_n21827_, new_n21828_, new_n21829_, new_n21830_,
    new_n21831_, new_n21832_, new_n21833_, new_n21834_, new_n21835_,
    new_n21836_, new_n21837_, new_n21838_, new_n21839_, new_n21840_,
    new_n21841_, new_n21842_, new_n21843_, new_n21844_, new_n21845_,
    new_n21846_, new_n21847_, new_n21848_, new_n21849_, new_n21850_,
    new_n21851_, new_n21852_, new_n21853_, new_n21854_, new_n21855_,
    new_n21856_, new_n21857_, new_n21858_, new_n21859_, new_n21860_,
    new_n21861_, new_n21862_, new_n21863_, new_n21864_, new_n21865_,
    new_n21866_, new_n21867_, new_n21868_, new_n21869_, new_n21870_,
    new_n21871_, new_n21872_, new_n21873_, new_n21874_, new_n21875_,
    new_n21876_, new_n21877_, new_n21878_, new_n21879_, new_n21880_,
    new_n21881_, new_n21882_, new_n21883_, new_n21884_, new_n21885_,
    new_n21886_, new_n21887_, new_n21888_, new_n21889_, new_n21890_,
    new_n21891_, new_n21892_, new_n21893_, new_n21894_, new_n21895_,
    new_n21896_, new_n21897_, new_n21898_, new_n21899_, new_n21900_,
    new_n21901_, new_n21902_, new_n21903_, new_n21904_, new_n21905_,
    new_n21906_, new_n21907_, new_n21908_, new_n21909_, new_n21910_,
    new_n21911_, new_n21912_, new_n21913_, new_n21914_, new_n21915_,
    new_n21916_, new_n21917_, new_n21918_, new_n21919_, new_n21920_,
    new_n21921_, new_n21922_, new_n21923_, new_n21924_, new_n21925_,
    new_n21926_, new_n21927_, new_n21928_, new_n21929_, new_n21930_,
    new_n21931_, new_n21932_, new_n21933_, new_n21934_, new_n21935_,
    new_n21936_, new_n21937_, new_n21938_, new_n21939_, new_n21940_,
    new_n21941_, new_n21942_, new_n21943_, new_n21944_, new_n21945_,
    new_n21946_, new_n21947_, new_n21948_, new_n21949_, new_n21950_,
    new_n21951_, new_n21952_, new_n21953_, new_n21954_, new_n21955_,
    new_n21956_, new_n21957_, new_n21958_, new_n21959_, new_n21960_,
    new_n21961_, new_n21962_, new_n21963_, new_n21964_, new_n21965_,
    new_n21966_, new_n21967_, new_n21968_, new_n21969_, new_n21970_,
    new_n21971_, new_n21972_, new_n21973_, new_n21974_, new_n21975_,
    new_n21976_, new_n21977_, new_n21978_, new_n21979_, new_n21980_,
    new_n21981_, new_n21982_, new_n21983_, new_n21984_, new_n21985_,
    new_n21986_, new_n21987_, new_n21988_, new_n21989_, new_n21990_,
    new_n21991_, new_n21992_, new_n21993_, new_n21994_, new_n21995_,
    new_n21996_, new_n21997_, new_n21998_, new_n21999_, new_n22000_,
    new_n22001_, new_n22002_, new_n22003_, new_n22004_, new_n22005_,
    new_n22006_, new_n22007_, new_n22008_, new_n22009_, new_n22010_,
    new_n22011_, new_n22012_, new_n22013_, new_n22014_, new_n22015_,
    new_n22016_, new_n22017_, new_n22018_, new_n22019_, new_n22020_,
    new_n22021_, new_n22022_, new_n22023_, new_n22024_, new_n22025_,
    new_n22026_, new_n22027_, new_n22028_, new_n22029_, new_n22030_,
    new_n22031_, new_n22032_, new_n22033_, new_n22034_, new_n22035_,
    new_n22036_, new_n22037_, new_n22038_, new_n22039_, new_n22040_,
    new_n22041_, new_n22042_, new_n22043_, new_n22044_, new_n22045_,
    new_n22046_, new_n22047_, new_n22048_, new_n22049_, new_n22050_,
    new_n22051_, new_n22052_, new_n22053_, new_n22054_, new_n22055_,
    new_n22056_, new_n22057_, new_n22058_, new_n22059_, new_n22060_,
    new_n22061_, new_n22062_, new_n22063_, new_n22064_, new_n22065_,
    new_n22066_, new_n22067_, new_n22068_, new_n22069_, new_n22070_,
    new_n22071_, new_n22072_, new_n22073_, new_n22074_, new_n22075_,
    new_n22076_, new_n22077_, new_n22078_, new_n22079_, new_n22080_,
    new_n22081_, new_n22082_, new_n22083_, new_n22084_, new_n22085_,
    new_n22086_, new_n22087_, new_n22088_, new_n22089_, new_n22090_,
    new_n22091_, new_n22092_, new_n22093_, new_n22094_, new_n22095_,
    new_n22096_, new_n22097_, new_n22098_, new_n22099_, new_n22100_,
    new_n22101_, new_n22102_, new_n22103_, new_n22104_, new_n22105_,
    new_n22106_, new_n22107_, new_n22108_, new_n22109_, new_n22110_,
    new_n22111_, new_n22112_, new_n22113_, new_n22114_, new_n22115_,
    new_n22116_, new_n22117_, new_n22118_, new_n22119_, new_n22120_,
    new_n22121_, new_n22122_, new_n22123_, new_n22124_, new_n22125_,
    new_n22126_, new_n22127_, new_n22128_, new_n22129_, new_n22130_,
    new_n22131_, new_n22132_, new_n22133_, new_n22134_, new_n22135_,
    new_n22136_, new_n22137_, new_n22138_, new_n22139_, new_n22140_,
    new_n22141_, new_n22142_, new_n22143_, new_n22144_, new_n22145_,
    new_n22146_, new_n22147_, new_n22148_, new_n22149_, new_n22150_,
    new_n22151_, new_n22152_, new_n22153_, new_n22154_, new_n22155_,
    new_n22156_, new_n22157_, new_n22158_, new_n22159_, new_n22160_,
    new_n22161_, new_n22162_, new_n22163_, new_n22164_, new_n22165_,
    new_n22166_, new_n22167_, new_n22168_, new_n22169_, new_n22170_,
    new_n22171_, new_n22172_, new_n22173_, new_n22174_, new_n22175_,
    new_n22176_, new_n22177_, new_n22178_, new_n22179_, new_n22180_,
    new_n22181_, new_n22182_, new_n22183_, new_n22184_, new_n22185_,
    new_n22186_, new_n22187_, new_n22188_, new_n22189_, new_n22190_,
    new_n22191_, new_n22192_, new_n22193_, new_n22194_, new_n22195_,
    new_n22196_, new_n22197_, new_n22198_, new_n22199_, new_n22200_,
    new_n22201_, new_n22202_, new_n22203_, new_n22204_, new_n22205_,
    new_n22206_, new_n22207_, new_n22208_, new_n22209_, new_n22210_,
    new_n22211_, new_n22212_, new_n22213_, new_n22214_, new_n22215_,
    new_n22216_, new_n22217_, new_n22218_, new_n22219_, new_n22220_,
    new_n22221_, new_n22222_, new_n22223_, new_n22224_, new_n22225_,
    new_n22226_, new_n22227_, new_n22228_, new_n22229_, new_n22230_,
    new_n22231_, new_n22232_, new_n22233_, new_n22234_, new_n22235_,
    new_n22236_, new_n22237_, new_n22238_, new_n22239_, new_n22240_,
    new_n22241_, new_n22242_, new_n22243_, new_n22244_, new_n22245_,
    new_n22246_, new_n22247_, new_n22248_, new_n22249_, new_n22250_,
    new_n22251_, new_n22252_, new_n22253_, new_n22254_, new_n22255_,
    new_n22256_, new_n22257_, new_n22258_, new_n22259_, new_n22260_,
    new_n22261_, new_n22262_, new_n22263_, new_n22264_, new_n22265_,
    new_n22266_, new_n22267_, new_n22268_, new_n22269_, new_n22270_,
    new_n22271_, new_n22272_, new_n22273_, new_n22274_, new_n22275_,
    new_n22276_, new_n22277_, new_n22278_, new_n22279_, new_n22280_,
    new_n22281_, new_n22282_, new_n22283_, new_n22284_, new_n22285_,
    new_n22286_, new_n22287_, new_n22288_, new_n22289_, new_n22290_,
    new_n22291_, new_n22292_, new_n22293_, new_n22294_, new_n22295_,
    new_n22296_, new_n22297_, new_n22298_, new_n22299_, new_n22300_,
    new_n22301_, new_n22302_, new_n22303_, new_n22304_, new_n22305_,
    new_n22306_, new_n22307_, new_n22308_, new_n22309_, new_n22310_,
    new_n22311_, new_n22312_, new_n22313_, new_n22314_, new_n22315_,
    new_n22316_, new_n22317_, new_n22318_, new_n22319_, new_n22320_,
    new_n22321_, new_n22322_, new_n22323_, new_n22324_, new_n22325_,
    new_n22326_, new_n22327_, new_n22328_, new_n22329_, new_n22330_,
    new_n22331_, new_n22332_, new_n22333_, new_n22334_, new_n22335_,
    new_n22336_, new_n22337_, new_n22338_, new_n22339_, new_n22340_,
    new_n22341_, new_n22342_, new_n22343_, new_n22344_, new_n22345_,
    new_n22346_, new_n22347_, new_n22348_, new_n22349_, new_n22350_,
    new_n22351_, new_n22352_, new_n22353_, new_n22354_, new_n22355_,
    new_n22356_, new_n22357_, new_n22358_, new_n22359_, new_n22360_,
    new_n22361_, new_n22362_, new_n22363_, new_n22364_, new_n22365_,
    new_n22366_, new_n22367_, new_n22368_, new_n22369_, new_n22370_,
    new_n22371_, new_n22372_, new_n22373_, new_n22374_, new_n22375_,
    new_n22376_, new_n22377_, new_n22378_, new_n22379_, new_n22380_,
    new_n22381_, new_n22382_, new_n22383_, new_n22384_, new_n22385_,
    new_n22386_, new_n22387_, new_n22388_, new_n22389_, new_n22390_,
    new_n22391_, new_n22392_, new_n22393_, new_n22394_, new_n22395_,
    new_n22396_, new_n22397_, new_n22398_, new_n22399_, new_n22400_,
    new_n22401_, new_n22402_, new_n22403_, new_n22404_, new_n22405_,
    new_n22406_, new_n22407_, new_n22408_, new_n22409_, new_n22410_,
    new_n22411_, new_n22412_, new_n22413_, new_n22414_, new_n22415_,
    new_n22416_, new_n22417_, new_n22418_, new_n22419_, new_n22420_,
    new_n22421_, new_n22422_, new_n22423_, new_n22424_, new_n22425_,
    new_n22426_, new_n22427_, new_n22428_, new_n22429_, new_n22430_,
    new_n22431_, new_n22432_, new_n22433_, new_n22434_, new_n22435_,
    new_n22436_, new_n22437_, new_n22438_, new_n22439_, new_n22440_,
    new_n22441_, new_n22442_, new_n22443_, new_n22444_, new_n22445_,
    new_n22446_, new_n22447_, new_n22448_, new_n22449_, new_n22450_,
    new_n22451_, new_n22452_, new_n22453_, new_n22454_, new_n22455_,
    new_n22456_, new_n22457_, new_n22458_, new_n22459_, new_n22460_,
    new_n22461_, new_n22462_, new_n22463_, new_n22464_, new_n22465_,
    new_n22466_, new_n22467_, new_n22468_, new_n22469_, new_n22470_,
    new_n22471_, new_n22472_, new_n22473_, new_n22474_, new_n22475_,
    new_n22476_, new_n22477_, new_n22478_, new_n22479_, new_n22480_,
    new_n22481_, new_n22482_, new_n22483_, new_n22484_, new_n22485_,
    new_n22486_, new_n22487_, new_n22488_, new_n22489_, new_n22490_,
    new_n22491_, new_n22492_, new_n22493_, new_n22494_, new_n22495_,
    new_n22496_, new_n22497_, new_n22498_, new_n22499_, new_n22500_,
    new_n22501_, new_n22502_, new_n22503_, new_n22504_, new_n22505_,
    new_n22506_, new_n22507_, new_n22508_, new_n22509_, new_n22510_,
    new_n22511_, new_n22512_, new_n22513_, new_n22514_, new_n22515_,
    new_n22516_, new_n22517_, new_n22518_, new_n22519_, new_n22520_,
    new_n22521_, new_n22522_, new_n22523_, new_n22524_, new_n22525_,
    new_n22526_, new_n22527_, new_n22528_, new_n22529_, new_n22530_,
    new_n22531_, new_n22532_, new_n22533_, new_n22534_, new_n22535_,
    new_n22536_, new_n22537_, new_n22538_, new_n22539_, new_n22540_,
    new_n22541_, new_n22542_, new_n22543_, new_n22544_, new_n22545_,
    new_n22546_, new_n22547_, new_n22548_, new_n22549_, new_n22550_,
    new_n22551_, new_n22552_, new_n22553_, new_n22554_, new_n22555_,
    new_n22556_, new_n22557_, new_n22558_, new_n22559_, new_n22560_,
    new_n22561_, new_n22562_, new_n22563_, new_n22564_, new_n22565_,
    new_n22566_, new_n22567_, new_n22568_, new_n22569_, new_n22570_,
    new_n22571_, new_n22572_, new_n22573_, new_n22574_, new_n22575_,
    new_n22576_, new_n22577_, new_n22578_, new_n22579_, new_n22580_,
    new_n22581_, new_n22582_, new_n22583_, new_n22584_, new_n22585_,
    new_n22586_, new_n22587_, new_n22588_, new_n22589_, new_n22590_,
    new_n22591_, new_n22592_, new_n22593_, new_n22594_, new_n22595_,
    new_n22596_, new_n22597_, new_n22598_, new_n22599_, new_n22600_,
    new_n22601_, new_n22602_, new_n22603_, new_n22604_, new_n22605_,
    new_n22606_, new_n22607_, new_n22608_, new_n22609_, new_n22610_,
    new_n22611_, new_n22612_, new_n22613_, new_n22614_, new_n22615_,
    new_n22616_, new_n22617_, new_n22618_, new_n22619_, new_n22620_,
    new_n22621_, new_n22622_, new_n22623_, new_n22624_, new_n22625_,
    new_n22626_, new_n22627_, new_n22628_, new_n22629_, new_n22630_,
    new_n22631_, new_n22632_, new_n22633_, new_n22634_, new_n22635_,
    new_n22636_, new_n22637_, new_n22638_, new_n22639_, new_n22640_,
    new_n22641_, new_n22642_, new_n22643_, new_n22644_, new_n22645_,
    new_n22646_, new_n22647_, new_n22648_, new_n22649_, new_n22650_,
    new_n22651_, new_n22652_, new_n22653_, new_n22654_, new_n22655_,
    new_n22656_, new_n22657_, new_n22658_, new_n22659_, new_n22660_,
    new_n22661_, new_n22662_, new_n22663_, new_n22664_, new_n22665_,
    new_n22666_, new_n22667_, new_n22668_, new_n22669_, new_n22670_,
    new_n22671_, new_n22672_, new_n22673_, new_n22674_, new_n22675_,
    new_n22676_, new_n22677_, new_n22678_, new_n22679_, new_n22680_,
    new_n22681_, new_n22682_, new_n22683_, new_n22684_, new_n22685_,
    new_n22686_, new_n22687_, new_n22688_, new_n22689_, new_n22690_,
    new_n22691_, new_n22692_, new_n22693_, new_n22694_, new_n22695_,
    new_n22696_, new_n22697_, new_n22698_, new_n22699_, new_n22700_,
    new_n22701_, new_n22702_, new_n22703_, new_n22704_, new_n22705_,
    new_n22706_, new_n22707_, new_n22708_, new_n22709_, new_n22710_,
    new_n22711_, new_n22712_, new_n22713_, new_n22714_, new_n22715_,
    new_n22716_, new_n22717_, new_n22718_, new_n22719_, new_n22720_,
    new_n22721_, new_n22722_, new_n22723_, new_n22724_, new_n22725_,
    new_n22726_, new_n22727_, new_n22728_, new_n22729_, new_n22730_,
    new_n22731_, new_n22732_, new_n22733_, new_n22734_, new_n22735_,
    new_n22736_, new_n22737_, new_n22738_, new_n22739_, new_n22740_,
    new_n22741_, new_n22742_, new_n22743_, new_n22744_, new_n22745_,
    new_n22746_, new_n22747_, new_n22748_, new_n22749_, new_n22750_,
    new_n22751_, new_n22752_, new_n22753_, new_n22754_, new_n22755_,
    new_n22756_, new_n22757_, new_n22758_, new_n22759_, new_n22760_,
    new_n22761_, new_n22762_, new_n22763_, new_n22764_, new_n22765_,
    new_n22766_, new_n22767_, new_n22768_, new_n22769_, new_n22770_,
    new_n22771_, new_n22772_, new_n22773_, new_n22774_, new_n22775_,
    new_n22776_, new_n22777_, new_n22778_, new_n22779_, new_n22780_,
    new_n22781_, new_n22782_, new_n22783_, new_n22784_, new_n22785_,
    new_n22786_, new_n22787_, new_n22788_, new_n22789_, new_n22790_,
    new_n22791_, new_n22792_, new_n22793_, new_n22794_, new_n22795_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22891_, new_n22892_, new_n22893_, new_n22894_, new_n22895_,
    new_n22896_, new_n22897_, new_n22898_, new_n22899_, new_n22900_,
    new_n22901_, new_n22902_, new_n22903_, new_n22904_, new_n22905_,
    new_n22906_, new_n22907_, new_n22908_, new_n22909_, new_n22910_,
    new_n22911_, new_n22912_, new_n22913_, new_n22914_, new_n22915_,
    new_n22916_, new_n22917_, new_n22918_, new_n22919_, new_n22920_,
    new_n22921_, new_n22922_, new_n22923_, new_n22924_, new_n22925_,
    new_n22926_, new_n22927_, new_n22928_, new_n22929_, new_n22930_,
    new_n22931_, new_n22932_, new_n22933_, new_n22934_, new_n22935_,
    new_n22936_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22942_, new_n22943_, new_n22944_, new_n22945_,
    new_n22946_, new_n22947_, new_n22948_, new_n22949_, new_n22950_,
    new_n22951_, new_n22952_, new_n22953_, new_n22954_, new_n22955_,
    new_n22956_, new_n22957_, new_n22958_, new_n22959_, new_n22960_,
    new_n22961_, new_n22962_, new_n22963_, new_n22964_, new_n22965_,
    new_n22966_, new_n22967_, new_n22968_, new_n22969_, new_n22970_,
    new_n22971_, new_n22972_, new_n22973_, new_n22974_, new_n22975_,
    new_n22976_, new_n22977_, new_n22978_, new_n22979_, new_n22980_,
    new_n22981_, new_n22982_, new_n22983_, new_n22984_, new_n22985_,
    new_n22986_, new_n22987_, new_n22988_, new_n22989_, new_n22990_,
    new_n22991_, new_n22992_, new_n22993_, new_n22994_, new_n22995_,
    new_n22996_, new_n22997_, new_n22998_, new_n22999_, new_n23000_,
    new_n23001_, new_n23002_, new_n23003_, new_n23004_, new_n23005_,
    new_n23006_, new_n23007_, new_n23008_, new_n23009_, new_n23010_,
    new_n23011_, new_n23012_, new_n23013_, new_n23014_, new_n23015_,
    new_n23016_, new_n23017_, new_n23018_, new_n23019_, new_n23020_,
    new_n23021_, new_n23022_, new_n23023_, new_n23024_, new_n23025_,
    new_n23026_, new_n23027_, new_n23028_, new_n23029_, new_n23030_,
    new_n23031_, new_n23032_, new_n23033_, new_n23034_, new_n23035_,
    new_n23036_, new_n23037_, new_n23038_, new_n23039_, new_n23040_,
    new_n23041_, new_n23042_, new_n23043_, new_n23044_, new_n23045_,
    new_n23046_, new_n23047_, new_n23048_, new_n23049_, new_n23050_,
    new_n23051_, new_n23052_, new_n23053_, new_n23054_, new_n23055_,
    new_n23056_, new_n23057_, new_n23058_, new_n23059_, new_n23060_,
    new_n23061_, new_n23062_, new_n23063_, new_n23064_, new_n23065_,
    new_n23066_, new_n23067_, new_n23068_, new_n23069_, new_n23070_,
    new_n23071_, new_n23072_, new_n23073_, new_n23074_, new_n23075_,
    new_n23076_, new_n23077_, new_n23078_, new_n23079_, new_n23080_,
    new_n23081_, new_n23082_, new_n23083_, new_n23084_, new_n23085_,
    new_n23086_, new_n23087_, new_n23088_, new_n23089_, new_n23090_,
    new_n23091_, new_n23092_, new_n23093_, new_n23094_, new_n23095_,
    new_n23096_, new_n23097_, new_n23098_, new_n23099_, new_n23100_,
    new_n23101_, new_n23102_, new_n23103_, new_n23104_, new_n23105_,
    new_n23106_, new_n23107_, new_n23108_, new_n23109_, new_n23110_,
    new_n23111_, new_n23112_, new_n23113_, new_n23114_, new_n23115_,
    new_n23116_, new_n23117_, new_n23118_, new_n23119_, new_n23120_,
    new_n23121_, new_n23122_, new_n23123_, new_n23124_, new_n23125_,
    new_n23126_, new_n23127_, new_n23128_, new_n23129_, new_n23130_,
    new_n23131_, new_n23132_, new_n23133_, new_n23134_, new_n23135_,
    new_n23136_, new_n23137_, new_n23138_, new_n23139_, new_n23140_,
    new_n23141_, new_n23142_, new_n23143_, new_n23144_, new_n23145_,
    new_n23146_, new_n23147_, new_n23148_, new_n23149_, new_n23150_,
    new_n23151_, new_n23152_, new_n23153_, new_n23154_, new_n23155_,
    new_n23156_, new_n23157_, new_n23158_, new_n23159_, new_n23160_,
    new_n23161_, new_n23162_, new_n23163_, new_n23164_, new_n23165_,
    new_n23166_, new_n23167_, new_n23168_, new_n23169_, new_n23170_,
    new_n23171_, new_n23172_, new_n23173_, new_n23174_, new_n23175_,
    new_n23176_, new_n23177_, new_n23178_, new_n23179_, new_n23180_,
    new_n23181_, new_n23182_, new_n23183_, new_n23184_, new_n23185_,
    new_n23186_, new_n23187_, new_n23188_, new_n23189_, new_n23190_,
    new_n23191_, new_n23192_, new_n23193_, new_n23194_, new_n23195_,
    new_n23196_, new_n23197_, new_n23198_, new_n23199_, new_n23200_,
    new_n23201_, new_n23202_, new_n23203_, new_n23204_, new_n23205_,
    new_n23206_, new_n23207_, new_n23208_, new_n23209_, new_n23210_,
    new_n23211_, new_n23212_, new_n23213_, new_n23214_, new_n23215_,
    new_n23216_, new_n23217_, new_n23218_, new_n23219_, new_n23220_,
    new_n23221_, new_n23222_, new_n23223_, new_n23224_, new_n23225_,
    new_n23226_, new_n23227_, new_n23228_, new_n23229_, new_n23230_,
    new_n23231_, new_n23232_, new_n23233_, new_n23234_, new_n23235_,
    new_n23236_, new_n23237_, new_n23238_, new_n23239_, new_n23240_,
    new_n23241_, new_n23242_, new_n23243_, new_n23244_, new_n23245_,
    new_n23246_, new_n23247_, new_n23248_, new_n23249_, new_n23250_,
    new_n23251_, new_n23252_, new_n23253_, new_n23254_, new_n23255_,
    new_n23256_, new_n23257_, new_n23258_, new_n23259_, new_n23260_,
    new_n23261_, new_n23262_, new_n23263_, new_n23264_, new_n23265_,
    new_n23266_, new_n23267_, new_n23268_, new_n23269_, new_n23270_,
    new_n23271_, new_n23272_, new_n23273_, new_n23274_, new_n23275_,
    new_n23276_, new_n23277_, new_n23278_, new_n23279_, new_n23280_,
    new_n23281_, new_n23282_, new_n23283_, new_n23284_, new_n23285_,
    new_n23286_, new_n23287_, new_n23288_, new_n23289_, new_n23290_,
    new_n23291_, new_n23292_, new_n23293_, new_n23294_, new_n23295_,
    new_n23296_, new_n23297_, new_n23298_, new_n23299_, new_n23300_,
    new_n23301_, new_n23302_, new_n23303_, new_n23304_, new_n23305_,
    new_n23306_, new_n23307_, new_n23308_, new_n23309_, new_n23310_,
    new_n23311_, new_n23312_, new_n23313_, new_n23314_, new_n23315_,
    new_n23316_, new_n23317_, new_n23318_, new_n23319_, new_n23320_,
    new_n23321_, new_n23322_, new_n23323_, new_n23324_, new_n23325_,
    new_n23326_, new_n23327_, new_n23328_, new_n23329_, new_n23330_,
    new_n23331_, new_n23332_, new_n23333_, new_n23334_, new_n23335_,
    new_n23336_, new_n23337_, new_n23338_, new_n23339_, new_n23340_,
    new_n23341_, new_n23342_, new_n23343_, new_n23344_, new_n23345_,
    new_n23346_, new_n23347_, new_n23348_, new_n23349_, new_n23350_,
    new_n23351_, new_n23352_, new_n23353_, new_n23354_, new_n23355_,
    new_n23356_, new_n23357_, new_n23358_, new_n23359_, new_n23360_,
    new_n23361_, new_n23362_, new_n23363_, new_n23364_, new_n23365_,
    new_n23366_, new_n23367_, new_n23368_, new_n23369_, new_n23370_,
    new_n23371_, new_n23372_, new_n23373_, new_n23374_, new_n23375_,
    new_n23376_, new_n23377_, new_n23378_, new_n23379_, new_n23380_,
    new_n23381_, new_n23382_, new_n23383_, new_n23384_, new_n23385_,
    new_n23386_, new_n23387_, new_n23388_, new_n23389_, new_n23390_,
    new_n23391_, new_n23392_, new_n23393_, new_n23394_, new_n23395_,
    new_n23396_, new_n23397_, new_n23398_, new_n23399_, new_n23400_,
    new_n23401_, new_n23402_, new_n23403_, new_n23404_, new_n23405_,
    new_n23406_, new_n23407_, new_n23408_, new_n23409_, new_n23410_,
    new_n23411_, new_n23412_, new_n23413_, new_n23414_, new_n23415_,
    new_n23416_, new_n23417_, new_n23418_, new_n23419_, new_n23420_,
    new_n23421_, new_n23422_, new_n23423_, new_n23424_, new_n23425_,
    new_n23426_, new_n23427_, new_n23428_, new_n23429_, new_n23430_,
    new_n23431_, new_n23432_, new_n23433_, new_n23434_, new_n23435_,
    new_n23436_, new_n23437_, new_n23438_, new_n23439_, new_n23440_,
    new_n23441_, new_n23442_, new_n23443_, new_n23444_, new_n23445_,
    new_n23446_, new_n23447_, new_n23448_, new_n23449_, new_n23450_,
    new_n23451_, new_n23452_, new_n23453_, new_n23454_, new_n23455_,
    new_n23456_, new_n23457_, new_n23458_, new_n23459_, new_n23460_,
    new_n23461_, new_n23462_, new_n23463_, new_n23464_, new_n23465_,
    new_n23466_, new_n23467_, new_n23468_, new_n23469_, new_n23470_,
    new_n23471_, new_n23472_, new_n23473_, new_n23474_, new_n23475_,
    new_n23476_, new_n23477_, new_n23478_, new_n23479_, new_n23480_,
    new_n23481_, new_n23482_, new_n23483_, new_n23484_, new_n23485_,
    new_n23486_, new_n23487_, new_n23488_, new_n23489_, new_n23490_,
    new_n23491_, new_n23492_, new_n23493_, new_n23494_, new_n23495_,
    new_n23496_, new_n23497_, new_n23498_, new_n23499_, new_n23500_,
    new_n23501_, new_n23502_, new_n23503_, new_n23504_, new_n23505_,
    new_n23506_, new_n23507_, new_n23508_, new_n23509_, new_n23510_,
    new_n23511_, new_n23512_, new_n23513_, new_n23514_, new_n23515_,
    new_n23516_, new_n23517_, new_n23518_, new_n23519_, new_n23520_,
    new_n23521_, new_n23522_, new_n23523_, new_n23524_, new_n23525_,
    new_n23526_, new_n23527_, new_n23528_, new_n23529_, new_n23530_,
    new_n23531_, new_n23532_, new_n23533_, new_n23534_, new_n23535_,
    new_n23536_, new_n23537_, new_n23538_, new_n23539_, new_n23540_,
    new_n23541_, new_n23542_, new_n23543_, new_n23544_, new_n23545_,
    new_n23546_, new_n23547_, new_n23548_, new_n23549_, new_n23550_,
    new_n23551_, new_n23552_, new_n23553_, new_n23554_, new_n23555_,
    new_n23556_, new_n23557_, new_n23558_, new_n23559_, new_n23560_,
    new_n23561_, new_n23562_, new_n23563_, new_n23564_, new_n23565_,
    new_n23566_, new_n23567_, new_n23568_, new_n23569_, new_n23570_,
    new_n23571_, new_n23572_, new_n23573_, new_n23574_, new_n23575_,
    new_n23576_, new_n23577_, new_n23578_, new_n23579_, new_n23580_,
    new_n23581_, new_n23582_, new_n23583_, new_n23584_, new_n23585_,
    new_n23586_, new_n23587_, new_n23588_, new_n23589_, new_n23590_,
    new_n23591_, new_n23592_, new_n23593_, new_n23594_, new_n23595_,
    new_n23596_, new_n23597_, new_n23598_, new_n23599_, new_n23600_,
    new_n23601_, new_n23602_, new_n23603_, new_n23604_, new_n23605_,
    new_n23606_, new_n23607_, new_n23608_, new_n23609_, new_n23610_,
    new_n23611_, new_n23612_, new_n23613_, new_n23614_, new_n23615_,
    new_n23616_, new_n23617_, new_n23618_, new_n23619_, new_n23620_,
    new_n23621_, new_n23622_, new_n23623_, new_n23624_, new_n23625_,
    new_n23626_, new_n23627_, new_n23628_, new_n23629_, new_n23630_,
    new_n23631_, new_n23632_, new_n23633_, new_n23634_, new_n23635_,
    new_n23636_, new_n23637_, new_n23638_, new_n23639_, new_n23640_,
    new_n23641_, new_n23642_, new_n23643_, new_n23644_, new_n23645_,
    new_n23646_, new_n23647_, new_n23648_, new_n23649_, new_n23650_,
    new_n23651_, new_n23652_, new_n23653_, new_n23654_, new_n23655_,
    new_n23656_, new_n23657_, new_n23658_, new_n23659_, new_n23660_,
    new_n23661_, new_n23662_, new_n23663_, new_n23664_, new_n23665_,
    new_n23666_, new_n23667_, new_n23668_, new_n23669_, new_n23670_,
    new_n23671_, new_n23672_, new_n23673_, new_n23674_, new_n23675_,
    new_n23676_, new_n23677_, new_n23678_, new_n23679_, new_n23680_,
    new_n23681_, new_n23682_, new_n23683_, new_n23684_, new_n23685_,
    new_n23686_, new_n23687_, new_n23688_, new_n23689_, new_n23690_,
    new_n23691_, new_n23692_, new_n23693_, new_n23694_, new_n23695_,
    new_n23696_, new_n23697_, new_n23698_, new_n23699_, new_n23700_,
    new_n23701_, new_n23702_, new_n23703_, new_n23704_, new_n23705_,
    new_n23706_, new_n23707_, new_n23708_, new_n23709_, new_n23710_,
    new_n23711_, new_n23712_, new_n23713_, new_n23714_, new_n23715_,
    new_n23716_, new_n23717_, new_n23718_, new_n23719_, new_n23720_,
    new_n23721_, new_n23722_, new_n23723_, new_n23724_, new_n23725_,
    new_n23726_, new_n23727_, new_n23728_, new_n23729_, new_n23730_,
    new_n23731_, new_n23732_, new_n23733_, new_n23734_, new_n23735_,
    new_n23736_, new_n23737_, new_n23738_, new_n23739_, new_n23740_,
    new_n23741_, new_n23742_, new_n23743_, new_n23744_, new_n23745_,
    new_n23746_, new_n23747_, new_n23748_, new_n23749_, new_n23750_,
    new_n23751_, new_n23752_, new_n23753_, new_n23754_, new_n23755_,
    new_n23756_, new_n23757_, new_n23758_, new_n23759_, new_n23760_,
    new_n23761_, new_n23762_, new_n23763_, new_n23764_, new_n23765_,
    new_n23766_, new_n23767_, new_n23768_, new_n23769_, new_n23770_,
    new_n23771_, new_n23772_, new_n23773_, new_n23774_, new_n23775_,
    new_n23776_, new_n23777_, new_n23778_, new_n23779_, new_n23780_,
    new_n23781_, new_n23782_, new_n23783_, new_n23784_, new_n23785_,
    new_n23786_, new_n23787_, new_n23788_, new_n23789_, new_n23790_,
    new_n23791_, new_n23792_, new_n23793_, new_n23794_, new_n23795_,
    new_n23796_, new_n23797_, new_n23798_, new_n23799_, new_n23800_,
    new_n23801_, new_n23802_, new_n23803_, new_n23804_, new_n23805_,
    new_n23806_, new_n23807_, new_n23808_, new_n23809_, new_n23810_,
    new_n23811_, new_n23812_, new_n23813_, new_n23814_, new_n23815_,
    new_n23816_, new_n23817_, new_n23818_, new_n23819_, new_n23820_,
    new_n23821_, new_n23822_, new_n23823_, new_n23824_, new_n23825_,
    new_n23826_, new_n23827_, new_n23828_, new_n23829_, new_n23830_,
    new_n23831_, new_n23832_, new_n23833_, new_n23834_, new_n23835_,
    new_n23836_, new_n23837_, new_n23838_, new_n23839_, new_n23840_,
    new_n23841_, new_n23842_, new_n23843_, new_n23844_, new_n23845_,
    new_n23846_, new_n23847_, new_n23848_, new_n23849_, new_n23850_,
    new_n23851_, new_n23852_, new_n23853_, new_n23854_, new_n23855_,
    new_n23856_, new_n23857_, new_n23858_, new_n23859_, new_n23860_,
    new_n23861_, new_n23862_, new_n23863_, new_n23864_, new_n23865_,
    new_n23866_, new_n23867_, new_n23868_, new_n23869_, new_n23870_,
    new_n23871_, new_n23872_, new_n23873_, new_n23874_, new_n23875_,
    new_n23876_, new_n23877_, new_n23878_, new_n23879_, new_n23880_,
    new_n23881_, new_n23882_, new_n23883_, new_n23884_, new_n23885_,
    new_n23886_, new_n23887_, new_n23888_, new_n23889_, new_n23890_,
    new_n23891_, new_n23892_, new_n23893_, new_n23894_, new_n23895_,
    new_n23896_, new_n23897_, new_n23898_, new_n23899_, new_n23900_,
    new_n23901_, new_n23902_, new_n23903_, new_n23904_, new_n23905_,
    new_n23906_, new_n23907_, new_n23908_, new_n23909_, new_n23910_,
    new_n23911_, new_n23912_, new_n23913_, new_n23914_, new_n23915_,
    new_n23916_, new_n23917_, new_n23918_, new_n23919_, new_n23920_,
    new_n23921_, new_n23922_, new_n23923_, new_n23924_, new_n23925_,
    new_n23926_, new_n23927_, new_n23928_, new_n23929_, new_n23930_,
    new_n23931_, new_n23932_, new_n23933_, new_n23934_, new_n23935_,
    new_n23936_, new_n23937_, new_n23938_, new_n23939_, new_n23940_,
    new_n23941_, new_n23942_, new_n23943_, new_n23944_, new_n23945_,
    new_n23946_, new_n23947_, new_n23948_, new_n23949_, new_n23950_,
    new_n23951_, new_n23952_, new_n23953_, new_n23954_, new_n23955_,
    new_n23956_, new_n23957_, new_n23958_, new_n23959_, new_n23960_,
    new_n23961_, new_n23962_, new_n23963_, new_n23964_, new_n23965_,
    new_n23966_, new_n23967_, new_n23968_, new_n23969_, new_n23970_,
    new_n23971_, new_n23972_, new_n23973_, new_n23974_, new_n23975_,
    new_n23976_, new_n23977_, new_n23978_, new_n23979_, new_n23980_,
    new_n23981_, new_n23982_, new_n23983_, new_n23984_, new_n23985_,
    new_n23986_, new_n23987_, new_n23988_, new_n23989_, new_n23990_,
    new_n23991_, new_n23992_, new_n23993_, new_n23994_, new_n23995_,
    new_n23996_, new_n23997_, new_n23998_, new_n23999_, new_n24000_,
    new_n24001_, new_n24002_, new_n24003_, new_n24004_, new_n24005_,
    new_n24006_, new_n24007_, new_n24008_, new_n24009_, new_n24010_,
    new_n24011_, new_n24012_, new_n24013_, new_n24014_, new_n24015_,
    new_n24016_, new_n24017_, new_n24018_, new_n24019_, new_n24020_,
    new_n24021_, new_n24022_, new_n24023_, new_n24024_, new_n24025_,
    new_n24026_, new_n24027_, new_n24028_, new_n24029_, new_n24030_,
    new_n24031_, new_n24032_, new_n24033_, new_n24034_, new_n24035_,
    new_n24036_, new_n24037_, new_n24038_, new_n24039_, new_n24040_,
    new_n24041_, new_n24042_, new_n24043_, new_n24044_, new_n24045_,
    new_n24046_, new_n24047_, new_n24048_, new_n24049_, new_n24050_,
    new_n24051_, new_n24052_, new_n24053_, new_n24054_, new_n24055_,
    new_n24056_, new_n24057_, new_n24058_, new_n24059_, new_n24060_,
    new_n24061_, new_n24062_, new_n24063_, new_n24064_, new_n24065_,
    new_n24066_, new_n24067_, new_n24068_, new_n24069_, new_n24070_,
    new_n24071_, new_n24072_, new_n24073_, new_n24074_, new_n24075_,
    new_n24076_, new_n24077_, new_n24078_, new_n24079_, new_n24080_,
    new_n24081_, new_n24082_, new_n24083_, new_n24084_, new_n24085_,
    new_n24086_, new_n24087_, new_n24088_, new_n24089_, new_n24090_,
    new_n24091_, new_n24092_, new_n24093_, new_n24094_, new_n24095_,
    new_n24096_, new_n24097_, new_n24098_, new_n24099_, new_n24100_,
    new_n24101_, new_n24102_, new_n24103_, new_n24104_, new_n24105_,
    new_n24106_, new_n24107_, new_n24108_, new_n24109_, new_n24110_,
    new_n24111_, new_n24112_, new_n24113_, new_n24114_, new_n24115_,
    new_n24116_, new_n24117_, new_n24118_, new_n24119_, new_n24120_,
    new_n24121_, new_n24122_, new_n24123_, new_n24124_, new_n24125_,
    new_n24126_, new_n24127_, new_n24128_, new_n24129_, new_n24130_,
    new_n24131_, new_n24132_, new_n24133_, new_n24134_, new_n24135_,
    new_n24136_, new_n24137_, new_n24138_, new_n24139_, new_n24140_,
    new_n24141_, new_n24142_, new_n24143_, new_n24144_, new_n24145_,
    new_n24146_, new_n24147_, new_n24148_, new_n24149_, new_n24150_,
    new_n24151_, new_n24152_, new_n24153_, new_n24154_, new_n24155_,
    new_n24156_, new_n24157_, new_n24158_, new_n24159_, new_n24160_,
    new_n24161_, new_n24162_, new_n24163_, new_n24164_, new_n24165_,
    new_n24166_, new_n24167_, new_n24168_, new_n24169_, new_n24170_,
    new_n24171_, new_n24172_, new_n24173_, new_n24174_, new_n24175_,
    new_n24176_, new_n24177_, new_n24178_, new_n24179_, new_n24180_,
    new_n24181_, new_n24182_, new_n24183_, new_n24184_, new_n24185_,
    new_n24186_, new_n24187_, new_n24188_, new_n24189_, new_n24190_,
    new_n24191_, new_n24192_, new_n24193_, new_n24194_, new_n24195_,
    new_n24196_, new_n24197_, new_n24198_, new_n24199_, new_n24200_,
    new_n24201_, new_n24202_, new_n24203_, new_n24204_, new_n24205_,
    new_n24206_, new_n24207_, new_n24208_, new_n24209_, new_n24210_,
    new_n24211_, new_n24212_, new_n24213_, new_n24214_, new_n24215_,
    new_n24216_, new_n24217_, new_n24218_, new_n24219_, new_n24220_,
    new_n24221_, new_n24222_, new_n24223_, new_n24224_, new_n24225_,
    new_n24226_, new_n24227_, new_n24228_, new_n24229_, new_n24230_,
    new_n24231_, new_n24232_, new_n24233_, new_n24234_, new_n24235_,
    new_n24236_, new_n24237_, new_n24238_, new_n24239_, new_n24240_,
    new_n24241_, new_n24242_, new_n24243_, new_n24244_, new_n24245_,
    new_n24246_, new_n24247_, new_n24248_, new_n24249_, new_n24250_,
    new_n24251_, new_n24252_, new_n24253_, new_n24254_, new_n24255_,
    new_n24256_, new_n24257_, new_n24258_, new_n24259_, new_n24260_,
    new_n24261_, new_n24262_, new_n24263_, new_n24264_, new_n24265_,
    new_n24266_, new_n24267_, new_n24268_, new_n24269_, new_n24270_,
    new_n24271_, new_n24272_, new_n24273_, new_n24274_, new_n24275_,
    new_n24276_, new_n24277_, new_n24278_, new_n24279_, new_n24280_,
    new_n24281_, new_n24282_, new_n24283_, new_n24284_, new_n24285_,
    new_n24286_, new_n24287_, new_n24288_, new_n24289_, new_n24290_,
    new_n24291_, new_n24292_, new_n24293_, new_n24294_, new_n24295_,
    new_n24296_, new_n24297_, new_n24298_, new_n24299_, new_n24300_,
    new_n24301_, new_n24302_, new_n24303_, new_n24304_, new_n24305_,
    new_n24306_, new_n24307_, new_n24308_, new_n24309_, new_n24310_,
    new_n24311_, new_n24312_, new_n24313_, new_n24314_, new_n24315_,
    new_n24316_, new_n24317_, new_n24318_, new_n24319_, new_n24320_,
    new_n24321_, new_n24322_, new_n24323_, new_n24324_, new_n24325_,
    new_n24326_, new_n24327_, new_n24328_, new_n24329_, new_n24330_,
    new_n24331_, new_n24332_, new_n24333_, new_n24334_, new_n24335_,
    new_n24336_, new_n24337_, new_n24338_, new_n24339_, new_n24340_,
    new_n24341_, new_n24342_, new_n24343_, new_n24344_, new_n24345_,
    new_n24346_, new_n24347_, new_n24348_, new_n24349_, new_n24350_,
    new_n24351_, new_n24352_, new_n24353_, new_n24354_, new_n24355_,
    new_n24356_, new_n24357_, new_n24358_, new_n24359_, new_n24360_,
    new_n24361_, new_n24362_, new_n24363_, new_n24364_, new_n24365_,
    new_n24366_, new_n24367_, new_n24368_, new_n24369_, new_n24370_,
    new_n24371_, new_n24372_, new_n24373_, new_n24374_, new_n24375_,
    new_n24376_, new_n24377_, new_n24378_, new_n24379_, new_n24380_,
    new_n24381_, new_n24382_, new_n24383_, new_n24384_, new_n24385_,
    new_n24386_, new_n24387_, new_n24388_, new_n24389_, new_n24390_,
    new_n24391_, new_n24392_, new_n24393_, new_n24394_, new_n24395_,
    new_n24396_, new_n24397_, new_n24398_, new_n24399_, new_n24400_,
    new_n24401_, new_n24402_, new_n24403_, new_n24404_, new_n24405_,
    new_n24406_, new_n24407_, new_n24408_, new_n24409_, new_n24410_,
    new_n24411_, new_n24412_, new_n24413_, new_n24414_, new_n24415_,
    new_n24416_, new_n24417_, new_n24418_, new_n24419_, new_n24420_,
    new_n24421_, new_n24422_, new_n24423_, new_n24424_, new_n24425_,
    new_n24426_, new_n24427_, new_n24428_, new_n24429_, new_n24430_,
    new_n24431_, new_n24432_, new_n24433_, new_n24434_, new_n24435_,
    new_n24436_, new_n24437_, new_n24438_, new_n24439_, new_n24440_,
    new_n24441_, new_n24442_, new_n24443_, new_n24444_, new_n24445_,
    new_n24446_, new_n24447_, new_n24448_, new_n24449_, new_n24450_,
    new_n24451_, new_n24452_, new_n24453_, new_n24454_, new_n24455_,
    new_n24456_, new_n24457_, new_n24458_, new_n24459_, new_n24460_,
    new_n24461_, new_n24462_, new_n24463_, new_n24464_, new_n24465_,
    new_n24466_, new_n24467_, new_n24468_, new_n24469_, new_n24470_,
    new_n24471_, new_n24472_, new_n24473_, new_n24474_, new_n24475_,
    new_n24476_, new_n24477_, new_n24478_, new_n24479_, new_n24480_,
    new_n24481_, new_n24482_, new_n24483_, new_n24484_, new_n24485_,
    new_n24486_, new_n24487_, new_n24488_, new_n24489_, new_n24490_,
    new_n24491_, new_n24492_, new_n24493_, new_n24494_, new_n24495_,
    new_n24496_, new_n24497_, new_n24498_, new_n24499_, new_n24500_,
    new_n24501_, new_n24502_, new_n24503_, new_n24504_, new_n24505_,
    new_n24506_, new_n24507_, new_n24508_, new_n24509_, new_n24510_,
    new_n24511_, new_n24512_, new_n24513_, new_n24514_, new_n24515_,
    new_n24516_, new_n24517_, new_n24518_, new_n24519_, new_n24520_,
    new_n24521_, new_n24522_, new_n24523_, new_n24524_, new_n24525_,
    new_n24526_, new_n24527_, new_n24528_, new_n24529_, new_n24530_,
    new_n24531_, new_n24532_, new_n24533_, new_n24534_, new_n24535_,
    new_n24536_, new_n24537_, new_n24538_, new_n24539_, new_n24540_,
    new_n24541_, new_n24542_, new_n24543_, new_n24544_, new_n24545_,
    new_n24546_, new_n24547_, new_n24548_, new_n24549_, new_n24550_,
    new_n24551_, new_n24552_, new_n24553_, new_n24554_, new_n24555_,
    new_n24556_, new_n24557_, new_n24558_, new_n24559_, new_n24560_,
    new_n24561_, new_n24562_, new_n24563_, new_n24564_, new_n24565_,
    new_n24566_, new_n24567_, new_n24568_, new_n24569_, new_n24570_,
    new_n24571_, new_n24572_, new_n24573_, new_n24574_, new_n24575_,
    new_n24576_, new_n24577_, new_n24578_, new_n24579_, new_n24580_,
    new_n24581_, new_n24582_, new_n24583_, new_n24584_, new_n24585_,
    new_n24586_, new_n24587_, new_n24588_, new_n24589_, new_n24590_,
    new_n24591_, new_n24592_, new_n24593_, new_n24594_, new_n24595_,
    new_n24596_, new_n24597_, new_n24598_, new_n24599_, new_n24600_,
    new_n24601_, new_n24602_, new_n24603_, new_n24604_, new_n24605_,
    new_n24606_, new_n24607_, new_n24608_, new_n24609_, new_n24610_,
    new_n24611_, new_n24612_, new_n24613_, new_n24614_, new_n24615_,
    new_n24616_, new_n24617_, new_n24618_, new_n24619_, new_n24620_,
    new_n24621_, new_n24622_, new_n24623_, new_n24624_, new_n24625_,
    new_n24626_, new_n24627_, new_n24628_, new_n24629_, new_n24630_,
    new_n24631_, new_n24632_, new_n24633_, new_n24634_, new_n24635_,
    new_n24636_, new_n24637_, new_n24638_, new_n24639_, new_n24640_,
    new_n24641_, new_n24642_, new_n24643_, new_n24644_, new_n24645_,
    new_n24646_, new_n24647_, new_n24648_, new_n24649_, new_n24650_,
    new_n24651_, new_n24652_, new_n24653_, new_n24654_, new_n24655_,
    new_n24656_, new_n24657_, new_n24658_, new_n24659_, new_n24660_,
    new_n24661_, new_n24662_, new_n24663_, new_n24664_, new_n24665_,
    new_n24666_, new_n24667_, new_n24668_, new_n24669_, new_n24670_,
    new_n24671_, new_n24672_, new_n24673_, new_n24674_, new_n24675_,
    new_n24676_, new_n24677_, new_n24678_, new_n24679_, new_n24680_,
    new_n24681_, new_n24682_, new_n24683_, new_n24684_, new_n24685_,
    new_n24686_, new_n24687_, new_n24688_, new_n24689_, new_n24690_,
    new_n24691_, new_n24692_, new_n24693_, new_n24694_, new_n24695_,
    new_n24696_, new_n24697_, new_n24698_, new_n24699_, new_n24700_,
    new_n24701_, new_n24702_, new_n24703_, new_n24704_, new_n24705_,
    new_n24706_, new_n24707_, new_n24708_, new_n24709_, new_n24710_,
    new_n24711_, new_n24712_, new_n24713_, new_n24714_, new_n24715_,
    new_n24716_, new_n24717_, new_n24718_, new_n24719_, new_n24720_,
    new_n24721_, new_n24722_, new_n24723_, new_n24724_, new_n24725_,
    new_n24726_, new_n24727_, new_n24728_, new_n24729_, new_n24730_,
    new_n24731_, new_n24732_, new_n24733_, new_n24734_, new_n24735_,
    new_n24736_, new_n24737_, new_n24738_, new_n24739_, new_n24740_,
    new_n24741_, new_n24742_, new_n24743_, new_n24744_, new_n24745_,
    new_n24746_, new_n24747_, new_n24748_, new_n24749_, new_n24750_,
    new_n24751_, new_n24752_, new_n24753_, new_n24754_, new_n24755_,
    new_n24756_, new_n24757_, new_n24758_, new_n24759_, new_n24760_,
    new_n24761_, new_n24762_, new_n24763_, new_n24764_, new_n24765_,
    new_n24766_, new_n24767_, new_n24768_, new_n24769_, new_n24770_,
    new_n24771_, new_n24772_, new_n24773_, new_n24774_, new_n24775_,
    new_n24776_, new_n24777_, new_n24778_, new_n24779_, new_n24780_,
    new_n24781_, new_n24782_, new_n24783_, new_n24784_, new_n24785_,
    new_n24786_, new_n24787_, new_n24788_, new_n24789_, new_n24790_,
    new_n24791_, new_n24792_, new_n24793_, new_n24794_, new_n24795_,
    new_n24796_, new_n24797_, new_n24798_, new_n24799_, new_n24800_,
    new_n24801_, new_n24802_, new_n24803_, new_n24804_, new_n24805_,
    new_n24806_, new_n24807_, new_n24808_, new_n24809_, new_n24810_,
    new_n24811_, new_n24812_, new_n24813_, new_n24814_, new_n24815_,
    new_n24816_, new_n24817_, new_n24818_, new_n24819_, new_n24820_,
    new_n24821_, new_n24822_, new_n24823_, new_n24824_, new_n24825_,
    new_n24826_, new_n24827_, new_n24828_, new_n24829_, new_n24830_,
    new_n24831_, new_n24832_, new_n24833_, new_n24834_, new_n24835_,
    new_n24836_, new_n24837_, new_n24838_, new_n24839_, new_n24840_,
    new_n24841_, new_n24842_, new_n24843_, new_n24844_, new_n24845_,
    new_n24846_, new_n24847_, new_n24848_, new_n24849_, new_n24850_,
    new_n24851_, new_n24852_, new_n24853_, new_n24854_, new_n24855_,
    new_n24856_, new_n24857_, new_n24858_, new_n24859_, new_n24860_,
    new_n24861_, new_n24862_, new_n24863_, new_n24864_, new_n24865_,
    new_n24866_, new_n24867_, new_n24868_, new_n24869_, new_n24870_,
    new_n24871_, new_n24872_, new_n24873_, new_n24874_, new_n24875_,
    new_n24876_, new_n24877_, new_n24878_, new_n24879_, new_n24880_,
    new_n24881_, new_n24882_, new_n24883_, new_n24884_, new_n24885_,
    new_n24886_, new_n24887_, new_n24888_, new_n24889_, new_n24890_,
    new_n24891_, new_n24892_, new_n24893_, new_n24894_, new_n24895_,
    new_n24896_, new_n24897_, new_n24898_, new_n24899_, new_n24900_,
    new_n24901_, new_n24902_, new_n24903_, new_n24904_, new_n24905_,
    new_n24906_, new_n24907_, new_n24908_, new_n24909_, new_n24910_,
    new_n24911_, new_n24912_, new_n24913_, new_n24914_, new_n24915_,
    new_n24916_, new_n24917_, new_n24918_, new_n24919_, new_n24920_,
    new_n24921_, new_n24922_, new_n24923_, new_n24924_, new_n24925_,
    new_n24926_, new_n24927_, new_n24928_, new_n24929_, new_n24930_,
    new_n24931_, new_n24932_, new_n24933_, new_n24934_, new_n24935_,
    new_n24936_, new_n24937_, new_n24938_, new_n24939_, new_n24940_,
    new_n24941_, new_n24942_, new_n24943_, new_n24944_, new_n24945_,
    new_n24946_, new_n24947_, new_n24948_, new_n24949_, new_n24950_,
    new_n24951_, new_n24952_, new_n24953_, new_n24954_, new_n24955_,
    new_n24956_, new_n24957_, new_n24958_, new_n24959_, new_n24960_,
    new_n24961_, new_n24962_, new_n24963_, new_n24964_, new_n24965_,
    new_n24966_, new_n24967_, new_n24968_, new_n24969_, new_n24970_,
    new_n24971_, new_n24972_, new_n24973_, new_n24974_, new_n24975_,
    new_n24976_, new_n24977_, new_n24978_, new_n24979_, new_n24980_,
    new_n24981_, new_n24982_, new_n24983_, new_n24984_, new_n24985_,
    new_n24986_, new_n24987_, new_n24988_, new_n24989_, new_n24990_,
    new_n24991_, new_n24992_, new_n24993_, new_n24994_, new_n24995_,
    new_n24996_, new_n24997_, new_n24998_, new_n24999_, new_n25000_,
    new_n25001_, new_n25002_, new_n25003_, new_n25004_, new_n25005_,
    new_n25006_, new_n25007_, new_n25008_, new_n25009_, new_n25010_,
    new_n25011_, new_n25012_, new_n25013_, new_n25014_, new_n25015_,
    new_n25016_, new_n25017_, new_n25018_, new_n25019_, new_n25020_,
    new_n25021_, new_n25022_, new_n25023_, new_n25024_, new_n25025_,
    new_n25026_, new_n25027_, new_n25028_, new_n25029_, new_n25030_,
    new_n25031_, new_n25032_, new_n25033_, new_n25034_, new_n25035_,
    new_n25036_, new_n25037_, new_n25038_, new_n25039_, new_n25040_,
    new_n25041_, new_n25042_, new_n25043_, new_n25044_, new_n25045_,
    new_n25046_, new_n25047_, new_n25048_, new_n25049_, new_n25050_,
    new_n25051_, new_n25052_, new_n25053_, new_n25054_, new_n25055_,
    new_n25056_, new_n25057_, new_n25058_, new_n25059_, new_n25060_,
    new_n25061_, new_n25062_, new_n25063_, new_n25064_, new_n25065_,
    new_n25066_, new_n25067_, new_n25068_, new_n25069_, new_n25070_,
    new_n25071_, new_n25072_, new_n25073_, new_n25074_, new_n25075_,
    new_n25076_, new_n25077_, new_n25078_, new_n25079_, new_n25080_,
    new_n25081_, new_n25082_, new_n25083_, new_n25084_, new_n25085_,
    new_n25086_, new_n25087_, new_n25088_, new_n25089_, new_n25090_,
    new_n25091_, new_n25092_, new_n25093_, new_n25094_, new_n25095_,
    new_n25096_, new_n25097_, new_n25098_, new_n25099_, new_n25100_,
    new_n25101_, new_n25102_, new_n25103_, new_n25104_, new_n25105_,
    new_n25106_, new_n25107_, new_n25108_, new_n25109_, new_n25110_,
    new_n25111_, new_n25112_, new_n25113_, new_n25114_, new_n25115_,
    new_n25116_, new_n25117_, new_n25118_, new_n25119_, new_n25120_,
    new_n25121_, new_n25122_, new_n25123_, new_n25124_, new_n25125_,
    new_n25126_, new_n25127_, new_n25128_, new_n25129_, new_n25130_,
    new_n25131_, new_n25132_, new_n25133_, new_n25134_, new_n25135_,
    new_n25136_, new_n25137_, new_n25138_, new_n25139_, new_n25140_,
    new_n25141_, new_n25142_, new_n25143_, new_n25144_, new_n25145_,
    new_n25146_, new_n25147_, new_n25148_, new_n25149_, new_n25150_,
    new_n25151_, new_n25152_, new_n25153_, new_n25154_, new_n25155_,
    new_n25156_, new_n25157_, new_n25158_, new_n25159_, new_n25160_,
    new_n25161_, new_n25162_, new_n25163_, new_n25164_, new_n25165_,
    new_n25166_, new_n25167_, new_n25168_, new_n25169_, new_n25170_,
    new_n25171_, new_n25172_, new_n25173_, new_n25174_, new_n25175_,
    new_n25176_, new_n25177_, new_n25178_, new_n25179_, new_n25180_,
    new_n25181_, new_n25182_, new_n25183_, new_n25184_, new_n25185_,
    new_n25186_, new_n25187_, new_n25188_, new_n25189_, new_n25190_,
    new_n25191_, new_n25192_, new_n25193_, new_n25194_, new_n25195_,
    new_n25196_, new_n25197_, new_n25198_, new_n25199_, new_n25200_,
    new_n25201_, new_n25202_, new_n25203_, new_n25204_, new_n25205_,
    new_n25206_, new_n25207_, new_n25208_, new_n25209_, new_n25210_,
    new_n25211_, new_n25212_, new_n25213_, new_n25214_, new_n25215_,
    new_n25216_, new_n25217_, new_n25218_, new_n25219_, new_n25220_,
    new_n25221_, new_n25222_, new_n25223_, new_n25224_, new_n25225_,
    new_n25226_, new_n25227_, new_n25228_, new_n25229_, new_n25230_,
    new_n25231_, new_n25232_, new_n25233_, new_n25234_, new_n25235_,
    new_n25236_, new_n25237_, new_n25238_, new_n25239_, new_n25240_,
    new_n25241_, new_n25242_, new_n25243_, new_n25244_, new_n25245_,
    new_n25246_, new_n25247_, new_n25248_, new_n25249_, new_n25250_,
    new_n25251_, new_n25252_, new_n25253_, new_n25254_, new_n25255_,
    new_n25256_, new_n25257_, new_n25258_, new_n25259_, new_n25260_,
    new_n25261_, new_n25262_, new_n25263_, new_n25264_, new_n25265_,
    new_n25266_, new_n25267_, new_n25268_, new_n25269_, new_n25270_,
    new_n25271_, new_n25272_, new_n25273_, new_n25274_, new_n25275_,
    new_n25276_, new_n25277_, new_n25278_, new_n25279_, new_n25280_,
    new_n25281_, new_n25282_, new_n25283_, new_n25284_, new_n25285_,
    new_n25286_, new_n25287_, new_n25288_, new_n25289_, new_n25290_,
    new_n25291_, new_n25292_, new_n25293_, new_n25294_, new_n25295_,
    new_n25296_, new_n25297_, new_n25298_, new_n25299_, new_n25300_,
    new_n25301_, new_n25302_, new_n25303_, new_n25304_, new_n25305_,
    new_n25306_, new_n25307_, new_n25308_, new_n25309_, new_n25310_,
    new_n25311_, new_n25312_, new_n25313_, new_n25314_, new_n25315_,
    new_n25316_, new_n25317_, new_n25318_, new_n25319_, new_n25320_,
    new_n25321_, new_n25322_, new_n25323_, new_n25324_, new_n25325_,
    new_n25326_, new_n25327_, new_n25328_, new_n25329_, new_n25330_,
    new_n25331_, new_n25332_, new_n25333_, new_n25334_, new_n25335_,
    new_n25336_, new_n25337_, new_n25338_, new_n25339_, new_n25340_,
    new_n25341_, new_n25342_, new_n25343_, new_n25344_, new_n25345_,
    new_n25346_, new_n25347_, new_n25348_, new_n25349_, new_n25350_,
    new_n25351_, new_n25352_, new_n25353_, new_n25354_, new_n25355_,
    new_n25356_, new_n25357_, new_n25358_, new_n25359_, new_n25360_,
    new_n25361_, new_n25362_, new_n25363_, new_n25364_, new_n25365_,
    new_n25366_, new_n25367_, new_n25368_, new_n25369_, new_n25370_,
    new_n25371_, new_n25372_, new_n25373_, new_n25374_, new_n25375_,
    new_n25376_, new_n25377_, new_n25378_, new_n25379_, new_n25380_,
    new_n25381_, new_n25382_, new_n25383_, new_n25384_, new_n25385_,
    new_n25386_, new_n25387_, new_n25388_, new_n25389_, new_n25390_,
    new_n25391_, new_n25392_, new_n25393_, new_n25394_, new_n25395_,
    new_n25396_, new_n25397_, new_n25398_, new_n25399_, new_n25400_,
    new_n25401_, new_n25402_, new_n25403_, new_n25404_, new_n25405_,
    new_n25406_, new_n25407_, new_n25408_, new_n25409_, new_n25410_,
    new_n25411_, new_n25412_, new_n25413_, new_n25414_, new_n25415_,
    new_n25416_, new_n25417_, new_n25418_, new_n25419_, new_n25420_,
    new_n25421_, new_n25422_, new_n25423_, new_n25424_, new_n25425_,
    new_n25426_, new_n25427_, new_n25428_, new_n25429_, new_n25430_,
    new_n25431_, new_n25432_, new_n25433_, new_n25434_, new_n25435_,
    new_n25436_, new_n25437_, new_n25438_, new_n25439_, new_n25440_,
    new_n25441_, new_n25442_, new_n25443_, new_n25444_, new_n25445_,
    new_n25446_, new_n25447_, new_n25448_, new_n25449_, new_n25450_,
    new_n25451_, new_n25452_, new_n25453_, new_n25454_, new_n25455_,
    new_n25456_, new_n25457_, new_n25458_, new_n25459_, new_n25460_,
    new_n25461_, new_n25462_, new_n25463_, new_n25464_, new_n25465_,
    new_n25466_, new_n25467_, new_n25468_, new_n25469_, new_n25470_,
    new_n25471_, new_n25472_, new_n25473_, new_n25474_, new_n25475_,
    new_n25476_, new_n25477_, new_n25478_, new_n25479_, new_n25480_,
    new_n25481_, new_n25482_, new_n25483_, new_n25484_, new_n25485_,
    new_n25486_, new_n25487_, new_n25488_, new_n25489_, new_n25490_,
    new_n25491_, new_n25492_, new_n25493_, new_n25494_, new_n25495_,
    new_n25496_, new_n25497_, new_n25498_, new_n25499_, new_n25500_,
    new_n25501_, new_n25502_, new_n25503_, new_n25504_, new_n25505_,
    new_n25506_, new_n25507_, new_n25508_, new_n25509_, new_n25510_,
    new_n25511_, new_n25512_, new_n25513_, new_n25514_, new_n25515_,
    new_n25516_, new_n25517_, new_n25518_, new_n25519_, new_n25520_,
    new_n25521_, new_n25522_, new_n25523_, new_n25524_, new_n25525_,
    new_n25526_, new_n25527_, new_n25528_, new_n25529_, new_n25530_,
    new_n25531_, new_n25532_, new_n25533_, new_n25534_, new_n25535_,
    new_n25536_, new_n25537_, new_n25538_, new_n25539_, new_n25540_,
    new_n25541_, new_n25542_, new_n25543_, new_n25544_, new_n25545_,
    new_n25546_, new_n25547_, new_n25548_, new_n25549_, new_n25550_,
    new_n25551_, new_n25552_, new_n25553_, new_n25554_, new_n25555_,
    new_n25556_, new_n25557_, new_n25558_, new_n25559_, new_n25560_,
    new_n25561_, new_n25562_, new_n25563_, new_n25564_, new_n25565_,
    new_n25566_, new_n25567_, new_n25568_, new_n25569_, new_n25570_,
    new_n25571_, new_n25572_, new_n25573_, new_n25574_, new_n25575_,
    new_n25576_, new_n25577_, new_n25578_, new_n25579_, new_n25580_,
    new_n25581_, new_n25582_, new_n25583_, new_n25584_, new_n25585_,
    new_n25586_, new_n25587_, new_n25588_, new_n25589_, new_n25590_,
    new_n25591_, new_n25592_, new_n25593_, new_n25594_, new_n25595_,
    new_n25596_, new_n25597_, new_n25598_, new_n25599_, new_n25600_,
    new_n25601_, new_n25602_, new_n25603_, new_n25604_, new_n25605_,
    new_n25606_, new_n25607_, new_n25608_, new_n25609_, new_n25610_,
    new_n25611_, new_n25612_, new_n25613_, new_n25614_, new_n25615_,
    new_n25616_, new_n25617_, new_n25618_, new_n25619_, new_n25620_,
    new_n25621_, new_n25622_, new_n25623_, new_n25624_, new_n25625_,
    new_n25626_, new_n25627_, new_n25628_, new_n25629_, new_n25630_,
    new_n25631_, new_n25632_, new_n25633_, new_n25634_, new_n25635_,
    new_n25636_, new_n25637_, new_n25638_, new_n25639_, new_n25640_,
    new_n25641_, new_n25642_, new_n25643_, new_n25644_, new_n25645_,
    new_n25646_, new_n25647_, new_n25648_, new_n25649_, new_n25650_,
    new_n25651_, new_n25652_, new_n25653_, new_n25654_, new_n25655_,
    new_n25656_, new_n25657_, new_n25658_, new_n25659_, new_n25660_,
    new_n25661_, new_n25662_, new_n25663_, new_n25664_, new_n25665_,
    new_n25666_, new_n25667_, new_n25668_, new_n25669_, new_n25670_,
    new_n25671_, new_n25672_, new_n25673_, new_n25674_, new_n25675_,
    new_n25676_, new_n25677_, new_n25678_, new_n25679_, new_n25680_,
    new_n25681_, new_n25682_, new_n25683_, new_n25684_, new_n25685_,
    new_n25686_, new_n25687_, new_n25688_, new_n25689_, new_n25690_,
    new_n25691_, new_n25692_, new_n25693_, new_n25694_, new_n25695_,
    new_n25696_, new_n25697_, new_n25698_, new_n25699_, new_n25700_,
    new_n25701_, new_n25702_, new_n25703_, new_n25704_, new_n25705_,
    new_n25706_, new_n25707_, new_n25708_, new_n25709_, new_n25710_,
    new_n25711_, new_n25712_, new_n25713_, new_n25714_, new_n25715_,
    new_n25716_, new_n25717_, new_n25718_, new_n25719_, new_n25720_,
    new_n25721_, new_n25722_, new_n25723_, new_n25724_, new_n25725_,
    new_n25726_, new_n25727_, new_n25728_, new_n25729_, new_n25730_,
    new_n25731_, new_n25732_, new_n25733_, new_n25734_, new_n25735_,
    new_n25736_, new_n25737_, new_n25738_, new_n25739_, new_n25740_,
    new_n25741_, new_n25742_, new_n25743_, new_n25744_, new_n25745_,
    new_n25746_, new_n25747_, new_n25748_, new_n25749_, new_n25750_,
    new_n25751_, new_n25752_, new_n25753_, new_n25754_, new_n25755_,
    new_n25756_, new_n25757_, new_n25758_, new_n25759_, new_n25760_,
    new_n25761_, new_n25762_, new_n25763_, new_n25764_, new_n25765_,
    new_n25766_, new_n25767_, new_n25768_, new_n25769_, new_n25770_,
    new_n25771_, new_n25772_, new_n25773_, new_n25774_, new_n25775_,
    new_n25776_, new_n25777_, new_n25778_, new_n25779_, new_n25780_,
    new_n25781_, new_n25782_, new_n25783_, new_n25784_, new_n25785_,
    new_n25786_, new_n25787_, new_n25788_, new_n25789_, new_n25790_,
    new_n25791_, new_n25792_, new_n25793_, new_n25794_, new_n25795_,
    new_n25796_, new_n25797_, new_n25798_, new_n25799_, new_n25800_,
    new_n25801_, new_n25802_, new_n25803_, new_n25804_, new_n25805_,
    new_n25806_, new_n25807_, new_n25808_, new_n25809_, new_n25810_,
    new_n25811_, new_n25812_, new_n25813_, new_n25814_, new_n25815_,
    new_n25816_, new_n25817_, new_n25818_, new_n25819_, new_n25820_,
    new_n25821_, new_n25822_, new_n25823_, new_n25824_, new_n25825_,
    new_n25826_, new_n25827_, new_n25828_, new_n25829_, new_n25830_,
    new_n25831_, new_n25832_, new_n25833_, new_n25834_, new_n25835_,
    new_n25836_, new_n25837_, new_n25838_, new_n25839_, new_n25840_,
    new_n25841_, new_n25842_, new_n25843_, new_n25844_, new_n25845_,
    new_n25846_, new_n25847_, new_n25848_, new_n25849_, new_n25850_,
    new_n25851_, new_n25852_, new_n25853_, new_n25854_, new_n25855_,
    new_n25856_, new_n25857_, new_n25858_, new_n25859_, new_n25860_,
    new_n25861_, new_n25862_, new_n25863_, new_n25864_, new_n25865_,
    new_n25866_, new_n25867_, new_n25868_, new_n25869_, new_n25870_,
    new_n25871_, new_n25872_, new_n25873_, new_n25874_, new_n25875_,
    new_n25876_, new_n25877_, new_n25878_, new_n25879_, new_n25880_,
    new_n25881_, new_n25882_, new_n25883_, new_n25884_, new_n25885_,
    new_n25886_, new_n25887_, new_n25888_, new_n25889_, new_n25890_,
    new_n25891_, new_n25892_, new_n25893_, new_n25894_, new_n25895_,
    new_n25896_, new_n25897_, new_n25898_, new_n25899_, new_n25900_,
    new_n25901_, new_n25902_, new_n25903_, new_n25904_, new_n25905_,
    new_n25906_, new_n25907_, new_n25908_, new_n25909_, new_n25910_,
    new_n25911_, new_n25912_, new_n25913_, new_n25914_, new_n25915_,
    new_n25916_, new_n25917_, new_n25918_, new_n25919_, new_n25920_,
    new_n25921_, new_n25922_, new_n25923_, new_n25924_, new_n25925_,
    new_n25926_, new_n25927_, new_n25928_, new_n25929_, new_n25930_,
    new_n25931_, new_n25932_, new_n25933_, new_n25934_, new_n25935_,
    new_n25936_, new_n25937_, new_n25938_, new_n25939_, new_n25940_,
    new_n25941_, new_n25942_, new_n25943_, new_n25944_, new_n25945_,
    new_n25946_, new_n25947_, new_n25948_, new_n25949_, new_n25950_,
    new_n25951_, new_n25952_, new_n25953_, new_n25954_, new_n25955_,
    new_n25956_, new_n25957_, new_n25958_, new_n25959_, new_n25960_,
    new_n25961_, new_n25962_, new_n25963_, new_n25964_, new_n25965_,
    new_n25966_, new_n25967_, new_n25968_, new_n25969_, new_n25970_,
    new_n25971_, new_n25972_, new_n25973_, new_n25974_, new_n25975_,
    new_n25976_, new_n25977_, new_n25978_, new_n25979_, new_n25980_,
    new_n25981_, new_n25982_, new_n25983_, new_n25984_, new_n25985_,
    new_n25986_, new_n25987_, new_n25988_, new_n25989_, new_n25990_,
    new_n25991_, new_n25992_, new_n25993_, new_n25994_, new_n25995_,
    new_n25996_, new_n25997_, new_n25998_, new_n25999_, new_n26000_,
    new_n26001_, new_n26002_, new_n26003_, new_n26004_, new_n26005_,
    new_n26006_, new_n26007_, new_n26008_, new_n26009_, new_n26010_,
    new_n26011_, new_n26012_, new_n26013_, new_n26014_, new_n26015_,
    new_n26016_, new_n26017_, new_n26018_, new_n26019_, new_n26020_,
    new_n26021_, new_n26022_, new_n26023_, new_n26024_, new_n26025_,
    new_n26026_, new_n26027_, new_n26028_, new_n26029_, new_n26030_,
    new_n26031_, new_n26032_, new_n26033_, new_n26034_, new_n26035_,
    new_n26036_, new_n26037_, new_n26038_, new_n26039_, new_n26040_,
    new_n26041_, new_n26042_, new_n26043_, new_n26044_, new_n26045_,
    new_n26046_, new_n26047_, new_n26048_, new_n26049_, new_n26050_,
    new_n26051_, new_n26052_, new_n26053_, new_n26054_, new_n26055_,
    new_n26056_, new_n26057_, new_n26058_, new_n26059_, new_n26060_,
    new_n26061_, new_n26062_, new_n26063_, new_n26064_, new_n26065_,
    new_n26066_, new_n26067_, new_n26068_, new_n26069_, new_n26070_,
    new_n26071_, new_n26072_, new_n26073_, new_n26074_, new_n26075_,
    new_n26076_, new_n26077_, new_n26078_, new_n26079_, new_n26080_,
    new_n26081_, new_n26082_, new_n26083_, new_n26084_, new_n26085_,
    new_n26086_, new_n26087_, new_n26088_, new_n26089_, new_n26090_,
    new_n26091_, new_n26092_, new_n26093_, new_n26094_, new_n26095_,
    new_n26096_, new_n26097_, new_n26098_, new_n26099_, new_n26100_,
    new_n26101_, new_n26102_, new_n26103_, new_n26104_, new_n26105_,
    new_n26106_, new_n26107_, new_n26108_, new_n26109_, new_n26110_,
    new_n26111_, new_n26112_, new_n26113_, new_n26114_, new_n26115_,
    new_n26116_, new_n26117_, new_n26118_, new_n26119_, new_n26120_,
    new_n26121_, new_n26122_, new_n26123_, new_n26124_, new_n26125_,
    new_n26126_, new_n26127_, new_n26128_, new_n26129_, new_n26130_,
    new_n26131_, new_n26132_, new_n26133_, new_n26134_, new_n26135_,
    new_n26136_, new_n26137_, new_n26138_, new_n26139_, new_n26140_,
    new_n26141_, new_n26142_, new_n26143_, new_n26144_, new_n26145_,
    new_n26146_, new_n26147_, new_n26148_, new_n26149_, new_n26150_,
    new_n26151_, new_n26152_, new_n26153_, new_n26154_, new_n26155_,
    new_n26156_, new_n26157_, new_n26158_, new_n26159_, new_n26160_,
    new_n26161_, new_n26162_, new_n26163_, new_n26164_, new_n26165_,
    new_n26166_, new_n26167_, new_n26168_, new_n26169_, new_n26170_,
    new_n26171_, new_n26172_, new_n26173_, new_n26174_, new_n26175_,
    new_n26176_, new_n26177_, new_n26178_, new_n26179_, new_n26180_,
    new_n26181_, new_n26182_, new_n26183_, new_n26184_, new_n26185_,
    new_n26186_, new_n26187_, new_n26188_, new_n26189_, new_n26190_,
    new_n26191_, new_n26192_, new_n26193_, new_n26194_, new_n26195_,
    new_n26196_, new_n26197_, new_n26198_, new_n26199_, new_n26200_,
    new_n26201_, new_n26202_, new_n26203_, new_n26204_, new_n26205_,
    new_n26206_, new_n26207_, new_n26208_, new_n26209_, new_n26210_,
    new_n26211_, new_n26212_, new_n26213_, new_n26214_, new_n26215_,
    new_n26216_, new_n26217_, new_n26218_, new_n26219_, new_n26220_,
    new_n26221_, new_n26222_, new_n26223_, new_n26224_, new_n26225_,
    new_n26226_, new_n26227_, new_n26228_, new_n26229_, new_n26230_,
    new_n26231_, new_n26232_, new_n26233_, new_n26234_, new_n26235_,
    new_n26236_, new_n26237_, new_n26238_, new_n26239_, new_n26240_,
    new_n26241_, new_n26242_, new_n26243_, new_n26244_, new_n26245_,
    new_n26246_, new_n26247_, new_n26248_, new_n26249_, new_n26250_,
    new_n26251_, new_n26252_, new_n26253_, new_n26254_, new_n26255_,
    new_n26256_, new_n26257_, new_n26258_, new_n26259_, new_n26260_,
    new_n26261_, new_n26262_, new_n26263_, new_n26264_, new_n26265_,
    new_n26266_, new_n26267_, new_n26268_, new_n26269_, new_n26270_,
    new_n26271_, new_n26272_, new_n26273_, new_n26274_, new_n26275_,
    new_n26276_, new_n26277_, new_n26278_, new_n26279_, new_n26280_,
    new_n26281_, new_n26282_, new_n26283_, new_n26284_, new_n26285_,
    new_n26286_, new_n26287_, new_n26288_, new_n26289_, new_n26290_,
    new_n26291_, new_n26292_, new_n26293_, new_n26294_, new_n26295_,
    new_n26296_, new_n26297_, new_n26298_, new_n26299_, new_n26300_,
    new_n26301_, new_n26302_, new_n26303_, new_n26304_, new_n26305_,
    new_n26306_, new_n26307_, new_n26308_, new_n26309_, new_n26310_,
    new_n26311_, new_n26312_, new_n26313_, new_n26314_, new_n26315_,
    new_n26316_, new_n26317_, new_n26318_, new_n26319_, new_n26320_,
    new_n26321_, new_n26322_, new_n26323_, new_n26324_, new_n26325_,
    new_n26326_, new_n26327_, new_n26328_, new_n26329_, new_n26330_,
    new_n26331_, new_n26332_, new_n26333_, new_n26334_, new_n26335_,
    new_n26336_, new_n26337_, new_n26338_, new_n26339_, new_n26340_,
    new_n26341_, new_n26342_, new_n26343_, new_n26344_, new_n26345_,
    new_n26346_, new_n26347_, new_n26348_, new_n26349_, new_n26350_,
    new_n26351_, new_n26352_, new_n26353_, new_n26354_, new_n26355_,
    new_n26356_, new_n26357_, new_n26358_, new_n26359_, new_n26360_,
    new_n26361_, new_n26362_, new_n26363_, new_n26364_, new_n26365_,
    new_n26366_, new_n26367_, new_n26368_, new_n26369_, new_n26370_,
    new_n26371_, new_n26372_, new_n26373_, new_n26374_, new_n26375_,
    new_n26376_, new_n26377_, new_n26378_, new_n26379_, new_n26380_,
    new_n26381_, new_n26382_, new_n26383_, new_n26384_, new_n26385_,
    new_n26386_, new_n26387_, new_n26388_, new_n26389_, new_n26390_,
    new_n26391_, new_n26392_, new_n26393_, new_n26394_, new_n26395_,
    new_n26396_, new_n26397_, new_n26398_, new_n26399_, new_n26400_,
    new_n26401_, new_n26402_, new_n26403_, new_n26404_, new_n26405_,
    new_n26406_, new_n26407_, new_n26408_, new_n26409_, new_n26410_,
    new_n26411_, new_n26412_, new_n26413_, new_n26414_, new_n26415_,
    new_n26416_, new_n26417_, new_n26418_, new_n26419_, new_n26420_,
    new_n26421_, new_n26422_, new_n26423_, new_n26424_, new_n26425_,
    new_n26426_, new_n26427_, new_n26428_, new_n26429_, new_n26430_,
    new_n26431_, new_n26432_, new_n26433_, new_n26434_, new_n26435_,
    new_n26436_, new_n26437_, new_n26438_, new_n26439_, new_n26440_,
    new_n26441_, new_n26442_, new_n26443_, new_n26444_, new_n26445_,
    new_n26446_, new_n26447_, new_n26448_, new_n26449_, new_n26450_,
    new_n26451_, new_n26452_, new_n26453_, new_n26454_, new_n26455_,
    new_n26456_, new_n26457_, new_n26458_, new_n26459_, new_n26460_,
    new_n26461_, new_n26462_, new_n26463_, new_n26464_, new_n26465_,
    new_n26466_, new_n26467_, new_n26468_, new_n26469_, new_n26470_,
    new_n26471_, new_n26472_, new_n26473_, new_n26474_, new_n26475_,
    new_n26476_, new_n26477_, new_n26478_, new_n26479_, new_n26480_,
    new_n26481_, new_n26482_, new_n26483_, new_n26484_, new_n26485_,
    new_n26486_, new_n26487_, new_n26488_, new_n26489_, new_n26490_,
    new_n26491_, new_n26492_, new_n26493_, new_n26494_, new_n26495_,
    new_n26496_, new_n26497_, new_n26498_, new_n26499_, new_n26500_,
    new_n26501_, new_n26502_, new_n26503_, new_n26504_, new_n26505_,
    new_n26506_, new_n26507_, new_n26508_, new_n26509_, new_n26510_,
    new_n26511_, new_n26512_, new_n26513_, new_n26514_, new_n26515_,
    new_n26516_, new_n26517_, new_n26518_, new_n26519_, new_n26520_,
    new_n26521_, new_n26522_, new_n26523_, new_n26524_, new_n26525_,
    new_n26526_, new_n26527_, new_n26528_, new_n26529_, new_n26530_,
    new_n26531_, new_n26532_, new_n26533_, new_n26534_, new_n26535_,
    new_n26536_, new_n26537_, new_n26538_, new_n26539_, new_n26540_,
    new_n26541_, new_n26542_, new_n26543_, new_n26544_, new_n26545_,
    new_n26546_, new_n26547_, new_n26548_, new_n26549_, new_n26550_,
    new_n26551_, new_n26552_, new_n26553_, new_n26554_, new_n26555_,
    new_n26556_, new_n26557_, new_n26558_, new_n26559_, new_n26560_,
    new_n26561_, new_n26562_, new_n26563_, new_n26564_, new_n26565_,
    new_n26566_, new_n26567_, new_n26568_, new_n26569_, new_n26570_,
    new_n26571_, new_n26572_, new_n26573_, new_n26574_, new_n26575_,
    new_n26576_, new_n26577_, new_n26578_, new_n26579_, new_n26580_,
    new_n26581_, new_n26582_, new_n26583_, new_n26584_, new_n26585_,
    new_n26586_, new_n26587_, new_n26588_, new_n26589_, new_n26590_,
    new_n26591_, new_n26592_, new_n26593_, new_n26594_, new_n26595_,
    new_n26596_, new_n26597_, new_n26598_, new_n26599_, new_n26600_,
    new_n26601_, new_n26602_, new_n26603_, new_n26604_, new_n26605_,
    new_n26606_, new_n26607_, new_n26608_, new_n26609_, new_n26610_,
    new_n26611_, new_n26612_, new_n26613_, new_n26614_, new_n26615_,
    new_n26616_, new_n26617_, new_n26618_, new_n26619_, new_n26620_,
    new_n26621_, new_n26622_, new_n26623_, new_n26624_, new_n26625_,
    new_n26626_, new_n26627_, new_n26628_, new_n26629_, new_n26630_,
    new_n26631_, new_n26632_, new_n26633_, new_n26634_, new_n26635_,
    new_n26636_, new_n26637_, new_n26638_, new_n26639_, new_n26640_,
    new_n26641_, new_n26642_, new_n26643_, new_n26644_, new_n26645_,
    new_n26646_, new_n26647_, new_n26648_, new_n26649_, new_n26650_,
    new_n26651_, new_n26652_, new_n26653_, new_n26654_, new_n26655_,
    new_n26656_, new_n26657_, new_n26658_, new_n26659_, new_n26660_,
    new_n26661_, new_n26662_, new_n26663_, new_n26664_, new_n26665_,
    new_n26666_, new_n26667_, new_n26668_, new_n26669_, new_n26670_,
    new_n26671_, new_n26672_, new_n26673_, new_n26674_, new_n26675_,
    new_n26676_, new_n26677_, new_n26678_, new_n26679_, new_n26680_,
    new_n26681_, new_n26682_, new_n26683_, new_n26684_, new_n26685_,
    new_n26686_, new_n26687_, new_n26688_, new_n26689_, new_n26690_,
    new_n26691_, new_n26692_, new_n26693_, new_n26694_, new_n26695_,
    new_n26696_, new_n26697_, new_n26698_, new_n26699_, new_n26700_,
    new_n26701_, new_n26702_, new_n26703_, new_n26704_, new_n26705_,
    new_n26706_, new_n26707_, new_n26708_, new_n26709_, new_n26710_,
    new_n26711_, new_n26712_, new_n26713_, new_n26714_, new_n26715_,
    new_n26716_, new_n26717_, new_n26718_, new_n26719_, new_n26720_,
    new_n26721_, new_n26722_, new_n26723_, new_n26724_, new_n26725_,
    new_n26726_, new_n26727_, new_n26728_, new_n26729_, new_n26730_,
    new_n26731_, new_n26732_, new_n26733_, new_n26734_, new_n26735_,
    new_n26736_, new_n26737_, new_n26738_, new_n26739_, new_n26740_,
    new_n26741_, new_n26742_, new_n26743_, new_n26744_, new_n26745_,
    new_n26746_, new_n26747_, new_n26748_, new_n26749_, new_n26750_,
    new_n26751_, new_n26752_, new_n26753_, new_n26754_, new_n26755_,
    new_n26756_, new_n26757_, new_n26758_, new_n26759_, new_n26760_,
    new_n26761_, new_n26762_, new_n26763_, new_n26764_, new_n26765_,
    new_n26766_, new_n26767_, new_n26768_, new_n26769_, new_n26770_,
    new_n26771_, new_n26772_, new_n26773_, new_n26774_, new_n26775_,
    new_n26776_, new_n26777_, new_n26778_, new_n26779_, new_n26780_,
    new_n26781_, new_n26782_, new_n26783_, new_n26784_, new_n26785_,
    new_n26786_, new_n26787_, new_n26788_, new_n26789_, new_n26790_,
    new_n26791_, new_n26792_, new_n26793_, new_n26794_, new_n26795_,
    new_n26796_, new_n26797_, new_n26798_, new_n26799_, new_n26800_,
    new_n26801_, new_n26802_, new_n26803_, new_n26804_, new_n26805_,
    new_n26806_, new_n26807_, new_n26808_, new_n26809_, new_n26810_,
    new_n26811_, new_n26812_, new_n26813_, new_n26814_, new_n26815_,
    new_n26816_, new_n26817_, new_n26818_, new_n26819_, new_n26820_,
    new_n26821_, new_n26822_, new_n26823_, new_n26824_, new_n26825_,
    new_n26826_, new_n26827_, new_n26828_, new_n26829_, new_n26830_,
    new_n26831_, new_n26832_, new_n26833_, new_n26834_, new_n26835_,
    new_n26836_, new_n26837_, new_n26838_, new_n26839_, new_n26840_,
    new_n26841_, new_n26842_, new_n26843_, new_n26844_, new_n26845_,
    new_n26846_, new_n26847_, new_n26848_, new_n26849_, new_n26850_,
    new_n26851_, new_n26852_, new_n26853_, new_n26854_, new_n26855_,
    new_n26856_, new_n26857_, new_n26858_, new_n26859_, new_n26860_,
    new_n26861_, new_n26862_, new_n26863_, new_n26864_, new_n26865_,
    new_n26866_, new_n26867_, new_n26868_, new_n26869_, new_n26870_,
    new_n26871_, new_n26872_, new_n26873_, new_n26874_, new_n26875_,
    new_n26876_, new_n26877_, new_n26878_, new_n26879_, new_n26880_,
    new_n26881_, new_n26882_, new_n26883_, new_n26884_, new_n26885_,
    new_n26886_, new_n26887_, new_n26888_, new_n26889_, new_n26890_,
    new_n26891_, new_n26892_, new_n26893_, new_n26894_, new_n26895_,
    new_n26896_, new_n26897_, new_n26898_, new_n26899_, new_n26900_,
    new_n26901_, new_n26902_, new_n26903_, new_n26904_, new_n26905_,
    new_n26906_, new_n26907_, new_n26908_, new_n26909_, new_n26910_,
    new_n26911_, new_n26912_, new_n26913_, new_n26914_, new_n26915_,
    new_n26916_, new_n26917_, new_n26918_, new_n26919_, new_n26920_,
    new_n26921_, new_n26922_, new_n26923_, new_n26924_, new_n26925_,
    new_n26926_, new_n26927_, new_n26928_, new_n26929_, new_n26930_,
    new_n26931_, new_n26932_, new_n26933_, new_n26934_, new_n26935_,
    new_n26936_, new_n26937_, new_n26938_, new_n26939_, new_n26940_,
    new_n26941_, new_n26942_, new_n26943_, new_n26944_, new_n26945_,
    new_n26946_, new_n26947_, new_n26948_, new_n26949_, new_n26950_,
    new_n26951_, new_n26952_, new_n26953_, new_n26954_, new_n26955_,
    new_n26956_, new_n26957_, new_n26958_, new_n26959_, new_n26960_,
    new_n26961_, new_n26962_, new_n26963_, new_n26964_, new_n26965_,
    new_n26966_, new_n26967_, new_n26968_, new_n26969_, new_n26970_,
    new_n26971_, new_n26972_, new_n26973_, new_n26974_, new_n26975_,
    new_n26976_, new_n26977_, new_n26978_, new_n26979_, new_n26980_,
    new_n26981_, new_n26982_, new_n26983_, new_n26984_, new_n26985_,
    new_n26986_, new_n26987_, new_n26988_, new_n26989_, new_n26990_,
    new_n26991_, new_n26992_, new_n26993_, new_n26994_, new_n26995_,
    new_n26996_, new_n26997_, new_n26998_, new_n26999_, new_n27000_,
    new_n27001_, new_n27002_, new_n27003_, new_n27004_, new_n27005_,
    new_n27006_, new_n27007_, new_n27008_, new_n27009_, new_n27010_,
    new_n27011_, new_n27012_, new_n27013_, new_n27014_, new_n27015_,
    new_n27016_, new_n27017_, new_n27018_, new_n27019_, new_n27020_,
    new_n27021_, new_n27022_, new_n27023_, new_n27024_, new_n27025_,
    new_n27026_, new_n27027_, new_n27028_, new_n27029_, new_n27030_,
    new_n27031_, new_n27032_, new_n27033_, new_n27034_, new_n27035_,
    new_n27036_, new_n27037_, new_n27038_, new_n27039_, new_n27040_,
    new_n27041_, new_n27042_, new_n27043_, new_n27044_, new_n27045_,
    new_n27046_, new_n27047_, new_n27048_, new_n27049_, new_n27050_,
    new_n27051_, new_n27052_, new_n27053_, new_n27054_, new_n27055_,
    new_n27056_, new_n27057_, new_n27058_, new_n27059_, new_n27060_,
    new_n27061_, new_n27062_, new_n27063_, new_n27064_, new_n27065_,
    new_n27066_, new_n27067_, new_n27068_, new_n27069_, new_n27070_,
    new_n27071_, new_n27072_, new_n27073_, new_n27074_, new_n27075_,
    new_n27076_, new_n27077_, new_n27078_, new_n27079_, new_n27080_,
    new_n27081_, new_n27082_, new_n27083_, new_n27084_, new_n27085_,
    new_n27086_, new_n27087_, new_n27088_, new_n27089_, new_n27090_,
    new_n27091_, new_n27092_, new_n27093_, new_n27094_, new_n27095_,
    new_n27096_, new_n27097_, new_n27098_, new_n27099_, new_n27100_,
    new_n27101_, new_n27102_, new_n27103_, new_n27104_, new_n27105_,
    new_n27106_, new_n27107_, new_n27108_, new_n27109_, new_n27110_,
    new_n27111_, new_n27112_, new_n27113_, new_n27114_, new_n27115_,
    new_n27116_, new_n27117_, new_n27118_, new_n27119_, new_n27120_,
    new_n27121_, new_n27122_, new_n27123_, new_n27124_, new_n27125_,
    new_n27126_, new_n27127_, new_n27128_, new_n27129_, new_n27130_,
    new_n27131_, new_n27132_, new_n27133_, new_n27134_, new_n27135_,
    new_n27136_, new_n27137_, new_n27138_, new_n27139_, new_n27140_,
    new_n27141_, new_n27142_, new_n27143_, new_n27144_, new_n27145_,
    new_n27146_, new_n27147_, new_n27148_, new_n27149_, new_n27150_,
    new_n27151_, new_n27152_, new_n27153_, new_n27154_, new_n27155_,
    new_n27156_, new_n27157_, new_n27158_, new_n27159_, new_n27160_,
    new_n27161_, new_n27162_, new_n27163_, new_n27164_, new_n27165_,
    new_n27166_, new_n27167_, new_n27168_, new_n27169_, new_n27170_,
    new_n27171_, new_n27172_, new_n27173_, new_n27174_, new_n27175_,
    new_n27176_, new_n27177_, new_n27178_, new_n27179_, new_n27180_,
    new_n27181_, new_n27182_, new_n27183_, new_n27184_, new_n27185_,
    new_n27186_, new_n27187_, new_n27188_, new_n27189_, new_n27190_,
    new_n27191_, new_n27192_, new_n27193_, new_n27194_, new_n27195_,
    new_n27196_, new_n27197_, new_n27198_, new_n27199_, new_n27200_,
    new_n27201_, new_n27202_, new_n27203_, new_n27204_, new_n27205_,
    new_n27206_, new_n27207_, new_n27208_, new_n27209_, new_n27210_,
    new_n27211_, new_n27212_, new_n27213_, new_n27214_, new_n27215_,
    new_n27216_, new_n27217_, new_n27218_, new_n27219_, new_n27220_,
    new_n27221_, new_n27222_, new_n27223_, new_n27224_, new_n27225_,
    new_n27226_, new_n27227_, new_n27228_, new_n27229_, new_n27230_,
    new_n27231_, new_n27232_, new_n27233_, new_n27234_, new_n27235_,
    new_n27236_, new_n27237_, new_n27238_, new_n27239_, new_n27240_,
    new_n27241_, new_n27242_, new_n27243_, new_n27244_, new_n27245_,
    new_n27246_, new_n27247_, new_n27248_, new_n27249_, new_n27250_,
    new_n27251_, new_n27252_, new_n27253_, new_n27254_, new_n27255_,
    new_n27256_, new_n27257_, new_n27258_, new_n27259_, new_n27260_,
    new_n27261_, new_n27262_, new_n27263_, new_n27264_, new_n27265_,
    new_n27266_, new_n27267_, new_n27268_, new_n27269_, new_n27270_,
    new_n27271_, new_n27272_, new_n27273_, new_n27274_, new_n27275_,
    new_n27276_, new_n27277_, new_n27278_, new_n27279_, new_n27280_,
    new_n27281_, new_n27282_, new_n27283_, new_n27284_, new_n27285_,
    new_n27286_, new_n27287_, new_n27288_, new_n27289_, new_n27290_,
    new_n27291_, new_n27292_, new_n27293_, new_n27294_, new_n27295_,
    new_n27296_, new_n27297_, new_n27298_, new_n27299_, new_n27300_,
    new_n27301_, new_n27302_, new_n27303_, new_n27304_, new_n27305_,
    new_n27306_, new_n27307_, new_n27308_, new_n27309_, new_n27310_,
    new_n27311_, new_n27312_, new_n27313_, new_n27314_, new_n27315_,
    new_n27316_, new_n27317_, new_n27318_, new_n27319_, new_n27320_,
    new_n27321_, new_n27322_, new_n27323_, new_n27324_, new_n27325_,
    new_n27326_, new_n27327_, new_n27328_, new_n27329_, new_n27330_,
    new_n27331_, new_n27332_, new_n27333_, new_n27334_, new_n27335_,
    new_n27336_, new_n27337_, new_n27338_, new_n27339_, new_n27340_,
    new_n27341_, new_n27342_, new_n27343_, new_n27344_, new_n27345_,
    new_n27346_, new_n27347_, new_n27348_, new_n27349_, new_n27350_,
    new_n27351_, new_n27352_, new_n27353_, new_n27354_, new_n27355_,
    new_n27356_, new_n27357_, new_n27358_, new_n27359_, new_n27360_,
    new_n27361_, new_n27362_, new_n27363_, new_n27364_, new_n27365_,
    new_n27366_, new_n27367_, new_n27368_, new_n27369_, new_n27370_,
    new_n27371_, new_n27372_, new_n27373_, new_n27374_, new_n27375_,
    new_n27376_, new_n27377_, new_n27378_, new_n27379_, new_n27380_,
    new_n27381_, new_n27382_, new_n27383_, new_n27384_, new_n27385_,
    new_n27386_, new_n27387_, new_n27388_, new_n27389_, new_n27390_,
    new_n27391_, new_n27392_, new_n27393_, new_n27394_, new_n27395_,
    new_n27396_, new_n27397_, new_n27398_, new_n27399_, new_n27400_,
    new_n27401_, new_n27402_, new_n27403_, new_n27404_, new_n27405_,
    new_n27406_, new_n27407_, new_n27408_, new_n27409_, new_n27410_,
    new_n27411_, new_n27412_, new_n27413_, new_n27414_, new_n27415_,
    new_n27416_, new_n27417_, new_n27418_, new_n27419_, new_n27420_,
    new_n27421_, new_n27422_, new_n27423_, new_n27424_, new_n27425_,
    new_n27426_, new_n27427_, new_n27428_, new_n27429_, new_n27430_,
    new_n27431_, new_n27432_, new_n27433_, new_n27434_, new_n27435_,
    new_n27436_, new_n27437_, new_n27438_, new_n27439_, new_n27440_,
    new_n27441_, new_n27442_, new_n27443_, new_n27444_, new_n27445_,
    new_n27446_, new_n27447_, new_n27448_, new_n27449_, new_n27450_,
    new_n27451_, new_n27452_, new_n27453_, new_n27454_, new_n27455_,
    new_n27456_, new_n27457_, new_n27458_, new_n27459_, new_n27460_,
    new_n27461_, new_n27462_, new_n27463_, new_n27464_, new_n27465_,
    new_n27466_, new_n27467_, new_n27468_, new_n27469_, new_n27470_,
    new_n27471_, new_n27472_, new_n27473_, new_n27474_, new_n27475_,
    new_n27476_, new_n27477_, new_n27478_, new_n27479_, new_n27480_,
    new_n27481_, new_n27482_, new_n27483_, new_n27484_, new_n27485_,
    new_n27486_, new_n27487_, new_n27488_, new_n27489_, new_n27490_,
    new_n27491_, new_n27492_, new_n27493_, new_n27494_, new_n27495_,
    new_n27496_, new_n27497_, new_n27498_, new_n27499_, new_n27500_,
    new_n27501_, new_n27502_, new_n27503_, new_n27504_, new_n27505_,
    new_n27506_, new_n27507_, new_n27508_, new_n27509_, new_n27510_,
    new_n27511_, new_n27512_, new_n27513_, new_n27514_, new_n27515_,
    new_n27516_, new_n27517_, new_n27518_, new_n27519_, new_n27520_,
    new_n27521_, new_n27522_, new_n27523_, new_n27524_, new_n27525_,
    new_n27526_, new_n27527_, new_n27528_, new_n27529_, new_n27530_,
    new_n27531_, new_n27532_, new_n27533_, new_n27534_, new_n27535_,
    new_n27536_, new_n27537_, new_n27538_, new_n27539_, new_n27540_,
    new_n27541_, new_n27542_, new_n27543_, new_n27544_, new_n27545_,
    new_n27546_, new_n27547_, new_n27548_, new_n27549_, new_n27550_,
    new_n27551_, new_n27552_, new_n27553_, new_n27554_, new_n27555_,
    new_n27556_, new_n27557_, new_n27558_, new_n27559_, new_n27560_,
    new_n27561_, new_n27562_, new_n27563_, new_n27564_, new_n27565_,
    new_n27566_, new_n27567_, new_n27568_, new_n27569_, new_n27570_,
    new_n27571_, new_n27572_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27577_, new_n27578_, new_n27579_, new_n27580_,
    new_n27581_, new_n27582_, new_n27583_, new_n27584_, new_n27585_,
    new_n27586_, new_n27587_, new_n27588_, new_n27589_, new_n27590_,
    new_n27591_, new_n27592_, new_n27593_, new_n27594_, new_n27595_,
    new_n27596_, new_n27597_, new_n27598_, new_n27599_, new_n27600_,
    new_n27601_, new_n27602_, new_n27603_, new_n27604_, new_n27605_,
    new_n27606_, new_n27607_, new_n27608_, new_n27609_, new_n27610_,
    new_n27611_, new_n27612_, new_n27613_, new_n27614_, new_n27615_,
    new_n27616_, new_n27617_, new_n27618_, new_n27619_, new_n27620_,
    new_n27621_, new_n27622_, new_n27623_, new_n27624_, new_n27625_,
    new_n27626_, new_n27627_, new_n27628_, new_n27629_, new_n27630_,
    new_n27631_, new_n27632_, new_n27633_, new_n27634_, new_n27635_,
    new_n27636_, new_n27637_, new_n27638_, new_n27639_, new_n27640_,
    new_n27641_, new_n27642_, new_n27643_, new_n27644_, new_n27645_,
    new_n27646_, new_n27647_, new_n27648_, new_n27649_, new_n27650_,
    new_n27651_, new_n27652_, new_n27653_, new_n27654_, new_n27655_,
    new_n27656_, new_n27657_, new_n27658_, new_n27659_, new_n27660_,
    new_n27661_, new_n27662_, new_n27663_, new_n27664_, new_n27665_,
    new_n27666_, new_n27667_, new_n27668_, new_n27669_, new_n27670_,
    new_n27671_, new_n27672_, new_n27673_, new_n27674_, new_n27675_,
    new_n27676_, new_n27677_, new_n27678_, new_n27679_, new_n27680_,
    new_n27681_, new_n27682_, new_n27683_, new_n27684_, new_n27685_,
    new_n27686_, new_n27687_, new_n27688_, new_n27689_, new_n27690_,
    new_n27691_, new_n27692_, new_n27693_, new_n27694_, new_n27695_,
    new_n27696_, new_n27697_, new_n27698_, new_n27699_, new_n27700_,
    new_n27701_, new_n27702_, new_n27703_, new_n27704_, new_n27705_,
    new_n27706_, new_n27707_, new_n27708_, new_n27709_, new_n27710_,
    new_n27711_, new_n27712_, new_n27713_, new_n27714_, new_n27715_,
    new_n27716_, new_n27717_, new_n27718_, new_n27719_, new_n27720_,
    new_n27721_, new_n27722_, new_n27723_, new_n27724_, new_n27725_,
    new_n27726_, new_n27727_, new_n27728_, new_n27729_, new_n27730_,
    new_n27731_, new_n27732_, new_n27733_, new_n27734_, new_n27735_,
    new_n27736_, new_n27737_, new_n27738_, new_n27739_, new_n27740_,
    new_n27741_, new_n27742_, new_n27743_, new_n27744_, new_n27745_,
    new_n27746_, new_n27747_, new_n27748_, new_n27749_, new_n27750_,
    new_n27751_, new_n27752_, new_n27753_, new_n27754_, new_n27755_,
    new_n27756_, new_n27757_, new_n27758_, new_n27759_, new_n27760_,
    new_n27761_, new_n27762_, new_n27763_, new_n27764_, new_n27765_,
    new_n27766_, new_n27767_, new_n27768_, new_n27769_, new_n27770_,
    new_n27771_, new_n27772_, new_n27773_, new_n27774_, new_n27775_,
    new_n27776_, new_n27777_, new_n27778_, new_n27779_, new_n27780_,
    new_n27781_, new_n27782_, new_n27783_, new_n27784_, new_n27785_,
    new_n27786_, new_n27787_, new_n27788_, new_n27789_, new_n27790_,
    new_n27791_, new_n27792_, new_n27793_, new_n27794_, new_n27795_,
    new_n27796_, new_n27797_, new_n27798_, new_n27799_, new_n27800_,
    new_n27801_, new_n27802_, new_n27803_, new_n27804_, new_n27805_,
    new_n27806_, new_n27807_, new_n27808_, new_n27809_, new_n27810_,
    new_n27811_, new_n27812_, new_n27813_, new_n27814_, new_n27815_,
    new_n27816_, new_n27817_, new_n27818_, new_n27819_, new_n27820_,
    new_n27821_, new_n27822_, new_n27823_, new_n27824_, new_n27825_,
    new_n27826_, new_n27827_, new_n27828_, new_n27829_, new_n27830_,
    new_n27831_, new_n27832_, new_n27833_, new_n27834_, new_n27835_,
    new_n27836_, new_n27837_, new_n27838_, new_n27839_, new_n27840_,
    new_n27841_, new_n27842_, new_n27843_, new_n27844_, new_n27845_,
    new_n27846_, new_n27847_, new_n27848_, new_n27849_, new_n27850_,
    new_n27851_, new_n27852_, new_n27853_, new_n27854_, new_n27855_,
    new_n27856_, new_n27857_, new_n27858_, new_n27859_, new_n27860_,
    new_n27861_, new_n27862_, new_n27863_, new_n27864_, new_n27865_,
    new_n27866_, new_n27867_, new_n27868_, new_n27869_, new_n27870_,
    new_n27871_, new_n27872_, new_n27873_, new_n27874_, new_n27875_,
    new_n27876_, new_n27877_, new_n27878_, new_n27879_, new_n27880_,
    new_n27881_, new_n27882_, new_n27883_, new_n27884_, new_n27885_,
    new_n27886_, new_n27887_, new_n27888_, new_n27889_, new_n27890_,
    new_n27891_, new_n27892_, new_n27893_, new_n27894_, new_n27895_,
    new_n27896_, new_n27897_, new_n27898_, new_n27899_, new_n27900_,
    new_n27901_, new_n27902_, new_n27903_, new_n27904_, new_n27905_,
    new_n27906_, new_n27907_, new_n27908_, new_n27909_, new_n27910_,
    new_n27911_, new_n27912_, new_n27913_, new_n27914_, new_n27915_,
    new_n27916_, new_n27917_, new_n27918_, new_n27919_, new_n27920_,
    new_n27921_, new_n27922_, new_n27923_, new_n27924_, new_n27925_,
    new_n27926_, new_n27927_, new_n27928_, new_n27929_, new_n27930_,
    new_n27931_, new_n27932_, new_n27933_, new_n27934_, new_n27935_,
    new_n27936_, new_n27937_, new_n27938_, new_n27939_, new_n27940_,
    new_n27941_, new_n27942_, new_n27943_, new_n27944_, new_n27945_,
    new_n27946_, new_n27947_, new_n27948_, new_n27949_, new_n27950_,
    new_n27951_, new_n27952_, new_n27953_, new_n27954_, new_n27955_,
    new_n27956_, new_n27957_, new_n27958_, new_n27959_, new_n27960_,
    new_n27961_, new_n27962_, new_n27963_, new_n27964_, new_n27965_,
    new_n27966_, new_n27967_, new_n27968_, new_n27969_, new_n27970_,
    new_n27971_, new_n27972_, new_n27973_, new_n27974_, new_n27975_,
    new_n27976_, new_n27977_, new_n27978_, new_n27979_, new_n27980_,
    new_n27981_, new_n27982_, new_n27983_, new_n27984_, new_n27985_,
    new_n27986_, new_n27987_, new_n27988_, new_n27989_, new_n27990_,
    new_n27991_, new_n27992_, new_n27993_, new_n27994_, new_n27995_,
    new_n27996_, new_n27997_, new_n27998_, new_n27999_, new_n28000_,
    new_n28001_, new_n28002_, new_n28003_, new_n28004_, new_n28005_,
    new_n28006_, new_n28007_, new_n28008_, new_n28009_, new_n28010_,
    new_n28011_, new_n28012_, new_n28013_, new_n28014_, new_n28015_,
    new_n28016_, new_n28017_, new_n28018_, new_n28019_, new_n28020_,
    new_n28021_, new_n28022_, new_n28023_, new_n28024_, new_n28025_,
    new_n28026_, new_n28027_, new_n28028_, new_n28029_, new_n28030_,
    new_n28031_, new_n28032_, new_n28033_, new_n28034_, new_n28035_,
    new_n28036_, new_n28037_, new_n28038_, new_n28039_, new_n28040_,
    new_n28041_, new_n28042_, new_n28043_, new_n28044_, new_n28045_,
    new_n28046_, new_n28047_, new_n28048_, new_n28049_, new_n28050_,
    new_n28051_, new_n28052_, new_n28053_, new_n28054_, new_n28055_,
    new_n28056_, new_n28057_, new_n28058_, new_n28059_, new_n28060_,
    new_n28061_, new_n28062_, new_n28063_, new_n28064_, new_n28065_,
    new_n28066_, new_n28067_, new_n28068_, new_n28069_, new_n28070_,
    new_n28071_, new_n28072_, new_n28073_, new_n28074_, new_n28075_,
    new_n28076_, new_n28077_, new_n28078_, new_n28079_, new_n28080_,
    new_n28081_, new_n28082_, new_n28083_, new_n28084_, new_n28085_,
    new_n28086_, new_n28087_, new_n28088_, new_n28089_, new_n28090_,
    new_n28091_, new_n28092_, new_n28093_, new_n28094_, new_n28095_,
    new_n28096_, new_n28097_, new_n28098_, new_n28099_, new_n28100_,
    new_n28101_, new_n28102_, new_n28103_, new_n28104_, new_n28105_,
    new_n28106_, new_n28107_, new_n28108_, new_n28109_, new_n28110_,
    new_n28111_, new_n28112_, new_n28113_, new_n28114_, new_n28115_,
    new_n28116_, new_n28117_, new_n28118_, new_n28119_, new_n28120_,
    new_n28121_, new_n28122_, new_n28123_, new_n28124_, new_n28125_,
    new_n28126_, new_n28127_, new_n28128_, new_n28129_, new_n28130_,
    new_n28131_, new_n28132_, new_n28133_, new_n28134_, new_n28135_,
    new_n28136_, new_n28137_, new_n28138_, new_n28139_, new_n28140_,
    new_n28141_, new_n28142_, new_n28143_, new_n28144_, new_n28145_,
    new_n28146_, new_n28147_, new_n28148_, new_n28149_, new_n28150_,
    new_n28151_, new_n28152_, new_n28153_, new_n28154_, new_n28155_,
    new_n28156_, new_n28157_, new_n28158_, new_n28159_, new_n28160_,
    new_n28161_, new_n28162_, new_n28163_, new_n28164_, new_n28165_,
    new_n28166_, new_n28167_, new_n28168_, new_n28169_, new_n28170_,
    new_n28171_, new_n28172_, new_n28173_, new_n28174_, new_n28175_,
    new_n28176_, new_n28177_, new_n28178_, new_n28179_, new_n28180_,
    new_n28181_, new_n28182_, new_n28183_, new_n28184_, new_n28185_,
    new_n28186_, new_n28187_, new_n28188_, new_n28189_, new_n28190_,
    new_n28191_, new_n28192_, new_n28193_, new_n28194_, new_n28195_,
    new_n28196_, new_n28197_, new_n28198_, new_n28199_, new_n28200_,
    new_n28201_, new_n28202_, new_n28203_, new_n28204_, new_n28205_,
    new_n28206_, new_n28207_, new_n28208_, new_n28209_, new_n28210_,
    new_n28211_, new_n28212_, new_n28213_, new_n28214_, new_n28215_,
    new_n28216_, new_n28217_, new_n28218_, new_n28219_, new_n28220_,
    new_n28221_, new_n28222_, new_n28223_, new_n28224_, new_n28225_,
    new_n28226_, new_n28227_, new_n28228_, new_n28229_, new_n28230_,
    new_n28231_, new_n28232_, new_n28233_, new_n28234_, new_n28235_,
    new_n28236_, new_n28237_, new_n28238_, new_n28239_, new_n28240_,
    new_n28241_, new_n28242_, new_n28243_, new_n28244_, new_n28245_,
    new_n28246_, new_n28247_, new_n28248_, new_n28249_, new_n28250_,
    new_n28251_, new_n28252_, new_n28253_, new_n28254_, new_n28255_,
    new_n28256_, new_n28257_, new_n28258_, new_n28259_, new_n28260_,
    new_n28261_, new_n28262_, new_n28263_, new_n28264_, new_n28265_,
    new_n28266_, new_n28267_, new_n28268_, new_n28269_, new_n28270_,
    new_n28271_, new_n28272_, new_n28273_, new_n28274_, new_n28275_,
    new_n28276_, new_n28277_, new_n28278_, new_n28279_, new_n28280_,
    new_n28281_, new_n28282_, new_n28283_, new_n28284_, new_n28285_,
    new_n28286_, new_n28287_, new_n28288_, new_n28289_, new_n28290_,
    new_n28291_, new_n28292_, new_n28293_, new_n28294_, new_n28295_,
    new_n28296_, new_n28297_, new_n28298_, new_n28299_, new_n28300_,
    new_n28301_, new_n28302_, new_n28303_, new_n28304_, new_n28305_,
    new_n28306_, new_n28307_, new_n28308_, new_n28309_, new_n28310_,
    new_n28311_, new_n28312_, new_n28313_, new_n28314_, new_n28315_,
    new_n28316_, new_n28317_, new_n28318_, new_n28319_, new_n28320_,
    new_n28321_, new_n28322_, new_n28323_, new_n28324_, new_n28325_,
    new_n28326_, new_n28327_, new_n28328_, new_n28329_, new_n28330_,
    new_n28331_, new_n28332_, new_n28333_, new_n28334_, new_n28335_,
    new_n28336_, new_n28337_, new_n28338_, new_n28339_, new_n28340_,
    new_n28341_, new_n28342_, new_n28343_, new_n28344_, new_n28345_,
    new_n28346_, new_n28347_, new_n28348_, new_n28349_, new_n28350_,
    new_n28351_, new_n28352_, new_n28353_, new_n28354_, new_n28355_,
    new_n28356_, new_n28357_, new_n28358_, new_n28359_, new_n28360_,
    new_n28361_, new_n28362_, new_n28363_, new_n28364_, new_n28365_,
    new_n28366_, new_n28367_, new_n28368_, new_n28369_, new_n28370_,
    new_n28371_, new_n28372_, new_n28373_, new_n28374_, new_n28375_,
    new_n28376_, new_n28377_, new_n28378_, new_n28379_, new_n28380_,
    new_n28381_, new_n28382_, new_n28383_, new_n28384_, new_n28385_,
    new_n28386_, new_n28387_, new_n28388_, new_n28389_, new_n28390_,
    new_n28391_, new_n28392_, new_n28393_, new_n28394_, new_n28395_,
    new_n28396_, new_n28397_, new_n28398_, new_n28399_, new_n28400_,
    new_n28401_, new_n28402_, new_n28403_, new_n28404_, new_n28405_,
    new_n28406_, new_n28407_, new_n28408_, new_n28409_, new_n28410_,
    new_n28411_, new_n28412_, new_n28413_, new_n28414_, new_n28415_,
    new_n28416_, new_n28417_, new_n28418_, new_n28419_, new_n28420_,
    new_n28421_, new_n28422_, new_n28423_, new_n28424_, new_n28425_,
    new_n28426_, new_n28427_, new_n28428_, new_n28429_, new_n28430_,
    new_n28431_, new_n28432_, new_n28433_, new_n28434_, new_n28435_,
    new_n28436_, new_n28437_, new_n28438_, new_n28439_, new_n28440_,
    new_n28441_, new_n28442_, new_n28443_, new_n28444_, new_n28445_,
    new_n28446_, new_n28447_, new_n28448_, new_n28449_, new_n28450_,
    new_n28451_, new_n28452_, new_n28453_, new_n28454_, new_n28455_,
    new_n28456_, new_n28457_, new_n28458_, new_n28459_, new_n28460_,
    new_n28461_, new_n28462_, new_n28463_, new_n28464_, new_n28465_,
    new_n28466_, new_n28467_, new_n28468_, new_n28469_, new_n28470_,
    new_n28471_, new_n28472_, new_n28473_, new_n28474_, new_n28475_,
    new_n28476_, new_n28477_, new_n28478_, new_n28479_, new_n28480_,
    new_n28481_, new_n28482_, new_n28483_, new_n28484_, new_n28485_,
    new_n28486_, new_n28487_, new_n28488_, new_n28489_, new_n28490_,
    new_n28491_, new_n28492_, new_n28493_, new_n28494_, new_n28495_,
    new_n28496_, new_n28497_, new_n28498_, new_n28499_, new_n28500_,
    new_n28501_, new_n28502_, new_n28503_, new_n28504_, new_n28505_,
    new_n28506_, new_n28507_, new_n28508_, new_n28509_, new_n28510_,
    new_n28511_, new_n28512_, new_n28513_, new_n28514_, new_n28515_,
    new_n28516_, new_n28517_, new_n28518_, new_n28519_, new_n28520_,
    new_n28521_, new_n28522_, new_n28523_, new_n28524_, new_n28525_,
    new_n28526_, new_n28527_, new_n28528_, new_n28529_, new_n28530_,
    new_n28531_, new_n28532_, new_n28533_, new_n28534_, new_n28535_,
    new_n28536_, new_n28537_, new_n28538_, new_n28539_, new_n28540_,
    new_n28541_, new_n28542_, new_n28543_, new_n28544_, new_n28545_,
    new_n28546_, new_n28547_, new_n28548_, new_n28549_, new_n28550_,
    new_n28551_, new_n28552_, new_n28553_, new_n28554_, new_n28555_,
    new_n28556_, new_n28557_, new_n28558_, new_n28559_, new_n28560_,
    new_n28561_, new_n28562_, new_n28563_, new_n28564_, new_n28565_,
    new_n28566_, new_n28567_, new_n28568_, new_n28569_, new_n28570_,
    new_n28571_, new_n28572_, new_n28573_, new_n28574_, new_n28575_,
    new_n28576_, new_n28577_, new_n28578_, new_n28579_, new_n28580_,
    new_n28581_, new_n28582_, new_n28583_, new_n28584_, new_n28585_,
    new_n28586_, new_n28587_, new_n28588_, new_n28589_, new_n28590_,
    new_n28591_, new_n28592_, new_n28593_, new_n28594_, new_n28595_,
    new_n28596_, new_n28597_, new_n28598_, new_n28599_, new_n28600_,
    new_n28601_, new_n28602_, new_n28603_, new_n28604_, new_n28605_,
    new_n28606_, new_n28607_, new_n28608_, new_n28609_, new_n28610_,
    new_n28611_, new_n28612_, new_n28613_, new_n28614_, new_n28615_,
    new_n28616_, new_n28617_, new_n28618_, new_n28619_, new_n28620_,
    new_n28621_, new_n28622_, new_n28623_, new_n28624_, new_n28625_,
    new_n28626_, new_n28627_, new_n28628_, new_n28629_, new_n28630_,
    new_n28631_, new_n28632_, new_n28633_, new_n28634_, new_n28635_,
    new_n28636_, new_n28637_, new_n28638_, new_n28639_, new_n28640_,
    new_n28641_, new_n28642_, new_n28643_, new_n28644_, new_n28645_,
    new_n28646_, new_n28647_, new_n28648_, new_n28649_, new_n28650_,
    new_n28651_, new_n28652_, new_n28653_, new_n28654_, new_n28655_,
    new_n28656_, new_n28657_, new_n28658_, new_n28659_, new_n28660_,
    new_n28661_, new_n28662_, new_n28663_, new_n28664_, new_n28665_,
    new_n28666_, new_n28667_, new_n28668_, new_n28669_, new_n28670_,
    new_n28671_, new_n28672_, new_n28673_, new_n28674_, new_n28675_,
    new_n28676_, new_n28677_, new_n28678_, new_n28679_, new_n28680_,
    new_n28681_, new_n28682_, new_n28683_, new_n28684_, new_n28685_,
    new_n28686_, new_n28687_, new_n28688_, new_n28689_, new_n28690_,
    new_n28691_, new_n28692_, new_n28693_, new_n28694_, new_n28695_,
    new_n28696_, new_n28697_, new_n28698_, new_n28699_, new_n28700_,
    new_n28701_, new_n28702_, new_n28703_, new_n28704_, new_n28705_,
    new_n28706_, new_n28707_, new_n28708_, new_n28709_, new_n28710_,
    new_n28711_, new_n28712_, new_n28713_, new_n28714_, new_n28715_,
    new_n28716_, new_n28717_, new_n28718_, new_n28719_, new_n28720_,
    new_n28721_, new_n28722_, new_n28723_, new_n28724_, new_n28725_,
    new_n28726_, new_n28727_, new_n28728_, new_n28729_, new_n28730_,
    new_n28731_, new_n28732_, new_n28733_, new_n28734_, new_n28735_,
    new_n28736_, new_n28737_, new_n28738_, new_n28739_, new_n28740_,
    new_n28741_, new_n28742_, new_n28743_, new_n28744_, new_n28745_,
    new_n28746_, new_n28747_, new_n28748_, new_n28749_, new_n28750_,
    new_n28751_, new_n28752_, new_n28753_, new_n28754_, new_n28755_,
    new_n28756_, new_n28757_, new_n28758_, new_n28759_, new_n28760_,
    new_n28761_, new_n28762_, new_n28763_, new_n28764_, new_n28765_,
    new_n28766_, new_n28767_, new_n28768_, new_n28769_, new_n28770_,
    new_n28771_, new_n28772_, new_n28773_, new_n28774_, new_n28775_,
    new_n28776_, new_n28777_, new_n28778_, new_n28779_, new_n28780_,
    new_n28781_, new_n28782_, new_n28783_, new_n28784_, new_n28785_,
    new_n28786_, new_n28787_, new_n28788_, new_n28789_, new_n28790_,
    new_n28791_, new_n28792_, new_n28793_, new_n28794_, new_n28795_,
    new_n28796_, new_n28797_, new_n28798_, new_n28799_, new_n28800_,
    new_n28801_, new_n28802_, new_n28803_, new_n28804_, new_n28805_,
    new_n28806_, new_n28807_, new_n28808_, new_n28809_, new_n28810_,
    new_n28811_, new_n28812_, new_n28813_, new_n28814_, new_n28815_,
    new_n28816_, new_n28817_, new_n28818_, new_n28819_, new_n28820_,
    new_n28821_, new_n28822_, new_n28823_, new_n28824_, new_n28825_,
    new_n28826_, new_n28827_, new_n28828_, new_n28829_, new_n28830_,
    new_n28831_, new_n28832_, new_n28833_, new_n28834_, new_n28835_,
    new_n28836_, new_n28837_, new_n28838_, new_n28839_, new_n28840_,
    new_n28841_, new_n28842_, new_n28843_, new_n28844_, new_n28845_,
    new_n28846_, new_n28847_, new_n28848_, new_n28849_, new_n28850_,
    new_n28851_, new_n28852_, new_n28853_, new_n28854_, new_n28855_,
    new_n28856_, new_n28857_, new_n28858_, new_n28859_, new_n28860_,
    new_n28861_, new_n28862_, new_n28863_, new_n28864_, new_n28865_,
    new_n28866_, new_n28867_, new_n28868_, new_n28869_, new_n28870_,
    new_n28871_, new_n28872_, new_n28873_, new_n28874_, new_n28875_,
    new_n28876_, new_n28877_, new_n28878_, new_n28879_, new_n28880_,
    new_n28881_, new_n28882_, new_n28883_, new_n28884_, new_n28885_,
    new_n28886_, new_n28887_, new_n28888_, new_n28889_, new_n28890_,
    new_n28891_, new_n28892_, new_n28893_, new_n28894_, new_n28895_,
    new_n28896_, new_n28897_, new_n28898_, new_n28899_, new_n28900_,
    new_n28901_, new_n28902_, new_n28903_, new_n28904_, new_n28905_,
    new_n28906_, new_n28907_, new_n28908_, new_n28909_, new_n28910_,
    new_n28911_, new_n28912_, new_n28913_, new_n28914_, new_n28915_,
    new_n28916_, new_n28917_, new_n28918_, new_n28919_, new_n28920_,
    new_n28921_, new_n28922_, new_n28923_, new_n28924_, new_n28925_,
    new_n28926_, new_n28927_, new_n28928_, new_n28929_, new_n28930_,
    new_n28931_, new_n28932_, new_n28933_, new_n28934_, new_n28935_,
    new_n28936_, new_n28937_, new_n28938_, new_n28939_, new_n28940_,
    new_n28941_, new_n28942_, new_n28943_, new_n28944_, new_n28945_,
    new_n28946_, new_n28947_, new_n28948_, new_n28949_, new_n28950_,
    new_n28951_, new_n28952_, new_n28953_, new_n28954_, new_n28955_,
    new_n28956_, new_n28957_, new_n28958_, new_n28959_, new_n28960_,
    new_n28961_, new_n28962_, new_n28963_, new_n28964_, new_n28965_,
    new_n28966_, new_n28967_, new_n28968_, new_n28969_, new_n28970_,
    new_n28971_, new_n28972_, new_n28973_, new_n28974_, new_n28975_,
    new_n28976_, new_n28977_, new_n28978_, new_n28979_, new_n28980_,
    new_n28981_, new_n28982_, new_n28983_, new_n28984_, new_n28985_,
    new_n28986_, new_n28987_, new_n28988_, new_n28989_, new_n28990_,
    new_n28991_, new_n28992_, new_n28993_, new_n28994_, new_n28995_,
    new_n28996_, new_n28997_, new_n28998_, new_n28999_, new_n29000_,
    new_n29001_, new_n29002_, new_n29003_, new_n29004_, new_n29005_,
    new_n29006_, new_n29007_, new_n29008_, new_n29009_, new_n29010_,
    new_n29011_, new_n29012_, new_n29013_, new_n29014_, new_n29015_,
    new_n29016_, new_n29017_, new_n29018_, new_n29019_, new_n29020_,
    new_n29021_, new_n29022_, new_n29023_, new_n29024_, new_n29025_,
    new_n29026_, new_n29027_, new_n29028_, new_n29029_, new_n29030_,
    new_n29031_, new_n29032_, new_n29033_, new_n29034_, new_n29035_,
    new_n29036_, new_n29037_, new_n29038_, new_n29039_, new_n29040_,
    new_n29041_, new_n29042_, new_n29043_, new_n29044_, new_n29045_,
    new_n29046_, new_n29047_, new_n29048_, new_n29049_, new_n29050_,
    new_n29051_, new_n29052_, new_n29053_, new_n29054_, new_n29055_,
    new_n29056_, new_n29057_, new_n29058_, new_n29059_, new_n29060_,
    new_n29061_, new_n29062_, new_n29063_, new_n29064_, new_n29065_,
    new_n29066_, new_n29067_, new_n29068_, new_n29069_, new_n29070_,
    new_n29071_, new_n29072_, new_n29073_, new_n29074_, new_n29075_,
    new_n29076_, new_n29077_, new_n29078_, new_n29079_, new_n29080_,
    new_n29081_, new_n29082_, new_n29083_, new_n29084_, new_n29085_,
    new_n29086_, new_n29087_, new_n29088_, new_n29089_, new_n29090_,
    new_n29091_, new_n29092_, new_n29093_, new_n29094_, new_n29095_,
    new_n29096_, new_n29097_, new_n29098_, new_n29099_, new_n29100_,
    new_n29101_, new_n29102_, new_n29103_, new_n29104_, new_n29105_,
    new_n29106_, new_n29107_, new_n29108_, new_n29109_, new_n29110_,
    new_n29111_, new_n29112_, new_n29113_, new_n29114_, new_n29115_,
    new_n29116_, new_n29117_, new_n29118_, new_n29119_, new_n29120_,
    new_n29121_, new_n29122_, new_n29123_, new_n29124_, new_n29125_,
    new_n29126_, new_n29127_, new_n29128_, new_n29129_, new_n29130_,
    new_n29131_, new_n29132_, new_n29133_, new_n29134_, new_n29135_,
    new_n29136_, new_n29137_, new_n29138_, new_n29139_, new_n29140_,
    new_n29141_, new_n29142_, new_n29143_, new_n29144_, new_n29145_,
    new_n29146_, new_n29147_, new_n29148_, new_n29149_, new_n29150_,
    new_n29151_, new_n29152_, new_n29153_, new_n29154_, new_n29155_,
    new_n29156_, new_n29157_, new_n29158_, new_n29159_, new_n29160_,
    new_n29161_, new_n29162_, new_n29163_, new_n29164_, new_n29165_,
    new_n29166_, new_n29167_, new_n29168_, new_n29169_, new_n29170_,
    new_n29171_, new_n29172_, new_n29173_, new_n29174_, new_n29175_,
    new_n29176_, new_n29177_, new_n29178_, new_n29179_, new_n29180_,
    new_n29181_, new_n29182_, new_n29183_, new_n29184_, new_n29185_,
    new_n29186_, new_n29187_, new_n29188_, new_n29189_, new_n29190_,
    new_n29191_, new_n29192_, new_n29193_, new_n29194_, new_n29195_,
    new_n29196_, new_n29197_, new_n29198_, new_n29199_, new_n29200_,
    new_n29201_, new_n29202_, new_n29203_, new_n29204_, new_n29205_,
    new_n29206_, new_n29207_, new_n29208_, new_n29209_, new_n29210_,
    new_n29211_, new_n29212_, new_n29213_, new_n29214_, new_n29215_,
    new_n29216_, new_n29217_, new_n29218_, new_n29219_, new_n29220_,
    new_n29221_, new_n29222_, new_n29223_, new_n29224_, new_n29225_,
    new_n29226_, new_n29227_, new_n29228_, new_n29229_, new_n29230_,
    new_n29231_, new_n29232_, new_n29233_, new_n29234_, new_n29235_,
    new_n29236_, new_n29237_, new_n29238_, new_n29239_, new_n29240_,
    new_n29241_, new_n29242_, new_n29243_, new_n29244_, new_n29245_,
    new_n29246_, new_n29247_, new_n29248_, new_n29249_, new_n29250_,
    new_n29251_, new_n29252_, new_n29253_, new_n29254_, new_n29255_,
    new_n29256_, new_n29257_, new_n29258_, new_n29259_, new_n29260_,
    new_n29261_, new_n29262_, new_n29263_, new_n29264_, new_n29265_,
    new_n29266_, new_n29267_, new_n29268_, new_n29269_, new_n29270_,
    new_n29271_, new_n29272_, new_n29273_, new_n29274_, new_n29275_,
    new_n29276_, new_n29277_, new_n29278_, new_n29279_, new_n29280_,
    new_n29281_, new_n29282_, new_n29283_, new_n29284_, new_n29285_,
    new_n29286_, new_n29287_, new_n29288_, new_n29289_, new_n29290_,
    new_n29291_, new_n29292_, new_n29293_, new_n29294_, new_n29295_,
    new_n29296_, new_n29297_, new_n29298_, new_n29299_, new_n29300_,
    new_n29301_, new_n29302_, new_n29303_, new_n29304_, new_n29305_,
    new_n29306_, new_n29307_, new_n29308_, new_n29309_, new_n29310_,
    new_n29311_, new_n29312_, new_n29313_, new_n29314_, new_n29315_,
    new_n29316_, new_n29317_, new_n29318_, new_n29319_, new_n29320_,
    new_n29321_, new_n29322_, new_n29323_, new_n29324_, new_n29325_,
    new_n29326_, new_n29327_, new_n29328_, new_n29329_, new_n29330_,
    new_n29331_, new_n29332_, new_n29333_, new_n29334_, new_n29335_,
    new_n29336_, new_n29337_, new_n29338_, new_n29339_, new_n29340_,
    new_n29341_, new_n29342_, new_n29343_, new_n29344_, new_n29345_,
    new_n29346_, new_n29347_, new_n29348_, new_n29349_, new_n29350_,
    new_n29351_, new_n29352_, new_n29353_, new_n29354_, new_n29355_,
    new_n29356_, new_n29357_, new_n29358_, new_n29359_, new_n29360_,
    new_n29361_, new_n29362_, new_n29363_, new_n29364_, new_n29365_,
    new_n29366_, new_n29367_, new_n29368_, new_n29369_, new_n29370_,
    new_n29371_, new_n29372_, new_n29373_, new_n29374_, new_n29375_,
    new_n29376_, new_n29377_, new_n29378_, new_n29379_, new_n29380_,
    new_n29381_, new_n29382_, new_n29383_, new_n29384_, new_n29385_,
    new_n29386_, new_n29387_, new_n29388_, new_n29389_, new_n29390_,
    new_n29391_, new_n29392_, new_n29393_, new_n29394_, new_n29395_,
    new_n29396_, new_n29397_, new_n29398_, new_n29399_, new_n29400_,
    new_n29401_, new_n29402_, new_n29403_, new_n29404_, new_n29405_,
    new_n29406_, new_n29407_, new_n29408_, new_n29409_, new_n29410_,
    new_n29411_, new_n29412_, new_n29413_, new_n29414_, new_n29415_,
    new_n29416_, new_n29417_, new_n29418_, new_n29419_, new_n29420_,
    new_n29421_, new_n29422_, new_n29423_, new_n29424_, new_n29425_,
    new_n29426_, new_n29427_, new_n29428_, new_n29429_, new_n29430_,
    new_n29431_, new_n29432_, new_n29433_, new_n29434_, new_n29435_,
    new_n29436_, new_n29437_, new_n29438_, new_n29439_, new_n29440_,
    new_n29441_, new_n29442_, new_n29443_, new_n29444_, new_n29445_,
    new_n29446_, new_n29447_, new_n29448_, new_n29449_, new_n29450_,
    new_n29451_, new_n29452_, new_n29453_, new_n29454_, new_n29455_,
    new_n29456_, new_n29457_, new_n29458_, new_n29459_, new_n29460_,
    new_n29461_, new_n29462_, new_n29463_, new_n29464_, new_n29465_,
    new_n29466_, new_n29467_, new_n29468_, new_n29469_, new_n29470_,
    new_n29471_, new_n29472_, new_n29473_, new_n29474_, new_n29475_,
    new_n29476_, new_n29477_, new_n29478_, new_n29479_, new_n29480_,
    new_n29481_, new_n29482_, new_n29483_, new_n29484_, new_n29485_,
    new_n29486_, new_n29487_, new_n29488_, new_n29489_, new_n29490_,
    new_n29491_, new_n29492_, new_n29493_, new_n29494_, new_n29495_,
    new_n29496_, new_n29497_, new_n29498_, new_n29499_, new_n29500_,
    new_n29501_, new_n29502_, new_n29503_, new_n29504_, new_n29505_,
    new_n29506_, new_n29507_, new_n29508_, new_n29509_, new_n29510_,
    new_n29511_, new_n29512_, new_n29513_, new_n29514_, new_n29515_,
    new_n29516_, new_n29517_, new_n29518_, new_n29519_, new_n29520_,
    new_n29521_, new_n29522_, new_n29523_, new_n29524_, new_n29525_,
    new_n29526_, new_n29527_, new_n29528_, new_n29529_, new_n29530_,
    new_n29531_, new_n29532_, new_n29533_, new_n29534_, new_n29535_,
    new_n29536_, new_n29537_, new_n29538_, new_n29539_, new_n29540_,
    new_n29541_, new_n29542_, new_n29543_, new_n29544_, new_n29545_,
    new_n29546_, new_n29547_, new_n29548_, new_n29549_, new_n29550_,
    new_n29551_, new_n29552_, new_n29553_, new_n29554_, new_n29555_,
    new_n29556_, new_n29557_, new_n29558_, new_n29559_, new_n29560_,
    new_n29561_, new_n29562_, new_n29563_, new_n29564_, new_n29565_,
    new_n29566_, new_n29567_, new_n29568_, new_n29569_, new_n29570_,
    new_n29571_, new_n29572_, new_n29573_, new_n29574_, new_n29575_,
    new_n29576_, new_n29577_, new_n29578_, new_n29579_, new_n29580_,
    new_n29581_, new_n29582_, new_n29583_, new_n29584_, new_n29585_,
    new_n29586_, new_n29587_, new_n29588_, new_n29589_, new_n29590_,
    new_n29591_, new_n29592_, new_n29593_, new_n29594_, new_n29595_,
    new_n29596_, new_n29597_, new_n29598_, new_n29599_, new_n29600_,
    new_n29601_, new_n29602_, new_n29603_, new_n29604_, new_n29605_,
    new_n29606_, new_n29607_, new_n29608_, new_n29609_, new_n29610_,
    new_n29611_, new_n29612_, new_n29613_, new_n29614_, new_n29615_,
    new_n29616_, new_n29617_, new_n29618_, new_n29619_, new_n29620_,
    new_n29621_, new_n29622_, new_n29623_, new_n29624_, new_n29625_,
    new_n29626_, new_n29627_, new_n29628_, new_n29629_, new_n29630_,
    new_n29631_, new_n29632_, new_n29633_, new_n29634_, new_n29635_,
    new_n29636_, new_n29637_, new_n29638_, new_n29639_, new_n29640_,
    new_n29641_, new_n29642_, new_n29643_, new_n29644_, new_n29645_,
    new_n29646_, new_n29647_, new_n29648_, new_n29649_, new_n29650_,
    new_n29651_, new_n29652_, new_n29653_, new_n29654_, new_n29655_,
    new_n29656_, new_n29657_, new_n29658_, new_n29659_, new_n29660_,
    new_n29661_, new_n29662_, new_n29663_, new_n29664_, new_n29665_,
    new_n29666_, new_n29667_, new_n29668_, new_n29669_, new_n29670_,
    new_n29671_, new_n29672_, new_n29673_, new_n29674_, new_n29675_,
    new_n29676_, new_n29677_, new_n29678_, new_n29679_, new_n29680_,
    new_n29681_, new_n29682_, new_n29683_, new_n29684_, new_n29685_,
    new_n29686_, new_n29687_, new_n29688_, new_n29689_, new_n29690_,
    new_n29691_, new_n29692_, new_n29693_, new_n29694_, new_n29695_,
    new_n29696_, new_n29697_, new_n29698_, new_n29699_, new_n29700_,
    new_n29701_, new_n29702_, new_n29703_, new_n29704_, new_n29705_,
    new_n29706_, new_n29707_, new_n29708_, new_n29709_, new_n29710_,
    new_n29711_, new_n29712_, new_n29713_, new_n29714_, new_n29715_,
    new_n29716_, new_n29717_, new_n29718_, new_n29719_, new_n29720_,
    new_n29721_, new_n29722_, new_n29723_, new_n29724_, new_n29725_,
    new_n29726_, new_n29727_, new_n29728_, new_n29729_, new_n29730_,
    new_n29731_, new_n29732_, new_n29733_, new_n29734_, new_n29735_,
    new_n29736_, new_n29737_, new_n29738_, new_n29739_, new_n29740_,
    new_n29741_, new_n29742_, new_n29743_, new_n29744_, new_n29745_,
    new_n29746_, new_n29747_, new_n29748_, new_n29749_, new_n29750_,
    new_n29751_, new_n29752_, new_n29753_, new_n29754_, new_n29755_,
    new_n29756_, new_n29757_, new_n29758_, new_n29759_, new_n29760_,
    new_n29761_, new_n29762_, new_n29763_, new_n29764_, new_n29765_,
    new_n29766_, new_n29767_, new_n29768_, new_n29769_, new_n29770_,
    new_n29771_, new_n29772_, new_n29773_, new_n29774_, new_n29775_,
    new_n29776_, new_n29777_, new_n29778_, new_n29779_, new_n29780_,
    new_n29781_, new_n29782_, new_n29783_, new_n29784_, new_n29785_,
    new_n29786_, new_n29787_, new_n29788_, new_n29789_, new_n29790_,
    new_n29791_, new_n29792_, new_n29793_, new_n29794_, new_n29795_,
    new_n29796_, new_n29797_, new_n29798_, new_n29799_, new_n29800_,
    new_n29801_, new_n29802_, new_n29803_, new_n29804_, new_n29805_,
    new_n29806_, new_n29807_, new_n29808_, new_n29809_, new_n29810_,
    new_n29811_, new_n29812_, new_n29813_, new_n29814_, new_n29815_,
    new_n29816_, new_n29817_, new_n29818_, new_n29819_, new_n29820_,
    new_n29821_, new_n29822_, new_n29823_, new_n29824_, new_n29825_,
    new_n29826_, new_n29827_, new_n29828_, new_n29829_, new_n29830_,
    new_n29831_, new_n29832_, new_n29833_, new_n29834_, new_n29835_,
    new_n29836_, new_n29837_, new_n29838_, new_n29839_, new_n29840_,
    new_n29841_, new_n29842_, new_n29843_, new_n29844_, new_n29845_,
    new_n29846_, new_n29847_, new_n29848_, new_n29849_, new_n29850_,
    new_n29851_, new_n29852_, new_n29853_, new_n29854_, new_n29855_,
    new_n29856_, new_n29857_, new_n29858_, new_n29859_, new_n29860_,
    new_n29861_, new_n29862_, new_n29863_, new_n29864_, new_n29865_,
    new_n29866_, new_n29867_, new_n29868_, new_n29869_, new_n29870_,
    new_n29871_, new_n29872_, new_n29873_, new_n29874_, new_n29875_,
    new_n29876_, new_n29877_, new_n29878_, new_n29879_, new_n29880_,
    new_n29881_, new_n29882_, new_n29883_, new_n29884_, new_n29885_,
    new_n29886_, new_n29887_, new_n29888_, new_n29889_, new_n29890_,
    new_n29891_, new_n29892_, new_n29893_, new_n29894_, new_n29895_,
    new_n29896_, new_n29897_, new_n29898_, new_n29899_, new_n29900_,
    new_n29901_, new_n29902_, new_n29903_, new_n29904_, new_n29905_,
    new_n29906_, new_n29907_, new_n29908_, new_n29909_, new_n29910_,
    new_n29911_, new_n29912_, new_n29913_, new_n29914_, new_n29915_,
    new_n29916_, new_n29917_, new_n29918_, new_n29919_, new_n29920_,
    new_n29921_, new_n29922_, new_n29923_, new_n29924_, new_n29925_,
    new_n29926_, new_n29927_, new_n29928_, new_n29929_, new_n29930_,
    new_n29931_, new_n29932_, new_n29933_, new_n29934_, new_n29935_,
    new_n29936_, new_n29937_, new_n29938_, new_n29939_, new_n29940_,
    new_n29941_, new_n29942_, new_n29943_, new_n29944_, new_n29945_,
    new_n29946_, new_n29947_, new_n29948_, new_n29949_, new_n29950_,
    new_n29951_, new_n29952_, new_n29953_, new_n29954_, new_n29955_,
    new_n29956_, new_n29957_, new_n29958_, new_n29959_, new_n29960_,
    new_n29961_, new_n29962_, new_n29963_, new_n29964_, new_n29965_,
    new_n29966_, new_n29967_, new_n29968_, new_n29969_, new_n29970_,
    new_n29971_, new_n29972_, new_n29973_, new_n29974_, new_n29975_,
    new_n29976_, new_n29977_, new_n29978_, new_n29979_, new_n29980_,
    new_n29981_, new_n29982_, new_n29983_, new_n29984_, new_n29985_,
    new_n29986_, new_n29987_, new_n29988_, new_n29989_, new_n29990_,
    new_n29991_, new_n29992_, new_n29993_, new_n29994_, new_n29995_,
    new_n29996_, new_n29997_, new_n29998_, new_n29999_, new_n30000_,
    new_n30001_, new_n30002_, new_n30003_, new_n30004_, new_n30005_,
    new_n30006_, new_n30007_, new_n30008_, new_n30009_, new_n30010_,
    new_n30011_, new_n30012_, new_n30013_, new_n30014_, new_n30015_,
    new_n30016_, new_n30017_, new_n30018_, new_n30019_, new_n30020_,
    new_n30021_, new_n30022_, new_n30023_, new_n30024_, new_n30025_,
    new_n30026_, new_n30027_, new_n30028_, new_n30029_, new_n30030_,
    new_n30031_, new_n30032_, new_n30033_, new_n30034_, new_n30035_,
    new_n30036_, new_n30037_, new_n30038_, new_n30039_, new_n30040_,
    new_n30041_, new_n30042_, new_n30043_, new_n30044_, new_n30045_,
    new_n30046_, new_n30047_, new_n30048_, new_n30049_, new_n30050_,
    new_n30051_, new_n30052_, new_n30053_, new_n30054_, new_n30055_,
    new_n30056_, new_n30057_, new_n30058_, new_n30059_, new_n30060_,
    new_n30061_, new_n30062_, new_n30063_, new_n30064_, new_n30065_,
    new_n30066_, new_n30067_, new_n30068_, new_n30069_, new_n30070_,
    new_n30071_, new_n30072_, new_n30073_, new_n30074_, new_n30075_,
    new_n30076_, new_n30077_, new_n30078_, new_n30079_, new_n30080_,
    new_n30081_, new_n30082_, new_n30083_, new_n30084_, new_n30085_,
    new_n30086_, new_n30087_, new_n30088_, new_n30089_, new_n30090_,
    new_n30091_, new_n30092_, new_n30093_, new_n30094_, new_n30095_,
    new_n30096_, new_n30097_, new_n30098_, new_n30099_, new_n30100_,
    new_n30101_, new_n30102_, new_n30103_, new_n30104_, new_n30105_,
    new_n30106_, new_n30107_, new_n30108_, new_n30109_, new_n30110_,
    new_n30111_, new_n30112_, new_n30113_, new_n30114_, new_n30115_,
    new_n30116_, new_n30117_, new_n30118_, new_n30119_, new_n30120_,
    new_n30121_, new_n30122_, new_n30123_, new_n30124_, new_n30125_,
    new_n30126_, new_n30127_, new_n30128_, new_n30129_, new_n30130_,
    new_n30131_, new_n30132_, new_n30133_, new_n30134_, new_n30135_,
    new_n30136_, new_n30137_, new_n30138_, new_n30139_, new_n30140_,
    new_n30141_, new_n30142_, new_n30143_, new_n30144_, new_n30145_,
    new_n30146_, new_n30147_, new_n30148_, new_n30149_, new_n30150_,
    new_n30151_, new_n30152_, new_n30153_, new_n30154_, new_n30155_,
    new_n30156_, new_n30157_, new_n30158_, new_n30159_, new_n30160_,
    new_n30161_, new_n30162_, new_n30163_, new_n30164_, new_n30165_,
    new_n30166_, new_n30167_, new_n30168_, new_n30169_, new_n30170_,
    new_n30171_, new_n30172_, new_n30173_, new_n30174_, new_n30175_,
    new_n30176_, new_n30177_, new_n30178_, new_n30179_, new_n30180_,
    new_n30181_, new_n30182_, new_n30183_, new_n30184_, new_n30185_,
    new_n30186_, new_n30187_, new_n30188_, new_n30189_, new_n30190_,
    new_n30191_, new_n30192_, new_n30193_, new_n30194_, new_n30195_,
    new_n30196_, new_n30197_, new_n30198_, new_n30199_, new_n30200_,
    new_n30201_, new_n30202_, new_n30203_, new_n30204_, new_n30205_,
    new_n30206_, new_n30207_, new_n30208_, new_n30209_, new_n30210_,
    new_n30211_, new_n30212_, new_n30213_, new_n30214_, new_n30215_,
    new_n30216_, new_n30217_, new_n30218_, new_n30219_, new_n30220_,
    new_n30221_, new_n30222_, new_n30223_, new_n30224_, new_n30225_,
    new_n30226_, new_n30227_, new_n30228_, new_n30229_, new_n30230_,
    new_n30231_, new_n30232_, new_n30233_, new_n30234_, new_n30235_,
    new_n30236_, new_n30237_, new_n30238_, new_n30239_, new_n30240_,
    new_n30241_, new_n30242_, new_n30243_, new_n30244_, new_n30245_,
    new_n30246_, new_n30247_, new_n30248_, new_n30249_, new_n30250_,
    new_n30251_, new_n30252_, new_n30253_, new_n30254_, new_n30255_,
    new_n30256_, new_n30257_, new_n30258_, new_n30259_, new_n30260_,
    new_n30261_, new_n30262_, new_n30263_, new_n30264_, new_n30265_,
    new_n30266_, new_n30267_, new_n30268_, new_n30269_, new_n30270_,
    new_n30271_, new_n30272_, new_n30273_, new_n30274_, new_n30275_,
    new_n30276_, new_n30277_, new_n30278_, new_n30279_, new_n30280_,
    new_n30281_, new_n30282_, new_n30283_, new_n30284_, new_n30285_,
    new_n30286_, new_n30287_, new_n30288_, new_n30289_, new_n30290_,
    new_n30291_, new_n30292_, new_n30293_, new_n30294_, new_n30295_,
    new_n30296_, new_n30297_, new_n30298_, new_n30299_, new_n30300_,
    new_n30301_, new_n30302_, new_n30303_, new_n30304_, new_n30305_,
    new_n30306_, new_n30307_, new_n30308_, new_n30309_, new_n30310_,
    new_n30311_, new_n30312_, new_n30313_, new_n30314_, new_n30315_,
    new_n30316_, new_n30317_, new_n30318_, new_n30319_, new_n30320_,
    new_n30321_, new_n30322_, new_n30323_, new_n30324_, new_n30325_,
    new_n30326_, new_n30327_, new_n30328_, new_n30329_, new_n30330_,
    new_n30331_, new_n30332_, new_n30333_, new_n30334_, new_n30335_,
    new_n30336_, new_n30337_, new_n30338_, new_n30339_, new_n30340_,
    new_n30341_, new_n30342_, new_n30343_, new_n30344_, new_n30345_,
    new_n30346_, new_n30347_, new_n30348_, new_n30349_, new_n30350_,
    new_n30351_, new_n30352_, new_n30353_, new_n30354_, new_n30355_,
    new_n30356_, new_n30357_, new_n30358_, new_n30359_, new_n30360_,
    new_n30361_, new_n30362_, new_n30363_, new_n30364_, new_n30365_,
    new_n30366_, new_n30367_, new_n30368_, new_n30369_, new_n30370_,
    new_n30371_, new_n30372_, new_n30373_, new_n30374_, new_n30375_,
    new_n30376_, new_n30377_, new_n30378_, new_n30379_, new_n30380_,
    new_n30381_, new_n30382_, new_n30383_, new_n30384_, new_n30385_,
    new_n30386_, new_n30387_, new_n30388_, new_n30389_, new_n30390_,
    new_n30391_, new_n30392_, new_n30393_, new_n30394_, new_n30395_,
    new_n30396_, new_n30397_, new_n30398_, new_n30399_, new_n30400_,
    new_n30401_, new_n30402_, new_n30403_, new_n30404_, new_n30405_,
    new_n30406_, new_n30407_, new_n30408_, new_n30409_, new_n30410_,
    new_n30411_, new_n30412_, new_n30413_, new_n30414_, new_n30415_,
    new_n30416_, new_n30417_, new_n30418_, new_n30419_, new_n30420_,
    new_n30421_, new_n30422_, new_n30423_, new_n30424_, new_n30425_,
    new_n30426_, new_n30427_, new_n30428_, new_n30429_, new_n30430_,
    new_n30431_, new_n30432_, new_n30433_, new_n30434_, new_n30435_,
    new_n30436_, new_n30437_, new_n30438_, new_n30439_, new_n30440_,
    new_n30441_, new_n30442_, new_n30443_, new_n30444_, new_n30445_,
    new_n30446_, new_n30447_, new_n30448_, new_n30449_, new_n30450_,
    new_n30451_, new_n30452_, new_n30453_, new_n30454_, new_n30455_,
    new_n30456_, new_n30457_, new_n30458_, new_n30459_, new_n30460_,
    new_n30461_, new_n30462_, new_n30463_, new_n30464_, new_n30465_,
    new_n30466_, new_n30467_, new_n30468_, new_n30469_, new_n30470_,
    new_n30471_, new_n30472_, new_n30473_, new_n30474_, new_n30475_,
    new_n30476_, new_n30477_, new_n30478_, new_n30479_, new_n30480_,
    new_n30481_, new_n30482_, new_n30483_, new_n30484_, new_n30485_,
    new_n30486_, new_n30487_, new_n30488_, new_n30489_, new_n30490_,
    new_n30491_, new_n30492_, new_n30493_, new_n30494_, new_n30495_,
    new_n30496_, new_n30497_, new_n30498_, new_n30499_, new_n30500_,
    new_n30501_, new_n30502_, new_n30503_, new_n30504_, new_n30505_,
    new_n30506_, new_n30507_, new_n30508_, new_n30509_, new_n30510_,
    new_n30511_, new_n30512_, new_n30513_, new_n30514_, new_n30515_,
    new_n30516_, new_n30517_, new_n30518_, new_n30519_, new_n30520_,
    new_n30521_, new_n30522_, new_n30523_, new_n30524_, new_n30525_,
    new_n30526_, new_n30527_, new_n30528_, new_n30529_, new_n30530_,
    new_n30531_, new_n30532_, new_n30533_, new_n30534_, new_n30535_,
    new_n30536_, new_n30537_, new_n30538_, new_n30539_, new_n30540_,
    new_n30541_, new_n30542_, new_n30543_, new_n30544_, new_n30545_,
    new_n30546_, new_n30547_, new_n30548_, new_n30549_, new_n30550_,
    new_n30551_, new_n30552_, new_n30553_, new_n30554_, new_n30555_,
    new_n30556_, new_n30557_, new_n30558_, new_n30559_, new_n30560_,
    new_n30561_, new_n30562_, new_n30563_, new_n30564_, new_n30565_,
    new_n30566_, new_n30567_, new_n30568_, new_n30569_, new_n30570_,
    new_n30571_, new_n30572_, new_n30573_, new_n30574_, new_n30575_,
    new_n30576_, new_n30577_, new_n30578_, new_n30579_, new_n30580_,
    new_n30581_, new_n30582_, new_n30583_, new_n30584_, new_n30585_,
    new_n30586_, new_n30587_, new_n30588_, new_n30589_, new_n30590_,
    new_n30591_, new_n30592_, new_n30593_, new_n30594_, new_n30595_,
    new_n30596_, new_n30597_, new_n30598_, new_n30599_, new_n30600_,
    new_n30601_, new_n30602_, new_n30603_, new_n30604_, new_n30605_,
    new_n30606_, new_n30607_, new_n30608_, new_n30609_, new_n30610_,
    new_n30611_, new_n30612_, new_n30613_, new_n30614_, new_n30615_,
    new_n30616_, new_n30617_, new_n30618_, new_n30619_, new_n30620_,
    new_n30621_, new_n30622_, new_n30623_, new_n30624_, new_n30625_,
    new_n30626_, new_n30627_, new_n30628_, new_n30629_, new_n30630_,
    new_n30631_, new_n30632_, new_n30633_, new_n30634_, new_n30635_,
    new_n30636_, new_n30637_, new_n30638_, new_n30639_, new_n30640_,
    new_n30641_, new_n30642_, new_n30643_, new_n30644_, new_n30645_,
    new_n30646_, new_n30647_, new_n30648_, new_n30649_, new_n30650_,
    new_n30651_, new_n30652_, new_n30653_, new_n30654_, new_n30655_,
    new_n30656_, new_n30657_, new_n30658_, new_n30659_, new_n30660_,
    new_n30661_, new_n30662_, new_n30663_, new_n30664_, new_n30665_,
    new_n30666_, new_n30667_, new_n30668_, new_n30669_, new_n30670_,
    new_n30671_, new_n30672_, new_n30673_, new_n30674_, new_n30675_,
    new_n30676_, new_n30677_, new_n30678_, new_n30679_, new_n30680_,
    new_n30681_, new_n30682_, new_n30683_, new_n30684_, new_n30685_,
    new_n30686_, new_n30687_;
  assign new_n1526_ = ~new_n8765_ | ~new_n30288_;
  assign new_n1527_ = ~new_n8454_ | ~new_n30287_;
  assign new_n1528_ = ~new_n8797_ | ~new_n30320_;
  assign po021 = pi767 | new_n1661_;
  assign po020 = pi766 | new_n1664_;
  assign new_n1531_ = ~new_n1674_ | ~new_n1673_;
  assign new_n1532_ = ~new_n1676_ | ~new_n1675_;
  assign new_n1533_ = ~new_n1678_ | ~new_n1677_;
  assign new_n1534_ = ~new_n1680_ | ~new_n1679_;
  assign new_n1535_ = ~new_n1682_ | ~new_n1681_;
  assign new_n1536_ = ~new_n1684_ | ~new_n1683_;
  assign new_n1537_ = ~new_n1686_ | ~new_n1685_;
  assign new_n1538_ = ~new_n1688_ | ~new_n1687_;
  assign new_n1539_ = ~new_n1690_ | ~new_n1689_;
  assign new_n1540_ = ~new_n1692_ | ~new_n1691_;
  assign new_n1541_ = ~new_n1694_ | ~new_n1693_;
  assign new_n1542_ = ~new_n1696_ | ~new_n1695_;
  assign new_n1543_ = ~new_n1698_ | ~new_n1697_;
  assign new_n1544_ = ~new_n1700_ | ~new_n1699_;
  assign new_n1545_ = ~new_n1702_ | ~new_n1701_;
  assign new_n1546_ = ~new_n1704_ | ~new_n1703_;
  assign new_n1547_ = ~new_n1706_ | ~new_n1705_;
  assign new_n1548_ = ~new_n1708_ | ~new_n1707_;
  assign new_n1549_ = ~new_n1710_ | ~new_n1709_;
  assign new_n1550_ = ~new_n1712_ | ~new_n1711_;
  assign new_n1551_ = ~new_n1714_ | ~new_n1713_;
  assign new_n1552_ = ~new_n1716_ | ~new_n1715_;
  assign new_n1553_ = ~new_n1718_ | ~new_n1717_;
  assign new_n1554_ = ~new_n1720_ | ~new_n1719_;
  assign new_n1555_ = ~new_n1722_ | ~new_n1721_;
  assign new_n1556_ = ~new_n1724_ | ~new_n1723_;
  assign new_n1557_ = ~new_n1726_ | ~new_n1725_;
  assign new_n1558_ = ~new_n1728_ | ~new_n1727_;
  assign new_n1559_ = ~new_n1730_ | ~new_n1729_;
  assign new_n1560_ = ~new_n1732_ | ~new_n1731_;
  assign new_n1561_ = ~new_n1734_ | ~new_n1733_;
  assign new_n1562_ = ~new_n1736_ | ~new_n1735_;
  assign new_n1563_ = ~new_n1738_ | ~new_n1737_;
  assign new_n1564_ = ~new_n1740_ | ~new_n1739_;
  assign new_n1565_ = ~new_n1742_ | ~new_n1741_;
  assign new_n1566_ = ~new_n1744_ | ~new_n1743_;
  assign new_n1567_ = ~new_n1746_ | ~new_n1745_;
  assign new_n1568_ = ~new_n1748_ | ~new_n1747_;
  assign new_n1569_ = ~new_n1750_ | ~new_n1749_;
  assign new_n1570_ = ~new_n1752_ | ~new_n1751_;
  assign new_n1571_ = ~new_n1754_ | ~new_n1753_;
  assign new_n1572_ = ~new_n1756_ | ~new_n1755_;
  assign new_n1573_ = ~new_n1758_ | ~new_n1757_;
  assign new_n1574_ = ~new_n1760_ | ~new_n1759_;
  assign new_n1575_ = ~new_n1762_ | ~new_n1761_;
  assign new_n1576_ = ~new_n1764_ | ~new_n1763_;
  assign new_n1577_ = ~new_n1766_ | ~new_n1765_;
  assign new_n1578_ = ~new_n1768_ | ~new_n1767_;
  assign new_n1579_ = ~new_n1770_ | ~new_n1769_;
  assign new_n1580_ = ~new_n1772_ | ~new_n1771_;
  assign new_n1581_ = ~new_n1774_ | ~new_n1773_;
  assign new_n1582_ = ~new_n1776_ | ~new_n1775_;
  assign new_n1583_ = ~new_n1778_ | ~new_n1777_;
  assign new_n1584_ = ~new_n1780_ | ~new_n1779_;
  assign new_n1585_ = ~new_n1782_ | ~new_n1781_;
  assign new_n1586_ = ~new_n1784_ | ~new_n1783_;
  assign new_n1587_ = ~new_n1786_ | ~new_n1785_;
  assign new_n1588_ = ~new_n1788_ | ~new_n1787_;
  assign new_n1589_ = ~new_n1790_ | ~new_n1789_;
  assign new_n1590_ = ~new_n1792_ | ~new_n1791_;
  assign new_n1591_ = ~new_n1794_ | ~new_n1793_;
  assign new_n1592_ = ~new_n1796_ | ~new_n1795_;
  assign new_n1593_ = ~new_n1798_ | ~new_n1797_;
  assign new_n1594_ = ~new_n1800_ | ~new_n1799_;
  assign new_n1595_ = ~new_n1802_ | ~new_n1801_;
  assign new_n1596_ = ~new_n1804_ | ~new_n1803_;
  assign new_n1597_ = ~new_n1806_ | ~new_n1805_;
  assign new_n1598_ = ~new_n1808_ | ~new_n1807_;
  assign new_n1599_ = ~new_n1810_ | ~new_n1809_;
  assign new_n1600_ = ~new_n1812_ | ~new_n1811_;
  assign new_n1601_ = ~new_n1814_ | ~new_n1813_;
  assign new_n1602_ = ~new_n1816_ | ~new_n1815_;
  assign new_n1603_ = ~new_n1818_ | ~new_n1817_;
  assign new_n1604_ = ~new_n1820_ | ~new_n1819_;
  assign new_n1605_ = ~new_n1822_ | ~new_n1821_;
  assign new_n1606_ = ~new_n1824_ | ~new_n1823_;
  assign new_n1607_ = ~new_n1826_ | ~new_n1825_;
  assign new_n1608_ = ~new_n1828_ | ~new_n1827_;
  assign new_n1609_ = ~new_n1830_ | ~new_n1829_;
  assign new_n1610_ = ~new_n1832_ | ~new_n1831_;
  assign new_n1611_ = ~new_n1834_ | ~new_n1833_;
  assign new_n1612_ = ~new_n1836_ | ~new_n1835_;
  assign new_n1613_ = ~new_n1838_ | ~new_n1837_;
  assign new_n1614_ = ~new_n1840_ | ~new_n1839_;
  assign new_n1615_ = ~new_n1842_ | ~new_n1841_;
  assign new_n1616_ = ~new_n1844_ | ~new_n1843_;
  assign new_n1617_ = ~new_n1846_ | ~new_n1845_;
  assign new_n1618_ = ~new_n1848_ | ~new_n1847_;
  assign new_n1619_ = ~new_n1850_ | ~new_n1849_;
  assign new_n1620_ = ~new_n1852_ | ~new_n1851_;
  assign new_n1621_ = ~new_n1854_ | ~new_n1853_;
  assign new_n1622_ = ~new_n1856_ | ~new_n1855_;
  assign new_n1623_ = ~new_n1858_ | ~new_n1857_;
  assign new_n1624_ = ~new_n1860_ | ~new_n1859_;
  assign new_n1625_ = ~new_n1862_ | ~new_n1861_;
  assign new_n1626_ = ~new_n1864_ | ~new_n1863_;
  assign new_n1627_ = ~new_n1866_ | ~new_n1865_;
  assign new_n1628_ = ~new_n1868_ | ~new_n1867_;
  assign new_n1629_ = ~new_n1870_ | ~new_n1869_;
  assign new_n1630_ = ~new_n1872_ | ~new_n1871_;
  assign new_n1631_ = ~new_n1874_ | ~new_n1873_;
  assign new_n1632_ = ~new_n1876_ | ~new_n1875_;
  assign new_n1633_ = ~new_n1878_ | ~new_n1877_;
  assign new_n1634_ = ~new_n1880_ | ~new_n1879_;
  assign new_n1635_ = ~new_n1882_ | ~new_n1881_;
  assign new_n1636_ = ~new_n1884_ | ~new_n1883_;
  assign new_n1637_ = ~new_n1886_ | ~new_n1885_;
  assign new_n1638_ = ~new_n1888_ | ~new_n1887_;
  assign new_n1639_ = ~new_n1890_ | ~new_n1889_;
  assign new_n1640_ = ~new_n1892_ | ~new_n1891_;
  assign new_n1641_ = ~new_n1894_ | ~new_n1893_;
  assign new_n1642_ = ~new_n1896_ | ~new_n1895_;
  assign new_n1643_ = ~new_n1898_ | ~new_n1897_;
  assign new_n1644_ = ~new_n1900_ | ~new_n1899_;
  assign new_n1645_ = ~new_n1902_ | ~new_n1901_;
  assign new_n1646_ = ~new_n1904_ | ~new_n1903_;
  assign new_n1647_ = ~new_n1906_ | ~new_n1905_;
  assign new_n1648_ = ~new_n1908_ | ~new_n1907_;
  assign new_n1649_ = ~new_n1910_ | ~new_n1909_;
  assign new_n1650_ = ~new_n1912_ | ~new_n1911_;
  assign new_n1651_ = ~new_n1914_ | ~new_n1913_;
  assign new_n1652_ = ~new_n1916_ | ~new_n1915_;
  assign new_n1653_ = ~new_n1918_ | ~new_n1917_;
  assign new_n1654_ = ~new_n1920_ | ~new_n1919_;
  assign new_n1655_ = ~new_n1922_ | ~new_n1921_;
  assign new_n1656_ = ~new_n1924_ | ~new_n1923_;
  assign new_n1657_ = ~new_n1926_ | ~new_n1925_;
  assign new_n1658_ = ~new_n1928_ | ~new_n1927_;
  assign new_n1659_ = ~pi522;
  assign new_n1660_ = ~pi277;
  assign new_n1661_ = new_n1670_ & new_n1669_;
  assign new_n1662_ = ~pi521;
  assign new_n1663_ = ~pi276;
  assign new_n1664_ = new_n1672_ & new_n1671_;
  assign new_n1665_ = ~new_n1667_ | ~new_n1666_;
  assign new_n1666_ = ~pi438 | ~new_n1662_ | ~new_n12472_ | ~pi193;
  assign new_n1667_ = ~new_n13031_ | ~new_n1663_ | ~pi683 | ~new_n12473_;
  assign new_n1668_ = ~new_n1665_;
  assign new_n1669_ = ~pi522 | ~new_n1660_;
  assign new_n1670_ = ~pi277 | ~new_n1659_;
  assign new_n1671_ = ~pi521 | ~new_n1663_;
  assign new_n1672_ = ~pi276 | ~new_n1662_;
  assign new_n1673_ = ~new_n11519_ | ~new_n1665_;
  assign new_n1674_ = ~pi023 | ~new_n1668_;
  assign new_n1675_ = ~new_n11520_ | ~new_n1665_;
  assign new_n1676_ = ~pi024 | ~new_n1668_;
  assign new_n1677_ = ~new_n11521_ | ~new_n1665_;
  assign new_n1678_ = ~pi025 | ~new_n1668_;
  assign new_n1679_ = ~new_n11522_ | ~new_n1665_;
  assign new_n1680_ = ~pi026 | ~new_n1668_;
  assign new_n1681_ = ~new_n11523_ | ~new_n1665_;
  assign new_n1682_ = ~pi027 | ~new_n1668_;
  assign new_n1683_ = ~new_n11524_ | ~new_n1665_;
  assign new_n1684_ = ~pi028 | ~new_n1668_;
  assign new_n1685_ = ~new_n11525_ | ~new_n1665_;
  assign new_n1686_ = ~pi029 | ~new_n1668_;
  assign new_n1687_ = ~new_n11452_ | ~new_n1665_;
  assign new_n1688_ = ~pi001 | ~new_n1668_;
  assign new_n1689_ = ~new_n11526_ | ~new_n1665_;
  assign new_n1690_ = ~pi002 | ~new_n1668_;
  assign new_n1691_ = ~new_n11527_ | ~new_n1665_;
  assign new_n1692_ = ~pi030 | ~new_n1668_;
  assign new_n1693_ = ~new_n11528_ | ~new_n1665_;
  assign new_n1694_ = ~pi003 | ~new_n1668_;
  assign new_n1695_ = ~new_n11529_ | ~new_n1665_;
  assign new_n1696_ = ~pi004 | ~new_n1668_;
  assign new_n1697_ = ~new_n11530_ | ~new_n1665_;
  assign new_n1698_ = ~pi005 | ~new_n1668_;
  assign new_n1699_ = ~new_n11531_ | ~new_n1665_;
  assign new_n1700_ = ~pi006 | ~new_n1668_;
  assign new_n1701_ = ~new_n11532_ | ~new_n1665_;
  assign new_n1702_ = ~pi007 | ~new_n1668_;
  assign new_n1703_ = ~new_n11533_ | ~new_n1665_;
  assign new_n1704_ = ~pi008 | ~new_n1668_;
  assign new_n1705_ = ~new_n11534_ | ~new_n1665_;
  assign new_n1706_ = ~pi009 | ~new_n1668_;
  assign new_n1707_ = ~new_n11535_ | ~new_n1665_;
  assign new_n1708_ = ~pi010 | ~new_n1668_;
  assign new_n1709_ = ~new_n11536_ | ~new_n1665_;
  assign new_n1710_ = ~pi011 | ~new_n1668_;
  assign new_n1711_ = ~new_n11537_ | ~new_n1665_;
  assign new_n1712_ = ~pi012 | ~new_n1668_;
  assign new_n1713_ = ~new_n11538_ | ~new_n1665_;
  assign new_n1714_ = ~pi031 | ~new_n1668_;
  assign new_n1715_ = ~new_n11539_ | ~new_n1665_;
  assign new_n1716_ = ~pi013 | ~new_n1668_;
  assign new_n1717_ = ~new_n11540_ | ~new_n1665_;
  assign new_n1718_ = ~pi014 | ~new_n1668_;
  assign new_n1719_ = ~new_n11541_ | ~new_n1665_;
  assign new_n1720_ = ~pi015 | ~new_n1668_;
  assign new_n1721_ = ~new_n11542_ | ~new_n1665_;
  assign new_n1722_ = ~pi016 | ~new_n1668_;
  assign new_n1723_ = ~new_n11543_ | ~new_n1665_;
  assign new_n1724_ = ~pi017 | ~new_n1668_;
  assign new_n1725_ = ~new_n11544_ | ~new_n1665_;
  assign new_n1726_ = ~pi018 | ~new_n1668_;
  assign new_n1727_ = ~new_n11545_ | ~new_n1665_;
  assign new_n1728_ = ~pi019 | ~new_n1668_;
  assign new_n1729_ = ~new_n11546_ | ~new_n1665_;
  assign new_n1730_ = ~pi020 | ~new_n1668_;
  assign new_n1731_ = ~new_n11547_ | ~new_n1665_;
  assign new_n1732_ = ~pi021 | ~new_n1668_;
  assign new_n1733_ = ~new_n11548_ | ~new_n1665_;
  assign new_n1734_ = ~pi022 | ~new_n1668_;
  assign new_n1735_ = ~new_n11453_ | ~new_n1665_;
  assign new_n1736_ = ~pi032 | ~new_n1668_;
  assign new_n1737_ = ~pi222 | ~new_n1665_;
  assign new_n1738_ = ~new_n12002_ | ~new_n1668_;
  assign new_n1739_ = ~pi221 | ~new_n1665_;
  assign new_n1740_ = ~new_n12003_ | ~new_n1668_;
  assign new_n1741_ = ~pi220 | ~new_n1665_;
  assign new_n1742_ = ~new_n12004_ | ~new_n1668_;
  assign new_n1743_ = ~pi219 | ~new_n1665_;
  assign new_n1744_ = ~new_n12005_ | ~new_n1668_;
  assign new_n1745_ = ~pi218 | ~new_n1665_;
  assign new_n1746_ = ~new_n12006_ | ~new_n1668_;
  assign new_n1747_ = ~pi217 | ~new_n1665_;
  assign new_n1748_ = ~new_n12007_ | ~new_n1668_;
  assign new_n1749_ = ~pi216 | ~new_n1665_;
  assign new_n1750_ = ~new_n12008_ | ~new_n1668_;
  assign new_n1751_ = ~pi244 | ~new_n1665_;
  assign new_n1752_ = ~new_n11929_ | ~new_n1668_;
  assign new_n1753_ = ~pi243 | ~new_n1665_;
  assign new_n1754_ = ~new_n12009_ | ~new_n1668_;
  assign new_n1755_ = ~pi215 | ~new_n1665_;
  assign new_n1756_ = ~new_n12010_ | ~new_n1668_;
  assign new_n1757_ = ~pi242 | ~new_n1665_;
  assign new_n1758_ = ~new_n12011_ | ~new_n1668_;
  assign new_n1759_ = ~pi241 | ~new_n1665_;
  assign new_n1760_ = ~new_n12012_ | ~new_n1668_;
  assign new_n1761_ = ~pi240 | ~new_n1665_;
  assign new_n1762_ = ~new_n12013_ | ~new_n1668_;
  assign new_n1763_ = ~pi239 | ~new_n1665_;
  assign new_n1764_ = ~new_n12014_ | ~new_n1668_;
  assign new_n1765_ = ~pi238 | ~new_n1665_;
  assign new_n1766_ = ~new_n12015_ | ~new_n1668_;
  assign new_n1767_ = ~pi237 | ~new_n1665_;
  assign new_n1768_ = ~new_n12016_ | ~new_n1668_;
  assign new_n1769_ = ~pi236 | ~new_n1665_;
  assign new_n1770_ = ~new_n12017_ | ~new_n1668_;
  assign new_n1771_ = ~pi235 | ~new_n1665_;
  assign new_n1772_ = ~new_n12018_ | ~new_n1668_;
  assign new_n1773_ = ~pi234 | ~new_n1665_;
  assign new_n1774_ = ~new_n12019_ | ~new_n1668_;
  assign new_n1775_ = ~pi233 | ~new_n1665_;
  assign new_n1776_ = ~new_n12020_ | ~new_n1668_;
  assign new_n1777_ = ~pi214 | ~new_n1665_;
  assign new_n1778_ = ~new_n11930_ | ~new_n1668_;
  assign new_n1779_ = ~pi232 | ~new_n1665_;
  assign new_n1780_ = ~new_n12021_ | ~new_n1668_;
  assign new_n1781_ = ~pi231 | ~new_n1665_;
  assign new_n1782_ = ~new_n12022_ | ~new_n1668_;
  assign new_n1783_ = ~pi230 | ~new_n1665_;
  assign new_n1784_ = ~new_n12023_ | ~new_n1668_;
  assign new_n1785_ = ~pi229 | ~new_n1665_;
  assign new_n1786_ = ~new_n12024_ | ~new_n1668_;
  assign new_n1787_ = ~pi228 | ~new_n1665_;
  assign new_n1788_ = ~new_n12025_ | ~new_n1668_;
  assign new_n1789_ = ~pi227 | ~new_n1665_;
  assign new_n1790_ = ~new_n12026_ | ~new_n1668_;
  assign new_n1791_ = ~pi226 | ~new_n1665_;
  assign new_n1792_ = ~new_n12027_ | ~new_n1668_;
  assign new_n1793_ = ~pi225 | ~new_n1665_;
  assign new_n1794_ = ~new_n12028_ | ~new_n1668_;
  assign new_n1795_ = ~pi224 | ~new_n1665_;
  assign new_n1796_ = ~new_n12029_ | ~new_n1668_;
  assign new_n1797_ = ~pi223 | ~new_n1665_;
  assign new_n1798_ = ~new_n12030_ | ~new_n1668_;
  assign new_n1799_ = ~pi213 | ~new_n1665_;
  assign new_n1800_ = ~new_n12001_ | ~new_n1668_;
  assign new_n1801_ = ~new_n12002_ | ~new_n1665_;
  assign new_n1802_ = ~pi467 | ~new_n1668_;
  assign new_n1803_ = ~new_n12003_ | ~new_n1665_;
  assign new_n1804_ = ~pi466 | ~new_n1668_;
  assign new_n1805_ = ~new_n12004_ | ~new_n1665_;
  assign new_n1806_ = ~pi465 | ~new_n1668_;
  assign new_n1807_ = ~new_n12005_ | ~new_n1665_;
  assign new_n1808_ = ~pi464 | ~new_n1668_;
  assign new_n1809_ = ~new_n12006_ | ~new_n1665_;
  assign new_n1810_ = ~pi463 | ~new_n1668_;
  assign new_n1811_ = ~new_n12007_ | ~new_n1665_;
  assign new_n1812_ = ~pi462 | ~new_n1668_;
  assign new_n1813_ = ~new_n12008_ | ~new_n1665_;
  assign new_n1814_ = ~pi461 | ~new_n1668_;
  assign new_n1815_ = ~new_n11929_ | ~new_n1665_;
  assign new_n1816_ = ~pi489 | ~new_n1668_;
  assign new_n1817_ = ~new_n12009_ | ~new_n1665_;
  assign new_n1818_ = ~pi488 | ~new_n1668_;
  assign new_n1819_ = ~new_n12010_ | ~new_n1665_;
  assign new_n1820_ = ~pi460 | ~new_n1668_;
  assign new_n1821_ = ~new_n12011_ | ~new_n1665_;
  assign new_n1822_ = ~pi487 | ~new_n1668_;
  assign new_n1823_ = ~new_n12012_ | ~new_n1665_;
  assign new_n1824_ = ~pi486 | ~new_n1668_;
  assign new_n1825_ = ~new_n12013_ | ~new_n1665_;
  assign new_n1826_ = ~pi485 | ~new_n1668_;
  assign new_n1827_ = ~new_n12014_ | ~new_n1665_;
  assign new_n1828_ = ~pi484 | ~new_n1668_;
  assign new_n1829_ = ~new_n12015_ | ~new_n1665_;
  assign new_n1830_ = ~pi483 | ~new_n1668_;
  assign new_n1831_ = ~new_n12016_ | ~new_n1665_;
  assign new_n1832_ = ~pi482 | ~new_n1668_;
  assign new_n1833_ = ~new_n12017_ | ~new_n1665_;
  assign new_n1834_ = ~pi481 | ~new_n1668_;
  assign new_n1835_ = ~new_n12018_ | ~new_n1665_;
  assign new_n1836_ = ~pi480 | ~new_n1668_;
  assign new_n1837_ = ~new_n12019_ | ~new_n1665_;
  assign new_n1838_ = ~pi479 | ~new_n1668_;
  assign new_n1839_ = ~new_n12020_ | ~new_n1665_;
  assign new_n1840_ = ~pi478 | ~new_n1668_;
  assign new_n1841_ = ~new_n11930_ | ~new_n1665_;
  assign new_n1842_ = ~pi459 | ~new_n1668_;
  assign new_n1843_ = ~new_n12021_ | ~new_n1665_;
  assign new_n1844_ = ~pi477 | ~new_n1668_;
  assign new_n1845_ = ~new_n12022_ | ~new_n1665_;
  assign new_n1846_ = ~pi476 | ~new_n1668_;
  assign new_n1847_ = ~new_n12023_ | ~new_n1665_;
  assign new_n1848_ = ~pi475 | ~new_n1668_;
  assign new_n1849_ = ~new_n12024_ | ~new_n1665_;
  assign new_n1850_ = ~pi474 | ~new_n1668_;
  assign new_n1851_ = ~new_n12025_ | ~new_n1665_;
  assign new_n1852_ = ~pi473 | ~new_n1668_;
  assign new_n1853_ = ~new_n12026_ | ~new_n1665_;
  assign new_n1854_ = ~pi472 | ~new_n1668_;
  assign new_n1855_ = ~new_n12027_ | ~new_n1665_;
  assign new_n1856_ = ~pi471 | ~new_n1668_;
  assign new_n1857_ = ~new_n12028_ | ~new_n1665_;
  assign new_n1858_ = ~pi470 | ~new_n1668_;
  assign new_n1859_ = ~new_n12029_ | ~new_n1665_;
  assign new_n1860_ = ~pi469 | ~new_n1668_;
  assign new_n1861_ = ~new_n12030_ | ~new_n1665_;
  assign new_n1862_ = ~pi468 | ~new_n1668_;
  assign new_n1863_ = ~new_n12001_ | ~new_n1665_;
  assign new_n1864_ = ~pi458 | ~new_n1668_;
  assign new_n1865_ = ~pi467 | ~new_n1665_;
  assign new_n1866_ = ~pi222 | ~new_n1668_;
  assign new_n1867_ = ~pi466 | ~new_n1665_;
  assign new_n1868_ = ~pi221 | ~new_n1668_;
  assign new_n1869_ = ~pi465 | ~new_n1665_;
  assign new_n1870_ = ~pi220 | ~new_n1668_;
  assign new_n1871_ = ~pi464 | ~new_n1665_;
  assign new_n1872_ = ~pi219 | ~new_n1668_;
  assign new_n1873_ = ~pi463 | ~new_n1665_;
  assign new_n1874_ = ~pi218 | ~new_n1668_;
  assign new_n1875_ = ~pi462 | ~new_n1665_;
  assign new_n1876_ = ~pi217 | ~new_n1668_;
  assign new_n1877_ = ~pi489 | ~new_n1665_;
  assign new_n1878_ = ~pi244 | ~new_n1668_;
  assign new_n1879_ = ~pi488 | ~new_n1665_;
  assign new_n1880_ = ~pi243 | ~new_n1668_;
  assign new_n1881_ = ~pi461 | ~new_n1665_;
  assign new_n1882_ = ~pi216 | ~new_n1668_;
  assign new_n1883_ = ~pi487 | ~new_n1665_;
  assign new_n1884_ = ~pi242 | ~new_n1668_;
  assign new_n1885_ = ~pi486 | ~new_n1665_;
  assign new_n1886_ = ~pi241 | ~new_n1668_;
  assign new_n1887_ = ~pi485 | ~new_n1665_;
  assign new_n1888_ = ~pi240 | ~new_n1668_;
  assign new_n1889_ = ~pi484 | ~new_n1665_;
  assign new_n1890_ = ~pi239 | ~new_n1668_;
  assign new_n1891_ = ~pi483 | ~new_n1665_;
  assign new_n1892_ = ~pi238 | ~new_n1668_;
  assign new_n1893_ = ~pi482 | ~new_n1665_;
  assign new_n1894_ = ~pi237 | ~new_n1668_;
  assign new_n1895_ = ~pi481 | ~new_n1665_;
  assign new_n1896_ = ~pi236 | ~new_n1668_;
  assign new_n1897_ = ~pi480 | ~new_n1665_;
  assign new_n1898_ = ~pi235 | ~new_n1668_;
  assign new_n1899_ = ~pi479 | ~new_n1665_;
  assign new_n1900_ = ~pi234 | ~new_n1668_;
  assign new_n1901_ = ~pi478 | ~new_n1665_;
  assign new_n1902_ = ~pi233 | ~new_n1668_;
  assign new_n1903_ = ~pi460 | ~new_n1665_;
  assign new_n1904_ = ~pi215 | ~new_n1668_;
  assign new_n1905_ = ~pi477 | ~new_n1665_;
  assign new_n1906_ = ~pi232 | ~new_n1668_;
  assign new_n1907_ = ~pi476 | ~new_n1665_;
  assign new_n1908_ = ~pi231 | ~new_n1668_;
  assign new_n1909_ = ~pi475 | ~new_n1665_;
  assign new_n1910_ = ~pi230 | ~new_n1668_;
  assign new_n1911_ = ~pi474 | ~new_n1665_;
  assign new_n1912_ = ~pi229 | ~new_n1668_;
  assign new_n1913_ = ~pi473 | ~new_n1665_;
  assign new_n1914_ = ~pi228 | ~new_n1668_;
  assign new_n1915_ = ~pi472 | ~new_n1665_;
  assign new_n1916_ = ~pi227 | ~new_n1668_;
  assign new_n1917_ = ~pi471 | ~new_n1665_;
  assign new_n1918_ = ~pi226 | ~new_n1668_;
  assign new_n1919_ = ~pi470 | ~new_n1665_;
  assign new_n1920_ = ~pi225 | ~new_n1668_;
  assign new_n1921_ = ~pi469 | ~new_n1665_;
  assign new_n1922_ = ~pi224 | ~new_n1668_;
  assign new_n1923_ = ~pi468 | ~new_n1665_;
  assign new_n1924_ = ~pi223 | ~new_n1668_;
  assign new_n1925_ = ~pi459 | ~new_n1665_;
  assign new_n1926_ = ~pi214 | ~new_n1668_;
  assign new_n1927_ = ~pi458 | ~new_n1665_;
  assign new_n1928_ = ~pi213 | ~new_n1668_;
  assign new_n1929_ = ~new_n8439_ | ~new_n30319_;
  assign new_n1930_ = ~new_n30502_ | ~new_n1932_;
  assign new_n1931_ = ~new_n30621_ | ~new_n30425_;
  assign new_n1932_ = ~new_n1933_ | ~new_n1934_;
  assign new_n1933_ = ~new_n8800_ | ~new_n30325_;
  assign new_n1934_ = ~new_n8440_ | ~new_n30324_;
  assign new_n1935_ = ~new_n1937_ | ~new_n30596_;
  assign new_n1936_ = ~new_n30620_ | ~new_n30351_;
  assign new_n1937_ = ~new_n1938_ | ~new_n1939_;
  assign new_n1938_ = ~new_n8803_ | ~new_n30323_;
  assign new_n1939_ = ~new_n8449_ | ~new_n30322_;
  assign new_n1940_ = ~new_n8806_ | ~new_n30328_;
  assign new_n1941_ = new_n2929_ & new_n2378_;
  assign new_n1942_ = new_n2382_ & new_n2376_;
  assign new_n1943_ = new_n2532_ & new_n2527_;
  assign new_n1944_ = new_n2374_ & new_n2375_;
  assign new_n1945_ = new_n4735_ & new_n2374_;
  assign new_n1946_ = new_n4732_ & new_n2375_;
  assign new_n1947_ = new_n4732_ & new_n4735_;
  assign new_n1948_ = new_n4339_ & new_n2352_;
  assign new_n1949_ = new_n2519_ & new_n2352_;
  assign new_n1950_ = new_n2970_ & new_n2355_;
  assign new_n1951_ = new_n1975_ & new_n4720_;
  assign new_n1952_ = new_n2957_ & new_n4738_;
  assign new_n1953_ = new_n2778_ & new_n2942_;
  assign new_n1954_ = new_n15358_ & new_n2364_;
  assign new_n1955_ = new_n15358_ & new_n2367_;
  assign new_n1956_ = new_n2284_ & pi275;
  assign new_n1957_ = new_n2935_ & new_n2958_;
  assign new_n1958_ = new_n2958_ & new_n2353_;
  assign new_n1959_ = new_n2930_ & new_n2958_;
  assign new_n1960_ = new_n2936_ & new_n2958_;
  assign new_n1961_ = new_n2957_ & new_n2376_;
  assign new_n1962_ = new_n2942_ & new_n4738_;
  assign new_n1963_ = new_n2958_ & new_n1952_;
  assign new_n1964_ = new_n2942_ & new_n2376_;
  assign new_n1965_ = new_n4744_ & new_n3850_;
  assign new_n1966_ = new_n1950_ & new_n4744_;
  assign new_n1967_ = new_n4738_ & new_n3850_;
  assign new_n1968_ = new_n1950_ & new_n4738_;
  assign new_n1969_ = new_n1942_ & new_n3850_;
  assign new_n1970_ = new_n1950_ & new_n1942_;
  assign new_n1971_ = new_n1949_ & new_n2355_;
  assign new_n1972_ = new_n1949_ & new_n4086_;
  assign new_n1973_ = new_n2533_ & new_n1943_;
  assign new_n1974_ = new_n2379_ & new_n2380_;
  assign new_n1975_ = new_n4726_ & new_n2379_;
  assign new_n1976_ = new_n4729_ & new_n4723_;
  assign new_n1977_ = new_n2777_ & new_n4075_;
  assign new_n1978_ = new_n2346_ & new_n2294_;
  assign new_n1979_ = new_n2806_ & new_n4468_ & new_n2349_;
  assign new_n1980_ = ~new_n3608_ | ~new_n3609_ | ~new_n3606_ | ~new_n3607_;
  assign new_n1981_ = ~new_n3627_ | ~new_n3628_ | ~new_n3625_ | ~new_n3626_;
  assign new_n1982_ = ~new_n3646_ | ~new_n3644_ | ~new_n3645_ | ~new_n3647_;
  assign new_n1983_ = ~new_n3683_ | ~new_n3684_ | ~new_n3685_;
  assign new_n1984_ = ~new_n3589_ | ~new_n3590_ | ~new_n3587_ | ~new_n3588_;
  assign new_n1985_ = ~new_n3570_ | ~new_n3571_ | ~new_n3568_ | ~new_n3569_;
  assign new_n1986_ = ~new_n3663_ | ~new_n3664_ | ~new_n3665_;
  assign new_n1987_ = ~new_n3171_ | ~new_n3169_ | ~new_n3170_ | ~new_n3172_;
  assign new_n1988_ = ~new_n3513_ | ~new_n3514_ | ~new_n3511_ | ~new_n3512_;
  assign new_n1989_ = ~new_n3285_ | ~new_n3286_ | ~new_n3283_ | ~new_n3284_;
  assign new_n1990_ = ~new_n3304_ | ~new_n3305_ | ~new_n3302_ | ~new_n3303_;
  assign new_n1991_ = ~new_n3152_ | ~new_n3150_ | ~new_n3151_ | ~new_n3153_;
  assign new_n1992_ = ~new_n3551_ | ~new_n3552_ | ~new_n3549_ | ~new_n3550_;
  assign new_n1993_ = ~new_n3532_ | ~new_n3533_ | ~new_n3530_ | ~new_n3531_;
  assign new_n1994_ = ~new_n3190_ | ~new_n3188_ | ~new_n3189_ | ~new_n3191_;
  assign new_n1995_ = ~new_n3128_ | ~new_n3126_ | ~new_n3127_ | ~new_n3129_;
  assign new_n1996_ = ~new_n3418_ | ~new_n3419_ | ~new_n3416_ | ~new_n3417_;
  assign new_n1997_ = ~new_n3228_ | ~new_n3226_ | ~new_n3227_ | ~new_n3229_;
  assign new_n1998_ = ~new_n3209_ | ~new_n3207_ | ~new_n3208_ | ~new_n3210_;
  assign new_n1999_ = ~new_n3323_ | ~new_n3324_ | ~new_n3321_ | ~new_n3322_;
  assign new_n2000_ = ~new_n3399_ | ~new_n3400_ | ~new_n3397_ | ~new_n3398_;
  assign new_n2001_ = ~new_n3380_ | ~new_n3381_ | ~new_n3378_ | ~new_n3379_;
  assign new_n2002_ = ~new_n3494_ | ~new_n3495_ | ~new_n3492_ | ~new_n3493_;
  assign new_n2003_ = ~new_n3475_ | ~new_n3476_ | ~new_n3473_ | ~new_n3474_;
  assign new_n2004_ = ~new_n3133_ | ~new_n3131_ | ~new_n3132_ | ~new_n3134_;
  assign new_n2005_ = ~new_n3109_ | ~new_n3107_ | ~new_n3108_ | ~new_n3110_;
  assign new_n2006_ = ~new_n3361_ | ~new_n3362_ | ~new_n3359_ | ~new_n3360_;
  assign new_n2007_ = ~new_n3342_ | ~new_n3343_ | ~new_n3340_ | ~new_n3341_;
  assign new_n2008_ = ~new_n3456_ | ~new_n3457_ | ~new_n3454_ | ~new_n3455_;
  assign new_n2009_ = ~new_n3437_ | ~new_n3438_ | ~new_n3435_ | ~new_n3436_;
  assign new_n2010_ = ~new_n3266_ | ~new_n3267_ | ~new_n3264_ | ~new_n3265_;
  assign new_n2011_ = ~new_n3247_ | ~new_n3245_ | ~new_n3246_ | ~new_n3248_;
  assign po265 = ~new_n3857_ | ~pi275;
  assign po264 = ~pi275;
  assign new_n2014_ = ~new_n4594_ | ~new_n4595_ | ~new_n4593_;
  assign new_n2015_ = ~new_n4597_ | ~new_n4598_ | ~new_n4596_;
  assign new_n2016_ = ~new_n4606_ | ~new_n2856_ | ~new_n4605_;
  assign new_n2017_ = ~new_n2857_ | ~new_n4610_ | ~new_n4609_;
  assign new_n2018_ = ~new_n2858_ | ~new_n4614_ | ~new_n4613_;
  assign new_n2019_ = ~new_n2859_ | ~new_n4618_ | ~new_n4617_;
  assign new_n2020_ = ~new_n2860_ | ~new_n4622_ | ~new_n4621_;
  assign new_n2021_ = ~new_n2861_ | ~new_n4626_ | ~new_n4625_;
  assign new_n2022_ = ~new_n2862_ | ~new_n4630_ | ~new_n4629_;
  assign new_n2023_ = ~new_n2863_ | ~new_n4634_ | ~new_n4633_;
  assign new_n2024_ = ~new_n2864_ | ~new_n4638_ | ~new_n4637_;
  assign new_n2025_ = ~new_n2865_ | ~new_n4642_ | ~new_n4641_;
  assign new_n2026_ = ~new_n2867_ | ~new_n4650_ | ~new_n4649_;
  assign new_n2027_ = ~new_n2868_ | ~new_n4654_ | ~new_n4653_;
  assign new_n2028_ = ~new_n2869_ | ~new_n4658_ | ~new_n4657_;
  assign new_n2029_ = ~new_n2870_ | ~new_n4662_ | ~new_n4661_;
  assign new_n2030_ = ~new_n2871_ | ~new_n4666_ | ~new_n4665_;
  assign new_n2031_ = ~new_n2872_ | ~new_n4670_ | ~new_n4669_;
  assign new_n2032_ = ~new_n2873_ | ~new_n4674_ | ~new_n4673_;
  assign new_n2033_ = ~new_n2874_ | ~new_n4678_ | ~new_n4677_;
  assign new_n2034_ = ~new_n2875_ | ~new_n4682_ | ~new_n4681_;
  assign new_n2035_ = ~new_n2876_ | ~new_n4686_ | ~new_n4685_;
  assign new_n2036_ = ~new_n4570_ | ~new_n2849_ | ~new_n4571_;
  assign new_n2037_ = ~new_n4574_ | ~new_n2850_ | ~new_n4575_;
  assign new_n2038_ = ~new_n2851_ | ~new_n4580_ | ~new_n4579_;
  assign new_n2039_ = ~new_n2852_ | ~new_n4584_ | ~new_n4583_;
  assign new_n2040_ = ~new_n2853_ | ~new_n4588_ | ~new_n4587_;
  assign new_n2041_ = ~new_n2854_ | ~new_n4592_ | ~new_n4591_;
  assign new_n2042_ = ~new_n2855_ | ~new_n4601_;
  assign new_n2043_ = ~new_n2866_ | ~new_n4645_;
  assign new_n2044_ = ~new_n2877_ | ~new_n4689_;
  assign new_n2045_ = ~new_n2878_ | ~new_n4693_;
  assign new_n2046_ = ~new_n2819_ | ~new_n4490_;
  assign new_n2047_ = ~new_n2820_ | ~new_n4493_;
  assign new_n2048_ = ~new_n2823_ | ~new_n4499_ | ~new_n4498_;
  assign new_n2049_ = ~new_n2824_ | ~new_n4502_ | ~new_n4501_;
  assign new_n2050_ = ~new_n2825_ | ~new_n4505_ | ~new_n4504_;
  assign new_n2051_ = ~new_n2826_ | ~new_n4508_ | ~new_n4507_;
  assign new_n2052_ = ~new_n2827_ | ~new_n4511_ | ~new_n4510_;
  assign new_n2053_ = ~new_n2828_ | ~new_n4514_ | ~new_n4513_;
  assign new_n2054_ = ~new_n2829_ | ~new_n4517_ | ~new_n4516_;
  assign new_n2055_ = ~new_n2830_ | ~new_n4520_ | ~new_n4519_;
  assign new_n2056_ = ~new_n2831_ | ~new_n4523_ | ~new_n4522_;
  assign new_n2057_ = ~new_n2832_ | ~new_n4526_ | ~new_n4525_;
  assign new_n2058_ = ~new_n2835_ | ~new_n4532_ | ~new_n4531_;
  assign new_n2059_ = ~new_n2836_ | ~new_n4535_ | ~new_n4534_;
  assign new_n2060_ = ~new_n2837_ | ~new_n4538_ | ~new_n4537_;
  assign new_n2061_ = ~new_n2838_ | ~new_n4541_ | ~new_n4540_;
  assign new_n2062_ = ~new_n2839_ | ~new_n4544_ | ~new_n4543_;
  assign new_n2063_ = ~new_n2840_ | ~new_n4547_ | ~new_n4546_;
  assign new_n2064_ = ~new_n2841_ | ~new_n4550_ | ~new_n4549_;
  assign new_n2065_ = ~new_n2842_ | ~new_n4553_ | ~new_n4552_;
  assign new_n2066_ = ~new_n2843_ | ~new_n4556_ | ~new_n4555_;
  assign new_n2067_ = ~new_n2844_ | ~new_n4559_ | ~new_n4558_;
  assign new_n2068_ = ~new_n4472_ | ~new_n2807_;
  assign new_n2069_ = ~new_n4475_ | ~new_n2809_;
  assign new_n2070_ = ~new_n4478_ | ~new_n2811_;
  assign new_n2071_ = ~new_n4481_ | ~new_n2813_;
  assign new_n2072_ = ~new_n4484_ | ~new_n2815_;
  assign new_n2073_ = ~new_n4487_ | ~new_n2817_;
  assign new_n2074_ = ~new_n4496_ | ~new_n2821_;
  assign new_n2075_ = ~new_n4529_ | ~new_n2833_;
  assign new_n2076_ = ~new_n4562_ | ~new_n2845_;
  assign new_n2077_ = ~new_n4565_ | ~new_n2847_;
  assign new_n2078_ = ~new_n2804_ | ~new_n4464_;
  assign new_n2079_ = ~new_n1941_ | ~new_n4713_;
  assign new_n2080_ = ~new_n4419_ | ~new_n4418_;
  assign new_n2081_ = ~new_n4421_ | ~new_n4420_;
  assign new_n2082_ = ~new_n4423_ | ~new_n4422_;
  assign new_n2083_ = ~new_n4425_ | ~new_n4424_;
  assign new_n2084_ = ~new_n4427_ | ~new_n4426_;
  assign new_n2085_ = ~new_n4429_ | ~new_n4428_;
  assign new_n2086_ = ~new_n4431_ | ~new_n4430_;
  assign new_n2087_ = ~new_n4433_ | ~new_n4432_;
  assign new_n2088_ = ~new_n4435_ | ~new_n4434_;
  assign new_n2089_ = ~new_n4439_ | ~new_n4438_;
  assign new_n2090_ = ~new_n4441_ | ~new_n4440_;
  assign new_n2091_ = ~new_n4443_ | ~new_n4442_;
  assign new_n2092_ = ~new_n4445_ | ~new_n4444_;
  assign new_n2093_ = ~new_n4447_ | ~new_n4446_;
  assign new_n2094_ = ~new_n4449_ | ~new_n4448_;
  assign new_n2095_ = ~new_n4451_ | ~new_n4450_;
  assign new_n2096_ = ~new_n4453_ | ~new_n4452_;
  assign new_n2097_ = ~new_n4455_ | ~new_n4454_;
  assign new_n2098_ = ~new_n4457_ | ~new_n4456_;
  assign new_n2099_ = ~new_n4405_ | ~new_n4404_;
  assign new_n2100_ = ~new_n4407_ | ~new_n4406_;
  assign new_n2101_ = ~new_n4409_ | ~new_n4408_;
  assign new_n2102_ = ~new_n4411_ | ~new_n4410_;
  assign new_n2103_ = ~new_n4413_ | ~new_n4412_;
  assign new_n2104_ = ~new_n4415_ | ~new_n4414_;
  assign new_n2105_ = ~new_n4417_ | ~new_n4416_;
  assign new_n2106_ = ~new_n4437_ | ~new_n4436_;
  assign new_n2107_ = ~new_n4459_ | ~new_n4458_;
  assign new_n2108_ = ~new_n2803_ | ~new_n4461_;
  assign new_n2109_ = ~new_n4360_ | ~new_n4359_;
  assign new_n2110_ = ~new_n4362_ | ~new_n4361_;
  assign new_n2111_ = ~new_n4364_ | ~new_n4363_;
  assign new_n2112_ = ~new_n4366_ | ~new_n4365_;
  assign new_n2113_ = ~new_n4368_ | ~new_n4367_;
  assign new_n2114_ = ~new_n4370_ | ~new_n4369_;
  assign new_n2115_ = ~new_n4372_ | ~new_n4371_;
  assign new_n2116_ = ~new_n4374_ | ~new_n4373_;
  assign new_n2117_ = ~new_n4376_ | ~new_n4375_;
  assign new_n2118_ = ~new_n4380_ | ~new_n4379_;
  assign new_n2119_ = ~new_n4382_ | ~new_n4381_;
  assign new_n2120_ = ~new_n4384_ | ~new_n4383_;
  assign new_n2121_ = ~new_n4386_ | ~new_n4385_;
  assign new_n2122_ = ~new_n4388_ | ~new_n4387_;
  assign new_n2123_ = ~new_n4390_ | ~new_n4389_;
  assign new_n2124_ = ~new_n4392_ | ~new_n4391_;
  assign new_n2125_ = ~new_n4394_ | ~new_n4393_;
  assign new_n2126_ = ~new_n4396_ | ~new_n4395_;
  assign new_n2127_ = ~new_n4398_ | ~new_n4397_;
  assign new_n2128_ = ~new_n4346_ | ~new_n4345_;
  assign new_n2129_ = ~new_n4348_ | ~new_n4347_;
  assign new_n2130_ = ~new_n4350_ | ~new_n4349_;
  assign new_n2131_ = ~new_n4352_ | ~new_n4351_;
  assign new_n2132_ = ~new_n4354_ | ~new_n4353_;
  assign new_n2133_ = ~new_n4356_ | ~new_n4355_;
  assign new_n2134_ = ~new_n4358_ | ~new_n4357_;
  assign new_n2135_ = ~new_n4378_ | ~new_n4377_;
  assign new_n2136_ = ~new_n4400_ | ~new_n4399_;
  assign new_n2137_ = ~new_n2802_ | ~new_n4401_;
  assign new_n2138_ = new_n4338_ & new_n2352_;
  assign new_n2139_ = ~new_n4336_ | ~new_n5212_ | ~new_n5211_;
  assign po263 = ~new_n4329_ | ~new_n4331_ | ~new_n2799_ | ~new_n4330_;
  assign po262 = ~new_n4321_ | ~new_n4322_ | ~new_n4323_ | ~new_n4324_ | ~new_n4320_;
  assign po261 = ~new_n4312_ | ~new_n4313_ | ~new_n4314_ | ~new_n4315_ | ~new_n4311_;
  assign po260 = ~new_n4303_ | ~new_n4304_ | ~new_n4305_ | ~new_n4306_ | ~new_n4302_;
  assign po259 = ~new_n4293_ | ~new_n4295_ | ~new_n2798_ | ~new_n4294_;
  assign po258 = ~new_n2797_ | ~new_n2796_ | ~new_n4285_;
  assign po257 = ~new_n4276_ | ~new_n4277_ | ~new_n4278_ | ~new_n4279_ | ~new_n4275_;
  assign po256 = ~new_n4267_ | ~new_n4268_ | ~new_n4269_ | ~new_n4270_ | ~new_n4266_;
  assign po255 = ~new_n4257_ | ~new_n4259_ | ~new_n2795_ | ~new_n4258_;
  assign po254 = ~new_n2794_ | ~new_n2793_ | ~new_n4249_;
  assign po253 = ~new_n4240_ | ~new_n4241_ | ~new_n4242_ | ~new_n4243_ | ~new_n4239_;
  assign po252 = ~new_n4230_ | ~new_n4232_ | ~new_n2792_ | ~new_n4231_;
  assign po251 = ~new_n4222_ | ~new_n4223_ | ~new_n4224_ | ~new_n4225_ | ~new_n4221_;
  assign po250 = ~new_n4213_ | ~new_n4214_ | ~new_n4215_ | ~new_n4216_ | ~new_n4212_;
  assign po249 = ~new_n4203_ | ~new_n2791_ | ~new_n4205_ | ~new_n4204_;
  assign po248 = ~new_n4195_ | ~new_n4196_ | ~new_n4197_ | ~new_n4198_ | ~new_n4194_;
  assign po247 = ~new_n4186_ | ~new_n4187_ | ~new_n4188_ | ~new_n4189_ | ~new_n4185_;
  assign po246 = ~new_n2790_ | ~new_n2789_ | ~new_n4177_;
  assign po245 = ~new_n4167_ | ~new_n4169_ | ~new_n2788_ | ~new_n4168_;
  assign po244 = ~new_n4160_ | ~new_n2786_;
  assign po243 = ~new_n4151_ | ~new_n4152_ | ~new_n4153_ | ~new_n4154_ | ~new_n4150_;
  assign po242 = ~new_n4141_ | ~new_n4143_ | ~new_n2784_ | ~new_n4142_;
  assign po241 = ~new_n4133_ | ~new_n4134_ | ~new_n4135_ | ~new_n4136_ | ~new_n4132_;
  assign po240 = ~new_n4123_ | ~new_n4125_ | ~new_n2783_ | ~new_n4124_;
  assign po239 = ~new_n2782_ | ~new_n2781_ | ~new_n4115_;
  assign po238 = ~new_n4106_ | ~new_n4107_ | ~new_n4108_ | ~new_n4109_ | ~new_n4105_;
  assign po237 = ~new_n4096_ | ~new_n4098_ | ~new_n2780_ | ~new_n4097_;
  assign po236 = ~new_n4088_ | ~new_n4089_ | ~new_n4090_ | ~new_n4091_ | ~new_n4087_;
  assign po235 = ~new_n4077_ | ~new_n4078_ | ~new_n4079_ | ~new_n4080_ | ~new_n4076_;
  assign po234 = ~new_n2773_ | ~new_n4064_;
  assign po201 = ~new_n2758_ | ~new_n2757_ | ~new_n4050_;
  assign po200 = ~new_n2756_ | ~new_n2755_ | ~new_n4040_;
  assign po199 = ~new_n2754_ | ~new_n4030_ | ~new_n2752_;
  assign po198 = ~new_n2751_ | ~new_n2750_ | ~new_n4020_;
  assign po197 = ~new_n2749_ | ~new_n4010_ | ~new_n2747_;
  assign po196 = ~new_n2746_ | ~new_n2745_ | ~new_n4000_;
  assign po195 = ~new_n3990_ | ~new_n2743_ | ~new_n2744_;
  assign po194 = ~new_n3980_ | ~new_n2741_ | ~new_n2742_;
  assign po193 = ~new_n3970_ | ~new_n2739_ | ~new_n2740_;
  assign po192 = ~new_n3960_ | ~new_n2737_ | ~new_n2738_;
  assign po191 = ~new_n3950_ | ~new_n2735_ | ~new_n2736_;
  assign po190 = ~new_n3940_ | ~new_n2733_ | ~new_n2734_;
  assign po189 = ~new_n3930_ | ~new_n2731_ | ~new_n2732_;
  assign po188 = ~new_n3920_ | ~new_n2729_ | ~new_n2730_;
  assign po187 = ~new_n3910_ | ~new_n2727_ | ~new_n2728_;
  assign po186 = ~new_n3900_ | ~new_n2725_ | ~new_n2726_;
  assign po185 = ~new_n3890_ | ~new_n2723_ | ~new_n2724_;
  assign po184 = ~new_n3880_ | ~new_n2721_ | ~new_n2722_;
  assign po183 = ~new_n3870_ | ~new_n2719_ | ~new_n2720_;
  assign po182 = ~new_n3860_ | ~new_n2717_ | ~new_n2718_;
  assign po181 = ~new_n3849_ | ~new_n2916_ | ~new_n3848_;
  assign po180 = ~new_n3847_ | ~new_n2915_ | ~new_n3846_;
  assign po178 = ~new_n2712_ | ~new_n2912_ | ~new_n3839_ | ~new_n2711_;
  assign po177 = ~new_n2710_ | ~new_n2911_ | ~new_n3834_ | ~new_n2709_;
  assign po176 = ~new_n2708_ | ~new_n2910_ | ~new_n3829_ | ~new_n2707_;
  assign po175 = ~new_n2706_ | ~new_n2909_ | ~new_n3824_ | ~new_n2705_;
  assign po174 = ~new_n2704_ | ~new_n2908_ | ~new_n3819_ | ~new_n2703_;
  assign po173 = ~new_n2702_ | ~new_n2907_ | ~new_n3814_ | ~new_n2701_;
  assign po172 = ~new_n2700_ | ~new_n2906_ | ~new_n3809_ | ~new_n2699_;
  assign po171 = ~new_n2698_ | ~new_n2905_ | ~new_n3804_ | ~new_n2697_;
  assign po170 = ~new_n2696_ | ~new_n2904_ | ~new_n3799_ | ~new_n2695_;
  assign po169 = ~new_n2694_ | ~new_n2903_ | ~new_n3794_ | ~new_n2693_;
  assign po168 = ~new_n2902_ | ~new_n2692_ | ~new_n2691_;
  assign po167 = ~new_n2901_ | ~new_n2690_ | ~new_n2689_;
  assign po166 = ~new_n2688_ | ~new_n2900_ | ~new_n3779_ | ~new_n2687_;
  assign po165 = ~new_n2686_ | ~new_n2899_ | ~new_n3774_ | ~new_n2685_;
  assign po164 = ~new_n2898_ | ~new_n2684_ | ~new_n2683_;
  assign po163 = ~new_n2897_ | ~new_n2682_ | ~new_n2681_;
  assign po162 = ~new_n2896_ | ~new_n2680_ | ~new_n2679_;
  assign po161 = ~new_n2895_ | ~new_n2678_ | ~new_n2677_;
  assign po160 = ~new_n2676_ | ~new_n2894_ | ~new_n3749_ | ~new_n2675_;
  assign po159 = ~new_n2674_ | ~new_n2893_ | ~new_n3744_ | ~new_n2673_;
  assign po158 = ~new_n2892_ | ~new_n2672_ | ~new_n2671_;
  assign po157 = ~new_n2891_ | ~new_n2670_ | ~new_n2669_;
  assign po156 = ~new_n2890_ | ~new_n2668_ | ~new_n2667_;
  assign po155 = ~new_n2889_ | ~new_n2666_ | ~new_n2665_;
  assign po154 = ~new_n2664_ | ~new_n2663_;
  assign po153 = ~new_n2662_ | ~new_n2661_;
  assign po152 = ~new_n2660_ | ~new_n2659_;
  assign po151 = ~new_n2658_ | ~new_n2657_;
  assign po150 = ~new_n2656_ | ~new_n2655_;
  assign po085 = pi096 & new_n2880_;
  assign po084 = pi095 & new_n2880_;
  assign po083 = pi094 & new_n2880_;
  assign po082 = pi093 & new_n2880_;
  assign po081 = pi092 & new_n2880_;
  assign po080 = pi091 & new_n2880_;
  assign po079 = pi090 & new_n2880_;
  assign po078 = pi089 & new_n2880_;
  assign po077 = pi088 & new_n2880_;
  assign po076 = pi087 & new_n2880_;
  assign po075 = pi086 & new_n2880_;
  assign po074 = pi085 & new_n2880_;
  assign po073 = pi084 & new_n2880_;
  assign po072 = pi083 & new_n2880_;
  assign po071 = pi082 & new_n2880_;
  assign po070 = pi081 & new_n2880_;
  assign po069 = pi080 & new_n2880_;
  assign po068 = pi079 & new_n2880_;
  assign po067 = pi078 & new_n2880_;
  assign po066 = pi077 & new_n2880_;
  assign po065 = pi076 & new_n2880_;
  assign po064 = pi075 & new_n2880_;
  assign po063 = pi074 & new_n2880_;
  assign po062 = pi073 & new_n2880_;
  assign po061 = pi072 & new_n2880_;
  assign po060 = pi071 & new_n2880_;
  assign po059 = pi070 & new_n2880_;
  assign po058 = pi069 & new_n2880_;
  assign po057 = pi068 & new_n2880_;
  assign po056 = pi067 & new_n2880_;
  assign po053 = ~new_n3068_ | ~new_n3069_ | ~new_n3070_;
  assign po052 = ~new_n3065_ | ~new_n3066_ | ~new_n3067_;
  assign po051 = ~new_n3062_ | ~new_n3063_ | ~new_n3064_;
  assign po050 = ~new_n3059_ | ~new_n3060_ | ~new_n3061_;
  assign po049 = ~new_n3056_ | ~new_n3057_ | ~new_n3058_;
  assign po048 = ~new_n3053_ | ~new_n3054_ | ~new_n3055_;
  assign po047 = ~new_n3050_ | ~new_n3051_ | ~new_n3052_;
  assign po046 = ~new_n3047_ | ~new_n3048_ | ~new_n3049_;
  assign po045 = ~new_n3044_ | ~new_n3045_ | ~new_n3046_;
  assign po044 = ~new_n3041_ | ~new_n3042_ | ~new_n3043_;
  assign po043 = ~new_n3038_ | ~new_n3039_ | ~new_n3040_;
  assign po042 = ~new_n3035_ | ~new_n3036_ | ~new_n3037_;
  assign po041 = ~new_n3032_ | ~new_n3033_ | ~new_n3034_;
  assign po040 = ~new_n3029_ | ~new_n3030_ | ~new_n3031_;
  assign po039 = ~new_n3026_ | ~new_n3027_ | ~new_n3028_;
  assign po038 = ~new_n3023_ | ~new_n3024_ | ~new_n3025_;
  assign po037 = ~new_n3020_ | ~new_n3021_ | ~new_n3022_;
  assign po036 = ~new_n3017_ | ~new_n3018_ | ~new_n3019_;
  assign po035 = ~new_n3014_ | ~new_n3015_ | ~new_n3016_;
  assign po034 = ~new_n3011_ | ~new_n3012_ | ~new_n3013_;
  assign po033 = ~new_n3008_ | ~new_n3009_ | ~new_n3010_;
  assign po032 = ~new_n3005_ | ~new_n3006_ | ~new_n3007_;
  assign po031 = ~new_n3002_ | ~new_n3003_ | ~new_n3004_;
  assign po030 = ~new_n2999_ | ~new_n3000_ | ~new_n3001_;
  assign po029 = ~new_n2996_ | ~new_n2997_ | ~new_n2998_;
  assign po028 = ~new_n2993_ | ~new_n2994_ | ~new_n2995_;
  assign po027 = ~new_n2990_ | ~new_n2991_ | ~new_n2992_;
  assign po026 = ~new_n2987_ | ~new_n2988_ | ~new_n2989_;
  assign po025 = ~new_n2984_ | ~new_n2985_ | ~new_n2986_;
  assign po024 = ~new_n2981_ | ~new_n2982_ | ~new_n2983_;
  assign po023 = ~new_n2978_ | ~new_n2979_ | ~new_n2980_;
  assign po022 = ~new_n2975_ | ~new_n2976_ | ~new_n2977_;
  assign po179 = ~new_n3844_ | ~new_n2913_ | ~new_n3843_ | ~new_n3845_ | ~new_n3842_;
  assign new_n2284_ = ~pi275 | ~new_n2879_;
  assign new_n2285_ = ~new_n2370_ | ~new_n4705_;
  assign new_n2286_ = ~pi245;
  assign new_n2287_ = ~new_n2370_ | ~new_n4710_ | ~new_n4709_;
  assign new_n2288_ = ~new_n1975_ | ~new_n2378_;
  assign new_n2289_ = ~new_n1974_ | ~new_n2378_;
  assign new_n2290_ = ~new_n2380_ | ~new_n4723_;
  assign new_n2291_ = ~new_n2969_ | ~new_n2378_;
  assign new_n2292_ = ~new_n1974_ | ~new_n2377_;
  assign new_n2293_ = ~new_n2969_ | ~new_n2377_;
  assign new_n2294_ = ~new_n1976_ | ~new_n2378_;
  assign new_n2295_ = ~new_n2928_ | ~new_n4726_;
  assign new_n2296_ = ~new_n4726_ | ~new_n4723_;
  assign new_n2297_ = ~new_n2971_ | ~new_n2377_;
  assign new_n2298_ = ~new_n2929_ | ~new_n4720_;
  assign new_n2299_ = ~new_n2378_ | ~new_n2377_;
  assign new_n2300_ = ~new_n4729_ | ~new_n4726_ | ~new_n4720_;
  assign new_n2301_ = ~new_n1976_ | ~new_n4720_;
  assign new_n2302_ = ~new_n4729_ | ~new_n2379_;
  assign new_n2303_ = ~new_n3118_ | ~new_n2520_ | ~new_n2521_ | ~new_n3119_ | ~new_n3117_;
  assign new_n2304_ = ~pi161;
  assign new_n2305_ = ~new_n3136_ | ~new_n2537_ | ~new_n2535_ | ~new_n3137_;
  assign new_n2306_ = ~new_n3155_ | ~new_n2541_ | ~new_n2539_ | ~new_n3156_;
  assign new_n2307_ = ~new_n3174_ | ~new_n2545_ | ~new_n2543_ | ~new_n3175_;
  assign new_n2308_ = ~new_n3193_ | ~new_n2549_ | ~new_n2547_ | ~new_n3194_;
  assign new_n2309_ = ~new_n3212_ | ~new_n2553_ | ~new_n2551_ | ~new_n3213_;
  assign new_n2310_ = ~new_n3231_ | ~new_n2557_ | ~new_n2555_ | ~new_n3232_;
  assign new_n2311_ = ~new_n3250_ | ~new_n2561_ | ~new_n2559_ | ~new_n3251_;
  assign new_n2312_ = ~new_n3269_ | ~new_n2565_ | ~new_n2563_ | ~new_n3270_;
  assign new_n2313_ = ~new_n3288_ | ~new_n2569_ | ~new_n2567_ | ~new_n3289_;
  assign new_n2314_ = ~new_n3307_ | ~new_n2573_ | ~new_n2571_ | ~new_n3308_;
  assign new_n2315_ = ~new_n3326_ | ~new_n2577_ | ~new_n2575_ | ~new_n3327_;
  assign new_n2316_ = ~new_n3345_ | ~new_n2581_ | ~new_n2579_ | ~new_n3346_;
  assign new_n2317_ = ~new_n3364_ | ~new_n2585_ | ~new_n2583_ | ~new_n3365_;
  assign new_n2318_ = ~new_n3383_ | ~new_n2589_ | ~new_n2587_ | ~new_n3384_;
  assign new_n2319_ = ~new_n3402_ | ~new_n2593_ | ~new_n2591_ | ~new_n3403_;
  assign new_n2320_ = ~new_n3421_ | ~new_n2597_ | ~new_n2595_ | ~new_n3422_;
  assign new_n2321_ = ~new_n3440_ | ~new_n2601_ | ~new_n2599_ | ~new_n3441_;
  assign new_n2322_ = ~new_n3459_ | ~new_n2605_ | ~new_n2603_ | ~new_n3460_;
  assign new_n2323_ = ~new_n3478_ | ~new_n2609_ | ~new_n2607_ | ~new_n3479_;
  assign new_n2324_ = ~new_n1614_ | ~new_n2881_;
  assign new_n2325_ = ~new_n3497_ | ~new_n2613_ | ~new_n2611_ | ~new_n3498_;
  assign new_n2326_ = ~new_n1613_ | ~new_n2881_;
  assign new_n2327_ = ~new_n3516_ | ~new_n2617_ | ~new_n2615_ | ~new_n3517_;
  assign new_n2328_ = ~new_n1612_ | ~new_n2881_;
  assign new_n2329_ = ~new_n3535_ | ~new_n2621_ | ~new_n2619_ | ~new_n3536_;
  assign new_n2330_ = ~new_n1611_ | ~new_n2881_;
  assign new_n2331_ = ~new_n3554_ | ~new_n2625_ | ~new_n2623_ | ~new_n3555_;
  assign new_n2332_ = ~new_n1610_ | ~new_n2881_;
  assign new_n2333_ = ~new_n3573_ | ~new_n2629_ | ~new_n2627_ | ~new_n3574_;
  assign new_n2334_ = ~new_n1609_ | ~new_n2881_;
  assign new_n2335_ = ~new_n3592_ | ~new_n2633_ | ~new_n2631_ | ~new_n3593_;
  assign new_n2336_ = ~new_n1608_ | ~new_n2881_;
  assign new_n2337_ = ~new_n3611_ | ~new_n2637_ | ~new_n2635_ | ~new_n3612_;
  assign new_n2338_ = ~new_n1607_ | ~new_n2881_;
  assign new_n2339_ = ~new_n3630_ | ~new_n2641_ | ~new_n2639_ | ~new_n3631_;
  assign new_n2340_ = ~new_n1606_ | ~new_n2881_;
  assign new_n2341_ = ~new_n3649_ | ~new_n2645_ | ~new_n2643_ | ~new_n3650_;
  assign new_n2342_ = ~new_n1605_ | ~new_n2881_;
  assign new_n2343_ = ~new_n2650_ | ~new_n2648_;
  assign new_n2344_ = ~new_n1603_ | ~new_n2881_;
  assign new_n2345_ = ~new_n1602_ | ~new_n2881_;
  assign new_n2346_ = ~new_n2968_ | ~new_n4720_;
  assign new_n2347_ = ~new_n1949_ | ~new_n3694_;
  assign new_n2348_ = ~new_n2925_ | ~new_n4726_;
  assign new_n2349_ = ~new_n1975_ | ~new_n2377_;
  assign new_n2350_ = ~new_n1974_ | ~new_n4720_;
  assign new_n2351_ = ~new_n2920_ | ~new_n4726_;
  assign new_n2352_ = ~new_n2369_ | ~new_n2368_ | ~new_n2370_;
  assign new_n2353_ = ~new_n2937_ | ~new_n3695_;
  assign new_n2354_ = ~new_n2371_ | ~pi275;
  assign new_n2355_ = ~new_n2356_ | ~new_n3858_;
  assign new_n2356_ = ~new_n3072_ | ~new_n4713_;
  assign new_n2357_ = ~new_n2972_ | ~pi275;
  assign new_n2358_ = ~new_n1941_ | ~new_n1942_;
  assign new_n2359_ = ~new_n15169_;
  assign new_n2360_ = ~new_n1949_ | ~new_n2353_;
  assign new_n2361_ = ~new_n2774_ | ~new_n1943_;
  assign new_n2362_ = ~new_n2779_ | ~new_n4070_;
  assign new_n2363_ = ~new_n4342_ | ~new_n4341_;
  assign new_n2364_ = ~new_n2926_ | ~new_n2289_;
  assign new_n2365_ = ~new_n4463_ | ~new_n1978_;
  assign new_n2366_ = ~new_n15358_;
  assign new_n2367_ = ~new_n2291_ | ~new_n2350_;
  assign new_n2368_ = ~new_n4701_ | ~new_n4700_;
  assign new_n2369_ = ~new_n4704_ | ~new_n4703_;
  assign new_n2370_ = ~new_n4707_ | ~new_n4706_;
  assign new_n2371_ = ~new_n4712_ | ~new_n4711_;
  assign po054 = ~new_n4715_ | ~new_n4714_;
  assign po055 = ~new_n4717_ | ~new_n4716_;
  assign new_n2374_ = ~new_n4731_ | ~new_n4730_;
  assign new_n2375_ = ~new_n4734_ | ~new_n4733_;
  assign new_n2376_ = ~new_n4737_ | ~new_n4736_;
  assign new_n2377_ = ~new_n4728_ | ~new_n4727_;
  assign new_n2378_ = ~new_n4719_ | ~new_n4718_;
  assign new_n2379_ = ~new_n4722_ | ~new_n4721_;
  assign new_n2380_ = ~new_n4725_ | ~new_n4724_;
  assign new_n2381_ = ~new_n4740_ | ~new_n4739_;
  assign new_n2382_ = ~new_n4743_ | ~new_n4742_;
  assign new_n2383_ = ~new_n4746_ | ~new_n4745_;
  assign new_n2384_ = ~new_n4754_ | ~new_n4753_;
  assign new_n2385_ = ~new_n4751_ | ~new_n4750_;
  assign po086 = ~new_n4757_ | ~new_n4756_;
  assign new_n2387_ = ~new_n4759_ | ~new_n4758_;
  assign new_n2388_ = ~new_n4761_ | ~new_n4760_;
  assign po087 = ~new_n4764_ | ~new_n4763_;
  assign new_n2390_ = ~new_n4766_ | ~new_n4765_;
  assign new_n2391_ = ~new_n4768_ | ~new_n4767_;
  assign po088 = ~new_n4771_ | ~new_n4770_;
  assign new_n2393_ = ~new_n4773_ | ~new_n4772_;
  assign new_n2394_ = ~new_n4775_ | ~new_n4774_;
  assign po089 = ~new_n4778_ | ~new_n4777_;
  assign new_n2396_ = ~new_n4780_ | ~new_n4779_;
  assign new_n2397_ = ~new_n4782_ | ~new_n4781_;
  assign po090 = ~new_n4785_ | ~new_n4784_;
  assign new_n2399_ = ~new_n4787_ | ~new_n4786_;
  assign new_n2400_ = ~new_n4789_ | ~new_n4788_;
  assign po091 = ~new_n4792_ | ~new_n4791_;
  assign new_n2402_ = ~new_n4794_ | ~new_n4793_;
  assign new_n2403_ = ~new_n4796_ | ~new_n4795_;
  assign po092 = ~new_n4799_ | ~new_n4798_;
  assign new_n2405_ = ~new_n4801_ | ~new_n4800_;
  assign new_n2406_ = ~new_n4803_ | ~new_n4802_;
  assign po093 = ~new_n4806_ | ~new_n4805_;
  assign new_n2408_ = ~new_n4808_ | ~new_n4807_;
  assign new_n2409_ = ~new_n4810_ | ~new_n4809_;
  assign po094 = ~new_n4813_ | ~new_n4812_;
  assign new_n2411_ = ~new_n4815_ | ~new_n4814_;
  assign new_n2412_ = ~new_n4817_ | ~new_n4816_;
  assign po095 = ~new_n4820_ | ~new_n4819_;
  assign new_n2414_ = ~new_n4822_ | ~new_n4821_;
  assign new_n2415_ = ~new_n4824_ | ~new_n4823_;
  assign po096 = ~new_n4827_ | ~new_n4826_;
  assign new_n2417_ = ~new_n4829_ | ~new_n4828_;
  assign new_n2418_ = ~new_n4831_ | ~new_n4830_;
  assign po097 = ~new_n4834_ | ~new_n4833_;
  assign new_n2420_ = ~new_n4836_ | ~new_n4835_;
  assign new_n2421_ = ~new_n4838_ | ~new_n4837_;
  assign po098 = ~new_n4841_ | ~new_n4840_;
  assign new_n2423_ = ~new_n4843_ | ~new_n4842_;
  assign new_n2424_ = ~new_n4845_ | ~new_n4844_;
  assign po099 = ~new_n4848_ | ~new_n4847_;
  assign new_n2426_ = ~new_n4850_ | ~new_n4849_;
  assign new_n2427_ = ~new_n4852_ | ~new_n4851_;
  assign po100 = ~new_n4855_ | ~new_n4854_;
  assign new_n2429_ = ~new_n4857_ | ~new_n4856_;
  assign new_n2430_ = ~new_n4859_ | ~new_n4858_;
  assign po101 = ~new_n4862_ | ~new_n4861_;
  assign new_n2432_ = ~new_n4864_ | ~new_n4863_;
  assign new_n2433_ = ~new_n4866_ | ~new_n4865_;
  assign po102 = ~new_n4869_ | ~new_n4868_;
  assign new_n2435_ = ~new_n4871_ | ~new_n4870_;
  assign new_n2436_ = ~new_n4873_ | ~new_n4872_;
  assign po103 = ~new_n4876_ | ~new_n4875_;
  assign new_n2438_ = ~new_n4878_ | ~new_n4877_;
  assign new_n2439_ = ~new_n4880_ | ~new_n4879_;
  assign po104 = ~new_n4883_ | ~new_n4882_;
  assign new_n2441_ = ~new_n4885_ | ~new_n4884_;
  assign po105 = ~new_n4888_ | ~new_n4887_;
  assign po106 = ~new_n4890_ | ~new_n4889_;
  assign po107 = ~new_n4892_ | ~new_n4891_;
  assign po108 = ~new_n4894_ | ~new_n4893_;
  assign po109 = ~new_n4896_ | ~new_n4895_;
  assign po110 = ~new_n4898_ | ~new_n4897_;
  assign po111 = ~new_n4900_ | ~new_n4899_;
  assign po112 = ~new_n4902_ | ~new_n4901_;
  assign po113 = ~new_n4904_ | ~new_n4903_;
  assign po114 = ~new_n4906_ | ~new_n4905_;
  assign po115 = ~new_n4908_ | ~new_n4907_;
  assign po116 = ~new_n4910_ | ~new_n4909_;
  assign po117 = ~new_n4912_ | ~new_n4911_;
  assign po118 = ~new_n4914_ | ~new_n4913_;
  assign po119 = ~new_n4916_ | ~new_n4915_;
  assign po120 = ~new_n4918_ | ~new_n4917_;
  assign po121 = ~new_n4920_ | ~new_n4919_;
  assign po122 = ~new_n4922_ | ~new_n4921_;
  assign po123 = ~new_n4924_ | ~new_n4923_;
  assign po124 = ~new_n4926_ | ~new_n4925_;
  assign po125 = ~new_n4928_ | ~new_n4927_;
  assign po126 = ~new_n4930_ | ~new_n4929_;
  assign po127 = ~new_n4932_ | ~new_n4931_;
  assign po128 = ~new_n4934_ | ~new_n4933_;
  assign po129 = ~new_n4936_ | ~new_n4935_;
  assign po130 = ~new_n4938_ | ~new_n4937_;
  assign po131 = ~new_n4940_ | ~new_n4939_;
  assign po132 = ~new_n4942_ | ~new_n4941_;
  assign po133 = ~new_n4944_ | ~new_n4943_;
  assign po134 = ~new_n4946_ | ~new_n4945_;
  assign po135 = ~new_n4948_ | ~new_n4947_;
  assign po136 = ~new_n4950_ | ~new_n4949_;
  assign po137 = ~new_n4952_ | ~new_n4951_;
  assign po138 = ~new_n4954_ | ~new_n4953_;
  assign po139 = ~new_n4956_ | ~new_n4955_;
  assign po140 = ~new_n4958_ | ~new_n4957_;
  assign po141 = ~new_n4960_ | ~new_n4959_;
  assign po142 = ~new_n4962_ | ~new_n4961_;
  assign po143 = ~new_n4964_ | ~new_n4963_;
  assign po144 = ~new_n4966_ | ~new_n4965_;
  assign po145 = ~new_n4968_ | ~new_n4967_;
  assign po146 = ~new_n4970_ | ~new_n4969_;
  assign po147 = ~new_n4972_ | ~new_n4971_;
  assign po148 = ~new_n4974_ | ~new_n4973_;
  assign po149 = ~new_n4976_ | ~new_n4975_;
  assign po202 = ~new_n5042_ | ~new_n5041_;
  assign po203 = ~new_n5044_ | ~new_n5043_;
  assign po204 = ~new_n5046_ | ~new_n5045_;
  assign po205 = ~new_n5048_ | ~new_n5047_;
  assign po206 = ~new_n5050_ | ~new_n5049_;
  assign po207 = ~new_n5052_ | ~new_n5051_;
  assign po208 = ~new_n5054_ | ~new_n5053_;
  assign po209 = ~new_n5056_ | ~new_n5055_;
  assign po210 = ~new_n5058_ | ~new_n5057_;
  assign po211 = ~new_n5060_ | ~new_n5059_;
  assign po212 = ~new_n5062_ | ~new_n5061_;
  assign po213 = ~new_n5064_ | ~new_n5063_;
  assign po214 = ~new_n5066_ | ~new_n5065_;
  assign po215 = ~new_n5068_ | ~new_n5067_;
  assign po216 = ~new_n5070_ | ~new_n5069_;
  assign po217 = ~new_n5072_ | ~new_n5071_;
  assign po218 = ~new_n5074_ | ~new_n5073_;
  assign po219 = ~new_n5076_ | ~new_n5075_;
  assign po220 = ~new_n5078_ | ~new_n5077_;
  assign po221 = ~new_n5080_ | ~new_n5079_;
  assign po222 = ~new_n5082_ | ~new_n5081_;
  assign po223 = ~new_n5084_ | ~new_n5083_;
  assign po224 = ~new_n5086_ | ~new_n5085_;
  assign po225 = ~new_n5088_ | ~new_n5087_;
  assign po226 = ~new_n5090_ | ~new_n5089_;
  assign po227 = ~new_n5092_ | ~new_n5091_;
  assign po228 = ~new_n5094_ | ~new_n5093_;
  assign po229 = ~new_n5096_ | ~new_n5095_;
  assign po230 = ~new_n5098_ | ~new_n5097_;
  assign po231 = ~new_n5100_ | ~new_n5099_;
  assign po232 = ~new_n5102_ | ~new_n5101_;
  assign po233 = ~new_n5104_ | ~new_n5103_;
  assign new_n2519_ = new_n4713_ & pi275;
  assign new_n2520_ = new_n3114_ & new_n3113_;
  assign new_n2521_ = new_n3116_ & new_n3115_;
  assign new_n2522_ = new_n3122_ & new_n3123_;
  assign new_n2523_ = new_n3077_ & new_n3075_ & new_n3076_ & new_n3078_;
  assign new_n2524_ = new_n3081_ & new_n3079_ & new_n3080_ & new_n3082_;
  assign new_n2525_ = new_n3085_ & new_n3083_ & new_n3084_ & new_n3086_;
  assign new_n2526_ = new_n3089_ & new_n3088_ & new_n3087_;
  assign new_n2527_ = new_n2525_ & new_n2523_ & new_n2524_ & new_n2526_;
  assign new_n2528_ = new_n3092_ & new_n3090_ & new_n3091_ & new_n3093_;
  assign new_n2529_ = new_n3096_ & new_n3094_ & new_n3095_ & new_n3097_;
  assign new_n2530_ = new_n3100_ & new_n3098_ & new_n3099_ & new_n3101_;
  assign new_n2531_ = new_n3104_ & new_n3103_ & new_n3102_;
  assign new_n2532_ = new_n2530_ & new_n2528_ & new_n2529_ & new_n2531_;
  assign new_n2533_ = new_n4752_ & new_n3106_;
  assign new_n2534_ = new_n4755_ & new_n1949_;
  assign new_n2535_ = new_n3139_ & new_n3138_;
  assign new_n2536_ = new_n3141_ & new_n3140_;
  assign new_n2537_ = new_n2536_ & new_n3143_ & new_n3142_;
  assign new_n2538_ = new_n3145_ & new_n3146_ & new_n3148_ & new_n3147_;
  assign new_n2539_ = new_n3158_ & new_n3157_;
  assign new_n2540_ = new_n3160_ & new_n3159_;
  assign new_n2541_ = new_n2540_ & new_n3162_ & new_n3161_;
  assign new_n2542_ = new_n3164_ & new_n3165_ & new_n3167_ & new_n3166_;
  assign new_n2543_ = new_n3177_ & new_n3176_;
  assign new_n2544_ = new_n3179_ & new_n3178_;
  assign new_n2545_ = new_n2544_ & new_n3181_ & new_n3180_;
  assign new_n2546_ = new_n3183_ & new_n3184_ & new_n3186_ & new_n3185_;
  assign new_n2547_ = new_n3196_ & new_n3195_;
  assign new_n2548_ = new_n3198_ & new_n3197_;
  assign new_n2549_ = new_n2548_ & new_n3200_ & new_n3199_;
  assign new_n2550_ = new_n3202_ & new_n3203_ & new_n3205_ & new_n3204_;
  assign new_n2551_ = new_n3215_ & new_n3214_;
  assign new_n2552_ = new_n3217_ & new_n3216_;
  assign new_n2553_ = new_n2552_ & new_n3219_ & new_n3218_;
  assign new_n2554_ = new_n3221_ & new_n3222_ & new_n3224_ & new_n3223_;
  assign new_n2555_ = new_n3234_ & new_n3233_;
  assign new_n2556_ = new_n3236_ & new_n3235_;
  assign new_n2557_ = new_n2556_ & new_n3238_ & new_n3237_;
  assign new_n2558_ = new_n3240_ & new_n3241_ & new_n3243_ & new_n3242_;
  assign new_n2559_ = new_n3253_ & new_n3252_;
  assign new_n2560_ = new_n3255_ & new_n3254_;
  assign new_n2561_ = new_n2560_ & new_n3257_ & new_n3256_;
  assign new_n2562_ = new_n3259_ & new_n3260_ & new_n3262_ & new_n3261_;
  assign new_n2563_ = new_n3272_ & new_n3271_;
  assign new_n2564_ = new_n3274_ & new_n3273_;
  assign new_n2565_ = new_n2564_ & new_n3276_ & new_n3275_;
  assign new_n2566_ = new_n3278_ & new_n3279_ & new_n3281_ & new_n3280_;
  assign new_n2567_ = new_n3291_ & new_n3290_;
  assign new_n2568_ = new_n3293_ & new_n3292_;
  assign new_n2569_ = new_n2568_ & new_n3295_ & new_n3294_;
  assign new_n2570_ = new_n3297_ & new_n3298_ & new_n3300_ & new_n3299_;
  assign new_n2571_ = new_n3310_ & new_n3309_;
  assign new_n2572_ = new_n3312_ & new_n3311_;
  assign new_n2573_ = new_n2572_ & new_n3314_ & new_n3313_;
  assign new_n2574_ = new_n3316_ & new_n3317_ & new_n3319_ & new_n3318_;
  assign new_n2575_ = new_n3329_ & new_n3328_;
  assign new_n2576_ = new_n3331_ & new_n3330_;
  assign new_n2577_ = new_n2576_ & new_n3333_ & new_n3332_;
  assign new_n2578_ = new_n3337_ & new_n3335_ & new_n3336_ & new_n3338_;
  assign new_n2579_ = new_n3348_ & new_n3347_;
  assign new_n2580_ = new_n3350_ & new_n3349_;
  assign new_n2581_ = new_n2580_ & new_n3352_ & new_n3351_;
  assign new_n2582_ = new_n3355_ & new_n3354_ & new_n3356_ & new_n3357_;
  assign new_n2583_ = new_n3367_ & new_n3366_;
  assign new_n2584_ = new_n3369_ & new_n3368_;
  assign new_n2585_ = new_n2584_ & new_n3371_ & new_n3370_;
  assign new_n2586_ = new_n3375_ & new_n3373_ & new_n3374_ & new_n3376_;
  assign new_n2587_ = new_n3386_ & new_n3385_;
  assign new_n2588_ = new_n3388_ & new_n3387_;
  assign new_n2589_ = new_n2588_ & new_n3390_ & new_n3389_;
  assign new_n2590_ = new_n3393_ & new_n3392_ & new_n3394_ & new_n3395_;
  assign new_n2591_ = new_n3405_ & new_n3404_;
  assign new_n2592_ = new_n3407_ & new_n3406_;
  assign new_n2593_ = new_n2592_ & new_n3409_ & new_n3408_;
  assign new_n2594_ = new_n3411_ & new_n3412_ & new_n3414_ & new_n3413_;
  assign new_n2595_ = new_n3424_ & new_n3423_;
  assign new_n2596_ = new_n3426_ & new_n3425_;
  assign new_n2597_ = new_n2596_ & new_n3428_ & new_n3427_;
  assign new_n2598_ = new_n3430_ & new_n3431_ & new_n3433_ & new_n3432_;
  assign new_n2599_ = new_n3443_ & new_n3442_;
  assign new_n2600_ = new_n3445_ & new_n3444_;
  assign new_n2601_ = new_n2600_ & new_n3447_ & new_n3446_;
  assign new_n2602_ = new_n3450_ & new_n3449_ & new_n3451_ & new_n3452_;
  assign new_n2603_ = new_n3462_ & new_n3461_;
  assign new_n2604_ = new_n3464_ & new_n3463_;
  assign new_n2605_ = new_n2604_ & new_n3466_ & new_n3465_;
  assign new_n2606_ = new_n3469_ & new_n3468_ & new_n3470_ & new_n3471_;
  assign new_n2607_ = new_n3481_ & new_n3480_;
  assign new_n2608_ = new_n3483_ & new_n3482_;
  assign new_n2609_ = new_n2608_ & new_n3485_ & new_n3484_;
  assign new_n2610_ = new_n3487_ & new_n3488_ & new_n3490_ & new_n3489_;
  assign new_n2611_ = new_n3500_ & new_n3499_;
  assign new_n2612_ = new_n3502_ & new_n3501_;
  assign new_n2613_ = new_n2612_ & new_n3504_ & new_n3503_;
  assign new_n2614_ = new_n3506_ & new_n3507_ & new_n3509_ & new_n3508_;
  assign new_n2615_ = new_n3519_ & new_n3518_;
  assign new_n2616_ = new_n3521_ & new_n3520_;
  assign new_n2617_ = new_n2616_ & new_n3523_ & new_n3522_;
  assign new_n2618_ = new_n3525_ & new_n3526_ & new_n3528_ & new_n3527_;
  assign new_n2619_ = new_n3538_ & new_n3537_;
  assign new_n2620_ = new_n3540_ & new_n3539_;
  assign new_n2621_ = new_n2620_ & new_n3542_ & new_n3541_;
  assign new_n2622_ = new_n3544_ & new_n3545_ & new_n3547_ & new_n3546_;
  assign new_n2623_ = new_n3557_ & new_n3556_;
  assign new_n2624_ = new_n3559_ & new_n3558_;
  assign new_n2625_ = new_n2624_ & new_n3561_ & new_n3560_;
  assign new_n2626_ = new_n3563_ & new_n3564_ & new_n3566_ & new_n3565_;
  assign new_n2627_ = new_n3576_ & new_n3575_;
  assign new_n2628_ = new_n3578_ & new_n3577_;
  assign new_n2629_ = new_n2628_ & new_n3580_ & new_n3579_;
  assign new_n2630_ = new_n3582_ & new_n3583_ & new_n3585_ & new_n3584_;
  assign new_n2631_ = new_n3595_ & new_n3594_;
  assign new_n2632_ = new_n3597_ & new_n3596_;
  assign new_n2633_ = new_n2632_ & new_n3599_ & new_n3598_;
  assign new_n2634_ = new_n3601_ & new_n3602_ & new_n3604_ & new_n3603_;
  assign new_n2635_ = new_n3614_ & new_n3613_;
  assign new_n2636_ = new_n3616_ & new_n3615_;
  assign new_n2637_ = new_n2636_ & new_n3618_ & new_n3617_;
  assign new_n2638_ = new_n3620_ & new_n3621_ & new_n3623_ & new_n3622_;
  assign new_n2639_ = new_n3633_ & new_n3632_;
  assign new_n2640_ = new_n3635_ & new_n3634_;
  assign new_n2641_ = new_n2640_ & new_n3637_ & new_n3636_;
  assign new_n2642_ = new_n3639_ & new_n3640_ & new_n3642_ & new_n3641_;
  assign new_n2643_ = new_n3652_ & new_n3651_;
  assign new_n2644_ = new_n3654_ & new_n3653_;
  assign new_n2645_ = new_n2644_ & new_n3656_ & new_n3655_;
  assign new_n2646_ = new_n3658_ & new_n3659_ & new_n3661_ & new_n3660_;
  assign new_n2647_ = new_n3668_ & new_n2957_;
  assign new_n2648_ = new_n3670_ & new_n3673_ & new_n3672_ & new_n3671_ & new_n3669_;
  assign new_n2649_ = new_n3675_ & new_n3674_;
  assign new_n2650_ = new_n2649_ & new_n3677_ & new_n3676_;
  assign new_n2651_ = new_n3679_ & new_n3680_ & new_n3681_;
  assign new_n2652_ = new_n2957_ & new_n3668_;
  assign new_n2653_ = new_n1949_ & new_n2384_;
  assign new_n2654_ = new_n2385_ & new_n4755_ & new_n2939_;
  assign new_n2655_ = new_n3699_ & new_n3698_ & new_n3697_;
  assign new_n2656_ = new_n2884_ & new_n3701_ & new_n3700_;
  assign new_n2657_ = new_n3704_ & new_n3703_ & new_n3702_;
  assign new_n2658_ = new_n2885_ & new_n3706_ & new_n3705_;
  assign new_n2659_ = new_n3709_ & new_n3708_ & new_n3707_;
  assign new_n2660_ = new_n2886_ & new_n3711_ & new_n3710_;
  assign new_n2661_ = new_n3714_ & new_n3713_ & new_n3712_;
  assign new_n2662_ = new_n2887_ & new_n3716_ & new_n3715_;
  assign new_n2663_ = new_n3719_ & new_n3718_ & new_n3717_;
  assign new_n2664_ = new_n2888_ & new_n3721_ & new_n3720_;
  assign new_n2665_ = new_n3724_ & new_n3723_ & new_n3722_;
  assign new_n2666_ = new_n3726_ & new_n3725_;
  assign new_n2667_ = new_n3729_ & new_n3728_ & new_n3727_;
  assign new_n2668_ = new_n3731_ & new_n3730_;
  assign new_n2669_ = new_n3734_ & new_n3733_ & new_n3732_;
  assign new_n2670_ = new_n3736_ & new_n3735_;
  assign new_n2671_ = new_n3739_ & new_n3738_ & new_n3737_;
  assign new_n2672_ = new_n3741_ & new_n3740_;
  assign new_n2673_ = new_n3743_ & new_n3742_;
  assign new_n2674_ = new_n3746_ & new_n3745_;
  assign new_n2675_ = new_n3748_ & new_n3747_;
  assign new_n2676_ = new_n3751_ & new_n3750_;
  assign new_n2677_ = new_n3754_ & new_n3753_ & new_n3752_;
  assign new_n2678_ = new_n3756_ & new_n3755_;
  assign new_n2679_ = new_n3759_ & new_n3758_ & new_n3757_;
  assign new_n2680_ = new_n3761_ & new_n3760_;
  assign new_n2681_ = new_n3764_ & new_n3763_ & new_n3762_;
  assign new_n2682_ = new_n3766_ & new_n3765_;
  assign new_n2683_ = new_n3769_ & new_n3768_ & new_n3767_;
  assign new_n2684_ = new_n3771_ & new_n3770_;
  assign new_n2685_ = new_n3773_ & new_n3772_;
  assign new_n2686_ = new_n3776_ & new_n3775_;
  assign new_n2687_ = new_n3778_ & new_n3777_;
  assign new_n2688_ = new_n3781_ & new_n3780_;
  assign new_n2689_ = new_n3784_ & new_n3783_ & new_n3782_;
  assign new_n2690_ = new_n3786_ & new_n3785_;
  assign new_n2691_ = new_n3789_ & new_n3788_ & new_n3787_;
  assign new_n2692_ = new_n3791_ & new_n3790_;
  assign new_n2693_ = new_n3793_ & new_n3792_;
  assign new_n2694_ = new_n3796_ & new_n3795_;
  assign new_n2695_ = new_n3798_ & new_n3797_;
  assign new_n2696_ = new_n3801_ & new_n3800_;
  assign new_n2697_ = new_n3803_ & new_n3802_;
  assign new_n2698_ = new_n3806_ & new_n3805_;
  assign new_n2699_ = new_n3808_ & new_n3807_;
  assign new_n2700_ = new_n3811_ & new_n3810_;
  assign new_n2701_ = new_n3813_ & new_n3812_;
  assign new_n2702_ = new_n3816_ & new_n3815_;
  assign new_n2703_ = new_n3818_ & new_n3817_;
  assign new_n2704_ = new_n3821_ & new_n3820_;
  assign new_n2705_ = new_n3823_ & new_n3822_;
  assign new_n2706_ = new_n3826_ & new_n3825_;
  assign new_n2707_ = new_n3828_ & new_n3827_;
  assign new_n2708_ = new_n3831_ & new_n3830_;
  assign new_n2709_ = new_n3833_ & new_n3832_;
  assign new_n2710_ = new_n3836_ & new_n3835_;
  assign new_n2711_ = new_n3838_ & new_n3837_;
  assign new_n2712_ = new_n3841_ & new_n3840_;
  assign new_n2713_ = new_n2297_ & new_n2289_ & new_n2291_;
  assign new_n2714_ = new_n2292_ & new_n2293_ & new_n2349_;
  assign new_n2715_ = new_n2288_ & new_n2933_;
  assign new_n2716_ = new_n2715_ & new_n2351_;
  assign new_n2717_ = new_n3861_ & new_n3862_;
  assign new_n2718_ = new_n3864_ & new_n3865_ & new_n3863_;
  assign new_n2719_ = new_n3871_ & new_n3872_;
  assign new_n2720_ = new_n3874_ & new_n3875_ & new_n3873_;
  assign new_n2721_ = new_n3881_ & new_n3882_;
  assign new_n2722_ = new_n3884_ & new_n3885_ & new_n3883_;
  assign new_n2723_ = new_n3891_ & new_n3892_;
  assign new_n2724_ = new_n3894_ & new_n3895_ & new_n3893_;
  assign new_n2725_ = new_n3901_ & new_n3902_;
  assign new_n2726_ = new_n3904_ & new_n3905_ & new_n3903_;
  assign new_n2727_ = new_n3911_ & new_n3912_;
  assign new_n2728_ = new_n3914_ & new_n3915_ & new_n3913_;
  assign new_n2729_ = new_n3921_ & new_n3922_;
  assign new_n2730_ = new_n3924_ & new_n3925_ & new_n3923_;
  assign new_n2731_ = new_n3931_ & new_n3932_;
  assign new_n2732_ = new_n3934_ & new_n3935_ & new_n3933_;
  assign new_n2733_ = new_n3941_ & new_n3942_;
  assign new_n2734_ = new_n3944_ & new_n3945_ & new_n3943_;
  assign new_n2735_ = new_n3951_ & new_n3952_;
  assign new_n2736_ = new_n3954_ & new_n3955_ & new_n3953_;
  assign new_n2737_ = new_n3961_ & new_n3962_;
  assign new_n2738_ = new_n3964_ & new_n3965_ & new_n3963_;
  assign new_n2739_ = new_n3971_ & new_n3972_;
  assign new_n2740_ = new_n3974_ & new_n3975_ & new_n3973_;
  assign new_n2741_ = new_n3981_ & new_n3982_;
  assign new_n2742_ = new_n3984_ & new_n3985_ & new_n3983_;
  assign new_n2743_ = new_n3991_ & new_n3992_;
  assign new_n2744_ = new_n3995_ & new_n3994_ & new_n3993_;
  assign new_n2745_ = new_n4001_ & new_n4002_;
  assign new_n2746_ = new_n4005_ & new_n4004_ & new_n4003_;
  assign new_n2747_ = new_n2748_ & new_n4011_;
  assign new_n2748_ = new_n4012_ & new_n2967_;
  assign new_n2749_ = new_n4015_ & new_n4014_ & new_n4013_;
  assign new_n2750_ = new_n4021_ & new_n4022_;
  assign new_n2751_ = new_n4025_ & new_n4024_ & new_n4023_;
  assign new_n2752_ = new_n2753_ & new_n4031_;
  assign new_n2753_ = new_n4032_ & new_n2967_;
  assign new_n2754_ = new_n4035_ & new_n4034_ & new_n4033_;
  assign new_n2755_ = new_n4041_ & new_n4042_;
  assign new_n2756_ = new_n4045_ & new_n4044_ & new_n4043_;
  assign new_n2757_ = new_n4051_ & new_n4052_;
  assign new_n2758_ = new_n4055_ & new_n4054_ & new_n4053_;
  assign new_n2759_ = new_n5148_ & new_n5145_ & new_n5142_;
  assign new_n2760_ = new_n5160_ & new_n2761_ & new_n2759_;
  assign new_n2761_ = new_n5151_ & new_n5157_ & new_n5154_;
  assign new_n2762_ = new_n5172_ & new_n5169_ & new_n5166_;
  assign new_n2763_ = new_n5181_ & new_n5178_ & new_n5175_;
  assign new_n2764_ = new_n5163_ & new_n2763_ & new_n2762_;
  assign new_n2765_ = new_n5118_ & new_n5115_ & new_n5112_;
  assign new_n2766_ = new_n5130_ & new_n5133_ & new_n5121_ & new_n5124_ & new_n5127_;
  assign new_n2767_ = new_n5193_ & new_n5187_ & new_n5190_ & new_n5196_;
  assign new_n2768_ = new_n5202_ & new_n5199_;
  assign new_n2769_ = new_n2768_ & new_n2767_;
  assign new_n2770_ = new_n2764_ & new_n5136_ & new_n5184_ & new_n5139_ & new_n2760_;
  assign new_n2771_ = new_n5109_ & new_n2766_ & new_n2765_;
  assign new_n2772_ = new_n2356_ & pi275;
  assign new_n2773_ = new_n4065_ & new_n4063_;
  assign new_n2774_ = new_n2384_ & new_n2385_;
  assign new_n2775_ = new_n2923_ & new_n2924_ & new_n2298_;
  assign new_n2776_ = new_n2295_ & new_n2351_;
  assign new_n2777_ = new_n2354_ & new_n2357_;
  assign new_n2778_ = new_n1949_ & new_n4072_;
  assign new_n2779_ = new_n2352_ & pi275;
  assign new_n2780_ = new_n4100_ & new_n4099_;
  assign new_n2781_ = new_n4116_ & new_n4114_;
  assign new_n2782_ = new_n4118_ & new_n4117_;
  assign new_n2783_ = new_n4127_ & new_n4126_;
  assign new_n2784_ = new_n4145_ & new_n4144_;
  assign new_n2785_ = new_n2964_ & new_n2005_;
  assign new_n2786_ = new_n2787_ & new_n4159_ & new_n4158_;
  assign new_n2787_ = new_n4162_ & new_n4161_;
  assign new_n2788_ = new_n4171_ & new_n4170_;
  assign new_n2789_ = new_n4178_ & new_n4176_;
  assign new_n2790_ = new_n4180_ & new_n4179_;
  assign new_n2791_ = new_n4207_ & new_n4206_;
  assign new_n2792_ = new_n4234_ & new_n4233_;
  assign new_n2793_ = new_n4250_ & new_n4248_;
  assign new_n2794_ = new_n4252_ & new_n4251_;
  assign new_n2795_ = new_n4261_ & new_n4260_;
  assign new_n2796_ = new_n4286_ & new_n4284_;
  assign new_n2797_ = new_n4288_ & new_n4287_;
  assign new_n2798_ = new_n4297_ & new_n4296_;
  assign new_n2799_ = new_n4333_ & new_n4332_;
  assign new_n2800_ = new_n4729_ & new_n4720_;
  assign new_n2801_ = new_n2302_ & new_n4337_;
  assign new_n2802_ = new_n4402_ & new_n4403_;
  assign new_n2803_ = new_n4462_ & new_n4460_;
  assign new_n2804_ = new_n2371_ & new_n4465_;
  assign new_n2805_ = new_n2301_ & new_n2924_;
  assign new_n2806_ = new_n2805_ & new_n2298_;
  assign new_n2807_ = new_n2808_ & new_n4473_;
  assign new_n2808_ = new_n2371_ & new_n4471_;
  assign new_n2809_ = new_n2810_ & new_n4476_;
  assign new_n2810_ = new_n2371_ & new_n4474_;
  assign new_n2811_ = new_n2812_ & new_n4479_;
  assign new_n2812_ = new_n2371_ & new_n4477_;
  assign new_n2813_ = new_n2814_ & new_n4482_;
  assign new_n2814_ = new_n2371_ & new_n4480_;
  assign new_n2815_ = new_n2816_ & new_n4485_;
  assign new_n2816_ = new_n2371_ & new_n4483_;
  assign new_n2817_ = new_n2818_ & new_n4488_;
  assign new_n2818_ = new_n2371_ & new_n4486_;
  assign new_n2819_ = new_n4491_ & new_n4489_;
  assign new_n2820_ = new_n4494_ & new_n4492_;
  assign new_n2821_ = new_n2822_ & new_n4497_;
  assign new_n2822_ = new_n2371_ & new_n4495_;
  assign new_n2823_ = new_n2371_ & new_n4500_;
  assign new_n2824_ = new_n2371_ & new_n4503_;
  assign new_n2825_ = new_n2371_ & new_n4506_;
  assign new_n2826_ = new_n2371_ & new_n4509_;
  assign new_n2827_ = new_n2371_ & new_n4512_;
  assign new_n2828_ = new_n2371_ & new_n4515_;
  assign new_n2829_ = new_n2371_ & new_n4518_;
  assign new_n2830_ = new_n2371_ & new_n4521_;
  assign new_n2831_ = new_n2371_ & new_n4524_;
  assign new_n2832_ = new_n2371_ & new_n4527_;
  assign new_n2833_ = new_n2834_ & new_n4530_;
  assign new_n2834_ = new_n2371_ & new_n4528_;
  assign new_n2835_ = new_n2371_ & new_n4533_;
  assign new_n2836_ = new_n2371_ & new_n4536_;
  assign new_n2837_ = new_n2371_ & new_n4539_;
  assign new_n2838_ = new_n2371_ & new_n4542_;
  assign new_n2839_ = new_n2371_ & new_n4545_;
  assign new_n2840_ = new_n2371_ & new_n4548_;
  assign new_n2841_ = new_n2371_ & new_n4551_;
  assign new_n2842_ = new_n2371_ & new_n4554_;
  assign new_n2843_ = new_n2371_ & new_n4557_;
  assign new_n2844_ = new_n2371_ & new_n4560_;
  assign new_n2845_ = new_n2846_ & new_n4563_;
  assign new_n2846_ = new_n2371_ & new_n4561_;
  assign new_n2847_ = new_n2848_ & new_n4566_;
  assign new_n2848_ = new_n2371_ & new_n4564_;
  assign new_n2849_ = new_n4572_ & new_n4569_;
  assign new_n2850_ = new_n4576_ & new_n4573_;
  assign new_n2851_ = new_n4578_ & new_n4577_;
  assign new_n2852_ = new_n4582_ & new_n4581_;
  assign new_n2853_ = new_n4586_ & new_n4585_;
  assign new_n2854_ = new_n4590_ & new_n4589_;
  assign new_n2855_ = new_n4602_ & new_n4600_ & new_n4599_;
  assign new_n2856_ = new_n4604_ & new_n4603_;
  assign new_n2857_ = new_n4608_ & new_n4607_;
  assign new_n2858_ = new_n4612_ & new_n4611_;
  assign new_n2859_ = new_n4616_ & new_n4615_;
  assign new_n2860_ = new_n4620_ & new_n4619_;
  assign new_n2861_ = new_n4624_ & new_n4623_;
  assign new_n2862_ = new_n4628_ & new_n4627_;
  assign new_n2863_ = new_n4632_ & new_n4631_;
  assign new_n2864_ = new_n4636_ & new_n4635_;
  assign new_n2865_ = new_n4640_ & new_n4639_;
  assign new_n2866_ = new_n4646_ & new_n4644_ & new_n4643_;
  assign new_n2867_ = new_n4648_ & new_n4647_;
  assign new_n2868_ = new_n4652_ & new_n4651_;
  assign new_n2869_ = new_n4656_ & new_n4655_;
  assign new_n2870_ = new_n4660_ & new_n4659_;
  assign new_n2871_ = new_n4664_ & new_n4663_;
  assign new_n2872_ = new_n4668_ & new_n4667_;
  assign new_n2873_ = new_n4672_ & new_n4671_;
  assign new_n2874_ = new_n4676_ & new_n4675_;
  assign new_n2875_ = new_n4680_ & new_n4679_;
  assign new_n2876_ = new_n4684_ & new_n4683_;
  assign new_n2877_ = new_n4690_ & new_n4688_ & new_n4687_;
  assign new_n2878_ = new_n4692_ & new_n4691_;
  assign new_n2879_ = ~pi064;
  assign new_n2880_ = ~new_n1949_ | ~new_n2287_;
  assign new_n2881_ = ~new_n4744_ | ~new_n4738_;
  assign new_n2882_ = ~new_n2534_ | ~new_n1973_;
  assign new_n2883_ = ~new_n2653_ | ~new_n1973_;
  assign new_n2884_ = new_n4978_ & new_n4977_;
  assign new_n2885_ = new_n4980_ & new_n4979_;
  assign new_n2886_ = new_n4982_ & new_n4981_;
  assign new_n2887_ = new_n4984_ & new_n4983_;
  assign new_n2888_ = new_n4986_ & new_n4985_;
  assign new_n2889_ = new_n4988_ & new_n4987_;
  assign new_n2890_ = new_n4990_ & new_n4989_;
  assign new_n2891_ = new_n4992_ & new_n4991_;
  assign new_n2892_ = new_n4994_ & new_n4993_;
  assign new_n2893_ = new_n4996_ & new_n4995_;
  assign new_n2894_ = new_n4998_ & new_n4997_;
  assign new_n2895_ = new_n5000_ & new_n4999_;
  assign new_n2896_ = new_n5002_ & new_n5001_;
  assign new_n2897_ = new_n5004_ & new_n5003_;
  assign new_n2898_ = new_n5006_ & new_n5005_;
  assign new_n2899_ = new_n5008_ & new_n5007_;
  assign new_n2900_ = new_n5010_ & new_n5009_;
  assign new_n2901_ = new_n5012_ & new_n5011_;
  assign new_n2902_ = new_n5014_ & new_n5013_;
  assign new_n2903_ = new_n5016_ & new_n5015_;
  assign new_n2904_ = new_n5018_ & new_n5017_;
  assign new_n2905_ = new_n5020_ & new_n5019_;
  assign new_n2906_ = new_n5022_ & new_n5021_;
  assign new_n2907_ = new_n5024_ & new_n5023_;
  assign new_n2908_ = new_n5026_ & new_n5025_;
  assign new_n2909_ = new_n5028_ & new_n5027_;
  assign new_n2910_ = new_n5030_ & new_n5029_;
  assign new_n2911_ = new_n5032_ & new_n5031_;
  assign new_n2912_ = new_n5034_ & new_n5033_;
  assign new_n2913_ = new_n5036_ & new_n5035_;
  assign new_n2914_ = ~new_n2652_ | ~new_n1983_;
  assign new_n2915_ = new_n5038_ & new_n5037_;
  assign new_n2916_ = new_n5040_ & new_n5039_;
  assign new_n2917_ = new_n5106_ & new_n5105_;
  assign new_n2918_ = ~new_n2771_ | ~new_n2769_ | ~new_n2770_;
  assign new_n2919_ = ~new_n2298_;
  assign new_n2920_ = ~new_n2301_;
  assign new_n2921_ = ~new_n2291_;
  assign new_n2922_ = ~new_n2350_;
  assign new_n2923_ = ~new_n2930_ | ~new_n4720_;
  assign new_n2924_ = ~new_n2968_ | ~new_n2378_;
  assign new_n2925_ = ~new_n2346_;
  assign new_n2926_ = ~new_n2969_ | ~new_n4720_;
  assign new_n2927_ = ~new_n2289_;
  assign new_n2928_ = ~new_n2294_;
  assign new_n2929_ = ~new_n2297_;
  assign new_n2930_ = ~new_n2349_;
  assign new_n2931_ = ~new_n2293_;
  assign new_n2932_ = ~new_n2292_;
  assign new_n2933_ = ~new_n2971_ | ~new_n2378_;
  assign new_n2934_ = ~new_n2288_;
  assign new_n2935_ = ~new_n2351_;
  assign new_n2936_ = ~new_n2348_;
  assign new_n2937_ = ~new_n2920_ | ~new_n2380_;
  assign new_n2938_ = ~new_n2295_;
  assign new_n2939_ = ~new_n2957_ | ~new_n2296_;
  assign new_n2940_ = ~new_n2800_ | ~new_n2352_;
  assign new_n2941_ = ~new_n2881_;
  assign new_n2942_ = ~new_n2361_;
  assign po266 = ~new_n2357_;
  assign new_n2944_ = ~new_n2340_;
  assign new_n2945_ = ~new_n2338_;
  assign new_n2946_ = ~new_n2336_;
  assign new_n2947_ = ~new_n2334_;
  assign new_n2948_ = ~new_n2332_;
  assign new_n2949_ = ~new_n2330_;
  assign new_n2950_ = ~new_n2328_;
  assign new_n2951_ = ~new_n2326_;
  assign new_n2952_ = ~new_n2324_;
  assign new_n2953_ = ~new_n2345_;
  assign new_n2954_ = ~new_n2344_;
  assign new_n2955_ = ~new_n2342_;
  assign new_n2956_ = ~new_n2358_;
  assign new_n2957_ = ~new_n2299_;
  assign new_n2958_ = ~new_n2347_;
  assign new_n2959_ = ~new_n2883_;
  assign new_n2960_ = ~new_n2882_;
  assign new_n2961_ = ~new_n2880_;
  assign new_n2962_ = ~new_n2914_;
  assign new_n2963_ = ~new_n2300_;
  assign new_n2964_ = ~new_n2362_;
  assign new_n2965_ = ~new_n2360_;
  assign new_n2966_ = ~new_n2936_ | ~new_n1949_;
  assign new_n2967_ = ~po266 | ~new_n2139_;
  assign new_n2968_ = ~new_n2302_;
  assign new_n2969_ = ~new_n2290_;
  assign new_n2970_ = ~new_n2354_;
  assign new_n2971_ = ~new_n2296_;
  assign new_n2972_ = ~new_n2356_;
  assign new_n2973_ = ~new_n2285_;
  assign new_n2974_ = ~new_n2284_;
  assign new_n2975_ = ~new_n1626_ | ~po264;
  assign new_n2976_ = ~pi033 | ~new_n1956_;
  assign new_n2977_ = ~pi033 | ~new_n2974_;
  assign new_n2978_ = ~new_n1615_ | ~po264;
  assign new_n2979_ = ~new_n13521_ | ~new_n1956_;
  assign new_n2980_ = ~pi034 | ~new_n2974_;
  assign new_n2981_ = ~new_n1604_ | ~po264;
  assign new_n2982_ = ~new_n13502_ | ~new_n1956_;
  assign new_n2983_ = ~pi035 | ~new_n2974_;
  assign new_n2984_ = ~new_n1601_ | ~po264;
  assign new_n2985_ = ~new_n13503_ | ~new_n1956_;
  assign new_n2986_ = ~pi036 | ~new_n2974_;
  assign new_n2987_ = ~new_n1600_ | ~po264;
  assign new_n2988_ = ~new_n13504_ | ~new_n1956_;
  assign new_n2989_ = ~pi037 | ~new_n2974_;
  assign new_n2990_ = ~new_n1599_ | ~po264;
  assign new_n2991_ = ~new_n13643_ | ~new_n1956_;
  assign new_n2992_ = ~pi038 | ~new_n2974_;
  assign new_n2993_ = ~new_n1598_ | ~po264;
  assign new_n2994_ = ~new_n13505_ | ~new_n1956_;
  assign new_n2995_ = ~pi039 | ~new_n2974_;
  assign new_n2996_ = ~new_n1597_ | ~po264;
  assign new_n2997_ = ~new_n13506_ | ~new_n1956_;
  assign new_n2998_ = ~pi040 | ~new_n2974_;
  assign new_n2999_ = ~new_n1596_ | ~po264;
  assign new_n3000_ = ~new_n13507_ | ~new_n1956_;
  assign new_n3001_ = ~pi041 | ~new_n2974_;
  assign new_n3002_ = ~new_n1595_ | ~po264;
  assign new_n3003_ = ~new_n13641_ | ~new_n1956_;
  assign new_n3004_ = ~pi042 | ~new_n2974_;
  assign new_n3005_ = ~new_n1625_ | ~po264;
  assign new_n3006_ = ~new_n13487_ | ~new_n1956_;
  assign new_n3007_ = ~pi043 | ~new_n2974_;
  assign new_n3008_ = ~new_n1624_ | ~po264;
  assign new_n3009_ = ~new_n13488_ | ~new_n1956_;
  assign new_n3010_ = ~pi044 | ~new_n2974_;
  assign new_n3011_ = ~new_n1623_ | ~po264;
  assign new_n3012_ = ~new_n13489_ | ~new_n1956_;
  assign new_n3013_ = ~pi045 | ~new_n2974_;
  assign new_n3014_ = ~new_n1622_ | ~po264;
  assign new_n3015_ = ~new_n13660_ | ~new_n1956_;
  assign new_n3016_ = ~pi046 | ~new_n2974_;
  assign new_n3017_ = ~new_n1621_ | ~po264;
  assign new_n3018_ = ~new_n13490_ | ~new_n1956_;
  assign new_n3019_ = ~pi047 | ~new_n2974_;
  assign new_n3020_ = ~new_n1620_ | ~po264;
  assign new_n3021_ = ~new_n13491_ | ~new_n1956_;
  assign new_n3022_ = ~pi048 | ~new_n2974_;
  assign new_n3023_ = ~new_n1619_ | ~po264;
  assign new_n3024_ = ~new_n13492_ | ~new_n1956_;
  assign new_n3025_ = ~pi049 | ~new_n2974_;
  assign new_n3026_ = ~new_n1618_ | ~po264;
  assign new_n3027_ = ~new_n13658_ | ~new_n1956_;
  assign new_n3028_ = ~pi050 | ~new_n2974_;
  assign new_n3029_ = ~new_n1617_ | ~po264;
  assign new_n3030_ = ~new_n13493_ | ~new_n1956_;
  assign new_n3031_ = ~pi051 | ~new_n2974_;
  assign new_n3032_ = ~new_n1616_ | ~po264;
  assign new_n3033_ = ~new_n13494_ | ~new_n1956_;
  assign new_n3034_ = ~pi052 | ~new_n2974_;
  assign new_n3035_ = ~new_n1614_ | ~po264;
  assign new_n3036_ = ~new_n13495_ | ~new_n1956_;
  assign new_n3037_ = ~pi053 | ~new_n2974_;
  assign new_n3038_ = ~new_n1613_ | ~po264;
  assign new_n3039_ = ~new_n13654_ | ~new_n1956_;
  assign new_n3040_ = ~pi054 | ~new_n2974_;
  assign new_n3041_ = ~new_n1612_ | ~po264;
  assign new_n3042_ = ~new_n13496_ | ~new_n1956_;
  assign new_n3043_ = ~pi055 | ~new_n2974_;
  assign new_n3044_ = ~new_n1611_ | ~po264;
  assign new_n3045_ = ~new_n13497_ | ~new_n1956_;
  assign new_n3046_ = ~pi056 | ~new_n2974_;
  assign new_n3047_ = ~new_n1610_ | ~po264;
  assign new_n3048_ = ~new_n13498_ | ~new_n1956_;
  assign new_n3049_ = ~pi057 | ~new_n2974_;
  assign new_n3050_ = ~new_n1609_ | ~po264;
  assign new_n3051_ = ~new_n13651_ | ~new_n1956_;
  assign new_n3052_ = ~pi058 | ~new_n2974_;
  assign new_n3053_ = ~new_n1608_ | ~po264;
  assign new_n3054_ = ~new_n13499_ | ~new_n1956_;
  assign new_n3055_ = ~pi059 | ~new_n2974_;
  assign new_n3056_ = ~new_n1607_ | ~po264;
  assign new_n3057_ = ~new_n13523_ | ~new_n1956_;
  assign new_n3058_ = ~pi060 | ~new_n2974_;
  assign new_n3059_ = ~new_n1606_ | ~po264;
  assign new_n3060_ = ~new_n13500_ | ~new_n1956_;
  assign new_n3061_ = ~pi061 | ~new_n2974_;
  assign new_n3062_ = ~new_n1605_ | ~po264;
  assign new_n3063_ = ~new_n13501_ | ~new_n1956_;
  assign new_n3064_ = ~pi062 | ~new_n2974_;
  assign new_n3065_ = ~new_n1603_ | ~po264;
  assign new_n3066_ = ~new_n13646_ | ~new_n1956_;
  assign new_n3067_ = ~pi063 | ~new_n2974_;
  assign new_n3068_ = ~new_n1602_ | ~po264;
  assign new_n3069_ = ~new_n13522_ | ~new_n1956_;
  assign new_n3070_ = ~pi064 | ~new_n2974_;
  assign new_n3071_ = ~new_n2287_;
  assign new_n3072_ = ~new_n2352_;
  assign new_n3073_ = ~new_n2285_ | ~new_n4702_;
  assign new_n3074_ = ~new_n2285_ | ~new_n4705_;
  assign new_n3075_ = ~new_n3071_ | ~pi075;
  assign new_n3076_ = ~new_n3071_ | ~pi076;
  assign new_n3077_ = ~new_n3071_ | ~pi077;
  assign new_n3078_ = ~new_n3071_ | ~pi078;
  assign new_n3079_ = ~new_n3071_ | ~pi079;
  assign new_n3080_ = ~new_n3071_ | ~pi080;
  assign new_n3081_ = ~new_n3071_ | ~pi081;
  assign new_n3082_ = ~new_n3071_ | ~pi082;
  assign new_n3083_ = ~new_n3071_ | ~pi083;
  assign new_n3084_ = ~new_n3071_ | ~pi084;
  assign new_n3085_ = ~new_n3071_ | ~pi085;
  assign new_n3086_ = ~new_n3071_ | ~pi086;
  assign new_n3087_ = ~new_n3071_ | ~pi087;
  assign new_n3088_ = ~new_n3071_ | ~pi088;
  assign new_n3089_ = ~new_n3071_ | ~pi089;
  assign new_n3090_ = ~new_n3071_ | ~pi090;
  assign new_n3091_ = ~new_n3071_ | ~pi091;
  assign new_n3092_ = ~new_n3071_ | ~pi092;
  assign new_n3093_ = ~new_n3071_ | ~pi093;
  assign new_n3094_ = ~new_n3071_ | ~pi094;
  assign new_n3095_ = ~new_n3071_ | ~pi067;
  assign new_n3096_ = ~new_n3071_ | ~pi095;
  assign new_n3097_ = ~new_n3071_ | ~pi096;
  assign new_n3098_ = ~new_n3071_ | ~pi068;
  assign new_n3099_ = ~new_n3071_ | ~pi069;
  assign new_n3100_ = ~new_n3071_ | ~pi070;
  assign new_n3101_ = ~new_n3071_ | ~pi071;
  assign new_n3102_ = ~new_n3071_ | ~pi072;
  assign new_n3103_ = ~new_n3071_ | ~pi073;
  assign new_n3104_ = ~new_n3071_ | ~pi074;
  assign new_n3105_ = ~new_n4729_ | ~new_n4726_;
  assign new_n3106_ = ~new_n2296_ | ~new_n4749_ | ~new_n4748_;
  assign new_n3107_ = ~new_n1945_ | ~pi162;
  assign new_n3108_ = ~new_n1946_ | ~pi130;
  assign new_n3109_ = ~new_n1947_ | ~pi098;
  assign new_n3110_ = ~pi265 | ~new_n1944_;
  assign new_n3111_ = ~new_n2005_;
  assign new_n3112_ = ~new_n2346_ | ~new_n2937_;
  assign new_n3113_ = ~new_n2934_ | ~new_n16438_;
  assign new_n3114_ = ~new_n2927_ | ~new_n14710_;
  assign new_n3115_ = ~new_n2921_ | ~new_n17955_;
  assign new_n3116_ = ~new_n2932_ | ~new_n16909_;
  assign new_n3117_ = ~new_n2931_ | ~new_n15375_;
  assign new_n3118_ = ~new_n2938_ | ~new_n17457_;
  assign new_n3119_ = ~new_n2919_ | ~new_n13984_;
  assign new_n3120_ = ~new_n2303_;
  assign new_n3121_ = ~new_n1952_ | ~new_n2005_;
  assign new_n3122_ = ~new_n18453_ | ~new_n1951_;
  assign new_n3123_ = ~new_n2383_ | ~new_n2963_;
  assign new_n3124_ = ~new_n2383_ | ~new_n3112_;
  assign new_n3125_ = ~new_n3121_ | ~new_n3120_ | ~new_n2522_ | ~new_n3124_;
  assign new_n3126_ = ~pi163 | ~new_n1945_;
  assign new_n3127_ = ~pi131 | ~new_n1946_;
  assign new_n3128_ = ~pi099 | ~new_n1947_;
  assign new_n3129_ = ~pi250 | ~new_n1944_;
  assign new_n3130_ = ~new_n1995_;
  assign new_n3131_ = ~pi097 | ~new_n1947_;
  assign new_n3132_ = ~pi129 | ~new_n1946_;
  assign new_n3133_ = ~pi161 | ~new_n1945_;
  assign new_n3134_ = ~pi255 | ~new_n1944_;
  assign new_n3135_ = ~new_n2004_;
  assign new_n3136_ = ~new_n1961_ | ~new_n2004_;
  assign new_n3137_ = ~new_n16515_ | ~new_n2934_;
  assign new_n3138_ = ~new_n14787_ | ~new_n2927_;
  assign new_n3139_ = ~new_n17954_ | ~new_n2921_;
  assign new_n3140_ = ~new_n16986_ | ~new_n2932_;
  assign new_n3141_ = ~new_n15452_ | ~new_n2931_;
  assign new_n3142_ = ~new_n17456_ | ~new_n2938_;
  assign new_n3143_ = ~new_n13983_ | ~new_n2919_;
  assign new_n3144_ = ~new_n2305_;
  assign new_n3145_ = ~new_n1952_ | ~new_n1995_;
  assign new_n3146_ = ~new_n18452_ | ~new_n1951_;
  assign new_n3147_ = ~new_n13788_ | ~new_n2963_;
  assign new_n3148_ = ~new_n2388_ | ~new_n3112_;
  assign new_n3149_ = ~new_n2538_ | ~new_n3144_;
  assign new_n3150_ = ~pi164 | ~new_n1945_;
  assign new_n3151_ = ~pi132 | ~new_n1946_;
  assign new_n3152_ = ~pi100 | ~new_n1947_;
  assign new_n3153_ = ~new_n13032_ | ~new_n1944_;
  assign new_n3154_ = ~new_n1991_;
  assign new_n3155_ = ~new_n1961_ | ~new_n2005_;
  assign new_n3156_ = ~new_n16525_ | ~new_n2934_;
  assign new_n3157_ = ~new_n14797_ | ~new_n2927_;
  assign new_n3158_ = ~new_n17876_ | ~new_n2921_;
  assign new_n3159_ = ~new_n16996_ | ~new_n2932_;
  assign new_n3160_ = ~new_n15462_ | ~new_n2931_;
  assign new_n3161_ = ~new_n17378_ | ~new_n2938_;
  assign new_n3162_ = ~new_n13905_ | ~new_n2919_;
  assign new_n3163_ = ~new_n2306_;
  assign new_n3164_ = ~new_n1952_ | ~new_n1991_;
  assign new_n3165_ = ~new_n18374_ | ~new_n1951_;
  assign new_n3166_ = ~new_n13750_ | ~new_n2963_;
  assign new_n3167_ = ~new_n2391_ | ~new_n3112_;
  assign new_n3168_ = ~new_n2542_ | ~new_n3163_;
  assign new_n3169_ = ~pi165 | ~new_n1945_;
  assign new_n3170_ = ~pi133 | ~new_n1946_;
  assign new_n3171_ = ~pi101 | ~new_n1947_;
  assign new_n3172_ = ~new_n13087_ | ~new_n1944_;
  assign new_n3173_ = ~new_n1987_;
  assign new_n3174_ = ~new_n1961_ | ~new_n1995_;
  assign new_n3175_ = ~new_n16435_ | ~new_n2934_;
  assign new_n3176_ = ~new_n14707_ | ~new_n2927_;
  assign new_n3177_ = ~new_n17960_ | ~new_n2921_;
  assign new_n3178_ = ~new_n16906_ | ~new_n2932_;
  assign new_n3179_ = ~new_n15372_ | ~new_n2931_;
  assign new_n3180_ = ~new_n17462_ | ~new_n2938_;
  assign new_n3181_ = ~new_n13989_ | ~new_n2919_;
  assign new_n3182_ = ~new_n2307_;
  assign new_n3183_ = ~new_n1952_ | ~new_n1987_;
  assign new_n3184_ = ~new_n18458_ | ~new_n1951_;
  assign new_n3185_ = ~new_n13752_ | ~new_n2963_;
  assign new_n3186_ = ~new_n2394_ | ~new_n3112_;
  assign new_n3187_ = ~new_n2546_ | ~new_n3182_;
  assign new_n3188_ = ~pi166 | ~new_n1945_;
  assign new_n3189_ = ~pi134 | ~new_n1946_;
  assign new_n3190_ = ~pi102 | ~new_n1947_;
  assign new_n3191_ = ~new_n13086_ | ~new_n1944_;
  assign new_n3192_ = ~new_n1994_;
  assign new_n3193_ = ~new_n1961_ | ~new_n1991_;
  assign new_n3194_ = ~new_n16524_ | ~new_n2934_;
  assign new_n3195_ = ~new_n14796_ | ~new_n2927_;
  assign new_n3196_ = ~new_n17959_ | ~new_n2921_;
  assign new_n3197_ = ~new_n16995_ | ~new_n2932_;
  assign new_n3198_ = ~new_n15461_ | ~new_n2931_;
  assign new_n3199_ = ~new_n17461_ | ~new_n2938_;
  assign new_n3200_ = ~new_n13988_ | ~new_n2919_;
  assign new_n3201_ = ~new_n2308_;
  assign new_n3202_ = ~new_n1952_ | ~new_n1994_;
  assign new_n3203_ = ~new_n18457_ | ~new_n1951_;
  assign new_n3204_ = ~new_n13753_ | ~new_n2963_;
  assign new_n3205_ = ~new_n2397_ | ~new_n3112_;
  assign new_n3206_ = ~new_n2550_ | ~new_n3201_;
  assign new_n3207_ = ~pi167 | ~new_n1945_;
  assign new_n3208_ = ~pi135 | ~new_n1946_;
  assign new_n3209_ = ~pi103 | ~new_n1947_;
  assign new_n3210_ = ~new_n13085_ | ~new_n1944_;
  assign new_n3211_ = ~new_n1998_;
  assign new_n3212_ = ~new_n1961_ | ~new_n1987_;
  assign new_n3213_ = ~new_n16523_ | ~new_n2934_;
  assign new_n3214_ = ~new_n14795_ | ~new_n2927_;
  assign new_n3215_ = ~new_n17877_ | ~new_n2921_;
  assign new_n3216_ = ~new_n16994_ | ~new_n2932_;
  assign new_n3217_ = ~new_n15460_ | ~new_n2931_;
  assign new_n3218_ = ~new_n17379_ | ~new_n2938_;
  assign new_n3219_ = ~new_n13906_ | ~new_n2919_;
  assign new_n3220_ = ~new_n2309_;
  assign new_n3221_ = ~new_n1952_ | ~new_n1998_;
  assign new_n3222_ = ~new_n18375_ | ~new_n1951_;
  assign new_n3223_ = ~new_n13797_ | ~new_n2963_;
  assign new_n3224_ = ~new_n2400_ | ~new_n3112_;
  assign new_n3225_ = ~new_n2554_ | ~new_n3220_;
  assign new_n3226_ = ~pi168 | ~new_n1945_;
  assign new_n3227_ = ~pi136 | ~new_n1946_;
  assign new_n3228_ = ~pi104 | ~new_n1947_;
  assign new_n3229_ = ~new_n13084_ | ~new_n1944_;
  assign new_n3230_ = ~new_n1997_;
  assign new_n3231_ = ~new_n1961_ | ~new_n1994_;
  assign new_n3232_ = ~new_n16436_ | ~new_n2934_;
  assign new_n3233_ = ~new_n14708_ | ~new_n2927_;
  assign new_n3234_ = ~new_n17958_ | ~new_n2921_;
  assign new_n3235_ = ~new_n16907_ | ~new_n2932_;
  assign new_n3236_ = ~new_n15373_ | ~new_n2931_;
  assign new_n3237_ = ~new_n17460_ | ~new_n2938_;
  assign new_n3238_ = ~new_n13987_ | ~new_n2919_;
  assign new_n3239_ = ~new_n2310_;
  assign new_n3240_ = ~new_n1952_ | ~new_n1997_;
  assign new_n3241_ = ~new_n18456_ | ~new_n1951_;
  assign new_n3242_ = ~new_n13754_ | ~new_n2963_;
  assign new_n3243_ = ~new_n2403_ | ~new_n3112_;
  assign new_n3244_ = ~new_n2558_ | ~new_n3239_;
  assign new_n3245_ = ~pi169 | ~new_n1945_;
  assign new_n3246_ = ~pi137 | ~new_n1946_;
  assign new_n3247_ = ~pi105 | ~new_n1947_;
  assign new_n3248_ = ~new_n13083_ | ~new_n1944_;
  assign new_n3249_ = ~new_n2011_;
  assign new_n3250_ = ~new_n1961_ | ~new_n1998_;
  assign new_n3251_ = ~new_n16522_ | ~new_n2934_;
  assign new_n3252_ = ~new_n14794_ | ~new_n2927_;
  assign new_n3253_ = ~new_n17878_ | ~new_n2921_;
  assign new_n3254_ = ~new_n16993_ | ~new_n2932_;
  assign new_n3255_ = ~new_n15459_ | ~new_n2931_;
  assign new_n3256_ = ~new_n17380_ | ~new_n2938_;
  assign new_n3257_ = ~new_n13907_ | ~new_n2919_;
  assign new_n3258_ = ~new_n2311_;
  assign new_n3259_ = ~new_n1952_ | ~new_n2011_;
  assign new_n3260_ = ~new_n18376_ | ~new_n1951_;
  assign new_n3261_ = ~new_n13755_ | ~new_n2963_;
  assign new_n3262_ = ~new_n2406_ | ~new_n3112_;
  assign new_n3263_ = ~new_n2562_ | ~new_n3258_;
  assign new_n3264_ = ~pi170 | ~new_n1945_;
  assign new_n3265_ = ~pi138 | ~new_n1946_;
  assign new_n3266_ = ~pi106 | ~new_n1947_;
  assign new_n3267_ = ~new_n13082_ | ~new_n1944_;
  assign new_n3268_ = ~new_n2010_;
  assign new_n3269_ = ~new_n1961_ | ~new_n1997_;
  assign new_n3270_ = ~new_n16437_ | ~new_n2934_;
  assign new_n3271_ = ~new_n14709_ | ~new_n2927_;
  assign new_n3272_ = ~new_n17957_ | ~new_n2921_;
  assign new_n3273_ = ~new_n16908_ | ~new_n2932_;
  assign new_n3274_ = ~new_n15374_ | ~new_n2931_;
  assign new_n3275_ = ~new_n17459_ | ~new_n2938_;
  assign new_n3276_ = ~new_n13986_ | ~new_n2919_;
  assign new_n3277_ = ~new_n2312_;
  assign new_n3278_ = ~new_n1952_ | ~new_n2010_;
  assign new_n3279_ = ~new_n18455_ | ~new_n1951_;
  assign new_n3280_ = ~new_n13756_ | ~new_n2963_;
  assign new_n3281_ = ~new_n2409_ | ~new_n3112_;
  assign new_n3282_ = ~new_n2566_ | ~new_n3277_;
  assign new_n3283_ = ~pi171 | ~new_n1945_;
  assign new_n3284_ = ~pi139 | ~new_n1946_;
  assign new_n3285_ = ~pi107 | ~new_n1947_;
  assign new_n3286_ = ~new_n13106_ | ~new_n1944_;
  assign new_n3287_ = ~new_n1989_;
  assign new_n3288_ = ~new_n1961_ | ~new_n2011_;
  assign new_n3289_ = ~new_n16521_ | ~new_n2934_;
  assign new_n3290_ = ~new_n14793_ | ~new_n2927_;
  assign new_n3291_ = ~new_n17956_ | ~new_n2921_;
  assign new_n3292_ = ~new_n16992_ | ~new_n2932_;
  assign new_n3293_ = ~new_n15458_ | ~new_n2931_;
  assign new_n3294_ = ~new_n17458_ | ~new_n2938_;
  assign new_n3295_ = ~new_n13985_ | ~new_n2919_;
  assign new_n3296_ = ~new_n2313_;
  assign new_n3297_ = ~new_n1952_ | ~new_n1989_;
  assign new_n3298_ = ~new_n18454_ | ~new_n1951_;
  assign new_n3299_ = ~new_n13795_ | ~new_n2963_;
  assign new_n3300_ = ~new_n2412_ | ~new_n3112_;
  assign new_n3301_ = ~new_n2570_ | ~new_n3296_;
  assign new_n3302_ = ~pi172 | ~new_n1945_;
  assign new_n3303_ = ~pi140 | ~new_n1946_;
  assign new_n3304_ = ~pi108 | ~new_n1947_;
  assign new_n3305_ = ~new_n13105_ | ~new_n1944_;
  assign new_n3306_ = ~new_n1990_;
  assign new_n3307_ = ~new_n1961_ | ~new_n2010_;
  assign new_n3308_ = ~new_n16531_ | ~new_n2934_;
  assign new_n3309_ = ~new_n14803_ | ~new_n2927_;
  assign new_n3310_ = ~new_n17870_ | ~new_n2921_;
  assign new_n3311_ = ~new_n17002_ | ~new_n2932_;
  assign new_n3312_ = ~new_n15468_ | ~new_n2931_;
  assign new_n3313_ = ~new_n17372_ | ~new_n2938_;
  assign new_n3314_ = ~new_n13899_ | ~new_n2919_;
  assign new_n3315_ = ~new_n2314_;
  assign new_n3316_ = ~new_n1952_ | ~new_n1990_;
  assign new_n3317_ = ~new_n18368_ | ~new_n1951_;
  assign new_n3318_ = ~new_n13738_ | ~new_n2963_;
  assign new_n3319_ = ~new_n2415_ | ~new_n3112_;
  assign new_n3320_ = ~new_n2574_ | ~new_n3315_;
  assign new_n3321_ = ~pi173 | ~new_n1945_;
  assign new_n3322_ = ~pi141 | ~new_n1946_;
  assign new_n3323_ = ~pi109 | ~new_n1947_;
  assign new_n3324_ = ~new_n13104_ | ~new_n1944_;
  assign new_n3325_ = ~new_n1999_;
  assign new_n3326_ = ~new_n1961_ | ~new_n1989_;
  assign new_n3327_ = ~new_n16430_ | ~new_n2934_;
  assign new_n3328_ = ~new_n14702_ | ~new_n2927_;
  assign new_n3329_ = ~new_n17974_ | ~new_n2921_;
  assign new_n3330_ = ~new_n16901_ | ~new_n2932_;
  assign new_n3331_ = ~new_n15367_ | ~new_n2931_;
  assign new_n3332_ = ~new_n17476_ | ~new_n2938_;
  assign new_n3333_ = ~new_n14003_ | ~new_n2919_;
  assign new_n3334_ = ~new_n2315_;
  assign new_n3335_ = ~new_n1952_ | ~new_n1999_;
  assign new_n3336_ = ~new_n18472_ | ~new_n1951_;
  assign new_n3337_ = ~new_n13739_ | ~new_n2963_;
  assign new_n3338_ = ~new_n2418_ | ~new_n3112_;
  assign new_n3339_ = ~new_n2578_ | ~new_n3334_;
  assign new_n3340_ = ~pi174 | ~new_n1945_;
  assign new_n3341_ = ~pi142 | ~new_n1946_;
  assign new_n3342_ = ~pi110 | ~new_n1947_;
  assign new_n3343_ = ~new_n13103_ | ~new_n1944_;
  assign new_n3344_ = ~new_n2007_;
  assign new_n3345_ = ~new_n1961_ | ~new_n1990_;
  assign new_n3346_ = ~new_n16520_ | ~new_n2934_;
  assign new_n3347_ = ~new_n14792_ | ~new_n2927_;
  assign new_n3348_ = ~new_n17973_ | ~new_n2921_;
  assign new_n3349_ = ~new_n16991_ | ~new_n2932_;
  assign new_n3350_ = ~new_n15457_ | ~new_n2931_;
  assign new_n3351_ = ~new_n17475_ | ~new_n2938_;
  assign new_n3352_ = ~new_n14002_ | ~new_n2919_;
  assign new_n3353_ = ~new_n2316_;
  assign new_n3354_ = ~new_n1952_ | ~new_n2007_;
  assign new_n3355_ = ~new_n18471_ | ~new_n1951_;
  assign new_n3356_ = ~new_n13740_ | ~new_n2963_;
  assign new_n3357_ = ~new_n2421_ | ~new_n3112_;
  assign new_n3358_ = ~new_n2582_ | ~new_n3353_;
  assign new_n3359_ = ~pi175 | ~new_n1945_;
  assign new_n3360_ = ~pi143 | ~new_n1946_;
  assign new_n3361_ = ~pi111 | ~new_n1947_;
  assign new_n3362_ = ~new_n13102_ | ~new_n1944_;
  assign new_n3363_ = ~new_n2006_;
  assign new_n3364_ = ~new_n1961_ | ~new_n1999_;
  assign new_n3365_ = ~new_n16519_ | ~new_n2934_;
  assign new_n3366_ = ~new_n14791_ | ~new_n2927_;
  assign new_n3367_ = ~new_n17871_ | ~new_n2921_;
  assign new_n3368_ = ~new_n16990_ | ~new_n2932_;
  assign new_n3369_ = ~new_n15456_ | ~new_n2931_;
  assign new_n3370_ = ~new_n17373_ | ~new_n2938_;
  assign new_n3371_ = ~new_n13900_ | ~new_n2919_;
  assign new_n3372_ = ~new_n2317_;
  assign new_n3373_ = ~new_n1952_ | ~new_n2006_;
  assign new_n3374_ = ~new_n18369_ | ~new_n1951_;
  assign new_n3375_ = ~new_n13818_ | ~new_n2963_;
  assign new_n3376_ = ~new_n2424_ | ~new_n3112_;
  assign new_n3377_ = ~new_n2586_ | ~new_n3372_;
  assign new_n3378_ = ~pi176 | ~new_n1945_;
  assign new_n3379_ = ~pi144 | ~new_n1946_;
  assign new_n3380_ = ~pi112 | ~new_n1947_;
  assign new_n3381_ = ~new_n13101_ | ~new_n1944_;
  assign new_n3382_ = ~new_n2001_;
  assign new_n3383_ = ~new_n1961_ | ~new_n2007_;
  assign new_n3384_ = ~new_n16530_ | ~new_n2934_;
  assign new_n3385_ = ~new_n14802_ | ~new_n2927_;
  assign new_n3386_ = ~new_n17972_ | ~new_n2921_;
  assign new_n3387_ = ~new_n17001_ | ~new_n2932_;
  assign new_n3388_ = ~new_n15467_ | ~new_n2931_;
  assign new_n3389_ = ~new_n17474_ | ~new_n2938_;
  assign new_n3390_ = ~new_n14001_ | ~new_n2919_;
  assign new_n3391_ = ~new_n2318_;
  assign new_n3392_ = ~new_n1952_ | ~new_n2001_;
  assign new_n3393_ = ~new_n18470_ | ~new_n1951_;
  assign new_n3394_ = ~new_n13741_ | ~new_n2963_;
  assign new_n3395_ = ~new_n2427_ | ~new_n3112_;
  assign new_n3396_ = ~new_n2590_ | ~new_n3391_;
  assign new_n3397_ = ~pi177 | ~new_n1945_;
  assign new_n3398_ = ~pi145 | ~new_n1946_;
  assign new_n3399_ = ~pi113 | ~new_n1947_;
  assign new_n3400_ = ~new_n13100_ | ~new_n1944_;
  assign new_n3401_ = ~new_n2000_;
  assign new_n3402_ = ~new_n1961_ | ~new_n2006_;
  assign new_n3403_ = ~new_n16529_ | ~new_n2934_;
  assign new_n3404_ = ~new_n14801_ | ~new_n2927_;
  assign new_n3405_ = ~new_n17971_ | ~new_n2921_;
  assign new_n3406_ = ~new_n17000_ | ~new_n2932_;
  assign new_n3407_ = ~new_n15466_ | ~new_n2931_;
  assign new_n3408_ = ~new_n17473_ | ~new_n2938_;
  assign new_n3409_ = ~new_n14000_ | ~new_n2919_;
  assign new_n3410_ = ~new_n2319_;
  assign new_n3411_ = ~new_n1952_ | ~new_n2000_;
  assign new_n3412_ = ~new_n18469_ | ~new_n1951_;
  assign new_n3413_ = ~new_n13742_ | ~new_n2963_;
  assign new_n3414_ = ~new_n2430_ | ~new_n3112_;
  assign new_n3415_ = ~new_n2594_ | ~new_n3410_;
  assign new_n3416_ = ~pi178 | ~new_n1945_;
  assign new_n3417_ = ~pi146 | ~new_n1946_;
  assign new_n3418_ = ~pi114 | ~new_n1947_;
  assign new_n3419_ = ~new_n13099_ | ~new_n1944_;
  assign new_n3420_ = ~new_n1996_;
  assign new_n3421_ = ~new_n1961_ | ~new_n2001_;
  assign new_n3422_ = ~new_n16431_ | ~new_n2934_;
  assign new_n3423_ = ~new_n14703_ | ~new_n2927_;
  assign new_n3424_ = ~new_n17970_ | ~new_n2921_;
  assign new_n3425_ = ~new_n16902_ | ~new_n2932_;
  assign new_n3426_ = ~new_n15368_ | ~new_n2931_;
  assign new_n3427_ = ~new_n17472_ | ~new_n2938_;
  assign new_n3428_ = ~new_n13999_ | ~new_n2919_;
  assign new_n3429_ = ~new_n2320_;
  assign new_n3430_ = ~new_n1952_ | ~new_n1996_;
  assign new_n3431_ = ~new_n18468_ | ~new_n1951_;
  assign new_n3432_ = ~new_n13743_ | ~new_n2963_;
  assign new_n3433_ = ~new_n2433_ | ~new_n3112_;
  assign new_n3434_ = ~new_n2598_ | ~new_n3429_;
  assign new_n3435_ = ~pi179 | ~new_n1945_;
  assign new_n3436_ = ~pi147 | ~new_n1946_;
  assign new_n3437_ = ~pi115 | ~new_n1947_;
  assign new_n3438_ = ~new_n13098_ | ~new_n1944_;
  assign new_n3439_ = ~new_n2009_;
  assign new_n3440_ = ~new_n1961_ | ~new_n2000_;
  assign new_n3441_ = ~new_n16518_ | ~new_n2934_;
  assign new_n3442_ = ~new_n14790_ | ~new_n2927_;
  assign new_n3443_ = ~new_n17872_ | ~new_n2921_;
  assign new_n3444_ = ~new_n16989_ | ~new_n2932_;
  assign new_n3445_ = ~new_n15455_ | ~new_n2931_;
  assign new_n3446_ = ~new_n17374_ | ~new_n2938_;
  assign new_n3447_ = ~new_n13901_ | ~new_n2919_;
  assign new_n3448_ = ~new_n2321_;
  assign new_n3449_ = ~new_n1952_ | ~new_n2009_;
  assign new_n3450_ = ~new_n18370_ | ~new_n1951_;
  assign new_n3451_ = ~new_n13816_ | ~new_n2963_;
  assign new_n3452_ = ~new_n2436_ | ~new_n3112_;
  assign new_n3453_ = ~new_n2602_ | ~new_n3448_;
  assign new_n3454_ = ~pi180 | ~new_n1945_;
  assign new_n3455_ = ~pi148 | ~new_n1946_;
  assign new_n3456_ = ~pi116 | ~new_n1947_;
  assign new_n3457_ = ~new_n13097_ | ~new_n1944_;
  assign new_n3458_ = ~new_n2008_;
  assign new_n3459_ = ~new_n1961_ | ~new_n1996_;
  assign new_n3460_ = ~new_n16517_ | ~new_n2934_;
  assign new_n3461_ = ~new_n14789_ | ~new_n2927_;
  assign new_n3462_ = ~new_n17969_ | ~new_n2921_;
  assign new_n3463_ = ~new_n16988_ | ~new_n2932_;
  assign new_n3464_ = ~new_n15454_ | ~new_n2931_;
  assign new_n3465_ = ~new_n17471_ | ~new_n2938_;
  assign new_n3466_ = ~new_n13998_ | ~new_n2919_;
  assign new_n3467_ = ~new_n2322_;
  assign new_n3468_ = ~new_n1952_ | ~new_n2008_;
  assign new_n3469_ = ~new_n18467_ | ~new_n1951_;
  assign new_n3470_ = ~new_n13744_ | ~new_n2963_;
  assign new_n3471_ = ~new_n2439_ | ~new_n3112_;
  assign new_n3472_ = ~new_n2606_ | ~new_n3467_;
  assign new_n3473_ = ~pi181 | ~new_n1945_;
  assign new_n3474_ = ~pi149 | ~new_n1946_;
  assign new_n3475_ = ~pi117 | ~new_n1947_;
  assign new_n3476_ = ~new_n13096_ | ~new_n1944_;
  assign new_n3477_ = ~new_n2003_;
  assign new_n3478_ = ~new_n1961_ | ~new_n2009_;
  assign new_n3479_ = ~new_n16516_ | ~new_n2934_;
  assign new_n3480_ = ~new_n14788_ | ~new_n2927_;
  assign new_n3481_ = ~new_n17968_ | ~new_n2921_;
  assign new_n3482_ = ~new_n16987_ | ~new_n2932_;
  assign new_n3483_ = ~new_n15453_ | ~new_n2931_;
  assign new_n3484_ = ~new_n17470_ | ~new_n2938_;
  assign new_n3485_ = ~new_n13997_ | ~new_n2919_;
  assign new_n3486_ = ~new_n2323_;
  assign new_n3487_ = ~new_n1952_ | ~new_n2003_;
  assign new_n3488_ = ~new_n18466_ | ~new_n1951_;
  assign new_n3489_ = ~new_n13814_ | ~new_n2963_;
  assign new_n3490_ = ~new_n2441_ | ~new_n3112_;
  assign new_n3491_ = ~new_n2610_ | ~new_n3486_;
  assign new_n3492_ = ~pi182 | ~new_n1945_;
  assign new_n3493_ = ~pi150 | ~new_n1946_;
  assign new_n3494_ = ~pi118 | ~new_n1947_;
  assign new_n3495_ = ~new_n13095_ | ~new_n1944_;
  assign new_n3496_ = ~new_n2002_;
  assign new_n3497_ = ~new_n1961_ | ~new_n2008_;
  assign new_n3498_ = ~new_n16514_ | ~new_n2934_;
  assign new_n3499_ = ~new_n14786_ | ~new_n2927_;
  assign new_n3500_ = ~new_n17873_ | ~new_n2921_;
  assign new_n3501_ = ~new_n16985_ | ~new_n2932_;
  assign new_n3502_ = ~new_n15451_ | ~new_n2931_;
  assign new_n3503_ = ~new_n17375_ | ~new_n2938_;
  assign new_n3504_ = ~new_n13902_ | ~new_n2919_;
  assign new_n3505_ = ~new_n2325_;
  assign new_n3506_ = ~new_n1952_ | ~new_n2002_;
  assign new_n3507_ = ~new_n18371_ | ~new_n1951_;
  assign new_n3508_ = ~new_n13745_ | ~new_n2963_;
  assign new_n3509_ = ~new_n2952_ | ~new_n3112_;
  assign new_n3510_ = ~new_n2614_ | ~new_n3505_;
  assign new_n3511_ = ~pi183 | ~new_n1945_;
  assign new_n3512_ = ~pi151 | ~new_n1946_;
  assign new_n3513_ = ~pi119 | ~new_n1947_;
  assign new_n3514_ = ~new_n13094_ | ~new_n1944_;
  assign new_n3515_ = ~new_n1988_;
  assign new_n3516_ = ~new_n1961_ | ~new_n2003_;
  assign new_n3517_ = ~new_n16528_ | ~new_n2934_;
  assign new_n3518_ = ~new_n14800_ | ~new_n2927_;
  assign new_n3519_ = ~new_n17874_ | ~new_n2921_;
  assign new_n3520_ = ~new_n16999_ | ~new_n2932_;
  assign new_n3521_ = ~new_n15465_ | ~new_n2931_;
  assign new_n3522_ = ~new_n17376_ | ~new_n2938_;
  assign new_n3523_ = ~new_n13903_ | ~new_n2919_;
  assign new_n3524_ = ~new_n2327_;
  assign new_n3525_ = ~new_n1952_ | ~new_n1988_;
  assign new_n3526_ = ~new_n18372_ | ~new_n1951_;
  assign new_n3527_ = ~new_n13810_ | ~new_n2963_;
  assign new_n3528_ = ~new_n2951_ | ~new_n3112_;
  assign new_n3529_ = ~new_n2618_ | ~new_n3524_;
  assign new_n3530_ = ~pi184 | ~new_n1945_;
  assign new_n3531_ = ~pi152 | ~new_n1946_;
  assign new_n3532_ = ~pi120 | ~new_n1947_;
  assign new_n3533_ = ~new_n13093_ | ~new_n1944_;
  assign new_n3534_ = ~new_n1993_;
  assign new_n3535_ = ~new_n1961_ | ~new_n2002_;
  assign new_n3536_ = ~new_n16527_ | ~new_n2934_;
  assign new_n3537_ = ~new_n14799_ | ~new_n2927_;
  assign new_n3538_ = ~new_n17967_ | ~new_n2921_;
  assign new_n3539_ = ~new_n16998_ | ~new_n2932_;
  assign new_n3540_ = ~new_n15464_ | ~new_n2931_;
  assign new_n3541_ = ~new_n17469_ | ~new_n2938_;
  assign new_n3542_ = ~new_n13996_ | ~new_n2919_;
  assign new_n3543_ = ~new_n2329_;
  assign new_n3544_ = ~new_n1952_ | ~new_n1993_;
  assign new_n3545_ = ~new_n18465_ | ~new_n1951_;
  assign new_n3546_ = ~new_n13746_ | ~new_n2963_;
  assign new_n3547_ = ~new_n2950_ | ~new_n3112_;
  assign new_n3548_ = ~new_n2622_ | ~new_n3543_;
  assign new_n3549_ = ~pi185 | ~new_n1945_;
  assign new_n3550_ = ~pi153 | ~new_n1946_;
  assign new_n3551_ = ~pi121 | ~new_n1947_;
  assign new_n3552_ = ~new_n13092_ | ~new_n1944_;
  assign new_n3553_ = ~new_n1992_;
  assign new_n3554_ = ~new_n1961_ | ~new_n1988_;
  assign new_n3555_ = ~new_n16432_ | ~new_n2934_;
  assign new_n3556_ = ~new_n14704_ | ~new_n2927_;
  assign new_n3557_ = ~new_n17966_ | ~new_n2921_;
  assign new_n3558_ = ~new_n16903_ | ~new_n2932_;
  assign new_n3559_ = ~new_n15369_ | ~new_n2931_;
  assign new_n3560_ = ~new_n17468_ | ~new_n2938_;
  assign new_n3561_ = ~new_n13995_ | ~new_n2919_;
  assign new_n3562_ = ~new_n2331_;
  assign new_n3563_ = ~new_n1952_ | ~new_n1992_;
  assign new_n3564_ = ~new_n18464_ | ~new_n1951_;
  assign new_n3565_ = ~new_n13808_ | ~new_n2963_;
  assign new_n3566_ = ~new_n2949_ | ~new_n3112_;
  assign new_n3567_ = ~new_n2626_ | ~new_n3562_;
  assign new_n3568_ = ~pi186 | ~new_n1945_;
  assign new_n3569_ = ~pi154 | ~new_n1946_;
  assign new_n3570_ = ~pi122 | ~new_n1947_;
  assign new_n3571_ = ~new_n13091_ | ~new_n1944_;
  assign new_n3572_ = ~new_n1985_;
  assign new_n3573_ = ~new_n1961_ | ~new_n1993_;
  assign new_n3574_ = ~new_n16513_ | ~new_n2934_;
  assign new_n3575_ = ~new_n14785_ | ~new_n2927_;
  assign new_n3576_ = ~new_n17965_ | ~new_n2921_;
  assign new_n3577_ = ~new_n16984_ | ~new_n2932_;
  assign new_n3578_ = ~new_n15450_ | ~new_n2931_;
  assign new_n3579_ = ~new_n17467_ | ~new_n2938_;
  assign new_n3580_ = ~new_n13994_ | ~new_n2919_;
  assign new_n3581_ = ~new_n2333_;
  assign new_n3582_ = ~new_n1952_ | ~new_n1985_;
  assign new_n3583_ = ~new_n18463_ | ~new_n1951_;
  assign new_n3584_ = ~new_n13747_ | ~new_n2963_;
  assign new_n3585_ = ~new_n2948_ | ~new_n3112_;
  assign new_n3586_ = ~new_n2630_ | ~new_n3581_;
  assign new_n3587_ = ~pi187 | ~new_n1945_;
  assign new_n3588_ = ~pi155 | ~new_n1946_;
  assign new_n3589_ = ~pi123 | ~new_n1947_;
  assign new_n3590_ = ~new_n13090_ | ~new_n1944_;
  assign new_n3591_ = ~new_n1984_;
  assign new_n3592_ = ~new_n1961_ | ~new_n1992_;
  assign new_n3593_ = ~new_n16512_ | ~new_n2934_;
  assign new_n3594_ = ~new_n14784_ | ~new_n2927_;
  assign new_n3595_ = ~new_n17964_ | ~new_n2921_;
  assign new_n3596_ = ~new_n16983_ | ~new_n2932_;
  assign new_n3597_ = ~new_n15449_ | ~new_n2931_;
  assign new_n3598_ = ~new_n17466_ | ~new_n2938_;
  assign new_n3599_ = ~new_n13993_ | ~new_n2919_;
  assign new_n3600_ = ~new_n2335_;
  assign new_n3601_ = ~new_n1952_ | ~new_n1984_;
  assign new_n3602_ = ~new_n18462_ | ~new_n1951_;
  assign new_n3603_ = ~new_n13806_ | ~new_n2963_;
  assign new_n3604_ = ~new_n2947_ | ~new_n3112_;
  assign new_n3605_ = ~new_n2634_ | ~new_n3600_;
  assign new_n3606_ = ~pi188 | ~new_n1945_;
  assign new_n3607_ = ~pi156 | ~new_n1946_;
  assign new_n3608_ = ~pi124 | ~new_n1947_;
  assign new_n3609_ = ~new_n13089_ | ~new_n1944_;
  assign new_n3610_ = ~new_n1980_;
  assign new_n3611_ = ~new_n1961_ | ~new_n1985_;
  assign new_n3612_ = ~new_n16526_ | ~new_n2934_;
  assign new_n3613_ = ~new_n14798_ | ~new_n2927_;
  assign new_n3614_ = ~new_n17875_ | ~new_n2921_;
  assign new_n3615_ = ~new_n16997_ | ~new_n2932_;
  assign new_n3616_ = ~new_n15463_ | ~new_n2931_;
  assign new_n3617_ = ~new_n17377_ | ~new_n2938_;
  assign new_n3618_ = ~new_n13904_ | ~new_n2919_;
  assign new_n3619_ = ~new_n2337_;
  assign new_n3620_ = ~new_n1952_ | ~new_n1980_;
  assign new_n3621_ = ~new_n18373_ | ~new_n1951_;
  assign new_n3622_ = ~new_n13748_ | ~new_n2963_;
  assign new_n3623_ = ~new_n2946_ | ~new_n3112_;
  assign new_n3624_ = ~new_n2638_ | ~new_n3619_;
  assign new_n3625_ = ~pi189 | ~new_n1945_;
  assign new_n3626_ = ~pi157 | ~new_n1946_;
  assign new_n3627_ = ~pi125 | ~new_n1947_;
  assign new_n3628_ = ~new_n13088_ | ~new_n1944_;
  assign new_n3629_ = ~new_n1981_;
  assign new_n3630_ = ~new_n1961_ | ~new_n1984_;
  assign new_n3631_ = ~new_n16433_ | ~new_n2934_;
  assign new_n3632_ = ~new_n14705_ | ~new_n2927_;
  assign new_n3633_ = ~new_n17963_ | ~new_n2921_;
  assign new_n3634_ = ~new_n16904_ | ~new_n2932_;
  assign new_n3635_ = ~new_n15370_ | ~new_n2931_;
  assign new_n3636_ = ~new_n17465_ | ~new_n2938_;
  assign new_n3637_ = ~new_n13992_ | ~new_n2919_;
  assign new_n3638_ = ~new_n2339_;
  assign new_n3639_ = ~new_n1952_ | ~new_n1981_;
  assign new_n3640_ = ~new_n18461_ | ~new_n1951_;
  assign new_n3641_ = ~new_n13804_ | ~new_n2963_;
  assign new_n3642_ = ~new_n2945_ | ~new_n3112_;
  assign new_n3643_ = ~new_n2642_ | ~new_n3638_;
  assign new_n3644_ = ~new_n13033_ | ~new_n1944_;
  assign new_n3645_ = ~pi190 | ~new_n1945_;
  assign new_n3646_ = ~pi158 | ~new_n1946_;
  assign new_n3647_ = ~pi126 | ~new_n1947_;
  assign new_n3648_ = ~new_n1982_;
  assign new_n3649_ = ~new_n1961_ | ~new_n1980_;
  assign new_n3650_ = ~new_n16511_ | ~new_n2934_;
  assign new_n3651_ = ~new_n14783_ | ~new_n2927_;
  assign new_n3652_ = ~new_n17962_ | ~new_n2921_;
  assign new_n3653_ = ~new_n16982_ | ~new_n2932_;
  assign new_n3654_ = ~new_n15448_ | ~new_n2931_;
  assign new_n3655_ = ~new_n17464_ | ~new_n2938_;
  assign new_n3656_ = ~new_n13991_ | ~new_n2919_;
  assign new_n3657_ = ~new_n2341_;
  assign new_n3658_ = ~new_n1952_ | ~new_n1982_;
  assign new_n3659_ = ~new_n18460_ | ~new_n1951_;
  assign new_n3660_ = ~new_n13749_ | ~new_n2963_;
  assign new_n3661_ = ~new_n2944_ | ~new_n3112_;
  assign new_n3662_ = ~new_n2646_ | ~new_n3657_;
  assign new_n3663_ = ~pi191 | ~new_n1945_;
  assign new_n3664_ = ~pi159 | ~new_n1946_;
  assign new_n3665_ = ~pi127 | ~new_n1947_;
  assign new_n3666_ = ~new_n1986_;
  assign new_n3667_ = ~new_n4738_ | ~new_n2286_;
  assign new_n3668_ = ~new_n2881_ | ~new_n3667_;
  assign new_n3669_ = ~new_n2647_ | ~new_n1986_;
  assign new_n3670_ = ~new_n1961_ | ~new_n1981_;
  assign new_n3671_ = ~new_n16434_ | ~new_n2934_;
  assign new_n3672_ = ~new_n14706_ | ~new_n2927_;
  assign new_n3673_ = ~new_n17961_ | ~new_n2921_;
  assign new_n3674_ = ~new_n16905_ | ~new_n2932_;
  assign new_n3675_ = ~new_n15371_ | ~new_n2931_;
  assign new_n3676_ = ~new_n17463_ | ~new_n2938_;
  assign new_n3677_ = ~new_n13990_ | ~new_n2919_;
  assign new_n3678_ = ~new_n2343_;
  assign new_n3679_ = ~new_n18459_ | ~new_n1951_;
  assign new_n3680_ = ~new_n13802_ | ~new_n2963_;
  assign new_n3681_ = ~new_n2955_ | ~new_n3112_;
  assign new_n3682_ = ~new_n2651_ | ~new_n3678_;
  assign new_n3683_ = ~pi192 | ~new_n1945_;
  assign new_n3684_ = ~pi160 | ~new_n1946_;
  assign new_n3685_ = ~pi128 | ~new_n1947_;
  assign new_n3686_ = ~new_n1983_;
  assign new_n3687_ = ~new_n13751_ | ~new_n2963_;
  assign new_n3688_ = ~new_n2954_ | ~new_n3112_;
  assign new_n3689_ = ~new_n3687_ | ~new_n3688_ | ~new_n2914_;
  assign new_n3690_ = ~new_n13800_ | ~new_n2963_;
  assign new_n3691_ = ~new_n2953_ | ~new_n3112_;
  assign new_n3692_ = ~new_n3690_ | ~new_n3691_ | ~new_n2914_;
  assign new_n3693_ = ~new_n2654_ | ~new_n1943_;
  assign new_n3694_ = ~new_n2348_ | ~new_n3693_;
  assign new_n3695_ = ~new_n2922_ | ~new_n4729_;
  assign new_n3696_ = ~new_n2353_;
  assign new_n3697_ = ~new_n1963_ | ~new_n2005_;
  assign new_n3698_ = ~new_n1960_ | ~pi255;
  assign new_n3699_ = ~new_n1959_ | ~new_n18453_;
  assign new_n3700_ = ~new_n1958_ | ~new_n2383_;
  assign new_n3701_ = ~new_n1957_ | ~new_n2383_;
  assign new_n3702_ = ~new_n1963_ | ~new_n1995_;
  assign new_n3703_ = ~new_n1960_ | ~pi265;
  assign new_n3704_ = ~new_n1959_ | ~new_n18452_;
  assign new_n3705_ = ~new_n1958_ | ~new_n2388_;
  assign new_n3706_ = ~new_n1957_ | ~new_n13788_;
  assign new_n3707_ = ~new_n1963_ | ~new_n1991_;
  assign new_n3708_ = ~new_n1960_ | ~pi250;
  assign new_n3709_ = ~new_n1959_ | ~new_n18374_;
  assign new_n3710_ = ~new_n1958_ | ~new_n2391_;
  assign new_n3711_ = ~new_n1957_ | ~new_n13750_;
  assign new_n3712_ = ~new_n1963_ | ~new_n1987_;
  assign new_n3713_ = ~new_n1960_ | ~new_n13032_;
  assign new_n3714_ = ~new_n1959_ | ~new_n18458_;
  assign new_n3715_ = ~new_n1958_ | ~new_n2394_;
  assign new_n3716_ = ~new_n1957_ | ~new_n13752_;
  assign new_n3717_ = ~new_n1963_ | ~new_n1994_;
  assign new_n3718_ = ~new_n1960_ | ~new_n13087_;
  assign new_n3719_ = ~new_n1959_ | ~new_n18457_;
  assign new_n3720_ = ~new_n1958_ | ~new_n2397_;
  assign new_n3721_ = ~new_n1957_ | ~new_n13753_;
  assign new_n3722_ = ~new_n1963_ | ~new_n1998_;
  assign new_n3723_ = ~new_n1960_ | ~new_n13086_;
  assign new_n3724_ = ~new_n1959_ | ~new_n18375_;
  assign new_n3725_ = ~new_n1958_ | ~new_n2400_;
  assign new_n3726_ = ~new_n1957_ | ~new_n13797_;
  assign new_n3727_ = ~new_n1963_ | ~new_n1997_;
  assign new_n3728_ = ~new_n1960_ | ~new_n13085_;
  assign new_n3729_ = ~new_n1959_ | ~new_n18456_;
  assign new_n3730_ = ~new_n1958_ | ~new_n2403_;
  assign new_n3731_ = ~new_n1957_ | ~new_n13754_;
  assign new_n3732_ = ~new_n1963_ | ~new_n2011_;
  assign new_n3733_ = ~new_n1960_ | ~new_n13084_;
  assign new_n3734_ = ~new_n1959_ | ~new_n18376_;
  assign new_n3735_ = ~new_n1958_ | ~new_n2406_;
  assign new_n3736_ = ~new_n1957_ | ~new_n13755_;
  assign new_n3737_ = ~new_n1963_ | ~new_n2010_;
  assign new_n3738_ = ~new_n1960_ | ~new_n13083_;
  assign new_n3739_ = ~new_n1959_ | ~new_n18455_;
  assign new_n3740_ = ~new_n1958_ | ~new_n2409_;
  assign new_n3741_ = ~new_n1957_ | ~new_n13756_;
  assign new_n3742_ = ~new_n1963_ | ~new_n1989_;
  assign new_n3743_ = ~new_n1960_ | ~new_n13082_;
  assign new_n3744_ = ~new_n1959_ | ~new_n18454_;
  assign new_n3745_ = ~new_n1958_ | ~new_n2412_;
  assign new_n3746_ = ~new_n1957_ | ~new_n13795_;
  assign new_n3747_ = ~new_n1963_ | ~new_n1990_;
  assign new_n3748_ = ~new_n1960_ | ~new_n13106_;
  assign new_n3749_ = ~new_n1959_ | ~new_n18368_;
  assign new_n3750_ = ~new_n1958_ | ~new_n2415_;
  assign new_n3751_ = ~new_n1957_ | ~new_n13738_;
  assign new_n3752_ = ~new_n1963_ | ~new_n1999_;
  assign new_n3753_ = ~new_n1960_ | ~new_n13105_;
  assign new_n3754_ = ~new_n1959_ | ~new_n18472_;
  assign new_n3755_ = ~new_n1958_ | ~new_n2418_;
  assign new_n3756_ = ~new_n1957_ | ~new_n13739_;
  assign new_n3757_ = ~new_n1963_ | ~new_n2007_;
  assign new_n3758_ = ~new_n1960_ | ~new_n13104_;
  assign new_n3759_ = ~new_n1959_ | ~new_n18471_;
  assign new_n3760_ = ~new_n1958_ | ~new_n2421_;
  assign new_n3761_ = ~new_n1957_ | ~new_n13740_;
  assign new_n3762_ = ~new_n1963_ | ~new_n2006_;
  assign new_n3763_ = ~new_n1960_ | ~new_n13103_;
  assign new_n3764_ = ~new_n1959_ | ~new_n18369_;
  assign new_n3765_ = ~new_n1958_ | ~new_n2424_;
  assign new_n3766_ = ~new_n1957_ | ~new_n13818_;
  assign new_n3767_ = ~new_n1963_ | ~new_n2001_;
  assign new_n3768_ = ~new_n1960_ | ~new_n13102_;
  assign new_n3769_ = ~new_n1959_ | ~new_n18470_;
  assign new_n3770_ = ~new_n1958_ | ~new_n2427_;
  assign new_n3771_ = ~new_n1957_ | ~new_n13741_;
  assign new_n3772_ = ~new_n1963_ | ~new_n2000_;
  assign new_n3773_ = ~new_n1960_ | ~new_n13101_;
  assign new_n3774_ = ~new_n1959_ | ~new_n18469_;
  assign new_n3775_ = ~new_n1958_ | ~new_n2430_;
  assign new_n3776_ = ~new_n1957_ | ~new_n13742_;
  assign new_n3777_ = ~new_n1963_ | ~new_n1996_;
  assign new_n3778_ = ~new_n1960_ | ~new_n13100_;
  assign new_n3779_ = ~new_n1959_ | ~new_n18468_;
  assign new_n3780_ = ~new_n1958_ | ~new_n2433_;
  assign new_n3781_ = ~new_n1957_ | ~new_n13743_;
  assign new_n3782_ = ~new_n1963_ | ~new_n2009_;
  assign new_n3783_ = ~new_n1960_ | ~new_n13099_;
  assign new_n3784_ = ~new_n1959_ | ~new_n18370_;
  assign new_n3785_ = ~new_n1958_ | ~new_n2436_;
  assign new_n3786_ = ~new_n1957_ | ~new_n13816_;
  assign new_n3787_ = ~new_n1963_ | ~new_n2008_;
  assign new_n3788_ = ~new_n1960_ | ~new_n13098_;
  assign new_n3789_ = ~new_n1959_ | ~new_n18467_;
  assign new_n3790_ = ~new_n1958_ | ~new_n2439_;
  assign new_n3791_ = ~new_n1957_ | ~new_n13744_;
  assign new_n3792_ = ~new_n1963_ | ~new_n2003_;
  assign new_n3793_ = ~new_n1960_ | ~new_n13097_;
  assign new_n3794_ = ~new_n1959_ | ~new_n18466_;
  assign new_n3795_ = ~new_n1958_ | ~new_n2441_;
  assign new_n3796_ = ~new_n1957_ | ~new_n13814_;
  assign new_n3797_ = ~new_n1963_ | ~new_n2002_;
  assign new_n3798_ = ~new_n1960_ | ~new_n13096_;
  assign new_n3799_ = ~new_n1959_ | ~new_n18371_;
  assign new_n3800_ = ~new_n1958_ | ~new_n2952_;
  assign new_n3801_ = ~new_n1957_ | ~new_n13745_;
  assign new_n3802_ = ~new_n1963_ | ~new_n1988_;
  assign new_n3803_ = ~new_n1960_ | ~new_n13095_;
  assign new_n3804_ = ~new_n1959_ | ~new_n18372_;
  assign new_n3805_ = ~new_n1958_ | ~new_n2951_;
  assign new_n3806_ = ~new_n1957_ | ~new_n13810_;
  assign new_n3807_ = ~new_n1963_ | ~new_n1993_;
  assign new_n3808_ = ~new_n1960_ | ~new_n13094_;
  assign new_n3809_ = ~new_n1959_ | ~new_n18465_;
  assign new_n3810_ = ~new_n1958_ | ~new_n2950_;
  assign new_n3811_ = ~new_n1957_ | ~new_n13746_;
  assign new_n3812_ = ~new_n1963_ | ~new_n1992_;
  assign new_n3813_ = ~new_n1960_ | ~new_n13093_;
  assign new_n3814_ = ~new_n1959_ | ~new_n18464_;
  assign new_n3815_ = ~new_n1958_ | ~new_n2949_;
  assign new_n3816_ = ~new_n1957_ | ~new_n13808_;
  assign new_n3817_ = ~new_n1963_ | ~new_n1985_;
  assign new_n3818_ = ~new_n1960_ | ~new_n13092_;
  assign new_n3819_ = ~new_n1959_ | ~new_n18463_;
  assign new_n3820_ = ~new_n1958_ | ~new_n2948_;
  assign new_n3821_ = ~new_n1957_ | ~new_n13747_;
  assign new_n3822_ = ~new_n1963_ | ~new_n1984_;
  assign new_n3823_ = ~new_n1960_ | ~new_n13091_;
  assign new_n3824_ = ~new_n1959_ | ~new_n18462_;
  assign new_n3825_ = ~new_n1958_ | ~new_n2947_;
  assign new_n3826_ = ~new_n1957_ | ~new_n13806_;
  assign new_n3827_ = ~new_n1963_ | ~new_n1980_;
  assign new_n3828_ = ~new_n1960_ | ~new_n13090_;
  assign new_n3829_ = ~new_n1959_ | ~new_n18373_;
  assign new_n3830_ = ~new_n1958_ | ~new_n2946_;
  assign new_n3831_ = ~new_n1957_ | ~new_n13748_;
  assign new_n3832_ = ~new_n1963_ | ~new_n1981_;
  assign new_n3833_ = ~new_n1960_ | ~new_n13089_;
  assign new_n3834_ = ~new_n1959_ | ~new_n18461_;
  assign new_n3835_ = ~new_n1958_ | ~new_n2945_;
  assign new_n3836_ = ~new_n1957_ | ~new_n13804_;
  assign new_n3837_ = ~new_n1963_ | ~new_n1982_;
  assign new_n3838_ = ~new_n1960_ | ~new_n13088_;
  assign new_n3839_ = ~new_n1959_ | ~new_n18460_;
  assign new_n3840_ = ~new_n1958_ | ~new_n2944_;
  assign new_n3841_ = ~new_n1957_ | ~new_n13749_;
  assign new_n3842_ = ~new_n1960_ | ~new_n13033_;
  assign new_n3843_ = ~new_n1959_ | ~new_n18459_;
  assign new_n3844_ = ~new_n1958_ | ~new_n2955_;
  assign new_n3845_ = ~new_n1957_ | ~new_n13802_;
  assign new_n3846_ = ~new_n1958_ | ~new_n2954_;
  assign new_n3847_ = ~new_n1957_ | ~new_n13751_;
  assign new_n3848_ = ~new_n1958_ | ~new_n2953_;
  assign new_n3849_ = ~new_n1957_ | ~new_n13800_;
  assign new_n3850_ = ~new_n2714_ | ~new_n2348_ | ~new_n3696_ | ~new_n2716_ | ~new_n2713_;
  assign new_n3851_ = ~new_n13191_ | ~new_n1969_;
  assign new_n3852_ = ~new_n1967_ | ~new_n2379_;
  assign new_n3853_ = ~new_n14399_ | ~new_n1965_;
  assign new_n3854_ = ~new_n3853_ | ~new_n3852_ | ~new_n3851_;
  assign new_n3855_ = ~new_n2352_ | ~new_n2299_;
  assign new_n3856_ = ~new_n4713_ | ~new_n3855_;
  assign new_n3857_ = ~new_n3856_ | ~new_n2881_;
  assign new_n3858_ = ~po265;
  assign new_n3859_ = ~new_n2355_;
  assign new_n3860_ = ~new_n1971_ | ~new_n3854_;
  assign new_n3861_ = ~new_n1970_ | ~new_n13191_;
  assign new_n3862_ = ~pi268 | ~po264;
  assign new_n3863_ = ~new_n1968_ | ~new_n2379_;
  assign new_n3864_ = ~new_n1966_ | ~new_n14399_;
  assign new_n3865_ = ~pi193 | ~new_n3859_;
  assign new_n3866_ = ~new_n13253_ | ~new_n1969_;
  assign new_n3867_ = ~new_n1967_ | ~new_n2438_;
  assign new_n3868_ = ~new_n14461_ | ~new_n1965_;
  assign new_n3869_ = ~new_n3868_ | ~new_n3867_ | ~new_n3866_;
  assign new_n3870_ = ~new_n1971_ | ~new_n3869_;
  assign new_n3871_ = ~new_n13253_ | ~new_n1970_;
  assign new_n3872_ = ~pi249 | ~po264;
  assign new_n3873_ = ~new_n1968_ | ~new_n2438_;
  assign new_n3874_ = ~new_n14461_ | ~new_n1966_;
  assign new_n3875_ = ~pi194 | ~new_n3859_;
  assign new_n3876_ = ~new_n13190_ | ~new_n1969_;
  assign new_n3877_ = ~new_n1967_ | ~new_n2435_;
  assign new_n3878_ = ~new_n14398_ | ~new_n1965_;
  assign new_n3879_ = ~new_n3878_ | ~new_n3877_ | ~new_n3876_;
  assign new_n3880_ = ~new_n1971_ | ~new_n3879_;
  assign new_n3881_ = ~new_n13190_ | ~new_n1970_;
  assign new_n3882_ = ~pi259 | ~po264;
  assign new_n3883_ = ~new_n1968_ | ~new_n2435_;
  assign new_n3884_ = ~new_n14398_ | ~new_n1966_;
  assign new_n3885_ = ~pi195 | ~new_n3859_;
  assign new_n3886_ = ~new_n13254_ | ~new_n1969_;
  assign new_n3887_ = ~new_n1967_ | ~new_n2432_;
  assign new_n3888_ = ~new_n14462_ | ~new_n1965_;
  assign new_n3889_ = ~new_n3888_ | ~new_n3887_ | ~new_n3886_;
  assign new_n3890_ = ~new_n1971_ | ~new_n3889_;
  assign new_n3891_ = ~new_n13254_ | ~new_n1970_;
  assign new_n3892_ = ~pi261 | ~po264;
  assign new_n3893_ = ~new_n1968_ | ~new_n2432_;
  assign new_n3894_ = ~new_n14462_ | ~new_n1966_;
  assign new_n3895_ = ~pi196 | ~new_n3859_;
  assign new_n3896_ = ~new_n13255_ | ~new_n1969_;
  assign new_n3897_ = ~new_n1967_ | ~new_n2429_;
  assign new_n3898_ = ~new_n14463_ | ~new_n1965_;
  assign new_n3899_ = ~new_n3898_ | ~new_n3897_ | ~new_n3896_;
  assign new_n3900_ = ~new_n1971_ | ~new_n3899_;
  assign new_n3901_ = ~new_n13255_ | ~new_n1970_;
  assign new_n3902_ = ~pi246 | ~po264;
  assign new_n3903_ = ~new_n1968_ | ~new_n2429_;
  assign new_n3904_ = ~new_n14463_ | ~new_n1966_;
  assign new_n3905_ = ~pi197 | ~new_n3859_;
  assign new_n3906_ = ~new_n13256_ | ~new_n1969_;
  assign new_n3907_ = ~new_n1967_ | ~new_n2426_;
  assign new_n3908_ = ~new_n14464_ | ~new_n1965_;
  assign new_n3909_ = ~new_n3908_ | ~new_n3907_ | ~new_n3906_;
  assign new_n3910_ = ~new_n1971_ | ~new_n3909_;
  assign new_n3911_ = ~new_n13256_ | ~new_n1970_;
  assign new_n3912_ = ~pi272 | ~po264;
  assign new_n3913_ = ~new_n1968_ | ~new_n2426_;
  assign new_n3914_ = ~new_n14464_ | ~new_n1966_;
  assign new_n3915_ = ~pi198 | ~new_n3859_;
  assign new_n3916_ = ~new_n13189_ | ~new_n1969_;
  assign new_n3917_ = ~new_n1967_ | ~new_n2423_;
  assign new_n3918_ = ~new_n14397_ | ~new_n1965_;
  assign new_n3919_ = ~new_n3918_ | ~new_n3917_ | ~new_n3916_;
  assign new_n3920_ = ~new_n1971_ | ~new_n3919_;
  assign new_n3921_ = ~new_n13189_ | ~new_n1970_;
  assign new_n3922_ = ~pi253 | ~po264;
  assign new_n3923_ = ~new_n1968_ | ~new_n2423_;
  assign new_n3924_ = ~new_n14397_ | ~new_n1966_;
  assign new_n3925_ = ~pi199 | ~new_n3859_;
  assign new_n3926_ = ~new_n13257_ | ~new_n1969_;
  assign new_n3927_ = ~new_n1967_ | ~new_n2420_;
  assign new_n3928_ = ~new_n14465_ | ~new_n1965_;
  assign new_n3929_ = ~new_n3928_ | ~new_n3927_ | ~new_n3926_;
  assign new_n3930_ = ~new_n1971_ | ~new_n3929_;
  assign new_n3931_ = ~new_n13257_ | ~new_n1970_;
  assign new_n3932_ = ~pi263 | ~po264;
  assign new_n3933_ = ~new_n1968_ | ~new_n2420_;
  assign new_n3934_ = ~new_n14465_ | ~new_n1966_;
  assign new_n3935_ = ~pi200 | ~new_n3859_;
  assign new_n3936_ = ~new_n13258_ | ~new_n1969_;
  assign new_n3937_ = ~new_n1967_ | ~new_n2417_;
  assign new_n3938_ = ~new_n14466_ | ~new_n1965_;
  assign new_n3939_ = ~new_n3938_ | ~new_n3937_ | ~new_n3936_;
  assign new_n3940_ = ~new_n1971_ | ~new_n3939_;
  assign new_n3941_ = ~new_n13258_ | ~new_n1970_;
  assign new_n3942_ = ~pi251 | ~po264;
  assign new_n3943_ = ~new_n1968_ | ~new_n2417_;
  assign new_n3944_ = ~new_n14466_ | ~new_n1966_;
  assign new_n3945_ = ~pi201 | ~new_n3859_;
  assign new_n3946_ = ~new_n13188_ | ~new_n1969_;
  assign new_n3947_ = ~new_n1967_ | ~new_n2414_;
  assign new_n3948_ = ~new_n14396_ | ~new_n1965_;
  assign new_n3949_ = ~new_n3948_ | ~new_n3947_ | ~new_n3946_;
  assign new_n3950_ = ~new_n1971_ | ~new_n3949_;
  assign new_n3951_ = ~new_n13188_ | ~new_n1970_;
  assign new_n3952_ = ~pi270 | ~po264;
  assign new_n3953_ = ~new_n1968_ | ~new_n2414_;
  assign new_n3954_ = ~new_n14396_ | ~new_n1966_;
  assign new_n3955_ = ~pi202 | ~new_n3859_;
  assign new_n3956_ = ~new_n13248_ | ~new_n1969_;
  assign new_n3957_ = ~new_n1967_ | ~new_n2411_;
  assign new_n3958_ = ~new_n14456_ | ~new_n1965_;
  assign new_n3959_ = ~new_n3958_ | ~new_n3957_ | ~new_n3956_;
  assign new_n3960_ = ~new_n1971_ | ~new_n3959_;
  assign new_n3961_ = ~new_n13248_ | ~new_n1970_;
  assign new_n3962_ = ~pi256 | ~po264;
  assign new_n3963_ = ~new_n1968_ | ~new_n2411_;
  assign new_n3964_ = ~new_n14456_ | ~new_n1966_;
  assign new_n3965_ = ~pi203 | ~new_n3859_;
  assign new_n3966_ = ~new_n13249_ | ~new_n1969_;
  assign new_n3967_ = ~new_n1967_ | ~new_n2408_;
  assign new_n3968_ = ~new_n14457_ | ~new_n1965_;
  assign new_n3969_ = ~new_n3968_ | ~new_n3967_ | ~new_n3966_;
  assign new_n3970_ = ~new_n1971_ | ~new_n3969_;
  assign new_n3971_ = ~new_n13249_ | ~new_n1970_;
  assign new_n3972_ = ~pi266 | ~po264;
  assign new_n3973_ = ~new_n1968_ | ~new_n2408_;
  assign new_n3974_ = ~new_n14457_ | ~new_n1966_;
  assign new_n3975_ = ~pi204 | ~new_n3859_;
  assign new_n3976_ = ~new_n13194_ | ~new_n1969_;
  assign new_n3977_ = ~new_n1967_ | ~new_n2405_;
  assign new_n3978_ = ~new_n14402_ | ~new_n1965_;
  assign new_n3979_ = ~new_n3978_ | ~new_n3977_ | ~new_n3976_;
  assign new_n3980_ = ~new_n1971_ | ~new_n3979_;
  assign new_n3981_ = ~new_n13194_ | ~new_n1970_;
  assign new_n3982_ = ~pi274 | ~po264;
  assign new_n3983_ = ~new_n1968_ | ~new_n2405_;
  assign new_n3984_ = ~new_n14402_ | ~new_n1966_;
  assign new_n3985_ = ~pi205 | ~new_n3859_;
  assign new_n3986_ = ~new_n13250_ | ~new_n1969_;
  assign new_n3987_ = ~new_n1967_ | ~new_n2402_;
  assign new_n3988_ = ~new_n14458_ | ~new_n1965_;
  assign new_n3989_ = ~new_n3988_ | ~new_n3987_ | ~new_n3986_;
  assign new_n3990_ = ~new_n1971_ | ~new_n3989_;
  assign new_n3991_ = ~new_n13250_ | ~new_n1970_;
  assign new_n3992_ = ~pi248 | ~po264;
  assign new_n3993_ = ~new_n1968_ | ~new_n2402_;
  assign new_n3994_ = ~new_n14458_ | ~new_n1966_;
  assign new_n3995_ = ~pi206 | ~new_n3859_;
  assign new_n3996_ = ~new_n13193_ | ~new_n1969_;
  assign new_n3997_ = ~new_n1967_ | ~new_n2399_;
  assign new_n3998_ = ~new_n14401_ | ~new_n1965_;
  assign new_n3999_ = ~new_n3998_ | ~new_n3997_ | ~new_n3996_;
  assign new_n4000_ = ~new_n1971_ | ~new_n3999_;
  assign new_n4001_ = ~new_n13193_ | ~new_n1970_;
  assign new_n4002_ = ~pi260 | ~po264;
  assign new_n4003_ = ~new_n1968_ | ~new_n2399_;
  assign new_n4004_ = ~new_n14401_ | ~new_n1966_;
  assign new_n4005_ = ~pi207 | ~new_n3859_;
  assign new_n4006_ = ~new_n13251_ | ~new_n1969_;
  assign new_n4007_ = ~new_n1967_ | ~new_n2396_;
  assign new_n4008_ = ~new_n14459_ | ~new_n1965_;
  assign new_n4009_ = ~new_n4008_ | ~new_n4007_ | ~new_n4006_;
  assign new_n4010_ = ~new_n1971_ | ~new_n4009_;
  assign new_n4011_ = ~new_n13251_ | ~new_n1970_;
  assign new_n4012_ = ~pi257 | ~po264;
  assign new_n4013_ = ~new_n1968_ | ~new_n2396_;
  assign new_n4014_ = ~new_n14459_ | ~new_n1966_;
  assign new_n4015_ = ~pi208 | ~new_n3859_;
  assign new_n4016_ = ~new_n13252_ | ~new_n1969_;
  assign new_n4017_ = ~new_n1967_ | ~new_n2393_;
  assign new_n4018_ = ~new_n14460_ | ~new_n1965_;
  assign new_n4019_ = ~new_n4018_ | ~new_n4017_ | ~new_n4016_;
  assign new_n4020_ = ~new_n1971_ | ~new_n4019_;
  assign new_n4021_ = ~new_n13252_ | ~new_n1970_;
  assign new_n4022_ = ~pi269 | ~po264;
  assign new_n4023_ = ~new_n1968_ | ~new_n2393_;
  assign new_n4024_ = ~new_n14460_ | ~new_n1966_;
  assign new_n4025_ = ~pi209 | ~new_n3859_;
  assign new_n4026_ = ~new_n13192_ | ~new_n1969_;
  assign new_n4027_ = ~new_n1967_ | ~new_n2390_;
  assign new_n4028_ = ~new_n14400_ | ~new_n1965_;
  assign new_n4029_ = ~new_n4028_ | ~new_n4027_ | ~new_n4026_;
  assign new_n4030_ = ~new_n1971_ | ~new_n4029_;
  assign new_n4031_ = ~new_n13192_ | ~new_n1970_;
  assign new_n4032_ = ~pi250 | ~po264;
  assign new_n4033_ = ~new_n1968_ | ~new_n2390_;
  assign new_n4034_ = ~new_n14400_ | ~new_n1966_;
  assign new_n4035_ = ~pi210 | ~new_n3859_;
  assign new_n4036_ = ~new_n13246_ | ~new_n1969_;
  assign new_n4037_ = ~new_n1967_ | ~new_n2387_;
  assign new_n4038_ = ~new_n14454_ | ~new_n1965_;
  assign new_n4039_ = ~new_n4038_ | ~new_n4037_ | ~new_n4036_;
  assign new_n4040_ = ~new_n1971_ | ~new_n4039_;
  assign new_n4041_ = ~new_n13246_ | ~new_n1970_;
  assign new_n4042_ = ~pi265 | ~po264;
  assign new_n4043_ = ~new_n1968_ | ~new_n2387_;
  assign new_n4044_ = ~new_n14454_ | ~new_n1966_;
  assign new_n4045_ = ~pi211 | ~new_n3859_;
  assign new_n4046_ = ~new_n13247_ | ~new_n1969_;
  assign new_n4047_ = ~new_n1967_ | ~new_n2381_;
  assign new_n4048_ = ~new_n14455_ | ~new_n1965_;
  assign new_n4049_ = ~new_n4048_ | ~new_n4047_ | ~new_n4046_;
  assign new_n4050_ = ~new_n1971_ | ~new_n4049_;
  assign new_n4051_ = ~new_n13247_ | ~new_n1970_;
  assign new_n4052_ = ~pi255 | ~po264;
  assign new_n4053_ = ~new_n1968_ | ~new_n2381_;
  assign new_n4054_ = ~new_n14455_ | ~new_n1966_;
  assign new_n4055_ = ~pi212 | ~new_n3859_;
  assign new_n4056_ = ~new_n2918_;
  assign new_n4057_ = ~new_n2917_ | ~new_n5204_ | ~new_n5203_;
  assign new_n4058_ = ~new_n2297_ | ~new_n2300_;
  assign new_n4059_ = ~new_n4729_ | ~new_n2378_;
  assign new_n4060_ = ~new_n2349_ | ~new_n4059_;
  assign new_n4061_ = ~new_n4699_ | ~new_n5206_ | ~new_n5205_;
  assign new_n4062_ = ~new_n2772_ | ~new_n5208_ | ~new_n5207_;
  assign new_n4063_ = ~new_n2359_ | ~new_n1949_ | ~new_n2956_;
  assign new_n4064_ = ~new_n2970_ | ~new_n4061_;
  assign new_n4065_ = ~pi245 | ~new_n4062_;
  assign new_n4066_ = ~new_n1964_ | ~new_n2006_;
  assign new_n4067_ = ~new_n1962_ | ~new_n2000_;
  assign new_n4068_ = ~new_n13101_ | ~new_n2361_;
  assign new_n4069_ = ~new_n4067_ | ~new_n4068_ | ~new_n4066_;
  assign new_n4070_ = ~new_n2079_;
  assign new_n4071_ = ~new_n2350_ | ~new_n2926_;
  assign new_n4072_ = ~new_n5209_ | ~new_n2775_ | ~new_n2776_ | ~new_n5210_;
  assign new_n4073_ = ~new_n4072_ | ~new_n2361_;
  assign new_n4074_ = ~new_n2939_ | ~new_n4073_;
  assign new_n4075_ = ~new_n1949_ | ~new_n4074_;
  assign new_n4076_ = ~new_n2430_ | ~new_n4697_;
  assign new_n4077_ = ~new_n13101_ | ~new_n4696_;
  assign new_n4078_ = ~new_n15932_ | ~new_n1953_;
  assign new_n4079_ = ~new_n2964_ | ~new_n4069_;
  assign new_n4080_ = ~pi246 | ~po264;
  assign new_n4081_ = ~new_n1964_ | ~new_n1985_;
  assign new_n4082_ = ~new_n1962_ | ~new_n1980_;
  assign new_n4083_ = ~new_n13090_ | ~new_n2361_;
  assign new_n4084_ = ~new_n4082_ | ~new_n4083_ | ~new_n4081_;
  assign new_n4085_ = ~new_n2942_ | ~new_n2353_;
  assign new_n4086_ = ~new_n2348_ | ~new_n4085_;
  assign new_n4087_ = ~new_n1972_ | ~new_n2946_;
  assign new_n4088_ = ~new_n13090_ | ~new_n4696_;
  assign new_n4089_ = ~new_n15839_ | ~new_n1953_;
  assign new_n4090_ = ~new_n2964_ | ~new_n4084_;
  assign new_n4091_ = ~pi247 | ~po264;
  assign new_n4092_ = ~new_n1964_ | ~new_n1994_;
  assign new_n4093_ = ~new_n1962_ | ~new_n1997_;
  assign new_n4094_ = ~new_n13085_ | ~new_n2361_;
  assign new_n4095_ = ~new_n4094_ | ~new_n4093_ | ~new_n4092_;
  assign new_n4096_ = ~new_n2403_ | ~new_n4697_;
  assign new_n4097_ = ~new_n13085_ | ~new_n4696_;
  assign new_n4098_ = ~new_n15917_ | ~new_n1953_;
  assign new_n4099_ = ~new_n2964_ | ~new_n4095_;
  assign new_n4100_ = ~pi248 | ~po264;
  assign new_n4101_ = ~new_n1964_ | ~new_n1996_;
  assign new_n4102_ = ~new_n1962_ | ~new_n2008_;
  assign new_n4103_ = ~new_n13098_ | ~new_n2361_;
  assign new_n4104_ = ~new_n4102_ | ~new_n4103_ | ~new_n4101_;
  assign new_n4105_ = ~new_n2439_ | ~new_n4697_;
  assign new_n4106_ = ~new_n13098_ | ~new_n4696_;
  assign new_n4107_ = ~new_n15930_ | ~new_n1953_;
  assign new_n4108_ = ~new_n2964_ | ~new_n4104_;
  assign new_n4109_ = ~pi249 | ~po264;
  assign new_n4110_ = ~new_n1964_ | ~new_n2005_;
  assign new_n4111_ = ~new_n1962_ | ~new_n1991_;
  assign new_n4112_ = ~pi250 | ~new_n2361_;
  assign new_n4113_ = ~new_n4112_ | ~new_n4111_ | ~new_n4110_;
  assign new_n4114_ = ~new_n2391_ | ~new_n4697_;
  assign new_n4115_ = ~pi250 | ~new_n4696_;
  assign new_n4116_ = ~new_n15920_ | ~new_n1953_;
  assign new_n4117_ = ~new_n2964_ | ~new_n4113_;
  assign new_n4118_ = ~pi250 | ~po264;
  assign new_n4119_ = ~new_n1964_ | ~new_n1989_;
  assign new_n4120_ = ~new_n1962_ | ~new_n1999_;
  assign new_n4121_ = ~new_n13105_ | ~new_n2361_;
  assign new_n4122_ = ~new_n4121_ | ~new_n4120_ | ~new_n4119_;
  assign new_n4123_ = ~new_n2418_ | ~new_n4697_;
  assign new_n4124_ = ~new_n13105_ | ~new_n4696_;
  assign new_n4125_ = ~new_n15935_ | ~new_n1953_;
  assign new_n4126_ = ~new_n2964_ | ~new_n4122_;
  assign new_n4127_ = ~pi251 | ~po264;
  assign new_n4128_ = ~new_n1964_ | ~new_n2002_;
  assign new_n4129_ = ~new_n1962_ | ~new_n1993_;
  assign new_n4130_ = ~new_n13094_ | ~new_n2361_;
  assign new_n4131_ = ~new_n4129_ | ~new_n4130_ | ~new_n4128_;
  assign new_n4132_ = ~new_n1972_ | ~new_n2950_;
  assign new_n4133_ = ~new_n13094_ | ~new_n4696_;
  assign new_n4134_ = ~new_n15926_ | ~new_n1953_;
  assign new_n4135_ = ~new_n2964_ | ~new_n4131_;
  assign new_n4136_ = ~pi252 | ~po264;
  assign new_n4137_ = ~new_n1964_ | ~new_n1999_;
  assign new_n4138_ = ~new_n1962_ | ~new_n2006_;
  assign new_n4139_ = ~new_n13103_ | ~new_n2361_;
  assign new_n4140_ = ~new_n4138_ | ~new_n4139_ | ~new_n4137_;
  assign new_n4141_ = ~new_n2424_ | ~new_n4697_;
  assign new_n4142_ = ~new_n13103_ | ~new_n4696_;
  assign new_n4143_ = ~new_n15836_ | ~new_n1953_;
  assign new_n4144_ = ~new_n2964_ | ~new_n4140_;
  assign new_n4145_ = ~pi253 | ~po264;
  assign new_n4146_ = ~new_n1964_ | ~new_n2008_;
  assign new_n4147_ = ~new_n1962_ | ~new_n2002_;
  assign new_n4148_ = ~new_n13096_ | ~new_n2361_;
  assign new_n4149_ = ~new_n4147_ | ~new_n4148_ | ~new_n4146_;
  assign new_n4150_ = ~new_n1972_ | ~new_n2952_;
  assign new_n4151_ = ~new_n13096_ | ~new_n4696_;
  assign new_n4152_ = ~new_n15927_ | ~new_n1953_;
  assign new_n4153_ = ~new_n2964_ | ~new_n4149_;
  assign new_n4154_ = ~pi254 | ~po264;
  assign new_n4155_ = ~new_n2362_ | ~new_n2360_;
  assign new_n4156_ = ~new_n4155_ | ~new_n2361_;
  assign new_n4157_ = ~new_n1977_ | ~new_n4156_;
  assign new_n4158_ = ~new_n2785_ | ~new_n1962_;
  assign new_n4159_ = ~new_n2383_ | ~new_n4697_;
  assign new_n4160_ = ~pi255 | ~new_n4157_;
  assign new_n4161_ = ~new_n15914_ | ~new_n1953_;
  assign new_n4162_ = ~pi255 | ~po264;
  assign new_n4163_ = ~new_n1964_ | ~new_n2011_;
  assign new_n4164_ = ~new_n1962_ | ~new_n1989_;
  assign new_n4165_ = ~new_n13082_ | ~new_n2361_;
  assign new_n4166_ = ~new_n4165_ | ~new_n4164_ | ~new_n4163_;
  assign new_n4167_ = ~new_n2412_ | ~new_n4697_;
  assign new_n4168_ = ~new_n13082_ | ~new_n4696_;
  assign new_n4169_ = ~new_n15915_ | ~new_n1953_;
  assign new_n4170_ = ~new_n2964_ | ~new_n4166_;
  assign new_n4171_ = ~pi256 | ~po264;
  assign new_n4172_ = ~new_n1964_ | ~new_n1991_;
  assign new_n4173_ = ~new_n1962_ | ~new_n1994_;
  assign new_n4174_ = ~new_n13087_ | ~new_n2361_;
  assign new_n4175_ = ~new_n4174_ | ~new_n4173_ | ~new_n4172_;
  assign new_n4176_ = ~new_n2397_ | ~new_n4697_;
  assign new_n4177_ = ~new_n13087_ | ~new_n4696_;
  assign new_n4178_ = ~new_n15919_ | ~new_n1953_;
  assign new_n4179_ = ~new_n2964_ | ~new_n4175_;
  assign new_n4180_ = ~pi257 | ~po264;
  assign new_n4181_ = ~new_n1964_ | ~new_n1993_;
  assign new_n4182_ = ~new_n1962_ | ~new_n1985_;
  assign new_n4183_ = ~new_n13092_ | ~new_n2361_;
  assign new_n4184_ = ~new_n4182_ | ~new_n4183_ | ~new_n4181_;
  assign new_n4185_ = ~new_n1972_ | ~new_n2948_;
  assign new_n4186_ = ~new_n13092_ | ~new_n4696_;
  assign new_n4187_ = ~new_n15924_ | ~new_n1953_;
  assign new_n4188_ = ~new_n2964_ | ~new_n4184_;
  assign new_n4189_ = ~pi258 | ~po264;
  assign new_n4190_ = ~new_n1964_ | ~new_n2000_;
  assign new_n4191_ = ~new_n1962_ | ~new_n2009_;
  assign new_n4192_ = ~new_n13099_ | ~new_n2361_;
  assign new_n4193_ = ~new_n4191_ | ~new_n4192_ | ~new_n4190_;
  assign new_n4194_ = ~new_n2436_ | ~new_n4697_;
  assign new_n4195_ = ~new_n13099_ | ~new_n4696_;
  assign new_n4196_ = ~new_n15837_ | ~new_n1953_;
  assign new_n4197_ = ~new_n2964_ | ~new_n4193_;
  assign new_n4198_ = ~pi259 | ~po264;
  assign new_n4199_ = ~new_n1964_ | ~new_n1987_;
  assign new_n4200_ = ~new_n1962_ | ~new_n1998_;
  assign new_n4201_ = ~new_n13086_ | ~new_n2361_;
  assign new_n4202_ = ~new_n4201_ | ~new_n4200_ | ~new_n4199_;
  assign new_n4203_ = ~new_n2400_ | ~new_n4697_;
  assign new_n4204_ = ~new_n13086_ | ~new_n4696_;
  assign new_n4205_ = ~new_n15918_ | ~new_n1953_;
  assign new_n4206_ = ~new_n2964_ | ~new_n4202_;
  assign new_n4207_ = ~pi260 | ~po264;
  assign new_n4208_ = ~new_n1964_ | ~new_n2001_;
  assign new_n4209_ = ~new_n1962_ | ~new_n1996_;
  assign new_n4210_ = ~new_n13100_ | ~new_n2361_;
  assign new_n4211_ = ~new_n4209_ | ~new_n4210_ | ~new_n4208_;
  assign new_n4212_ = ~new_n2433_ | ~new_n4697_;
  assign new_n4213_ = ~new_n13100_ | ~new_n4696_;
  assign new_n4214_ = ~new_n15931_ | ~new_n1953_;
  assign new_n4215_ = ~new_n2964_ | ~new_n4211_;
  assign new_n4216_ = ~pi261 | ~po264;
  assign new_n4217_ = ~new_n1964_ | ~new_n1992_;
  assign new_n4218_ = ~new_n1962_ | ~new_n1984_;
  assign new_n4219_ = ~new_n13091_ | ~new_n2361_;
  assign new_n4220_ = ~new_n4218_ | ~new_n4219_ | ~new_n4217_;
  assign new_n4221_ = ~new_n1972_ | ~new_n2947_;
  assign new_n4222_ = ~new_n13091_ | ~new_n4696_;
  assign new_n4223_ = ~new_n15923_ | ~new_n1953_;
  assign new_n4224_ = ~new_n2964_ | ~new_n4220_;
  assign new_n4225_ = ~pi262 | ~po264;
  assign new_n4226_ = ~new_n1964_ | ~new_n1990_;
  assign new_n4227_ = ~new_n1962_ | ~new_n2007_;
  assign new_n4228_ = ~new_n13104_ | ~new_n2361_;
  assign new_n4229_ = ~new_n4227_ | ~new_n4228_ | ~new_n4226_;
  assign new_n4230_ = ~new_n2421_ | ~new_n4697_;
  assign new_n4231_ = ~new_n13104_ | ~new_n4696_;
  assign new_n4232_ = ~new_n15934_ | ~new_n1953_;
  assign new_n4233_ = ~new_n2964_ | ~new_n4229_;
  assign new_n4234_ = ~pi263 | ~po264;
  assign new_n4235_ = ~new_n1964_ | ~new_n2003_;
  assign new_n4236_ = ~new_n1962_ | ~new_n1988_;
  assign new_n4237_ = ~new_n13095_ | ~new_n2361_;
  assign new_n4238_ = ~new_n4236_ | ~new_n4237_ | ~new_n4235_;
  assign new_n4239_ = ~new_n1972_ | ~new_n2951_;
  assign new_n4240_ = ~new_n13095_ | ~new_n4696_;
  assign new_n4241_ = ~new_n15838_ | ~new_n1953_;
  assign new_n4242_ = ~new_n2964_ | ~new_n4238_;
  assign new_n4243_ = ~pi264 | ~po264;
  assign new_n4244_ = ~new_n1964_ | ~new_n2004_;
  assign new_n4245_ = ~new_n1962_ | ~new_n1995_;
  assign new_n4246_ = ~pi265 | ~new_n2361_;
  assign new_n4247_ = ~new_n4246_ | ~new_n4245_ | ~new_n4244_;
  assign new_n4248_ = ~new_n2388_ | ~new_n4697_;
  assign new_n4249_ = ~pi265 | ~new_n4696_;
  assign new_n4250_ = ~new_n15928_ | ~new_n1953_;
  assign new_n4251_ = ~new_n2964_ | ~new_n4247_;
  assign new_n4252_ = ~pi265 | ~po264;
  assign new_n4253_ = ~new_n1964_ | ~new_n1997_;
  assign new_n4254_ = ~new_n1962_ | ~new_n2010_;
  assign new_n4255_ = ~new_n13083_ | ~new_n2361_;
  assign new_n4256_ = ~new_n4255_ | ~new_n4254_ | ~new_n4253_;
  assign new_n4257_ = ~new_n2409_ | ~new_n4697_;
  assign new_n4258_ = ~new_n13083_ | ~new_n4696_;
  assign new_n4259_ = ~new_n15916_ | ~new_n1953_;
  assign new_n4260_ = ~new_n2964_ | ~new_n4256_;
  assign new_n4261_ = ~pi266 | ~po264;
  assign new_n4262_ = ~new_n1964_ | ~new_n1980_;
  assign new_n4263_ = ~new_n1962_ | ~new_n1982_;
  assign new_n4264_ = ~new_n13088_ | ~new_n2361_;
  assign new_n4265_ = ~new_n4264_ | ~new_n4263_ | ~new_n4262_;
  assign new_n4266_ = ~new_n1972_ | ~new_n2944_;
  assign new_n4267_ = ~new_n13088_ | ~new_n4696_;
  assign new_n4268_ = ~new_n15921_ | ~new_n1953_;
  assign new_n4269_ = ~new_n2964_ | ~new_n4265_;
  assign new_n4270_ = ~pi267 | ~po264;
  assign new_n4271_ = ~new_n1964_ | ~new_n2009_;
  assign new_n4272_ = ~new_n1962_ | ~new_n2003_;
  assign new_n4273_ = ~new_n13097_ | ~new_n2361_;
  assign new_n4274_ = ~new_n4272_ | ~new_n4273_ | ~new_n4271_;
  assign new_n4275_ = ~new_n2441_ | ~new_n4697_;
  assign new_n4276_ = ~new_n13097_ | ~new_n4696_;
  assign new_n4277_ = ~new_n15929_ | ~new_n1953_;
  assign new_n4278_ = ~new_n2964_ | ~new_n4274_;
  assign new_n4279_ = ~pi268 | ~po264;
  assign new_n4280_ = ~new_n1964_ | ~new_n1995_;
  assign new_n4281_ = ~new_n1962_ | ~new_n1987_;
  assign new_n4282_ = ~new_n13032_ | ~new_n2361_;
  assign new_n4283_ = ~new_n4282_ | ~new_n4281_ | ~new_n4280_;
  assign new_n4284_ = ~new_n2394_ | ~new_n4697_;
  assign new_n4285_ = ~new_n13032_ | ~new_n4696_;
  assign new_n4286_ = ~new_n15840_ | ~new_n1953_;
  assign new_n4287_ = ~new_n2964_ | ~new_n4283_;
  assign new_n4288_ = ~pi269 | ~po264;
  assign new_n4289_ = ~new_n1964_ | ~new_n2010_;
  assign new_n4290_ = ~new_n1962_ | ~new_n1990_;
  assign new_n4291_ = ~new_n13106_ | ~new_n2361_;
  assign new_n4292_ = ~new_n4291_ | ~new_n4290_ | ~new_n4289_;
  assign new_n4293_ = ~new_n2415_ | ~new_n4697_;
  assign new_n4294_ = ~new_n13106_ | ~new_n4696_;
  assign new_n4295_ = ~new_n15936_ | ~new_n1953_;
  assign new_n4296_ = ~new_n2964_ | ~new_n4292_;
  assign new_n4297_ = ~pi270 | ~po264;
  assign new_n4298_ = ~new_n1964_ | ~new_n1988_;
  assign new_n4299_ = ~new_n1962_ | ~new_n1992_;
  assign new_n4300_ = ~new_n13093_ | ~new_n2361_;
  assign new_n4301_ = ~new_n4299_ | ~new_n4300_ | ~new_n4298_;
  assign new_n4302_ = ~new_n1972_ | ~new_n2949_;
  assign new_n4303_ = ~new_n13093_ | ~new_n4696_;
  assign new_n4304_ = ~new_n15925_ | ~new_n1953_;
  assign new_n4305_ = ~new_n2964_ | ~new_n4301_;
  assign new_n4306_ = ~pi271 | ~po264;
  assign new_n4307_ = ~new_n1964_ | ~new_n2007_;
  assign new_n4308_ = ~new_n1962_ | ~new_n2001_;
  assign new_n4309_ = ~new_n13102_ | ~new_n2361_;
  assign new_n4310_ = ~new_n4308_ | ~new_n4309_ | ~new_n4307_;
  assign new_n4311_ = ~new_n2427_ | ~new_n4697_;
  assign new_n4312_ = ~new_n13102_ | ~new_n4696_;
  assign new_n4313_ = ~new_n15933_ | ~new_n1953_;
  assign new_n4314_ = ~new_n2964_ | ~new_n4310_;
  assign new_n4315_ = ~pi272 | ~po264;
  assign new_n4316_ = ~new_n1964_ | ~new_n1984_;
  assign new_n4317_ = ~new_n1962_ | ~new_n1981_;
  assign new_n4318_ = ~new_n13089_ | ~new_n2361_;
  assign new_n4319_ = ~new_n4317_ | ~new_n4318_ | ~new_n4316_;
  assign new_n4320_ = ~new_n1972_ | ~new_n2945_;
  assign new_n4321_ = ~new_n13089_ | ~new_n4696_;
  assign new_n4322_ = ~new_n15922_ | ~new_n1953_;
  assign new_n4323_ = ~new_n2964_ | ~new_n4319_;
  assign new_n4324_ = ~pi273 | ~po264;
  assign new_n4325_ = ~new_n1964_ | ~new_n1998_;
  assign new_n4326_ = ~new_n1962_ | ~new_n2011_;
  assign new_n4327_ = ~new_n13084_ | ~new_n2361_;
  assign new_n4328_ = ~new_n4327_ | ~new_n4326_ | ~new_n4325_;
  assign new_n4329_ = ~new_n2406_ | ~new_n4697_;
  assign new_n4330_ = ~new_n13084_ | ~new_n4696_;
  assign new_n4331_ = ~new_n15841_ | ~new_n1953_;
  assign new_n4332_ = ~new_n2964_ | ~new_n4328_;
  assign new_n4333_ = ~pi274 | ~po264;
  assign new_n4334_ = ~new_n2382_ | ~new_n2304_;
  assign new_n4335_ = ~new_n2376_ | ~new_n4334_;
  assign new_n4336_ = ~new_n15914_ | ~new_n4744_ | ~new_n2376_;
  assign new_n4337_ = ~new_n2377_ | ~new_n2380_;
  assign new_n4338_ = ~new_n2801_ | ~new_n2940_;
  assign new_n4339_ = ~new_n2297_ | ~new_n2349_;
  assign new_n4340_ = ~new_n2292_ | ~new_n2933_ | ~new_n2290_;
  assign new_n4341_ = ~new_n2968_ | ~new_n2352_;
  assign new_n4342_ = ~new_n4340_ | ~new_n2352_;
  assign new_n4343_ = ~new_n2363_;
  assign new_n4344_ = ~new_n4343_ | ~new_n2940_;
  assign new_n4345_ = ~new_n2412_ | ~new_n4344_;
  assign new_n4346_ = ~new_n1948_ | ~new_n2010_;
  assign new_n4347_ = ~new_n2409_ | ~new_n4344_;
  assign new_n4348_ = ~new_n1948_ | ~new_n2011_;
  assign new_n4349_ = ~new_n2406_ | ~new_n4344_;
  assign new_n4350_ = ~new_n1948_ | ~new_n1997_;
  assign new_n4351_ = ~new_n2403_ | ~new_n4344_;
  assign new_n4352_ = ~new_n1948_ | ~new_n1998_;
  assign new_n4353_ = ~new_n2400_ | ~new_n4344_;
  assign new_n4354_ = ~new_n1948_ | ~new_n1994_;
  assign new_n4355_ = ~new_n2397_ | ~new_n4344_;
  assign new_n4356_ = ~new_n1948_ | ~new_n1987_;
  assign new_n4357_ = ~new_n2394_ | ~new_n4344_;
  assign new_n4358_ = ~new_n1948_ | ~new_n1991_;
  assign new_n4359_ = ~new_n2944_ | ~new_n4344_;
  assign new_n4360_ = ~new_n1948_ | ~new_n1981_;
  assign new_n4361_ = ~new_n2945_ | ~new_n4344_;
  assign new_n4362_ = ~new_n1948_ | ~new_n1980_;
  assign new_n4363_ = ~new_n2946_ | ~new_n4344_;
  assign new_n4364_ = ~new_n1948_ | ~new_n1984_;
  assign new_n4365_ = ~new_n2947_ | ~new_n4344_;
  assign new_n4366_ = ~new_n1948_ | ~new_n1985_;
  assign new_n4367_ = ~new_n2948_ | ~new_n4344_;
  assign new_n4368_ = ~new_n1948_ | ~new_n1992_;
  assign new_n4369_ = ~new_n2949_ | ~new_n4344_;
  assign new_n4370_ = ~new_n1948_ | ~new_n1993_;
  assign new_n4371_ = ~new_n2950_ | ~new_n4344_;
  assign new_n4372_ = ~new_n1948_ | ~new_n1988_;
  assign new_n4373_ = ~new_n2951_ | ~new_n4344_;
  assign new_n4374_ = ~new_n1948_ | ~new_n2002_;
  assign new_n4375_ = ~new_n2952_ | ~new_n4344_;
  assign new_n4376_ = ~new_n1948_ | ~new_n2003_;
  assign new_n4377_ = ~new_n2391_ | ~new_n4344_;
  assign new_n4378_ = ~new_n1948_ | ~new_n1995_;
  assign new_n4379_ = ~new_n2441_ | ~new_n4344_;
  assign new_n4380_ = ~new_n1948_ | ~new_n2008_;
  assign new_n4381_ = ~new_n2439_ | ~new_n4344_;
  assign new_n4382_ = ~new_n1948_ | ~new_n2009_;
  assign new_n4383_ = ~new_n2436_ | ~new_n4344_;
  assign new_n4384_ = ~new_n1948_ | ~new_n1996_;
  assign new_n4385_ = ~new_n2433_ | ~new_n4344_;
  assign new_n4386_ = ~new_n1948_ | ~new_n2000_;
  assign new_n4387_ = ~new_n2430_ | ~new_n4344_;
  assign new_n4388_ = ~new_n1948_ | ~new_n2001_;
  assign new_n4389_ = ~new_n2427_ | ~new_n4344_;
  assign new_n4390_ = ~new_n1948_ | ~new_n2006_;
  assign new_n4391_ = ~new_n2424_ | ~new_n4344_;
  assign new_n4392_ = ~new_n1948_ | ~new_n2007_;
  assign new_n4393_ = ~new_n2421_ | ~new_n4344_;
  assign new_n4394_ = ~new_n1948_ | ~new_n1999_;
  assign new_n4395_ = ~new_n2418_ | ~new_n4344_;
  assign new_n4396_ = ~new_n1948_ | ~new_n1990_;
  assign new_n4397_ = ~new_n2415_ | ~new_n4344_;
  assign new_n4398_ = ~new_n1948_ | ~new_n1989_;
  assign new_n4399_ = ~new_n2388_ | ~new_n4344_;
  assign new_n4400_ = ~new_n1948_ | ~new_n2005_;
  assign new_n4401_ = ~new_n2383_ | ~new_n4344_;
  assign new_n4402_ = ~new_n1948_ | ~new_n2004_;
  assign new_n4403_ = ~new_n3072_ | ~pi129;
  assign new_n4404_ = ~new_n1948_ | ~new_n2412_;
  assign new_n4405_ = ~new_n2363_ | ~new_n2010_;
  assign new_n4406_ = ~new_n1948_ | ~new_n2409_;
  assign new_n4407_ = ~new_n2363_ | ~new_n2011_;
  assign new_n4408_ = ~new_n1948_ | ~new_n2406_;
  assign new_n4409_ = ~new_n2363_ | ~new_n1997_;
  assign new_n4410_ = ~new_n1948_ | ~new_n2403_;
  assign new_n4411_ = ~new_n2363_ | ~new_n1998_;
  assign new_n4412_ = ~new_n1948_ | ~new_n2400_;
  assign new_n4413_ = ~new_n2363_ | ~new_n1994_;
  assign new_n4414_ = ~new_n1948_ | ~new_n2397_;
  assign new_n4415_ = ~new_n2363_ | ~new_n1987_;
  assign new_n4416_ = ~new_n1948_ | ~new_n2394_;
  assign new_n4417_ = ~new_n2363_ | ~new_n1991_;
  assign new_n4418_ = ~new_n1948_ | ~new_n2944_;
  assign new_n4419_ = ~new_n2363_ | ~new_n1981_;
  assign new_n4420_ = ~new_n1948_ | ~new_n2945_;
  assign new_n4421_ = ~new_n2363_ | ~new_n1980_;
  assign new_n4422_ = ~new_n1948_ | ~new_n2946_;
  assign new_n4423_ = ~new_n2363_ | ~new_n1984_;
  assign new_n4424_ = ~new_n1948_ | ~new_n2947_;
  assign new_n4425_ = ~new_n2363_ | ~new_n1985_;
  assign new_n4426_ = ~new_n1948_ | ~new_n2948_;
  assign new_n4427_ = ~new_n2363_ | ~new_n1992_;
  assign new_n4428_ = ~new_n1948_ | ~new_n2949_;
  assign new_n4429_ = ~new_n2363_ | ~new_n1993_;
  assign new_n4430_ = ~new_n1948_ | ~new_n2950_;
  assign new_n4431_ = ~new_n2363_ | ~new_n1988_;
  assign new_n4432_ = ~new_n1948_ | ~new_n2951_;
  assign new_n4433_ = ~new_n2363_ | ~new_n2002_;
  assign new_n4434_ = ~new_n1948_ | ~new_n2952_;
  assign new_n4435_ = ~new_n2363_ | ~new_n2003_;
  assign new_n4436_ = ~new_n1948_ | ~new_n2391_;
  assign new_n4437_ = ~new_n2363_ | ~new_n1995_;
  assign new_n4438_ = ~new_n1948_ | ~new_n2441_;
  assign new_n4439_ = ~new_n2363_ | ~new_n2008_;
  assign new_n4440_ = ~new_n1948_ | ~new_n2439_;
  assign new_n4441_ = ~new_n2363_ | ~new_n2009_;
  assign new_n4442_ = ~new_n1948_ | ~new_n2436_;
  assign new_n4443_ = ~new_n2363_ | ~new_n1996_;
  assign new_n4444_ = ~new_n1948_ | ~new_n2433_;
  assign new_n4445_ = ~new_n2363_ | ~new_n2000_;
  assign new_n4446_ = ~new_n1948_ | ~new_n2430_;
  assign new_n4447_ = ~new_n2363_ | ~new_n2001_;
  assign new_n4448_ = ~new_n1948_ | ~new_n2427_;
  assign new_n4449_ = ~new_n2363_ | ~new_n2006_;
  assign new_n4450_ = ~new_n1948_ | ~new_n2424_;
  assign new_n4451_ = ~new_n2363_ | ~new_n2007_;
  assign new_n4452_ = ~new_n1948_ | ~new_n2421_;
  assign new_n4453_ = ~new_n2363_ | ~new_n1999_;
  assign new_n4454_ = ~new_n1948_ | ~new_n2418_;
  assign new_n4455_ = ~new_n2363_ | ~new_n1990_;
  assign new_n4456_ = ~new_n1948_ | ~new_n2415_;
  assign new_n4457_ = ~new_n2363_ | ~new_n1989_;
  assign new_n4458_ = ~new_n1948_ | ~new_n2388_;
  assign new_n4459_ = ~new_n2363_ | ~new_n2005_;
  assign new_n4460_ = ~new_n1948_ | ~new_n2383_;
  assign new_n4461_ = ~new_n2363_ | ~new_n2004_;
  assign new_n4462_ = ~new_n3072_ | ~new_n2381_;
  assign new_n4463_ = ~new_n2364_;
  assign new_n4464_ = ~new_n2365_;
  assign new_n4465_ = ~new_n4726_ | ~new_n2377_;
  assign new_n4466_ = ~new_n2364_ | ~new_n2366_;
  assign new_n4467_ = ~new_n1978_ | ~new_n4466_;
  assign new_n4468_ = ~new_n1941_ | ~new_n2371_;
  assign new_n4469_ = ~new_n2367_;
  assign new_n4470_ = ~new_n1979_ | ~new_n4469_;
  assign new_n4471_ = ~new_n2010_ | ~new_n1954_;
  assign new_n4472_ = ~new_n2412_ | ~new_n4470_;
  assign new_n4473_ = ~new_n4467_ | ~new_n2010_;
  assign new_n4474_ = ~new_n2011_ | ~new_n1954_;
  assign new_n4475_ = ~new_n2409_ | ~new_n4470_;
  assign new_n4476_ = ~new_n4467_ | ~new_n2011_;
  assign new_n4477_ = ~new_n1997_ | ~new_n1954_;
  assign new_n4478_ = ~new_n2406_ | ~new_n4470_;
  assign new_n4479_ = ~new_n4467_ | ~new_n1997_;
  assign new_n4480_ = ~new_n1998_ | ~new_n1954_;
  assign new_n4481_ = ~new_n2403_ | ~new_n4470_;
  assign new_n4482_ = ~new_n4467_ | ~new_n1998_;
  assign new_n4483_ = ~new_n1994_ | ~new_n1954_;
  assign new_n4484_ = ~new_n2400_ | ~new_n4470_;
  assign new_n4485_ = ~new_n4467_ | ~new_n1994_;
  assign new_n4486_ = ~new_n1987_ | ~new_n1954_;
  assign new_n4487_ = ~new_n2397_ | ~new_n4470_;
  assign new_n4488_ = ~new_n4467_ | ~new_n1987_;
  assign new_n4489_ = ~new_n13735_ | ~new_n1954_;
  assign new_n4490_ = ~new_n2953_ | ~new_n4470_;
  assign new_n4491_ = ~new_n4467_ | ~new_n1983_;
  assign new_n4492_ = ~new_n13733_ | ~new_n1954_;
  assign new_n4493_ = ~new_n2954_ | ~new_n4470_;
  assign new_n4494_ = ~new_n4467_ | ~new_n1986_;
  assign new_n4495_ = ~new_n1991_ | ~new_n1954_;
  assign new_n4496_ = ~new_n2394_ | ~new_n4470_;
  assign new_n4497_ = ~new_n4467_ | ~new_n1991_;
  assign new_n4498_ = ~new_n1982_ | ~new_n1954_;
  assign new_n4499_ = ~new_n2955_ | ~new_n4470_;
  assign new_n4500_ = ~new_n4467_ | ~new_n1982_;
  assign new_n4501_ = ~new_n1981_ | ~new_n1954_;
  assign new_n4502_ = ~new_n2944_ | ~new_n4470_;
  assign new_n4503_ = ~new_n4467_ | ~new_n1981_;
  assign new_n4504_ = ~new_n1980_ | ~new_n1954_;
  assign new_n4505_ = ~new_n2945_ | ~new_n4470_;
  assign new_n4506_ = ~new_n4467_ | ~new_n1980_;
  assign new_n4507_ = ~new_n1984_ | ~new_n1954_;
  assign new_n4508_ = ~new_n2946_ | ~new_n4470_;
  assign new_n4509_ = ~new_n4467_ | ~new_n1984_;
  assign new_n4510_ = ~new_n1985_ | ~new_n1954_;
  assign new_n4511_ = ~new_n2947_ | ~new_n4470_;
  assign new_n4512_ = ~new_n4467_ | ~new_n1985_;
  assign new_n4513_ = ~new_n1992_ | ~new_n1954_;
  assign new_n4514_ = ~new_n2948_ | ~new_n4470_;
  assign new_n4515_ = ~new_n4467_ | ~new_n1992_;
  assign new_n4516_ = ~new_n1993_ | ~new_n1954_;
  assign new_n4517_ = ~new_n2949_ | ~new_n4470_;
  assign new_n4518_ = ~new_n4467_ | ~new_n1993_;
  assign new_n4519_ = ~new_n1988_ | ~new_n1954_;
  assign new_n4520_ = ~new_n2950_ | ~new_n4470_;
  assign new_n4521_ = ~new_n4467_ | ~new_n1988_;
  assign new_n4522_ = ~new_n2002_ | ~new_n1954_;
  assign new_n4523_ = ~new_n2951_ | ~new_n4470_;
  assign new_n4524_ = ~new_n4467_ | ~new_n2002_;
  assign new_n4525_ = ~new_n2003_ | ~new_n1954_;
  assign new_n4526_ = ~new_n2952_ | ~new_n4470_;
  assign new_n4527_ = ~new_n4467_ | ~new_n2003_;
  assign new_n4528_ = ~new_n1995_ | ~new_n1954_;
  assign new_n4529_ = ~new_n2391_ | ~new_n4470_;
  assign new_n4530_ = ~new_n4467_ | ~new_n1995_;
  assign new_n4531_ = ~new_n2008_ | ~new_n1954_;
  assign new_n4532_ = ~new_n2441_ | ~new_n4470_;
  assign new_n4533_ = ~new_n4467_ | ~new_n2008_;
  assign new_n4534_ = ~new_n2009_ | ~new_n1954_;
  assign new_n4535_ = ~new_n2439_ | ~new_n4470_;
  assign new_n4536_ = ~new_n4467_ | ~new_n2009_;
  assign new_n4537_ = ~new_n1996_ | ~new_n1954_;
  assign new_n4538_ = ~new_n2436_ | ~new_n4470_;
  assign new_n4539_ = ~new_n4467_ | ~new_n1996_;
  assign new_n4540_ = ~new_n2000_ | ~new_n1954_;
  assign new_n4541_ = ~new_n2433_ | ~new_n4470_;
  assign new_n4542_ = ~new_n4467_ | ~new_n2000_;
  assign new_n4543_ = ~new_n2001_ | ~new_n1954_;
  assign new_n4544_ = ~new_n2430_ | ~new_n4470_;
  assign new_n4545_ = ~new_n4467_ | ~new_n2001_;
  assign new_n4546_ = ~new_n2006_ | ~new_n1954_;
  assign new_n4547_ = ~new_n2427_ | ~new_n4470_;
  assign new_n4548_ = ~new_n4467_ | ~new_n2006_;
  assign new_n4549_ = ~new_n2007_ | ~new_n1954_;
  assign new_n4550_ = ~new_n2424_ | ~new_n4470_;
  assign new_n4551_ = ~new_n4467_ | ~new_n2007_;
  assign new_n4552_ = ~new_n1999_ | ~new_n1954_;
  assign new_n4553_ = ~new_n2421_ | ~new_n4470_;
  assign new_n4554_ = ~new_n4467_ | ~new_n1999_;
  assign new_n4555_ = ~new_n1990_ | ~new_n1954_;
  assign new_n4556_ = ~new_n2418_ | ~new_n4470_;
  assign new_n4557_ = ~new_n4467_ | ~new_n1990_;
  assign new_n4558_ = ~new_n1989_ | ~new_n1954_;
  assign new_n4559_ = ~new_n2415_ | ~new_n4470_;
  assign new_n4560_ = ~new_n4467_ | ~new_n1989_;
  assign new_n4561_ = ~new_n2005_ | ~new_n1954_;
  assign new_n4562_ = ~new_n2388_ | ~new_n4470_;
  assign new_n4563_ = ~new_n4467_ | ~new_n2005_;
  assign new_n4564_ = ~new_n2004_ | ~new_n1954_;
  assign new_n4565_ = ~new_n2383_ | ~new_n4470_;
  assign new_n4566_ = ~new_n4467_ | ~new_n2004_;
  assign new_n4567_ = ~new_n2367_ | ~new_n2366_;
  assign new_n4568_ = ~new_n1979_ | ~new_n4567_;
  assign new_n4569_ = ~new_n1955_ | ~new_n2010_;
  assign new_n4570_ = ~new_n2412_ | ~new_n2365_;
  assign new_n4571_ = ~new_n4568_ | ~new_n2010_;
  assign new_n4572_ = ~new_n4713_ | ~new_n2011_;
  assign new_n4573_ = ~new_n1955_ | ~new_n2011_;
  assign new_n4574_ = ~new_n2409_ | ~new_n2365_;
  assign new_n4575_ = ~new_n4568_ | ~new_n2011_;
  assign new_n4576_ = ~new_n4713_ | ~new_n1997_;
  assign new_n4577_ = ~new_n1955_ | ~new_n1997_;
  assign new_n4578_ = ~new_n2406_ | ~new_n2365_;
  assign new_n4579_ = ~new_n4568_ | ~new_n1997_;
  assign new_n4580_ = ~new_n4713_ | ~new_n1998_;
  assign new_n4581_ = ~new_n1955_ | ~new_n1998_;
  assign new_n4582_ = ~new_n2403_ | ~new_n2365_;
  assign new_n4583_ = ~new_n4568_ | ~new_n1998_;
  assign new_n4584_ = ~new_n4713_ | ~new_n1994_;
  assign new_n4585_ = ~new_n1955_ | ~new_n1994_;
  assign new_n4586_ = ~new_n2400_ | ~new_n2365_;
  assign new_n4587_ = ~new_n4568_ | ~new_n1994_;
  assign new_n4588_ = ~new_n4713_ | ~new_n1987_;
  assign new_n4589_ = ~new_n1955_ | ~new_n1987_;
  assign new_n4590_ = ~new_n2397_ | ~new_n2365_;
  assign new_n4591_ = ~new_n4568_ | ~new_n1987_;
  assign new_n4592_ = ~new_n4713_ | ~new_n1991_;
  assign new_n4593_ = ~new_n1955_ | ~new_n13735_;
  assign new_n4594_ = ~new_n2953_ | ~new_n2365_;
  assign new_n4595_ = ~new_n4568_ | ~new_n1983_;
  assign new_n4596_ = ~new_n1955_ | ~new_n13733_;
  assign new_n4597_ = ~new_n2954_ | ~new_n2365_;
  assign new_n4598_ = ~new_n4568_ | ~new_n1986_;
  assign new_n4599_ = ~new_n1955_ | ~new_n1991_;
  assign new_n4600_ = ~new_n2394_ | ~new_n2365_;
  assign new_n4601_ = ~new_n4568_ | ~new_n1991_;
  assign new_n4602_ = ~new_n4713_ | ~new_n1995_;
  assign new_n4603_ = ~new_n1955_ | ~new_n1982_;
  assign new_n4604_ = ~new_n2955_ | ~new_n2365_;
  assign new_n4605_ = ~new_n4568_ | ~new_n1982_;
  assign new_n4606_ = ~new_n4713_ | ~new_n1981_;
  assign new_n4607_ = ~new_n1955_ | ~new_n1981_;
  assign new_n4608_ = ~new_n2944_ | ~new_n2365_;
  assign new_n4609_ = ~new_n4568_ | ~new_n1981_;
  assign new_n4610_ = ~new_n4713_ | ~new_n1980_;
  assign new_n4611_ = ~new_n1955_ | ~new_n1980_;
  assign new_n4612_ = ~new_n2945_ | ~new_n2365_;
  assign new_n4613_ = ~new_n4568_ | ~new_n1980_;
  assign new_n4614_ = ~new_n4713_ | ~new_n1984_;
  assign new_n4615_ = ~new_n1955_ | ~new_n1984_;
  assign new_n4616_ = ~new_n2946_ | ~new_n2365_;
  assign new_n4617_ = ~new_n4568_ | ~new_n1984_;
  assign new_n4618_ = ~new_n4713_ | ~new_n1985_;
  assign new_n4619_ = ~new_n1955_ | ~new_n1985_;
  assign new_n4620_ = ~new_n2947_ | ~new_n2365_;
  assign new_n4621_ = ~new_n4568_ | ~new_n1985_;
  assign new_n4622_ = ~new_n4713_ | ~new_n1992_;
  assign new_n4623_ = ~new_n1955_ | ~new_n1992_;
  assign new_n4624_ = ~new_n2948_ | ~new_n2365_;
  assign new_n4625_ = ~new_n4568_ | ~new_n1992_;
  assign new_n4626_ = ~new_n4713_ | ~new_n1993_;
  assign new_n4627_ = ~new_n1955_ | ~new_n1993_;
  assign new_n4628_ = ~new_n2949_ | ~new_n2365_;
  assign new_n4629_ = ~new_n4568_ | ~new_n1993_;
  assign new_n4630_ = ~new_n4713_ | ~new_n1988_;
  assign new_n4631_ = ~new_n1955_ | ~new_n1988_;
  assign new_n4632_ = ~new_n2950_ | ~new_n2365_;
  assign new_n4633_ = ~new_n4568_ | ~new_n1988_;
  assign new_n4634_ = ~new_n4713_ | ~new_n2002_;
  assign new_n4635_ = ~new_n1955_ | ~new_n2002_;
  assign new_n4636_ = ~new_n2951_ | ~new_n2365_;
  assign new_n4637_ = ~new_n4568_ | ~new_n2002_;
  assign new_n4638_ = ~new_n4713_ | ~new_n2003_;
  assign new_n4639_ = ~new_n1955_ | ~new_n2003_;
  assign new_n4640_ = ~new_n2952_ | ~new_n2365_;
  assign new_n4641_ = ~new_n4568_ | ~new_n2003_;
  assign new_n4642_ = ~new_n4713_ | ~new_n2008_;
  assign new_n4643_ = ~new_n1955_ | ~new_n1995_;
  assign new_n4644_ = ~new_n2391_ | ~new_n2365_;
  assign new_n4645_ = ~new_n4568_ | ~new_n1995_;
  assign new_n4646_ = ~new_n4713_ | ~new_n2005_;
  assign new_n4647_ = ~new_n1955_ | ~new_n2008_;
  assign new_n4648_ = ~new_n2441_ | ~new_n2365_;
  assign new_n4649_ = ~new_n4568_ | ~new_n2008_;
  assign new_n4650_ = ~new_n4713_ | ~new_n2009_;
  assign new_n4651_ = ~new_n1955_ | ~new_n2009_;
  assign new_n4652_ = ~new_n2439_ | ~new_n2365_;
  assign new_n4653_ = ~new_n4568_ | ~new_n2009_;
  assign new_n4654_ = ~new_n4713_ | ~new_n1996_;
  assign new_n4655_ = ~new_n1955_ | ~new_n1996_;
  assign new_n4656_ = ~new_n2436_ | ~new_n2365_;
  assign new_n4657_ = ~new_n4568_ | ~new_n1996_;
  assign new_n4658_ = ~new_n4713_ | ~new_n2000_;
  assign new_n4659_ = ~new_n1955_ | ~new_n2000_;
  assign new_n4660_ = ~new_n2433_ | ~new_n2365_;
  assign new_n4661_ = ~new_n4568_ | ~new_n2000_;
  assign new_n4662_ = ~new_n4713_ | ~new_n2001_;
  assign new_n4663_ = ~new_n1955_ | ~new_n2001_;
  assign new_n4664_ = ~new_n2430_ | ~new_n2365_;
  assign new_n4665_ = ~new_n4568_ | ~new_n2001_;
  assign new_n4666_ = ~new_n4713_ | ~new_n2006_;
  assign new_n4667_ = ~new_n1955_ | ~new_n2006_;
  assign new_n4668_ = ~new_n2427_ | ~new_n2365_;
  assign new_n4669_ = ~new_n4568_ | ~new_n2006_;
  assign new_n4670_ = ~new_n4713_ | ~new_n2007_;
  assign new_n4671_ = ~new_n1955_ | ~new_n2007_;
  assign new_n4672_ = ~new_n2424_ | ~new_n2365_;
  assign new_n4673_ = ~new_n4568_ | ~new_n2007_;
  assign new_n4674_ = ~new_n4713_ | ~new_n1999_;
  assign new_n4675_ = ~new_n1955_ | ~new_n1999_;
  assign new_n4676_ = ~new_n2421_ | ~new_n2365_;
  assign new_n4677_ = ~new_n4568_ | ~new_n1999_;
  assign new_n4678_ = ~new_n4713_ | ~new_n1990_;
  assign new_n4679_ = ~new_n1955_ | ~new_n1990_;
  assign new_n4680_ = ~new_n2418_ | ~new_n2365_;
  assign new_n4681_ = ~new_n4568_ | ~new_n1990_;
  assign new_n4682_ = ~new_n4713_ | ~new_n1989_;
  assign new_n4683_ = ~new_n1955_ | ~new_n1989_;
  assign new_n4684_ = ~new_n2415_ | ~new_n2365_;
  assign new_n4685_ = ~new_n4568_ | ~new_n1989_;
  assign new_n4686_ = ~new_n4713_ | ~new_n2010_;
  assign new_n4687_ = ~new_n1955_ | ~new_n2005_;
  assign new_n4688_ = ~new_n2388_ | ~new_n2365_;
  assign new_n4689_ = ~new_n4568_ | ~new_n2005_;
  assign new_n4690_ = ~new_n4713_ | ~new_n2004_;
  assign new_n4691_ = ~new_n1955_ | ~new_n2004_;
  assign new_n4692_ = ~new_n2383_ | ~new_n2365_;
  assign new_n4693_ = ~new_n4568_ | ~new_n2004_;
  assign new_n4694_ = ~new_n2965_ | ~new_n2361_;
  assign new_n4695_ = ~new_n2942_ | ~new_n2965_;
  assign new_n4696_ = ~new_n1977_ | ~new_n4694_;
  assign new_n4697_ = ~new_n4695_ | ~new_n2966_;
  assign new_n4698_ = ~new_n4702_ | ~new_n4708_;
  assign new_n4699_ = ~new_n15169_ | ~new_n4058_;
  assign new_n4700_ = ~pi057 | ~new_n2879_;
  assign new_n4701_ = ~pi064 | ~new_n13498_;
  assign new_n4702_ = ~new_n2368_;
  assign new_n4703_ = ~pi058 | ~new_n2879_;
  assign new_n4704_ = ~pi064 | ~new_n13651_;
  assign new_n4705_ = ~new_n2369_;
  assign new_n4706_ = ~pi059 | ~new_n2879_;
  assign new_n4707_ = ~pi064 | ~new_n13499_;
  assign new_n4708_ = ~new_n2370_;
  assign new_n4709_ = ~new_n2368_ | ~new_n2286_;
  assign new_n4710_ = ~pi245 | ~new_n2973_ | ~new_n4702_;
  assign new_n4711_ = ~pi056 | ~new_n2879_;
  assign new_n4712_ = ~pi064 | ~new_n13497_;
  assign new_n4713_ = ~new_n2371_;
  assign new_n4714_ = ~pi065 | ~new_n2880_;
  assign new_n4715_ = ~new_n2961_ | ~new_n3073_;
  assign new_n4716_ = ~pi066 | ~new_n2880_;
  assign new_n4717_ = ~new_n2961_ | ~new_n3074_;
  assign new_n4718_ = ~pi055 | ~new_n2879_;
  assign new_n4719_ = ~pi064 | ~new_n13496_;
  assign new_n4720_ = ~new_n2378_;
  assign new_n4721_ = ~pi052 | ~new_n2879_;
  assign new_n4722_ = ~pi064 | ~new_n13494_;
  assign new_n4723_ = ~new_n2379_;
  assign new_n4724_ = ~pi053 | ~new_n2879_;
  assign new_n4725_ = ~pi064 | ~new_n13495_;
  assign new_n4726_ = ~new_n2380_;
  assign new_n4727_ = ~pi054 | ~new_n2879_;
  assign new_n4728_ = ~pi064 | ~new_n13654_;
  assign new_n4729_ = ~new_n2377_;
  assign new_n4730_ = ~pi063 | ~new_n2879_;
  assign new_n4731_ = ~pi064 | ~new_n13646_;
  assign new_n4732_ = ~new_n2374_;
  assign new_n4733_ = ~pi062 | ~new_n2879_;
  assign new_n4734_ = ~pi064 | ~new_n13501_;
  assign new_n4735_ = ~new_n2375_;
  assign new_n4736_ = ~pi061 | ~new_n2879_;
  assign new_n4737_ = ~pi064 | ~new_n13500_;
  assign new_n4738_ = ~new_n2376_;
  assign new_n4739_ = ~pi033 | ~new_n2879_;
  assign new_n4740_ = ~pi064 | ~pi033;
  assign new_n4741_ = ~new_n2381_;
  assign new_n4742_ = ~pi060 | ~new_n2879_;
  assign new_n4743_ = ~pi064 | ~new_n13523_;
  assign new_n4744_ = ~new_n2382_;
  assign new_n4745_ = ~new_n1626_ | ~new_n2881_;
  assign new_n4746_ = ~new_n2941_ | ~new_n2381_;
  assign new_n4747_ = ~new_n2383_;
  assign new_n4748_ = ~new_n2378_ | ~new_n4729_;
  assign new_n4749_ = ~new_n4720_ | ~new_n3105_;
  assign new_n4750_ = ~pi066 | ~new_n3071_;
  assign new_n4751_ = ~new_n3074_ | ~new_n2287_;
  assign new_n4752_ = ~new_n2385_;
  assign new_n4753_ = ~new_n4698_ | ~new_n2287_;
  assign new_n4754_ = ~pi065 | ~new_n3071_;
  assign new_n4755_ = ~new_n2384_;
  assign new_n4756_ = ~pi097 | ~new_n2882_;
  assign new_n4757_ = ~new_n2960_ | ~new_n3125_;
  assign new_n4758_ = ~pi034 | ~new_n2879_;
  assign new_n4759_ = ~pi064 | ~new_n13521_;
  assign new_n4760_ = ~new_n1615_ | ~new_n2881_;
  assign new_n4761_ = ~new_n2387_ | ~new_n2941_;
  assign new_n4762_ = ~new_n2388_;
  assign new_n4763_ = ~pi098 | ~new_n2882_;
  assign new_n4764_ = ~new_n2960_ | ~new_n3149_;
  assign new_n4765_ = ~pi035 | ~new_n2879_;
  assign new_n4766_ = ~pi064 | ~new_n13502_;
  assign new_n4767_ = ~new_n1604_ | ~new_n2881_;
  assign new_n4768_ = ~new_n2390_ | ~new_n2941_;
  assign new_n4769_ = ~new_n2391_;
  assign new_n4770_ = ~pi099 | ~new_n2882_;
  assign new_n4771_ = ~new_n2960_ | ~new_n3168_;
  assign new_n4772_ = ~pi036 | ~new_n2879_;
  assign new_n4773_ = ~pi064 | ~new_n13503_;
  assign new_n4774_ = ~new_n1601_ | ~new_n2881_;
  assign new_n4775_ = ~new_n2393_ | ~new_n2941_;
  assign new_n4776_ = ~new_n2394_;
  assign new_n4777_ = ~pi100 | ~new_n2882_;
  assign new_n4778_ = ~new_n2960_ | ~new_n3187_;
  assign new_n4779_ = ~pi037 | ~new_n2879_;
  assign new_n4780_ = ~pi064 | ~new_n13504_;
  assign new_n4781_ = ~new_n1600_ | ~new_n2881_;
  assign new_n4782_ = ~new_n2396_ | ~new_n2941_;
  assign new_n4783_ = ~new_n2397_;
  assign new_n4784_ = ~pi101 | ~new_n2882_;
  assign new_n4785_ = ~new_n2960_ | ~new_n3206_;
  assign new_n4786_ = ~pi038 | ~new_n2879_;
  assign new_n4787_ = ~pi064 | ~new_n13643_;
  assign new_n4788_ = ~new_n1599_ | ~new_n2881_;
  assign new_n4789_ = ~new_n2399_ | ~new_n2941_;
  assign new_n4790_ = ~new_n2400_;
  assign new_n4791_ = ~pi102 | ~new_n2882_;
  assign new_n4792_ = ~new_n2960_ | ~new_n3225_;
  assign new_n4793_ = ~pi039 | ~new_n2879_;
  assign new_n4794_ = ~pi064 | ~new_n13505_;
  assign new_n4795_ = ~new_n1598_ | ~new_n2881_;
  assign new_n4796_ = ~new_n2402_ | ~new_n2941_;
  assign new_n4797_ = ~new_n2403_;
  assign new_n4798_ = ~pi103 | ~new_n2882_;
  assign new_n4799_ = ~new_n2960_ | ~new_n3244_;
  assign new_n4800_ = ~pi040 | ~new_n2879_;
  assign new_n4801_ = ~pi064 | ~new_n13506_;
  assign new_n4802_ = ~new_n1597_ | ~new_n2881_;
  assign new_n4803_ = ~new_n2405_ | ~new_n2941_;
  assign new_n4804_ = ~new_n2406_;
  assign new_n4805_ = ~pi104 | ~new_n2882_;
  assign new_n4806_ = ~new_n2960_ | ~new_n3263_;
  assign new_n4807_ = ~pi041 | ~new_n2879_;
  assign new_n4808_ = ~pi064 | ~new_n13507_;
  assign new_n4809_ = ~new_n1596_ | ~new_n2881_;
  assign new_n4810_ = ~new_n2408_ | ~new_n2941_;
  assign new_n4811_ = ~new_n2409_;
  assign new_n4812_ = ~pi105 | ~new_n2882_;
  assign new_n4813_ = ~new_n2960_ | ~new_n3282_;
  assign new_n4814_ = ~pi042 | ~new_n2879_;
  assign new_n4815_ = ~pi064 | ~new_n13641_;
  assign new_n4816_ = ~new_n1595_ | ~new_n2881_;
  assign new_n4817_ = ~new_n2411_ | ~new_n2941_;
  assign new_n4818_ = ~new_n2412_;
  assign new_n4819_ = ~pi106 | ~new_n2882_;
  assign new_n4820_ = ~new_n2960_ | ~new_n3301_;
  assign new_n4821_ = ~pi043 | ~new_n2879_;
  assign new_n4822_ = ~pi064 | ~new_n13487_;
  assign new_n4823_ = ~new_n1625_ | ~new_n2881_;
  assign new_n4824_ = ~new_n2414_ | ~new_n2941_;
  assign new_n4825_ = ~new_n2415_;
  assign new_n4826_ = ~pi107 | ~new_n2882_;
  assign new_n4827_ = ~new_n2960_ | ~new_n3320_;
  assign new_n4828_ = ~pi044 | ~new_n2879_;
  assign new_n4829_ = ~pi064 | ~new_n13488_;
  assign new_n4830_ = ~new_n1624_ | ~new_n2881_;
  assign new_n4831_ = ~new_n2417_ | ~new_n2941_;
  assign new_n4832_ = ~new_n2418_;
  assign new_n4833_ = ~pi108 | ~new_n2882_;
  assign new_n4834_ = ~new_n2960_ | ~new_n3339_;
  assign new_n4835_ = ~pi045 | ~new_n2879_;
  assign new_n4836_ = ~pi064 | ~new_n13489_;
  assign new_n4837_ = ~new_n1623_ | ~new_n2881_;
  assign new_n4838_ = ~new_n2420_ | ~new_n2941_;
  assign new_n4839_ = ~new_n2421_;
  assign new_n4840_ = ~pi109 | ~new_n2882_;
  assign new_n4841_ = ~new_n2960_ | ~new_n3358_;
  assign new_n4842_ = ~pi046 | ~new_n2879_;
  assign new_n4843_ = ~pi064 | ~new_n13660_;
  assign new_n4844_ = ~new_n1622_ | ~new_n2881_;
  assign new_n4845_ = ~new_n2423_ | ~new_n2941_;
  assign new_n4846_ = ~new_n2424_;
  assign new_n4847_ = ~pi110 | ~new_n2882_;
  assign new_n4848_ = ~new_n2960_ | ~new_n3377_;
  assign new_n4849_ = ~pi047 | ~new_n2879_;
  assign new_n4850_ = ~pi064 | ~new_n13490_;
  assign new_n4851_ = ~new_n1621_ | ~new_n2881_;
  assign new_n4852_ = ~new_n2426_ | ~new_n2941_;
  assign new_n4853_ = ~new_n2427_;
  assign new_n4854_ = ~pi111 | ~new_n2882_;
  assign new_n4855_ = ~new_n2960_ | ~new_n3396_;
  assign new_n4856_ = ~pi048 | ~new_n2879_;
  assign new_n4857_ = ~pi064 | ~new_n13491_;
  assign new_n4858_ = ~new_n1620_ | ~new_n2881_;
  assign new_n4859_ = ~new_n2429_ | ~new_n2941_;
  assign new_n4860_ = ~new_n2430_;
  assign new_n4861_ = ~pi112 | ~new_n2882_;
  assign new_n4862_ = ~new_n2960_ | ~new_n3415_;
  assign new_n4863_ = ~pi049 | ~new_n2879_;
  assign new_n4864_ = ~pi064 | ~new_n13492_;
  assign new_n4865_ = ~new_n1619_ | ~new_n2881_;
  assign new_n4866_ = ~new_n2432_ | ~new_n2941_;
  assign new_n4867_ = ~new_n2433_;
  assign new_n4868_ = ~pi113 | ~new_n2882_;
  assign new_n4869_ = ~new_n2960_ | ~new_n3434_;
  assign new_n4870_ = ~pi050 | ~new_n2879_;
  assign new_n4871_ = ~pi064 | ~new_n13658_;
  assign new_n4872_ = ~new_n1618_ | ~new_n2881_;
  assign new_n4873_ = ~new_n2435_ | ~new_n2941_;
  assign new_n4874_ = ~new_n2436_;
  assign new_n4875_ = ~pi114 | ~new_n2882_;
  assign new_n4876_ = ~new_n2960_ | ~new_n3453_;
  assign new_n4877_ = ~pi051 | ~new_n2879_;
  assign new_n4878_ = ~pi064 | ~new_n13493_;
  assign new_n4879_ = ~new_n1617_ | ~new_n2881_;
  assign new_n4880_ = ~new_n2438_ | ~new_n2941_;
  assign new_n4881_ = ~new_n2439_;
  assign new_n4882_ = ~pi115 | ~new_n2882_;
  assign new_n4883_ = ~new_n2960_ | ~new_n3472_;
  assign new_n4884_ = ~new_n1616_ | ~new_n2881_;
  assign new_n4885_ = ~new_n2941_ | ~new_n2379_;
  assign new_n4886_ = ~new_n2441_;
  assign new_n4887_ = ~pi116 | ~new_n2882_;
  assign new_n4888_ = ~new_n2960_ | ~new_n3491_;
  assign new_n4889_ = ~pi117 | ~new_n2882_;
  assign new_n4890_ = ~new_n2960_ | ~new_n3510_;
  assign new_n4891_ = ~pi118 | ~new_n2882_;
  assign new_n4892_ = ~new_n2960_ | ~new_n3529_;
  assign new_n4893_ = ~pi119 | ~new_n2882_;
  assign new_n4894_ = ~new_n2960_ | ~new_n3548_;
  assign new_n4895_ = ~pi120 | ~new_n2882_;
  assign new_n4896_ = ~new_n2960_ | ~new_n3567_;
  assign new_n4897_ = ~pi121 | ~new_n2882_;
  assign new_n4898_ = ~new_n2960_ | ~new_n3586_;
  assign new_n4899_ = ~pi122 | ~new_n2882_;
  assign new_n4900_ = ~new_n2960_ | ~new_n3605_;
  assign new_n4901_ = ~pi123 | ~new_n2882_;
  assign new_n4902_ = ~new_n2960_ | ~new_n3624_;
  assign new_n4903_ = ~pi124 | ~new_n2882_;
  assign new_n4904_ = ~new_n2960_ | ~new_n3643_;
  assign new_n4905_ = ~pi125 | ~new_n2882_;
  assign new_n4906_ = ~new_n2960_ | ~new_n3662_;
  assign new_n4907_ = ~pi126 | ~new_n2882_;
  assign new_n4908_ = ~new_n2960_ | ~new_n3682_;
  assign new_n4909_ = ~pi127 | ~new_n2882_;
  assign new_n4910_ = ~new_n2960_ | ~new_n3689_;
  assign new_n4911_ = ~pi128 | ~new_n2882_;
  assign new_n4912_ = ~new_n2960_ | ~new_n3692_;
  assign new_n4913_ = ~pi129 | ~new_n2883_;
  assign new_n4914_ = ~new_n2959_ | ~new_n3125_;
  assign new_n4915_ = ~pi130 | ~new_n2883_;
  assign new_n4916_ = ~new_n2959_ | ~new_n3149_;
  assign new_n4917_ = ~pi131 | ~new_n2883_;
  assign new_n4918_ = ~new_n2959_ | ~new_n3168_;
  assign new_n4919_ = ~pi132 | ~new_n2883_;
  assign new_n4920_ = ~new_n2959_ | ~new_n3187_;
  assign new_n4921_ = ~pi133 | ~new_n2883_;
  assign new_n4922_ = ~new_n2959_ | ~new_n3206_;
  assign new_n4923_ = ~pi134 | ~new_n2883_;
  assign new_n4924_ = ~new_n2959_ | ~new_n3225_;
  assign new_n4925_ = ~pi135 | ~new_n2883_;
  assign new_n4926_ = ~new_n2959_ | ~new_n3244_;
  assign new_n4927_ = ~pi136 | ~new_n2883_;
  assign new_n4928_ = ~new_n2959_ | ~new_n3263_;
  assign new_n4929_ = ~pi137 | ~new_n2883_;
  assign new_n4930_ = ~new_n2959_ | ~new_n3282_;
  assign new_n4931_ = ~pi138 | ~new_n2883_;
  assign new_n4932_ = ~new_n2959_ | ~new_n3301_;
  assign new_n4933_ = ~pi139 | ~new_n2883_;
  assign new_n4934_ = ~new_n2959_ | ~new_n3320_;
  assign new_n4935_ = ~pi140 | ~new_n2883_;
  assign new_n4936_ = ~new_n2959_ | ~new_n3339_;
  assign new_n4937_ = ~pi141 | ~new_n2883_;
  assign new_n4938_ = ~new_n2959_ | ~new_n3358_;
  assign new_n4939_ = ~pi142 | ~new_n2883_;
  assign new_n4940_ = ~new_n2959_ | ~new_n3377_;
  assign new_n4941_ = ~pi143 | ~new_n2883_;
  assign new_n4942_ = ~new_n2959_ | ~new_n3396_;
  assign new_n4943_ = ~pi144 | ~new_n2883_;
  assign new_n4944_ = ~new_n2959_ | ~new_n3415_;
  assign new_n4945_ = ~pi145 | ~new_n2883_;
  assign new_n4946_ = ~new_n2959_ | ~new_n3434_;
  assign new_n4947_ = ~pi146 | ~new_n2883_;
  assign new_n4948_ = ~new_n2959_ | ~new_n3453_;
  assign new_n4949_ = ~pi147 | ~new_n2883_;
  assign new_n4950_ = ~new_n2959_ | ~new_n3472_;
  assign new_n4951_ = ~pi148 | ~new_n2883_;
  assign new_n4952_ = ~new_n2959_ | ~new_n3491_;
  assign new_n4953_ = ~pi149 | ~new_n2883_;
  assign new_n4954_ = ~new_n2959_ | ~new_n3510_;
  assign new_n4955_ = ~pi150 | ~new_n2883_;
  assign new_n4956_ = ~new_n2959_ | ~new_n3529_;
  assign new_n4957_ = ~pi151 | ~new_n2883_;
  assign new_n4958_ = ~new_n2959_ | ~new_n3548_;
  assign new_n4959_ = ~pi152 | ~new_n2883_;
  assign new_n4960_ = ~new_n2959_ | ~new_n3567_;
  assign new_n4961_ = ~pi153 | ~new_n2883_;
  assign new_n4962_ = ~new_n2959_ | ~new_n3586_;
  assign new_n4963_ = ~pi154 | ~new_n2883_;
  assign new_n4964_ = ~new_n2959_ | ~new_n3605_;
  assign new_n4965_ = ~pi155 | ~new_n2883_;
  assign new_n4966_ = ~new_n2959_ | ~new_n3624_;
  assign new_n4967_ = ~pi156 | ~new_n2883_;
  assign new_n4968_ = ~new_n2959_ | ~new_n3643_;
  assign new_n4969_ = ~pi157 | ~new_n2883_;
  assign new_n4970_ = ~new_n2959_ | ~new_n3662_;
  assign new_n4971_ = ~pi158 | ~new_n2883_;
  assign new_n4972_ = ~new_n2959_ | ~new_n3682_;
  assign new_n4973_ = ~pi159 | ~new_n2883_;
  assign new_n4974_ = ~new_n2959_ | ~new_n3689_;
  assign new_n4975_ = ~pi160 | ~new_n2883_;
  assign new_n4976_ = ~new_n2959_ | ~new_n3692_;
  assign new_n4977_ = ~pi161 | ~new_n2347_;
  assign new_n4978_ = ~new_n2958_ | ~new_n2303_;
  assign new_n4979_ = ~pi162 | ~new_n2347_;
  assign new_n4980_ = ~new_n2958_ | ~new_n2305_;
  assign new_n4981_ = ~pi163 | ~new_n2347_;
  assign new_n4982_ = ~new_n2958_ | ~new_n2306_;
  assign new_n4983_ = ~pi164 | ~new_n2347_;
  assign new_n4984_ = ~new_n2958_ | ~new_n2307_;
  assign new_n4985_ = ~pi165 | ~new_n2347_;
  assign new_n4986_ = ~new_n2958_ | ~new_n2308_;
  assign new_n4987_ = ~pi166 | ~new_n2347_;
  assign new_n4988_ = ~new_n2958_ | ~new_n2309_;
  assign new_n4989_ = ~pi167 | ~new_n2347_;
  assign new_n4990_ = ~new_n2958_ | ~new_n2310_;
  assign new_n4991_ = ~pi168 | ~new_n2347_;
  assign new_n4992_ = ~new_n2958_ | ~new_n2311_;
  assign new_n4993_ = ~pi169 | ~new_n2347_;
  assign new_n4994_ = ~new_n2958_ | ~new_n2312_;
  assign new_n4995_ = ~pi170 | ~new_n2347_;
  assign new_n4996_ = ~new_n2958_ | ~new_n2313_;
  assign new_n4997_ = ~pi171 | ~new_n2347_;
  assign new_n4998_ = ~new_n2958_ | ~new_n2314_;
  assign new_n4999_ = ~pi172 | ~new_n2347_;
  assign new_n5000_ = ~new_n2958_ | ~new_n2315_;
  assign new_n5001_ = ~pi173 | ~new_n2347_;
  assign new_n5002_ = ~new_n2958_ | ~new_n2316_;
  assign new_n5003_ = ~pi174 | ~new_n2347_;
  assign new_n5004_ = ~new_n2958_ | ~new_n2317_;
  assign new_n5005_ = ~pi175 | ~new_n2347_;
  assign new_n5006_ = ~new_n2958_ | ~new_n2318_;
  assign new_n5007_ = ~pi176 | ~new_n2347_;
  assign new_n5008_ = ~new_n2958_ | ~new_n2319_;
  assign new_n5009_ = ~pi177 | ~new_n2347_;
  assign new_n5010_ = ~new_n2958_ | ~new_n2320_;
  assign new_n5011_ = ~pi178 | ~new_n2347_;
  assign new_n5012_ = ~new_n2958_ | ~new_n2321_;
  assign new_n5013_ = ~pi179 | ~new_n2347_;
  assign new_n5014_ = ~new_n2958_ | ~new_n2322_;
  assign new_n5015_ = ~pi180 | ~new_n2347_;
  assign new_n5016_ = ~new_n2958_ | ~new_n2323_;
  assign new_n5017_ = ~pi181 | ~new_n2347_;
  assign new_n5018_ = ~new_n2958_ | ~new_n2325_;
  assign new_n5019_ = ~pi182 | ~new_n2347_;
  assign new_n5020_ = ~new_n2958_ | ~new_n2327_;
  assign new_n5021_ = ~pi183 | ~new_n2347_;
  assign new_n5022_ = ~new_n2958_ | ~new_n2329_;
  assign new_n5023_ = ~pi184 | ~new_n2347_;
  assign new_n5024_ = ~new_n2958_ | ~new_n2331_;
  assign new_n5025_ = ~pi185 | ~new_n2347_;
  assign new_n5026_ = ~new_n2958_ | ~new_n2333_;
  assign new_n5027_ = ~pi186 | ~new_n2347_;
  assign new_n5028_ = ~new_n2958_ | ~new_n2335_;
  assign new_n5029_ = ~pi187 | ~new_n2347_;
  assign new_n5030_ = ~new_n2958_ | ~new_n2337_;
  assign new_n5031_ = ~pi188 | ~new_n2347_;
  assign new_n5032_ = ~new_n2958_ | ~new_n2339_;
  assign new_n5033_ = ~pi189 | ~new_n2347_;
  assign new_n5034_ = ~new_n2958_ | ~new_n2341_;
  assign new_n5035_ = ~pi190 | ~new_n2347_;
  assign new_n5036_ = ~new_n2958_ | ~new_n2343_;
  assign new_n5037_ = ~pi191 | ~new_n2347_;
  assign new_n5038_ = ~new_n2962_ | ~new_n2958_;
  assign new_n5039_ = ~pi192 | ~new_n2347_;
  assign new_n5040_ = ~new_n2962_ | ~new_n2958_;
  assign new_n5041_ = ~pi213 | ~new_n2357_;
  assign new_n5042_ = ~po266 | ~new_n2004_;
  assign new_n5043_ = ~pi214 | ~new_n2357_;
  assign new_n5044_ = ~po266 | ~new_n2005_;
  assign new_n5045_ = ~pi215 | ~new_n2357_;
  assign new_n5046_ = ~po266 | ~new_n1995_;
  assign new_n5047_ = ~pi216 | ~new_n2357_;
  assign new_n5048_ = ~po266 | ~new_n1991_;
  assign new_n5049_ = ~pi217 | ~new_n2357_;
  assign new_n5050_ = ~po266 | ~new_n1987_;
  assign new_n5051_ = ~pi218 | ~new_n2357_;
  assign new_n5052_ = ~po266 | ~new_n1994_;
  assign new_n5053_ = ~pi219 | ~new_n2357_;
  assign new_n5054_ = ~po266 | ~new_n1998_;
  assign new_n5055_ = ~pi220 | ~new_n2357_;
  assign new_n5056_ = ~po266 | ~new_n1997_;
  assign new_n5057_ = ~pi221 | ~new_n2357_;
  assign new_n5058_ = ~po266 | ~new_n2011_;
  assign new_n5059_ = ~pi222 | ~new_n2357_;
  assign new_n5060_ = ~po266 | ~new_n2010_;
  assign new_n5061_ = ~pi223 | ~new_n2357_;
  assign new_n5062_ = ~po266 | ~new_n1989_;
  assign new_n5063_ = ~pi224 | ~new_n2357_;
  assign new_n5064_ = ~po266 | ~new_n1990_;
  assign new_n5065_ = ~pi225 | ~new_n2357_;
  assign new_n5066_ = ~po266 | ~new_n1999_;
  assign new_n5067_ = ~pi226 | ~new_n2357_;
  assign new_n5068_ = ~po266 | ~new_n2007_;
  assign new_n5069_ = ~pi227 | ~new_n2357_;
  assign new_n5070_ = ~po266 | ~new_n2006_;
  assign new_n5071_ = ~pi228 | ~new_n2357_;
  assign new_n5072_ = ~po266 | ~new_n2001_;
  assign new_n5073_ = ~pi229 | ~new_n2357_;
  assign new_n5074_ = ~po266 | ~new_n2000_;
  assign new_n5075_ = ~pi230 | ~new_n2357_;
  assign new_n5076_ = ~po266 | ~new_n1996_;
  assign new_n5077_ = ~pi231 | ~new_n2357_;
  assign new_n5078_ = ~po266 | ~new_n2009_;
  assign new_n5079_ = ~pi232 | ~new_n2357_;
  assign new_n5080_ = ~po266 | ~new_n2008_;
  assign new_n5081_ = ~pi233 | ~new_n2357_;
  assign new_n5082_ = ~po266 | ~new_n2003_;
  assign new_n5083_ = ~pi234 | ~new_n2357_;
  assign new_n5084_ = ~po266 | ~new_n2002_;
  assign new_n5085_ = ~pi235 | ~new_n2357_;
  assign new_n5086_ = ~po266 | ~new_n1988_;
  assign new_n5087_ = ~pi236 | ~new_n2357_;
  assign new_n5088_ = ~po266 | ~new_n1993_;
  assign new_n5089_ = ~pi237 | ~new_n2357_;
  assign new_n5090_ = ~po266 | ~new_n1992_;
  assign new_n5091_ = ~pi238 | ~new_n2357_;
  assign new_n5092_ = ~po266 | ~new_n1985_;
  assign new_n5093_ = ~pi239 | ~new_n2357_;
  assign new_n5094_ = ~po266 | ~new_n1984_;
  assign new_n5095_ = ~pi240 | ~new_n2357_;
  assign new_n5096_ = ~po266 | ~new_n1980_;
  assign new_n5097_ = ~pi241 | ~new_n2357_;
  assign new_n5098_ = ~po266 | ~new_n1981_;
  assign new_n5099_ = ~pi242 | ~new_n2357_;
  assign new_n5100_ = ~po266 | ~new_n1982_;
  assign new_n5101_ = ~pi243 | ~new_n2357_;
  assign new_n5102_ = ~po266 | ~new_n1986_;
  assign new_n5103_ = ~pi244 | ~new_n2357_;
  assign new_n5104_ = ~po266 | ~new_n1983_;
  assign new_n5105_ = ~new_n2359_ | ~new_n2377_ | ~new_n4720_;
  assign new_n5106_ = ~new_n15169_ | ~new_n2957_;
  assign new_n5107_ = ~new_n2944_ | ~new_n1981_;
  assign new_n5108_ = ~new_n2340_ | ~new_n3629_;
  assign new_n5109_ = ~new_n5108_ | ~new_n5107_;
  assign new_n5110_ = ~new_n2953_ | ~new_n1983_;
  assign new_n5111_ = ~new_n2345_ | ~new_n3686_;
  assign new_n5112_ = ~new_n5111_ | ~new_n5110_;
  assign new_n5113_ = ~new_n2952_ | ~new_n2003_;
  assign new_n5114_ = ~new_n2324_ | ~new_n3477_;
  assign new_n5115_ = ~new_n5114_ | ~new_n5113_;
  assign new_n5116_ = ~new_n2954_ | ~new_n1986_;
  assign new_n5117_ = ~new_n2344_ | ~new_n3666_;
  assign new_n5118_ = ~new_n5117_ | ~new_n5116_;
  assign new_n5119_ = ~new_n4886_ | ~new_n3458_;
  assign new_n5120_ = ~new_n2441_ | ~new_n2008_;
  assign new_n5121_ = ~new_n5120_ | ~new_n5119_;
  assign new_n5122_ = ~new_n4832_ | ~new_n3306_;
  assign new_n5123_ = ~new_n2418_ | ~new_n1990_;
  assign new_n5124_ = ~new_n5123_ | ~new_n5122_;
  assign new_n5125_ = ~new_n4783_ | ~new_n3173_;
  assign new_n5126_ = ~new_n2397_ | ~new_n1987_;
  assign new_n5127_ = ~new_n5126_ | ~new_n5125_;
  assign new_n5128_ = ~new_n4825_ | ~new_n3287_;
  assign new_n5129_ = ~new_n2415_ | ~new_n1989_;
  assign new_n5130_ = ~new_n5129_ | ~new_n5128_;
  assign new_n5131_ = ~new_n2955_ | ~new_n1982_;
  assign new_n5132_ = ~new_n2342_ | ~new_n3648_;
  assign new_n5133_ = ~new_n5132_ | ~new_n5131_;
  assign new_n5134_ = ~new_n2945_ | ~new_n1980_;
  assign new_n5135_ = ~new_n2338_ | ~new_n3610_;
  assign new_n5136_ = ~new_n5135_ | ~new_n5134_;
  assign new_n5137_ = ~new_n4874_ | ~new_n3420_;
  assign new_n5138_ = ~new_n2436_ | ~new_n1996_;
  assign new_n5139_ = ~new_n5138_ | ~new_n5137_;
  assign new_n5140_ = ~new_n4811_ | ~new_n3249_;
  assign new_n5141_ = ~new_n2409_ | ~new_n2011_;
  assign new_n5142_ = ~new_n5141_ | ~new_n5140_;
  assign new_n5143_ = ~new_n4818_ | ~new_n3268_;
  assign new_n5144_ = ~new_n2412_ | ~new_n2010_;
  assign new_n5145_ = ~new_n5144_ | ~new_n5143_;
  assign new_n5146_ = ~new_n4846_ | ~new_n3344_;
  assign new_n5147_ = ~new_n2424_ | ~new_n2007_;
  assign new_n5148_ = ~new_n5147_ | ~new_n5146_;
  assign new_n5149_ = ~new_n4853_ | ~new_n3363_;
  assign new_n5150_ = ~new_n2427_ | ~new_n2006_;
  assign new_n5151_ = ~new_n5150_ | ~new_n5149_;
  assign new_n5152_ = ~new_n4747_ | ~new_n3135_;
  assign new_n5153_ = ~new_n2383_ | ~new_n2004_;
  assign new_n5154_ = ~new_n5153_ | ~new_n5152_;
  assign new_n5155_ = ~new_n4762_ | ~new_n3111_;
  assign new_n5156_ = ~new_n2388_ | ~new_n2005_;
  assign new_n5157_ = ~new_n5156_ | ~new_n5155_;
  assign new_n5158_ = ~new_n4860_ | ~new_n3382_;
  assign new_n5159_ = ~new_n2430_ | ~new_n2001_;
  assign new_n5160_ = ~new_n5159_ | ~new_n5158_;
  assign new_n5161_ = ~new_n4867_ | ~new_n3401_;
  assign new_n5162_ = ~new_n2433_ | ~new_n2000_;
  assign new_n5163_ = ~new_n5162_ | ~new_n5161_;
  assign new_n5164_ = ~new_n4797_ | ~new_n3211_;
  assign new_n5165_ = ~new_n2403_ | ~new_n1998_;
  assign new_n5166_ = ~new_n5165_ | ~new_n5164_;
  assign new_n5167_ = ~new_n4804_ | ~new_n3230_;
  assign new_n5168_ = ~new_n2406_ | ~new_n1997_;
  assign new_n5169_ = ~new_n5168_ | ~new_n5167_;
  assign new_n5170_ = ~new_n4839_ | ~new_n3325_;
  assign new_n5171_ = ~new_n2421_ | ~new_n1999_;
  assign new_n5172_ = ~new_n5171_ | ~new_n5170_;
  assign new_n5173_ = ~new_n4769_ | ~new_n3130_;
  assign new_n5174_ = ~new_n2391_ | ~new_n1995_;
  assign new_n5175_ = ~new_n5174_ | ~new_n5173_;
  assign new_n5176_ = ~new_n4776_ | ~new_n3154_;
  assign new_n5177_ = ~new_n2394_ | ~new_n1991_;
  assign new_n5178_ = ~new_n5177_ | ~new_n5176_;
  assign new_n5179_ = ~new_n4790_ | ~new_n3192_;
  assign new_n5180_ = ~new_n2400_ | ~new_n1994_;
  assign new_n5181_ = ~new_n5180_ | ~new_n5179_;
  assign new_n5182_ = ~new_n4881_ | ~new_n3439_;
  assign new_n5183_ = ~new_n2439_ | ~new_n2009_;
  assign new_n5184_ = ~new_n5183_ | ~new_n5182_;
  assign new_n5185_ = ~new_n2948_ | ~new_n1992_;
  assign new_n5186_ = ~new_n2332_ | ~new_n3553_;
  assign new_n5187_ = ~new_n5186_ | ~new_n5185_;
  assign new_n5188_ = ~new_n2949_ | ~new_n1993_;
  assign new_n5189_ = ~new_n2330_ | ~new_n3534_;
  assign new_n5190_ = ~new_n5189_ | ~new_n5188_;
  assign new_n5191_ = ~new_n2951_ | ~new_n2002_;
  assign new_n5192_ = ~new_n2326_ | ~new_n3496_;
  assign new_n5193_ = ~new_n5192_ | ~new_n5191_;
  assign new_n5194_ = ~new_n2950_ | ~new_n1988_;
  assign new_n5195_ = ~new_n2328_ | ~new_n3515_;
  assign new_n5196_ = ~new_n5195_ | ~new_n5194_;
  assign new_n5197_ = ~new_n2947_ | ~new_n1985_;
  assign new_n5198_ = ~new_n2334_ | ~new_n3572_;
  assign new_n5199_ = ~new_n5198_ | ~new_n5197_;
  assign new_n5200_ = ~new_n2946_ | ~new_n1984_;
  assign new_n5201_ = ~new_n2336_ | ~new_n3591_;
  assign new_n5202_ = ~new_n5201_ | ~new_n5200_;
  assign new_n5203_ = ~new_n2968_ | ~new_n2918_;
  assign new_n5204_ = ~new_n4056_ | ~new_n1976_;
  assign new_n5205_ = ~new_n4726_ | ~new_n4060_ | ~new_n2359_;
  assign new_n5206_ = ~new_n2380_ | ~new_n4057_;
  assign new_n5207_ = ~new_n4713_ | ~new_n2358_;
  assign new_n5208_ = ~new_n2378_ | ~new_n2371_;
  assign new_n5209_ = ~new_n2377_ | ~new_n4071_;
  assign new_n5210_ = ~new_n4729_ | ~new_n2921_;
  assign new_n5211_ = ~new_n2381_ | ~new_n4335_;
  assign new_n5212_ = ~new_n4741_ | ~new_n1942_ | ~pi161;
  assign new_n5213_ = ~new_n8457_ | ~new_n30327_;
  assign new_n5214_ = ~new_n30512_ | ~new_n5216_;
  assign new_n5215_ = ~new_n30423_ | ~new_n30424_;
  assign new_n5216_ = ~new_n5217_ | ~new_n5218_;
  assign new_n5217_ = ~new_n8809_ | ~new_n30330_;
  assign new_n5218_ = ~new_n8456_ | ~new_n30329_;
  assign new_n5219_ = ~new_n8809_ | ~new_n30330_;
  assign new_n5220_ = ~new_n8456_ | ~new_n30329_;
  assign new_n5221_ = ~new_n30516_ | ~new_n5223_;
  assign new_n5222_ = ~new_n30421_ | ~new_n30422_;
  assign new_n5223_ = ~new_n5224_ | ~new_n5225_;
  assign new_n5224_ = ~new_n8812_ | ~new_n30332_;
  assign new_n5225_ = ~new_n8451_ | ~new_n30331_;
  assign new_n5226_ = ~new_n8812_ | ~new_n30332_;
  assign new_n5227_ = ~new_n8451_ | ~new_n30331_;
  assign new_n5228_ = ~new_n5230_ | ~new_n30520_;
  assign new_n5229_ = ~new_n30619_ | ~new_n30350_;
  assign new_n5230_ = ~new_n5231_ | ~new_n5232_;
  assign new_n5231_ = ~new_n8815_ | ~new_n30315_;
  assign new_n5232_ = ~new_n8450_ | ~new_n30314_;
  assign new_n5233_ = ~new_n8818_ | ~new_n30316_;
  assign new_n5234_ = new_n6144_ & new_n7891_;
  assign new_n5235_ = new_n6157_ & new_n5639_;
  assign new_n5236_ = new_n5795_ & new_n5790_;
  assign new_n5237_ = new_n7908_ & new_n5643_;
  assign new_n5238_ = new_n5646_ & new_n5643_;
  assign new_n5239_ = new_n5641_ & new_n5642_;
  assign new_n5240_ = new_n7900_ & new_n5641_;
  assign new_n5241_ = new_n7897_ & new_n5642_;
  assign new_n5242_ = new_n7897_ & new_n7900_;
  assign new_n5243_ = new_n5268_ & pi520;
  assign new_n5244_ = new_n5977_ & new_n5621_;
  assign new_n5245_ = new_n6196_ & new_n7891_;
  assign new_n5246_ = new_n6183_ & new_n7903_;
  assign new_n5247_ = new_n6164_ & new_n7891_;
  assign new_n5248_ = new_n6023_ & new_n6166_;
  assign new_n5249_ = new_n19210_ & new_n5631_;
  assign new_n5250_ = new_n5549_ & pi520;
  assign new_n5251_ = new_n6152_ & new_n6184_;
  assign new_n5252_ = new_n6184_ & new_n5618_;
  assign new_n5253_ = new_n6153_ & new_n6184_;
  assign new_n5254_ = new_n6158_ & new_n6184_;
  assign new_n5255_ = new_n6183_ & new_n5643_;
  assign new_n5256_ = new_n6166_ & new_n7903_;
  assign new_n5257_ = new_n6184_ & new_n5246_;
  assign new_n5258_ = new_n6166_ & new_n5643_;
  assign new_n5259_ = new_n7908_ & new_n7074_;
  assign new_n5260_ = new_n5244_ & new_n7908_;
  assign new_n5261_ = new_n7903_ & new_n7074_;
  assign new_n5262_ = new_n5244_ & new_n7903_;
  assign new_n5263_ = new_n5238_ & new_n7074_;
  assign new_n5264_ = new_n5244_ & new_n5238_;
  assign new_n5265_ = new_n5243_ & new_n5621_;
  assign new_n5266_ = new_n7404_ & pi520;
  assign new_n5267_ = new_n5243_ & new_n7406_;
  assign new_n5268_ = new_n7878_ & new_n5616_;
  assign new_n5269_ = new_n5638_ & new_n7888_;
  assign new_n5270_ = new_n5796_ & new_n5236_;
  assign new_n5271_ = new_n5561_ & new_n5557_ & new_n5558_ & new_n5612_ & new_n5622_;
  assign new_n5272_ = new_n5619_ & pi520;
  assign new_n5273_ = new_n6039_ & new_n6040_ & new_n7659_;
  assign new_n5274_ = new_n7681_ & new_n7680_;
  assign new_n5275_ = ~new_n6832_ | ~new_n6833_ | ~new_n6830_ | ~new_n6831_;
  assign new_n5276_ = ~new_n6851_ | ~new_n6852_ | ~new_n6849_ | ~new_n6850_;
  assign new_n5277_ = ~new_n6870_ | ~new_n6868_ | ~new_n6869_ | ~new_n6871_;
  assign new_n5278_ = ~new_n6907_ | ~new_n6908_ | ~new_n6909_;
  assign new_n5279_ = ~new_n6813_ | ~new_n6814_ | ~new_n6811_ | ~new_n6812_;
  assign new_n5280_ = ~new_n6794_ | ~new_n6795_ | ~new_n6792_ | ~new_n6793_;
  assign new_n5281_ = ~new_n6887_ | ~new_n6888_ | ~new_n6889_;
  assign new_n5282_ = ~new_n6395_ | ~new_n6393_ | ~new_n6394_ | ~new_n6396_;
  assign new_n5283_ = ~new_n6737_ | ~new_n6738_ | ~new_n6735_ | ~new_n6736_;
  assign new_n5284_ = ~new_n6509_ | ~new_n6507_ | ~new_n6508_ | ~new_n6510_;
  assign new_n5285_ = ~new_n6528_ | ~new_n6526_ | ~new_n6527_ | ~new_n6529_;
  assign new_n5286_ = ~new_n6376_ | ~new_n6374_ | ~new_n6375_ | ~new_n6377_;
  assign new_n5287_ = ~new_n6775_ | ~new_n6776_ | ~new_n6773_ | ~new_n6774_;
  assign new_n5288_ = ~new_n6756_ | ~new_n6757_ | ~new_n6754_ | ~new_n6755_;
  assign new_n5289_ = ~new_n6414_ | ~new_n6412_ | ~new_n6413_ | ~new_n6415_;
  assign new_n5290_ = ~new_n6352_ | ~new_n6350_ | ~new_n6351_ | ~new_n6353_;
  assign new_n5291_ = ~new_n6642_ | ~new_n6643_ | ~new_n6640_ | ~new_n6641_;
  assign new_n5292_ = ~new_n6452_ | ~new_n6450_ | ~new_n6451_ | ~new_n6453_;
  assign new_n5293_ = ~new_n6433_ | ~new_n6431_ | ~new_n6432_ | ~new_n6434_;
  assign new_n5294_ = ~new_n6547_ | ~new_n6545_ | ~new_n6546_ | ~new_n6548_;
  assign new_n5295_ = ~new_n6623_ | ~new_n6621_ | ~new_n6622_ | ~new_n6624_;
  assign new_n5296_ = ~new_n6604_ | ~new_n6602_ | ~new_n6603_ | ~new_n6605_;
  assign new_n5297_ = ~new_n6718_ | ~new_n6719_ | ~new_n6716_ | ~new_n6717_;
  assign new_n5298_ = ~new_n6699_ | ~new_n6700_ | ~new_n6697_ | ~new_n6698_;
  assign new_n5299_ = ~new_n6357_ | ~new_n6355_ | ~new_n6356_ | ~new_n6358_;
  assign new_n5300_ = ~new_n6333_ | ~new_n6331_ | ~new_n6332_ | ~new_n6334_;
  assign new_n5301_ = ~new_n6585_ | ~new_n6583_ | ~new_n6584_ | ~new_n6586_;
  assign new_n5302_ = ~new_n6566_ | ~new_n6564_ | ~new_n6565_ | ~new_n6567_;
  assign new_n5303_ = ~new_n6680_ | ~new_n6681_ | ~new_n6678_ | ~new_n6679_;
  assign new_n5304_ = ~new_n6661_ | ~new_n6662_ | ~new_n6659_ | ~new_n6660_;
  assign new_n5305_ = ~new_n6490_ | ~new_n6488_ | ~new_n6489_ | ~new_n6491_;
  assign new_n5306_ = ~new_n6471_ | ~new_n6469_ | ~new_n6470_ | ~new_n6472_;
  assign po510 = ~new_n6035_ | ~new_n7654_;
  assign po509 = ~pi520;
  assign new_n5309_ = ~new_n7777_ | ~new_n7776_;
  assign new_n5310_ = ~new_n7779_ | ~new_n7778_;
  assign new_n5311_ = ~new_n6079_ | ~new_n7783_;
  assign new_n5312_ = ~new_n6080_ | ~new_n7786_;
  assign new_n5313_ = ~new_n6081_ | ~new_n7789_;
  assign new_n5314_ = ~new_n6082_ | ~new_n7792_;
  assign new_n5315_ = ~new_n6083_ | ~new_n7795_;
  assign new_n5316_ = ~new_n6084_ | ~new_n7798_;
  assign new_n5317_ = ~new_n6085_ | ~new_n7801_;
  assign new_n5318_ = ~new_n6086_ | ~new_n7804_;
  assign new_n5319_ = ~new_n6087_ | ~new_n7807_;
  assign new_n5320_ = ~new_n6088_ | ~new_n7810_;
  assign new_n5321_ = ~new_n6089_ | ~new_n7816_;
  assign new_n5322_ = ~new_n6090_ | ~new_n7819_;
  assign new_n5323_ = ~new_n6091_ | ~new_n7822_;
  assign new_n5324_ = ~new_n6092_ | ~new_n7825_;
  assign new_n5325_ = ~new_n6093_ | ~new_n7828_;
  assign new_n5326_ = ~new_n6094_ | ~new_n7831_;
  assign new_n5327_ = ~new_n6095_ | ~new_n7834_;
  assign new_n5328_ = ~new_n6096_ | ~new_n7837_;
  assign new_n5329_ = ~new_n6097_ | ~new_n7840_;
  assign new_n5330_ = ~new_n6098_ | ~new_n7843_;
  assign new_n5331_ = ~new_n6077_ | ~new_n7758_;
  assign new_n5332_ = ~new_n6078_ | ~new_n7761_;
  assign new_n5333_ = ~new_n7766_ | ~new_n7765_ | ~new_n7764_;
  assign new_n5334_ = ~new_n7769_ | ~new_n7768_ | ~new_n7767_;
  assign new_n5335_ = ~new_n7772_ | ~new_n7771_ | ~new_n7770_;
  assign new_n5336_ = ~new_n7775_ | ~new_n7774_ | ~new_n7773_;
  assign new_n5337_ = ~new_n7782_ | ~new_n7781_ | ~new_n7780_;
  assign new_n5338_ = ~new_n7815_ | ~new_n7814_ | ~new_n7813_;
  assign new_n5339_ = ~new_n7848_ | ~new_n7847_ | ~new_n7846_;
  assign new_n5340_ = ~new_n7850_ | ~new_n7849_;
  assign new_n5341_ = new_n7858_ & new_n7857_ & new_n7852_;
  assign new_n5342_ = ~new_n7684_ | ~new_n7683_ | ~new_n7682_;
  assign new_n5343_ = ~new_n7690_ | ~new_n7689_ | ~new_n6051_;
  assign new_n5344_ = ~new_n7693_ | ~new_n7692_ | ~new_n6052_;
  assign new_n5345_ = ~new_n7696_ | ~new_n7695_ | ~new_n6053_;
  assign new_n5346_ = ~new_n7699_ | ~new_n7698_ | ~new_n6054_;
  assign new_n5347_ = ~new_n7702_ | ~new_n7701_ | ~new_n6055_;
  assign new_n5348_ = ~new_n7705_ | ~new_n7704_ | ~new_n6056_;
  assign new_n5349_ = ~new_n7708_ | ~new_n7707_ | ~new_n6057_;
  assign new_n5350_ = ~new_n7711_ | ~new_n7710_ | ~new_n6058_;
  assign new_n5351_ = ~new_n7714_ | ~new_n7713_ | ~new_n6059_;
  assign new_n5352_ = ~new_n7717_ | ~new_n7716_ | ~new_n6060_;
  assign new_n5353_ = ~new_n7723_ | ~new_n7722_ | ~new_n6063_;
  assign new_n5354_ = ~new_n7726_ | ~new_n7725_ | ~new_n6064_;
  assign new_n5355_ = ~new_n7729_ | ~new_n7728_ | ~new_n6065_;
  assign new_n5356_ = ~new_n7732_ | ~new_n7731_ | ~new_n6066_;
  assign new_n5357_ = ~new_n7735_ | ~new_n7734_ | ~new_n6067_;
  assign new_n5358_ = ~new_n7738_ | ~new_n7737_ | ~new_n6068_;
  assign new_n5359_ = ~new_n7741_ | ~new_n7740_ | ~new_n6069_;
  assign new_n5360_ = ~new_n7744_ | ~new_n7743_ | ~new_n6070_;
  assign new_n5361_ = ~new_n6071_ | ~new_n7746_ | ~new_n7745_;
  assign new_n5362_ = ~new_n6072_ | ~new_n7749_ | ~new_n7748_;
  assign new_n5363_ = ~new_n6041_ | ~new_n7663_ | ~new_n7662_;
  assign new_n5364_ = ~new_n6042_ | ~new_n7666_ | ~new_n7665_;
  assign new_n5365_ = ~new_n6043_ | ~new_n7669_ | ~new_n7668_;
  assign new_n5366_ = ~new_n6044_ | ~new_n7672_ | ~new_n7671_;
  assign new_n5367_ = ~new_n6045_ | ~new_n7675_ | ~new_n7674_;
  assign new_n5368_ = ~new_n7678_ | ~new_n6046_;
  assign new_n5369_ = ~new_n7686_ | ~new_n6049_;
  assign new_n5370_ = ~new_n7719_ | ~new_n6061_;
  assign new_n5371_ = ~new_n7752_ | ~new_n6073_;
  assign new_n5372_ = ~new_n7755_ | ~new_n6075_;
  assign new_n5373_ = ~new_n5635_ | ~new_n6037_ | ~new_n5565_;
  assign new_n5374_ = ~new_n5235_ | ~new_n7878_;
  assign new_n5375_ = new_n7657_ & new_n5276_;
  assign new_n5376_ = new_n7657_ & new_n5275_;
  assign new_n5377_ = new_n7657_ & new_n5279_;
  assign new_n5378_ = new_n7657_ & new_n5280_;
  assign new_n5379_ = new_n7657_ & new_n5287_;
  assign new_n5380_ = new_n7657_ & new_n5288_;
  assign new_n5381_ = new_n7657_ & new_n5283_;
  assign new_n5382_ = new_n7657_ & new_n5297_;
  assign new_n5383_ = new_n7657_ & new_n5298_;
  assign new_n5384_ = new_n7657_ & new_n5303_;
  assign new_n5385_ = new_n7657_ & new_n5304_;
  assign new_n5386_ = new_n7657_ & new_n5291_;
  assign new_n5387_ = new_n7657_ & new_n5295_;
  assign new_n5388_ = new_n7657_ & new_n5296_;
  assign new_n5389_ = new_n7657_ & new_n5301_;
  assign new_n5390_ = new_n7657_ & new_n5302_;
  assign new_n5391_ = new_n7657_ & new_n5294_;
  assign new_n5392_ = new_n7657_ & new_n5285_;
  assign new_n5393_ = new_n7657_ & new_n5284_;
  assign new_n5394_ = new_n7657_ & new_n5305_;
  assign new_n5395_ = new_n7657_ & new_n5306_;
  assign new_n5396_ = new_n7657_ & new_n5292_;
  assign new_n5397_ = new_n7657_ & new_n5293_;
  assign new_n5398_ = new_n7657_ & new_n5289_;
  assign new_n5399_ = new_n7657_ & new_n5282_;
  assign new_n5400_ = new_n7657_ & new_n5286_;
  assign new_n5401_ = new_n7657_ & new_n5290_;
  assign new_n5402_ = new_n7657_ & new_n5300_;
  assign new_n5403_ = new_n7657_ & new_n5299_;
  assign new_n5404_ = ~new_n5563_ | ~new_n5624_ | ~new_n7656_;
  assign po508 = ~new_n7652_ | ~new_n7650_ | ~new_n6034_ | ~new_n7653_;
  assign po507 = ~new_n7644_ | ~new_n7642_ | ~new_n7640_ | ~new_n7641_ | ~new_n7643_;
  assign po506 = ~new_n7632_ | ~new_n7633_ | ~new_n7634_ | ~new_n7635_ | ~new_n7631_;
  assign po505 = ~new_n7626_ | ~new_n7624_ | ~new_n7622_ | ~new_n7623_ | ~new_n7625_;
  assign po504 = ~new_n7614_ | ~new_n7616_ | ~new_n7617_ | ~new_n7615_ | ~new_n7613_;
  assign po503 = ~new_n7607_ | ~new_n7605_ | ~new_n6033_ | ~new_n7608_;
  assign po502 = ~new_n7596_ | ~new_n7597_ | ~new_n7598_ | ~new_n7599_ | ~new_n7595_;
  assign po501 = ~new_n7590_ | ~new_n7588_ | ~new_n7586_ | ~new_n7587_ | ~new_n7589_;
  assign po500 = ~new_n7580_ | ~new_n7578_ | ~new_n6032_ | ~new_n7581_;
  assign po499 = ~new_n7571_ | ~new_n7569_ | ~new_n6031_ | ~new_n7572_;
  assign po498 = ~new_n7560_ | ~new_n7561_ | ~new_n7562_ | ~new_n7563_ | ~new_n7559_;
  assign po497 = ~new_n7551_ | ~new_n7552_ | ~new_n7553_ | ~new_n7554_ | ~new_n7550_;
  assign po496 = ~new_n7545_ | ~new_n7543_ | ~new_n7541_ | ~new_n7542_ | ~new_n7544_;
  assign po495 = ~new_n7533_ | ~new_n7534_ | ~new_n7535_ | ~new_n7536_ | ~new_n7532_;
  assign po494 = ~new_n7526_ | ~new_n7524_ | ~new_n6030_ | ~new_n7527_;
  assign po493 = ~new_n7515_ | ~new_n7516_ | ~new_n7517_ | ~new_n7518_ | ~new_n7514_;
  assign po492 = ~new_n7509_ | ~new_n7507_ | ~new_n7505_ | ~new_n7506_ | ~new_n7508_;
  assign po491 = ~new_n7499_ | ~new_n7497_ | ~new_n6029_ | ~new_n7500_;
  assign po490 = ~new_n7488_ | ~new_n7490_ | ~new_n7491_ | ~new_n7489_ | ~new_n7487_;
  assign po489 = ~new_n6027_ | ~new_n6028_ | ~new_n7480_;
  assign po488 = ~new_n7471_ | ~new_n7472_ | ~new_n7473_ | ~new_n7474_ | ~new_n7470_;
  assign po487 = ~new_n7462_ | ~new_n7463_ | ~new_n7464_ | ~new_n7465_ | ~new_n7461_;
  assign po486 = ~new_n7456_ | ~new_n7454_ | ~new_n7452_ | ~new_n7453_ | ~new_n7455_;
  assign po485 = ~new_n7444_ | ~new_n7446_ | ~new_n7447_ | ~new_n7445_ | ~new_n7443_;
  assign po484 = ~new_n7437_ | ~new_n7435_ | ~new_n6025_ | ~new_n7438_;
  assign po483 = ~new_n7426_ | ~new_n7427_ | ~new_n7428_ | ~new_n7429_ | ~new_n7425_;
  assign po482 = ~new_n7419_ | ~new_n7417_ | ~new_n6024_ | ~new_n7420_;
  assign po481 = ~new_n7411_ | ~new_n7409_ | ~new_n7407_ | ~new_n7408_ | ~new_n7410_;
  assign po480 = ~new_n7395_ | ~new_n7396_ | ~new_n7397_ | ~new_n7398_ | ~new_n7394_;
  assign po446 = ~new_n7369_ | ~new_n6006_ | ~new_n6005_ | ~new_n7370_;
  assign po445 = ~new_n7354_ | ~new_n6004_ | ~new_n6003_ | ~new_n7355_;
  assign po444 = ~new_n7339_ | ~new_n6002_ | ~new_n6001_ | ~new_n7340_;
  assign po443 = ~new_n7324_ | ~new_n6000_ | ~new_n5999_ | ~new_n7325_;
  assign po442 = ~new_n7309_ | ~new_n5998_ | ~new_n5997_ | ~new_n7310_;
  assign po441 = ~new_n7294_ | ~new_n5996_ | ~new_n5995_ | ~new_n7295_;
  assign po440 = ~new_n7279_ | ~new_n5994_ | ~new_n5993_ | ~new_n7280_;
  assign po439 = ~new_n7264_ | ~new_n5992_ | ~new_n5991_ | ~new_n7265_;
  assign po438 = ~new_n7249_ | ~new_n5990_ | ~new_n5989_ | ~new_n7250_;
  assign po437 = ~new_n5988_ | ~new_n7235_ | ~new_n7234_;
  assign po436 = ~new_n5987_ | ~new_n7220_ | ~new_n7219_;
  assign po435 = ~new_n5986_ | ~new_n7205_ | ~new_n7204_;
  assign po434 = ~new_n5985_ | ~new_n7190_ | ~new_n7189_;
  assign po433 = ~new_n5984_ | ~new_n7175_ | ~new_n7174_;
  assign po432 = ~new_n5983_ | ~new_n7160_ | ~new_n7159_;
  assign po431 = ~new_n5982_ | ~new_n7145_ | ~new_n7144_;
  assign po430 = ~new_n5981_ | ~new_n7130_ | ~new_n7129_;
  assign po429 = ~new_n5980_ | ~new_n7115_ | ~new_n7114_;
  assign po428 = ~new_n5979_ | ~new_n7100_ | ~new_n7099_;
  assign po427 = ~new_n5978_ | ~new_n7085_ | ~new_n7084_;
  assign po426 = ~new_n7073_ | ~new_n6135_ | ~new_n7072_;
  assign po425 = ~new_n7071_ | ~new_n6134_ | ~new_n7070_;
  assign po424 = ~new_n7067_ | ~new_n6132_ | ~new_n7066_ | ~new_n7069_ | ~new_n7068_;
  assign po423 = ~new_n5974_ | ~new_n6131_ | ~new_n7062_ | ~new_n5973_;
  assign po422 = ~new_n5972_ | ~new_n6130_ | ~new_n7057_ | ~new_n5971_;
  assign po421 = ~new_n5970_ | ~new_n6129_ | ~new_n7052_ | ~new_n5969_;
  assign po420 = ~new_n5968_ | ~new_n6128_ | ~new_n7047_ | ~new_n5967_;
  assign po419 = ~new_n5966_ | ~new_n6127_ | ~new_n7042_ | ~new_n5965_;
  assign po418 = ~new_n5964_ | ~new_n6126_ | ~new_n7037_ | ~new_n5963_;
  assign po417 = ~new_n5962_ | ~new_n6125_ | ~new_n7032_ | ~new_n5961_;
  assign po416 = ~new_n5960_ | ~new_n6124_ | ~new_n7027_ | ~new_n5959_;
  assign po415 = ~new_n5958_ | ~new_n6123_ | ~new_n7022_ | ~new_n5957_;
  assign po414 = ~new_n5956_ | ~new_n6122_ | ~new_n7017_ | ~new_n5955_;
  assign po413 = ~new_n5954_ | ~new_n6121_ | ~new_n7012_ | ~new_n5953_;
  assign po412 = ~new_n5952_ | ~new_n6120_ | ~new_n7007_ | ~new_n5951_;
  assign po411 = ~new_n5950_ | ~new_n6119_ | ~new_n7002_ | ~new_n5949_;
  assign po410 = ~new_n6118_ | ~new_n5948_ | ~new_n5947_;
  assign po409 = ~new_n6117_ | ~new_n5946_ | ~new_n5945_;
  assign po408 = ~new_n6116_ | ~new_n5944_ | ~new_n5943_;
  assign po407 = ~new_n6115_ | ~new_n5942_ | ~new_n5941_;
  assign po406 = ~new_n6114_ | ~new_n5940_ | ~new_n5939_;
  assign po405 = ~new_n6113_ | ~new_n5938_ | ~new_n5937_;
  assign po404 = ~new_n5936_ | ~new_n5935_;
  assign po403 = ~new_n5934_ | ~new_n5933_;
  assign po402 = ~new_n5932_ | ~new_n5931_;
  assign po401 = ~new_n5930_ | ~new_n5929_;
  assign po400 = ~new_n5928_ | ~new_n5927_;
  assign po399 = ~new_n5926_ | ~new_n5925_;
  assign po398 = ~new_n5924_ | ~new_n5923_;
  assign po397 = ~new_n5922_ | ~new_n5921_;
  assign po396 = ~new_n5920_ | ~new_n5919_;
  assign po395 = ~new_n5918_ | ~new_n5917_;
  assign po330 = pi341 & new_n6100_;
  assign po329 = pi340 & new_n6100_;
  assign po328 = pi339 & new_n6100_;
  assign po327 = pi338 & new_n6100_;
  assign po326 = pi337 & new_n6100_;
  assign po325 = pi336 & new_n6100_;
  assign po324 = pi335 & new_n6100_;
  assign po323 = pi334 & new_n6100_;
  assign po322 = pi333 & new_n6100_;
  assign po321 = pi332 & new_n6100_;
  assign po320 = pi331 & new_n6100_;
  assign po319 = pi330 & new_n6100_;
  assign po318 = pi329 & new_n6100_;
  assign po317 = pi328 & new_n6100_;
  assign po316 = pi327 & new_n6100_;
  assign po315 = pi326 & new_n6100_;
  assign po314 = pi325 & new_n6100_;
  assign po313 = pi324 & new_n6100_;
  assign po312 = pi323 & new_n6100_;
  assign po311 = pi322 & new_n6100_;
  assign po310 = pi321 & new_n6100_;
  assign po309 = pi320 & new_n6100_;
  assign po308 = pi319 & new_n6100_;
  assign po307 = pi318 & new_n6100_;
  assign po306 = pi317 & new_n6100_;
  assign po305 = pi316 & new_n6100_;
  assign po304 = pi315 & new_n6100_;
  assign po303 = pi314 & new_n6100_;
  assign po302 = pi313 & new_n6100_;
  assign po301 = pi312 & new_n6100_;
  assign po298 = ~new_n6292_ | ~new_n6293_ | ~new_n6294_;
  assign po297 = ~new_n6289_ | ~new_n6290_ | ~new_n6291_;
  assign po296 = ~new_n6286_ | ~new_n6287_ | ~new_n6288_;
  assign po295 = ~new_n6283_ | ~new_n6284_ | ~new_n6285_;
  assign po294 = ~new_n6280_ | ~new_n6281_ | ~new_n6282_;
  assign po293 = ~new_n6277_ | ~new_n6278_ | ~new_n6279_;
  assign po292 = ~new_n6274_ | ~new_n6275_ | ~new_n6276_;
  assign po291 = ~new_n6271_ | ~new_n6272_ | ~new_n6273_;
  assign po290 = ~new_n6268_ | ~new_n6269_ | ~new_n6270_;
  assign po289 = ~new_n6265_ | ~new_n6266_ | ~new_n6267_;
  assign po288 = ~new_n6262_ | ~new_n6263_ | ~new_n6264_;
  assign po287 = ~new_n6259_ | ~new_n6260_ | ~new_n6261_;
  assign po286 = ~new_n6256_ | ~new_n6257_ | ~new_n6258_;
  assign po285 = ~new_n6253_ | ~new_n6254_ | ~new_n6255_;
  assign po284 = ~new_n6250_ | ~new_n6251_ | ~new_n6252_;
  assign po283 = ~new_n6247_ | ~new_n6248_ | ~new_n6249_;
  assign po282 = ~new_n6244_ | ~new_n6245_ | ~new_n6246_;
  assign po281 = ~new_n6241_ | ~new_n6242_ | ~new_n6243_;
  assign po280 = ~new_n6238_ | ~new_n6239_ | ~new_n6240_;
  assign po279 = ~new_n6235_ | ~new_n6236_ | ~new_n6237_;
  assign po278 = ~new_n6232_ | ~new_n6233_ | ~new_n6234_;
  assign po277 = ~new_n6229_ | ~new_n6230_ | ~new_n6231_;
  assign po276 = ~new_n6226_ | ~new_n6227_ | ~new_n6228_;
  assign po275 = ~new_n6223_ | ~new_n6224_ | ~new_n6225_;
  assign po274 = ~new_n6220_ | ~new_n6221_ | ~new_n6222_;
  assign po273 = ~new_n6217_ | ~new_n6218_ | ~new_n6219_;
  assign po272 = ~new_n6214_ | ~new_n6215_ | ~new_n6216_;
  assign po271 = ~new_n6211_ | ~new_n6212_ | ~new_n6213_;
  assign po270 = ~new_n6208_ | ~new_n6209_ | ~new_n6210_;
  assign po269 = ~new_n6205_ | ~new_n6206_ | ~new_n6207_;
  assign po268 = ~new_n6202_ | ~new_n6203_ | ~new_n6204_;
  assign po267 = ~new_n6199_ | ~new_n6200_ | ~new_n6201_;
  assign po479 = new_n6017_ & new_n7861_;
  assign new_n5549_ = ~pi520 | ~new_n6099_;
  assign new_n5550_ = ~new_n1570_;
  assign new_n5551_ = ~pi490;
  assign new_n5552_ = ~new_n5634_ | ~new_n7869_;
  assign new_n5553_ = ~new_n5634_ | ~new_n6295_;
  assign new_n5554_ = ~new_n5640_ | ~new_n7891_ | ~new_n5644_;
  assign new_n5555_ = ~new_n5640_ | ~new_n5638_ | ~new_n5644_;
  assign new_n5556_ = ~new_n5269_ | ~new_n5640_;
  assign new_n5557_ = ~new_n5639_ | ~new_n5638_ | ~new_n5644_;
  assign new_n5558_ = ~new_n5269_ | ~new_n5639_;
  assign new_n5559_ = ~new_n5640_ | ~new_n7888_ | ~new_n7894_;
  assign new_n5560_ = ~new_n7891_ | ~new_n7888_;
  assign new_n5561_ = ~new_n6194_ | ~new_n5639_;
  assign new_n5562_ = ~new_n6159_ | ~new_n7885_;
  assign new_n5563_ = ~new_n7885_ | ~new_n7894_;
  assign new_n5564_ = ~new_n5640_ | ~new_n5639_;
  assign new_n5565_ = ~new_n7885_ | ~new_n5644_;
  assign new_n5566_ = ~new_n5269_ | ~new_n7885_;
  assign new_n5567_ = ~new_n7908_ | ~new_n7903_;
  assign new_n5568_ = ~new_n5783_ | ~new_n5784_ | ~new_n6343_;
  assign new_n5569_ = ~new_n6360_ | ~new_n5800_ | ~new_n5798_ | ~new_n6361_;
  assign new_n5570_ = ~new_n6379_ | ~new_n5804_ | ~new_n5802_ | ~new_n6380_;
  assign new_n5571_ = ~new_n6398_ | ~new_n5808_ | ~new_n5806_ | ~new_n6399_;
  assign new_n5572_ = ~new_n6417_ | ~new_n5812_ | ~new_n5810_ | ~new_n6418_;
  assign new_n5573_ = ~new_n6436_ | ~new_n5816_ | ~new_n5814_ | ~new_n6437_;
  assign new_n5574_ = ~new_n6455_ | ~new_n5820_ | ~new_n5818_ | ~new_n6456_;
  assign new_n5575_ = ~new_n6474_ | ~new_n5824_ | ~new_n5822_ | ~new_n6475_;
  assign new_n5576_ = ~new_n6493_ | ~new_n5828_ | ~new_n5826_ | ~new_n6494_;
  assign new_n5577_ = ~new_n6512_ | ~new_n5832_ | ~new_n5830_ | ~new_n6513_;
  assign new_n5578_ = ~new_n6531_ | ~new_n5836_ | ~new_n5834_ | ~new_n6532_;
  assign new_n5579_ = ~new_n6550_ | ~new_n5840_ | ~new_n5838_ | ~new_n6551_;
  assign new_n5580_ = ~new_n6569_ | ~new_n5844_ | ~new_n5842_ | ~new_n6570_;
  assign new_n5581_ = ~new_n6588_ | ~new_n5848_ | ~new_n5846_ | ~new_n6589_;
  assign new_n5582_ = ~new_n6607_ | ~new_n5852_ | ~new_n5850_ | ~new_n6608_;
  assign new_n5583_ = ~new_n6626_ | ~new_n5856_ | ~new_n5854_ | ~new_n6627_;
  assign new_n5584_ = ~new_n6645_ | ~new_n5860_ | ~new_n5858_ | ~new_n6646_;
  assign new_n5585_ = ~new_n6664_ | ~new_n5864_ | ~new_n5862_ | ~new_n6665_;
  assign new_n5586_ = ~new_n6683_ | ~new_n5868_ | ~new_n5866_ | ~new_n6684_;
  assign new_n5587_ = ~new_n6702_ | ~new_n5872_ | ~new_n5870_ | ~new_n6703_;
  assign new_n5588_ = ~new_n1582_ | ~new_n5567_;
  assign new_n5589_ = ~new_n6721_ | ~new_n5876_ | ~new_n5874_ | ~new_n6722_;
  assign new_n5590_ = ~new_n1581_ | ~new_n5567_;
  assign new_n5591_ = ~new_n6740_ | ~new_n5880_ | ~new_n5878_ | ~new_n6741_;
  assign new_n5592_ = ~new_n1580_ | ~new_n5567_;
  assign new_n5593_ = ~new_n6759_ | ~new_n5884_ | ~new_n5882_ | ~new_n6760_;
  assign new_n5594_ = ~new_n1579_ | ~new_n5567_;
  assign new_n5595_ = ~new_n6778_ | ~new_n5888_ | ~new_n5886_ | ~new_n6779_;
  assign new_n5596_ = ~new_n1578_ | ~new_n5567_;
  assign new_n5597_ = ~new_n6797_ | ~new_n5892_ | ~new_n5890_ | ~new_n6798_;
  assign new_n5598_ = ~new_n1577_ | ~new_n5567_;
  assign new_n5599_ = ~new_n6816_ | ~new_n5896_ | ~new_n5894_ | ~new_n6817_;
  assign new_n5600_ = ~new_n1576_ | ~new_n5567_;
  assign new_n5601_ = ~new_n6835_ | ~new_n5900_ | ~new_n5898_ | ~new_n6836_;
  assign new_n5602_ = ~new_n1575_ | ~new_n5567_;
  assign new_n5603_ = ~new_n6854_ | ~new_n5904_ | ~new_n5902_ | ~new_n6855_;
  assign new_n5604_ = ~new_n1574_ | ~new_n5567_;
  assign new_n5605_ = ~new_n6874_ | ~new_n5907_ | ~new_n6876_ | ~new_n6875_ | ~new_n6873_;
  assign new_n5606_ = ~new_n1573_ | ~new_n5567_;
  assign new_n5607_ = ~new_n6894_ | ~new_n5912_ | ~new_n5910_ | ~new_n6895_ | ~new_n6893_;
  assign new_n5608_ = ~new_n1571_ | ~new_n5567_;
  assign new_n5609_ = ~new_n1570_ | ~new_n5567_;
  assign new_n5610_ = ~new_n6164_ | ~new_n5644_;
  assign new_n5611_ = ~new_n5243_ | ~new_n6918_;
  assign new_n5612_ = ~new_n5639_ | ~new_n7891_ | ~new_n5644_;
  assign new_n5613_ = ~new_n6141_ | ~new_n7891_;
  assign new_n5614_ = ~new_n6164_ | ~new_n7888_;
  assign new_n5615_ = ~new_n6147_ | ~new_n7891_;
  assign new_n5616_ = ~new_n5634_ | ~new_n5633_ | ~new_n5632_;
  assign new_n5617_ = ~new_n5564_ | ~new_n5567_;
  assign new_n5618_ = ~new_n6154_ | ~new_n6919_;
  assign new_n5619_ = ~new_n6182_ | ~new_n7878_;
  assign new_n5620_ = ~new_n6197_ | ~pi520;
  assign new_n5621_ = ~new_n5976_ | ~new_n5272_;
  assign new_n5622_ = ~new_n6194_ | ~new_n5640_;
  assign new_n5623_ = ~new_n5235_ | ~new_n5238_;
  assign new_n5624_ = ~new_n7894_ | ~new_n5644_;
  assign new_n5625_ = ~new_n5243_ | ~new_n5618_;
  assign new_n5626_ = ~new_n6018_ | ~new_n5236_;
  assign new_n5627_ = ~new_n5616_ | ~new_n7388_ | ~pi520;
  assign new_n5628_ = ~new_n6022_ | ~new_n7392_;
  assign new_n5629_ = ~new_n19210_;
  assign new_n5630_ = ~new_n6158_ | ~new_n7885_;
  assign new_n5631_ = ~new_n5556_ | ~new_n6143_ | ~new_n5566_ | ~new_n5555_;
  assign new_n5632_ = ~new_n7865_ | ~new_n7864_;
  assign new_n5633_ = ~new_n7868_ | ~new_n7867_;
  assign new_n5634_ = ~new_n7871_ | ~new_n7870_;
  assign new_n5635_ = ~new_n7877_ | ~new_n7876_;
  assign po299 = ~new_n7880_ | ~new_n7879_;
  assign po300 = ~new_n7882_ | ~new_n7881_;
  assign new_n5638_ = ~new_n7890_ | ~new_n7889_;
  assign new_n5639_ = ~new_n7893_ | ~new_n7892_;
  assign new_n5640_ = ~new_n7884_ | ~new_n7883_;
  assign new_n5641_ = ~new_n7896_ | ~new_n7895_;
  assign new_n5642_ = ~new_n7899_ | ~new_n7898_;
  assign new_n5643_ = ~new_n7902_ | ~new_n7901_;
  assign new_n5644_ = ~new_n7887_ | ~new_n7886_;
  assign new_n5645_ = ~new_n7905_ | ~new_n7904_;
  assign new_n5646_ = ~new_n7907_ | ~new_n7906_;
  assign new_n5647_ = ~new_n7910_ | ~new_n7909_;
  assign new_n5648_ = ~new_n7918_ | ~new_n7917_;
  assign new_n5649_ = ~new_n7915_ | ~new_n7914_;
  assign po331 = ~new_n7921_ | ~new_n7920_;
  assign new_n5651_ = ~new_n7923_ | ~new_n7922_;
  assign new_n5652_ = ~new_n7925_ | ~new_n7924_;
  assign po332 = ~new_n7928_ | ~new_n7927_;
  assign new_n5654_ = ~new_n7930_ | ~new_n7929_;
  assign new_n5655_ = ~new_n7932_ | ~new_n7931_;
  assign po333 = ~new_n7935_ | ~new_n7934_;
  assign new_n5657_ = ~new_n7937_ | ~new_n7936_;
  assign new_n5658_ = ~new_n7939_ | ~new_n7938_;
  assign po334 = ~new_n7942_ | ~new_n7941_;
  assign new_n5660_ = ~new_n7944_ | ~new_n7943_;
  assign new_n5661_ = ~new_n7946_ | ~new_n7945_;
  assign po335 = ~new_n7949_ | ~new_n7948_;
  assign new_n5663_ = ~new_n7951_ | ~new_n7950_;
  assign new_n5664_ = ~new_n7953_ | ~new_n7952_;
  assign po336 = ~new_n7956_ | ~new_n7955_;
  assign new_n5666_ = ~new_n7958_ | ~new_n7957_;
  assign new_n5667_ = ~new_n7960_ | ~new_n7959_;
  assign po337 = ~new_n7963_ | ~new_n7962_;
  assign new_n5669_ = ~new_n7965_ | ~new_n7964_;
  assign new_n5670_ = ~new_n7967_ | ~new_n7966_;
  assign po338 = ~new_n7970_ | ~new_n7969_;
  assign new_n5672_ = ~new_n7972_ | ~new_n7971_;
  assign new_n5673_ = ~new_n7974_ | ~new_n7973_;
  assign po339 = ~new_n7977_ | ~new_n7976_;
  assign new_n5675_ = ~new_n7979_ | ~new_n7978_;
  assign new_n5676_ = ~new_n7981_ | ~new_n7980_;
  assign po340 = ~new_n7984_ | ~new_n7983_;
  assign new_n5678_ = ~new_n7986_ | ~new_n7985_;
  assign new_n5679_ = ~new_n7988_ | ~new_n7987_;
  assign po341 = ~new_n7991_ | ~new_n7990_;
  assign new_n5681_ = ~new_n7993_ | ~new_n7992_;
  assign new_n5682_ = ~new_n7995_ | ~new_n7994_;
  assign po342 = ~new_n7998_ | ~new_n7997_;
  assign new_n5684_ = ~new_n8000_ | ~new_n7999_;
  assign new_n5685_ = ~new_n8002_ | ~new_n8001_;
  assign po343 = ~new_n8005_ | ~new_n8004_;
  assign new_n5687_ = ~new_n8007_ | ~new_n8006_;
  assign new_n5688_ = ~new_n8009_ | ~new_n8008_;
  assign po344 = ~new_n8012_ | ~new_n8011_;
  assign new_n5690_ = ~new_n8014_ | ~new_n8013_;
  assign new_n5691_ = ~new_n8016_ | ~new_n8015_;
  assign po345 = ~new_n8019_ | ~new_n8018_;
  assign new_n5693_ = ~new_n8021_ | ~new_n8020_;
  assign new_n5694_ = ~new_n8023_ | ~new_n8022_;
  assign po346 = ~new_n8026_ | ~new_n8025_;
  assign new_n5696_ = ~new_n8028_ | ~new_n8027_;
  assign new_n5697_ = ~new_n8030_ | ~new_n8029_;
  assign po347 = ~new_n8033_ | ~new_n8032_;
  assign new_n5699_ = ~new_n8035_ | ~new_n8034_;
  assign new_n5700_ = ~new_n8037_ | ~new_n8036_;
  assign po348 = ~new_n8040_ | ~new_n8039_;
  assign new_n5702_ = ~new_n8042_ | ~new_n8041_;
  assign new_n5703_ = ~new_n8044_ | ~new_n8043_;
  assign po349 = ~new_n8047_ | ~new_n8046_;
  assign new_n5705_ = ~new_n8049_ | ~new_n8048_;
  assign po350 = ~new_n8052_ | ~new_n8051_;
  assign po351 = ~new_n8054_ | ~new_n8053_;
  assign po352 = ~new_n8056_ | ~new_n8055_;
  assign po353 = ~new_n8058_ | ~new_n8057_;
  assign po354 = ~new_n8060_ | ~new_n8059_;
  assign po355 = ~new_n8062_ | ~new_n8061_;
  assign po356 = ~new_n8064_ | ~new_n8063_;
  assign po357 = ~new_n8066_ | ~new_n8065_;
  assign po358 = ~new_n8068_ | ~new_n8067_;
  assign po359 = ~new_n8070_ | ~new_n8069_;
  assign po360 = ~new_n8072_ | ~new_n8071_;
  assign po361 = ~new_n8074_ | ~new_n8073_;
  assign po362 = ~new_n8076_ | ~new_n8075_;
  assign po363 = ~new_n8078_ | ~new_n8077_;
  assign po364 = ~new_n8080_ | ~new_n8079_;
  assign po365 = ~new_n8082_ | ~new_n8081_;
  assign po366 = ~new_n8084_ | ~new_n8083_;
  assign po367 = ~new_n8086_ | ~new_n8085_;
  assign po368 = ~new_n8088_ | ~new_n8087_;
  assign po369 = ~new_n8090_ | ~new_n8089_;
  assign po370 = ~new_n8092_ | ~new_n8091_;
  assign po371 = ~new_n8094_ | ~new_n8093_;
  assign po372 = ~new_n8096_ | ~new_n8095_;
  assign po373 = ~new_n8098_ | ~new_n8097_;
  assign po374 = ~new_n8100_ | ~new_n8099_;
  assign po375 = ~new_n8102_ | ~new_n8101_;
  assign po376 = ~new_n8104_ | ~new_n8103_;
  assign po377 = ~new_n8106_ | ~new_n8105_;
  assign po378 = ~new_n8108_ | ~new_n8107_;
  assign po379 = ~new_n8110_ | ~new_n8109_;
  assign po380 = ~new_n8112_ | ~new_n8111_;
  assign po381 = ~new_n8114_ | ~new_n8113_;
  assign po382 = ~new_n8116_ | ~new_n8115_;
  assign po383 = ~new_n8118_ | ~new_n8117_;
  assign po384 = ~new_n8120_ | ~new_n8119_;
  assign po385 = ~new_n8122_ | ~new_n8121_;
  assign po386 = ~new_n8124_ | ~new_n8123_;
  assign po387 = ~new_n8126_ | ~new_n8125_;
  assign po388 = ~new_n8128_ | ~new_n8127_;
  assign po389 = ~new_n8130_ | ~new_n8129_;
  assign po390 = ~new_n8132_ | ~new_n8131_;
  assign po391 = ~new_n8134_ | ~new_n8133_;
  assign po392 = ~new_n8136_ | ~new_n8135_;
  assign po393 = ~new_n8138_ | ~new_n8137_;
  assign po394 = ~new_n8140_ | ~new_n8139_;
  assign po447 = ~new_n8206_ | ~new_n8205_;
  assign po448 = ~new_n8208_ | ~new_n8207_;
  assign po449 = ~new_n8210_ | ~new_n8209_;
  assign po450 = ~new_n8212_ | ~new_n8211_;
  assign po451 = ~new_n8214_ | ~new_n8213_;
  assign po452 = ~new_n8216_ | ~new_n8215_;
  assign po453 = ~new_n8218_ | ~new_n8217_;
  assign po454 = ~new_n8220_ | ~new_n8219_;
  assign po455 = ~new_n8222_ | ~new_n8221_;
  assign po456 = ~new_n8224_ | ~new_n8223_;
  assign po457 = ~new_n8226_ | ~new_n8225_;
  assign po458 = ~new_n8228_ | ~new_n8227_;
  assign po459 = ~new_n8230_ | ~new_n8229_;
  assign po460 = ~new_n8232_ | ~new_n8231_;
  assign po461 = ~new_n8234_ | ~new_n8233_;
  assign po462 = ~new_n8236_ | ~new_n8235_;
  assign po463 = ~new_n8238_ | ~new_n8237_;
  assign po464 = ~new_n8240_ | ~new_n8239_;
  assign po465 = ~new_n8242_ | ~new_n8241_;
  assign po466 = ~new_n8244_ | ~new_n8243_;
  assign po467 = ~new_n8246_ | ~new_n8245_;
  assign po468 = ~new_n8248_ | ~new_n8247_;
  assign po469 = ~new_n8250_ | ~new_n8249_;
  assign po470 = ~new_n8252_ | ~new_n8251_;
  assign po471 = ~new_n8254_ | ~new_n8253_;
  assign po472 = ~new_n8256_ | ~new_n8255_;
  assign po473 = ~new_n8258_ | ~new_n8257_;
  assign po474 = ~new_n8260_ | ~new_n8259_;
  assign po475 = ~new_n8262_ | ~new_n8261_;
  assign po476 = ~new_n8264_ | ~new_n8263_;
  assign po477 = ~new_n8266_ | ~new_n8265_;
  assign po478 = ~new_n8268_ | ~new_n8267_;
  assign new_n5783_ = new_n6339_ & new_n6337_ & new_n6338_ & new_n6340_;
  assign new_n5784_ = new_n6342_ & new_n6341_;
  assign new_n5785_ = new_n6347_ & new_n6345_;
  assign new_n5786_ = new_n6301_ & new_n6299_ & new_n6300_ & new_n6302_;
  assign new_n5787_ = new_n6305_ & new_n6303_ & new_n6304_ & new_n6306_;
  assign new_n5788_ = new_n6309_ & new_n6307_ & new_n6308_ & new_n6310_;
  assign new_n5789_ = new_n6313_ & new_n6312_ & new_n6311_;
  assign new_n5790_ = new_n5788_ & new_n5786_ & new_n5787_ & new_n5789_;
  assign new_n5791_ = new_n6316_ & new_n6314_ & new_n6315_ & new_n6317_;
  assign new_n5792_ = new_n6320_ & new_n6318_ & new_n6319_ & new_n6321_;
  assign new_n5793_ = new_n6324_ & new_n6322_ & new_n6323_ & new_n6325_;
  assign new_n5794_ = new_n6328_ & new_n6327_ & new_n6326_;
  assign new_n5795_ = new_n5793_ & new_n5791_ & new_n5792_ & new_n5794_;
  assign new_n5796_ = new_n7916_ & new_n6330_;
  assign new_n5797_ = new_n7919_ & new_n5243_;
  assign new_n5798_ = new_n6363_ & new_n6362_;
  assign new_n5799_ = new_n6365_ & new_n6364_;
  assign new_n5800_ = new_n5799_ & new_n6367_ & new_n6366_;
  assign new_n5801_ = new_n6369_ & new_n6371_ & new_n6372_ & new_n6370_;
  assign new_n5802_ = new_n6382_ & new_n6381_;
  assign new_n5803_ = new_n6384_ & new_n6383_;
  assign new_n5804_ = new_n5803_ & new_n6386_ & new_n6385_;
  assign new_n5805_ = new_n6388_ & new_n6390_ & new_n6391_ & new_n6389_;
  assign new_n5806_ = new_n6401_ & new_n6400_;
  assign new_n5807_ = new_n6403_ & new_n6402_;
  assign new_n5808_ = new_n5807_ & new_n6405_ & new_n6404_;
  assign new_n5809_ = new_n6407_ & new_n6409_ & new_n6410_ & new_n6408_;
  assign new_n5810_ = new_n6420_ & new_n6419_;
  assign new_n5811_ = new_n6422_ & new_n6421_;
  assign new_n5812_ = new_n5811_ & new_n6424_ & new_n6423_;
  assign new_n5813_ = new_n6426_ & new_n6428_ & new_n6429_ & new_n6427_;
  assign new_n5814_ = new_n6439_ & new_n6438_;
  assign new_n5815_ = new_n6441_ & new_n6440_;
  assign new_n5816_ = new_n5815_ & new_n6443_ & new_n6442_;
  assign new_n5817_ = new_n6445_ & new_n6447_ & new_n6448_ & new_n6446_;
  assign new_n5818_ = new_n6458_ & new_n6457_;
  assign new_n5819_ = new_n6460_ & new_n6459_;
  assign new_n5820_ = new_n5819_ & new_n6462_ & new_n6461_;
  assign new_n5821_ = new_n6464_ & new_n6466_ & new_n6467_ & new_n6465_;
  assign new_n5822_ = new_n6477_ & new_n6476_;
  assign new_n5823_ = new_n6479_ & new_n6478_;
  assign new_n5824_ = new_n5823_ & new_n6481_ & new_n6480_;
  assign new_n5825_ = new_n6483_ & new_n6485_ & new_n6486_ & new_n6484_;
  assign new_n5826_ = new_n6496_ & new_n6495_;
  assign new_n5827_ = new_n6498_ & new_n6497_;
  assign new_n5828_ = new_n5827_ & new_n6500_ & new_n6499_;
  assign new_n5829_ = new_n6502_ & new_n6504_ & new_n6505_ & new_n6503_;
  assign new_n5830_ = new_n6515_ & new_n6514_;
  assign new_n5831_ = new_n6517_ & new_n6516_;
  assign new_n5832_ = new_n5831_ & new_n6519_ & new_n6518_;
  assign new_n5833_ = new_n6521_ & new_n6523_ & new_n6524_ & new_n6522_;
  assign new_n5834_ = new_n6534_ & new_n6533_;
  assign new_n5835_ = new_n6536_ & new_n6535_;
  assign new_n5836_ = new_n5835_ & new_n6538_ & new_n6537_;
  assign new_n5837_ = new_n6540_ & new_n6542_ & new_n6543_ & new_n6541_;
  assign new_n5838_ = new_n6553_ & new_n6552_;
  assign new_n5839_ = new_n6555_ & new_n6554_;
  assign new_n5840_ = new_n5839_ & new_n6557_ & new_n6556_;
  assign new_n5841_ = new_n6559_ & new_n6561_ & new_n6562_ & new_n6560_;
  assign new_n5842_ = new_n6572_ & new_n6571_;
  assign new_n5843_ = new_n6574_ & new_n6573_;
  assign new_n5844_ = new_n5843_ & new_n6576_ & new_n6575_;
  assign new_n5845_ = new_n6578_ & new_n6580_ & new_n6581_ & new_n6579_;
  assign new_n5846_ = new_n6591_ & new_n6590_;
  assign new_n5847_ = new_n6593_ & new_n6592_;
  assign new_n5848_ = new_n5847_ & new_n6595_ & new_n6594_;
  assign new_n5849_ = new_n6597_ & new_n6599_ & new_n6600_ & new_n6598_;
  assign new_n5850_ = new_n6610_ & new_n6609_;
  assign new_n5851_ = new_n6612_ & new_n6611_;
  assign new_n5852_ = new_n5851_ & new_n6614_ & new_n6613_;
  assign new_n5853_ = new_n6616_ & new_n6618_ & new_n6619_ & new_n6617_;
  assign new_n5854_ = new_n6629_ & new_n6628_;
  assign new_n5855_ = new_n6631_ & new_n6630_;
  assign new_n5856_ = new_n5855_ & new_n6633_ & new_n6632_;
  assign new_n5857_ = new_n6635_ & new_n6637_ & new_n6638_ & new_n6636_;
  assign new_n5858_ = new_n6648_ & new_n6647_;
  assign new_n5859_ = new_n6650_ & new_n6649_;
  assign new_n5860_ = new_n5859_ & new_n6652_ & new_n6651_;
  assign new_n5861_ = new_n6654_ & new_n6656_ & new_n6657_ & new_n6655_;
  assign new_n5862_ = new_n6667_ & new_n6666_;
  assign new_n5863_ = new_n6669_ & new_n6668_;
  assign new_n5864_ = new_n5863_ & new_n6671_ & new_n6670_;
  assign new_n5865_ = new_n6673_ & new_n6675_ & new_n6676_ & new_n6674_;
  assign new_n5866_ = new_n6686_ & new_n6685_;
  assign new_n5867_ = new_n6688_ & new_n6687_;
  assign new_n5868_ = new_n5867_ & new_n6690_ & new_n6689_;
  assign new_n5869_ = new_n6692_ & new_n6694_ & new_n6695_ & new_n6693_;
  assign new_n5870_ = new_n6705_ & new_n6704_;
  assign new_n5871_ = new_n6707_ & new_n6706_;
  assign new_n5872_ = new_n5871_ & new_n6709_ & new_n6708_;
  assign new_n5873_ = new_n6711_ & new_n6713_ & new_n6714_ & new_n6712_;
  assign new_n5874_ = new_n6724_ & new_n6723_;
  assign new_n5875_ = new_n6726_ & new_n6725_;
  assign new_n5876_ = new_n5875_ & new_n6728_ & new_n6727_;
  assign new_n5877_ = new_n6730_ & new_n6732_ & new_n6733_ & new_n6731_;
  assign new_n5878_ = new_n6743_ & new_n6742_;
  assign new_n5879_ = new_n6745_ & new_n6744_;
  assign new_n5880_ = new_n5879_ & new_n6747_ & new_n6746_;
  assign new_n5881_ = new_n6749_ & new_n6751_ & new_n6752_ & new_n6750_;
  assign new_n5882_ = new_n6762_ & new_n6761_;
  assign new_n5883_ = new_n6764_ & new_n6763_;
  assign new_n5884_ = new_n5883_ & new_n6766_ & new_n6765_;
  assign new_n5885_ = new_n6768_ & new_n6770_ & new_n6771_ & new_n6769_;
  assign new_n5886_ = new_n6781_ & new_n6780_;
  assign new_n5887_ = new_n6783_ & new_n6782_;
  assign new_n5888_ = new_n5887_ & new_n6785_ & new_n6784_;
  assign new_n5889_ = new_n6787_ & new_n6789_ & new_n6790_ & new_n6788_;
  assign new_n5890_ = new_n6800_ & new_n6799_;
  assign new_n5891_ = new_n6802_ & new_n6801_;
  assign new_n5892_ = new_n5891_ & new_n6804_ & new_n6803_;
  assign new_n5893_ = new_n6806_ & new_n6808_ & new_n6809_ & new_n6807_;
  assign new_n5894_ = new_n6819_ & new_n6818_;
  assign new_n5895_ = new_n6821_ & new_n6820_;
  assign new_n5896_ = new_n5895_ & new_n6823_ & new_n6822_;
  assign new_n5897_ = new_n6825_ & new_n6827_ & new_n6828_ & new_n6826_;
  assign new_n5898_ = new_n6838_ & new_n6837_;
  assign new_n5899_ = new_n6840_ & new_n6839_;
  assign new_n5900_ = new_n5899_ & new_n6842_ & new_n6841_;
  assign new_n5901_ = new_n6844_ & new_n6846_ & new_n6847_ & new_n6845_;
  assign new_n5902_ = new_n6857_ & new_n6856_;
  assign new_n5903_ = new_n6859_ & new_n6858_;
  assign new_n5904_ = new_n5903_ & new_n6861_ & new_n6860_;
  assign new_n5905_ = new_n6863_ & new_n6865_ & new_n6866_ & new_n6864_;
  assign new_n5906_ = new_n6878_ & new_n6877_;
  assign new_n5907_ = new_n5906_ & new_n6880_ & new_n6879_;
  assign new_n5908_ = new_n6882_ & new_n6884_ & new_n6885_ & new_n6883_;
  assign new_n5909_ = new_n6892_ & new_n6183_;
  assign new_n5910_ = new_n6897_ & new_n6896_;
  assign new_n5911_ = new_n6899_ & new_n6898_;
  assign new_n5912_ = new_n5911_ & new_n6901_ & new_n6900_;
  assign new_n5913_ = new_n6904_ & new_n6905_ & new_n6903_;
  assign new_n5914_ = new_n6183_ & new_n6892_;
  assign new_n5915_ = new_n5243_ & new_n5648_;
  assign new_n5916_ = new_n5649_ & new_n7919_ & new_n6155_;
  assign new_n5917_ = new_n6923_ & new_n6922_ & new_n6921_;
  assign new_n5918_ = new_n6103_ & new_n6925_ & new_n6924_;
  assign new_n5919_ = new_n6928_ & new_n6927_ & new_n6926_;
  assign new_n5920_ = new_n6104_ & new_n6930_ & new_n6929_;
  assign new_n5921_ = new_n6933_ & new_n6932_ & new_n6931_;
  assign new_n5922_ = new_n6105_ & new_n6935_ & new_n6934_;
  assign new_n5923_ = new_n6938_ & new_n6937_ & new_n6936_;
  assign new_n5924_ = new_n6106_ & new_n6940_ & new_n6939_;
  assign new_n5925_ = new_n6943_ & new_n6942_ & new_n6941_;
  assign new_n5926_ = new_n6107_ & new_n6945_ & new_n6944_;
  assign new_n5927_ = new_n6948_ & new_n6947_ & new_n6946_;
  assign new_n5928_ = new_n6108_ & new_n6950_ & new_n6949_;
  assign new_n5929_ = new_n6953_ & new_n6952_ & new_n6951_;
  assign new_n5930_ = new_n6109_ & new_n6955_ & new_n6954_;
  assign new_n5931_ = new_n6958_ & new_n6957_ & new_n6956_;
  assign new_n5932_ = new_n6110_ & new_n6960_ & new_n6959_;
  assign new_n5933_ = new_n6963_ & new_n6962_ & new_n6961_;
  assign new_n5934_ = new_n6111_ & new_n6965_ & new_n6964_;
  assign new_n5935_ = new_n6968_ & new_n6967_ & new_n6966_;
  assign new_n5936_ = new_n6112_ & new_n6970_ & new_n6969_;
  assign new_n5937_ = new_n6973_ & new_n6972_ & new_n6971_;
  assign new_n5938_ = new_n6975_ & new_n6974_;
  assign new_n5939_ = new_n6978_ & new_n6977_ & new_n6976_;
  assign new_n5940_ = new_n6980_ & new_n6979_;
  assign new_n5941_ = new_n6983_ & new_n6982_ & new_n6981_;
  assign new_n5942_ = new_n6985_ & new_n6984_;
  assign new_n5943_ = new_n6987_ & new_n6988_ & new_n6986_;
  assign new_n5944_ = new_n6990_ & new_n6989_;
  assign new_n5945_ = new_n6993_ & new_n6992_ & new_n6991_;
  assign new_n5946_ = new_n6995_ & new_n6994_;
  assign new_n5947_ = new_n6997_ & new_n6998_ & new_n6996_;
  assign new_n5948_ = new_n7000_ & new_n6999_;
  assign new_n5949_ = new_n7003_ & new_n7001_;
  assign new_n5950_ = new_n7005_ & new_n7004_;
  assign new_n5951_ = new_n7008_ & new_n7006_;
  assign new_n5952_ = new_n7010_ & new_n7009_;
  assign new_n5953_ = new_n7013_ & new_n7011_;
  assign new_n5954_ = new_n7015_ & new_n7014_;
  assign new_n5955_ = new_n7018_ & new_n7016_;
  assign new_n5956_ = new_n7020_ & new_n7019_;
  assign new_n5957_ = new_n7023_ & new_n7021_;
  assign new_n5958_ = new_n7025_ & new_n7024_;
  assign new_n5959_ = new_n7028_ & new_n7026_;
  assign new_n5960_ = new_n7030_ & new_n7029_;
  assign new_n5961_ = new_n7033_ & new_n7031_;
  assign new_n5962_ = new_n7035_ & new_n7034_;
  assign new_n5963_ = new_n7038_ & new_n7036_;
  assign new_n5964_ = new_n7040_ & new_n7039_;
  assign new_n5965_ = new_n7043_ & new_n7041_;
  assign new_n5966_ = new_n7045_ & new_n7044_;
  assign new_n5967_ = new_n7048_ & new_n7046_;
  assign new_n5968_ = new_n7050_ & new_n7049_;
  assign new_n5969_ = new_n7053_ & new_n7051_;
  assign new_n5970_ = new_n7055_ & new_n7054_;
  assign new_n5971_ = new_n7058_ & new_n7056_;
  assign new_n5972_ = new_n7060_ & new_n7059_;
  assign new_n5973_ = new_n7063_ & new_n7061_;
  assign new_n5974_ = new_n7065_ & new_n7064_;
  assign new_n5975_ = new_n5554_ & new_n5555_ & new_n5556_;
  assign new_n5976_ = new_n7863_ & new_n5617_;
  assign new_n5977_ = new_n5635_ & pi520;
  assign new_n5978_ = new_n7090_ & new_n7086_ & new_n7087_ & new_n7089_ & new_n7088_;
  assign new_n5979_ = new_n7105_ & new_n7101_ & new_n7102_ & new_n7104_ & new_n7103_;
  assign new_n5980_ = new_n7120_ & new_n7116_ & new_n7117_ & new_n7119_ & new_n7118_;
  assign new_n5981_ = new_n7135_ & new_n7131_ & new_n7132_ & new_n7134_ & new_n7133_;
  assign new_n5982_ = new_n7150_ & new_n7146_ & new_n7147_ & new_n7149_ & new_n7148_;
  assign new_n5983_ = new_n7165_ & new_n7161_ & new_n7162_ & new_n7164_ & new_n7163_;
  assign new_n5984_ = new_n7180_ & new_n7176_ & new_n7177_ & new_n7179_ & new_n7178_;
  assign new_n5985_ = new_n7195_ & new_n7191_ & new_n7192_ & new_n7194_ & new_n7193_;
  assign new_n5986_ = new_n7209_ & new_n7206_ & new_n7207_ & new_n7210_ & new_n7208_;
  assign new_n5987_ = new_n7225_ & new_n7221_ & new_n7222_ & new_n7224_ & new_n7223_;
  assign new_n5988_ = new_n7239_ & new_n7236_ & new_n7237_ & new_n7240_ & new_n7238_;
  assign new_n5989_ = new_n7252_ & new_n7251_;
  assign new_n5990_ = new_n7255_ & new_n7254_ & new_n7253_;
  assign new_n5991_ = new_n7267_ & new_n7266_;
  assign new_n5992_ = new_n7270_ & new_n7269_ & new_n7268_;
  assign new_n5993_ = new_n7282_ & new_n7281_;
  assign new_n5994_ = new_n7285_ & new_n7284_ & new_n7283_;
  assign new_n5995_ = new_n7297_ & new_n7296_;
  assign new_n5996_ = new_n7300_ & new_n7299_ & new_n7298_;
  assign new_n5997_ = new_n7312_ & new_n7311_;
  assign new_n5998_ = new_n7315_ & new_n7314_ & new_n7313_;
  assign new_n5999_ = new_n7327_ & new_n7326_;
  assign new_n6000_ = new_n7330_ & new_n7329_ & new_n7328_;
  assign new_n6001_ = new_n7342_ & new_n7341_;
  assign new_n6002_ = new_n7345_ & new_n7344_ & new_n7343_;
  assign new_n6003_ = new_n7357_ & new_n7356_;
  assign new_n6004_ = new_n7360_ & new_n7359_ & new_n7358_;
  assign new_n6005_ = new_n7372_ & new_n7371_;
  assign new_n6006_ = new_n7375_ & new_n7374_ & new_n7373_;
  assign new_n6007_ = new_n7859_ & new_n7878_;
  assign new_n6008_ = new_n8326_ & new_n8323_ & new_n8320_;
  assign new_n6009_ = new_n8314_ & new_n8308_ & new_n8311_ & new_n8317_;
  assign new_n6010_ = new_n8338_ & new_n8332_ & new_n8335_ & new_n8341_;
  assign new_n6011_ = new_n8344_ & new_n8353_ & new_n8350_ & new_n8347_;
  assign new_n6012_ = new_n6008_ & new_n6010_ & new_n6011_ & new_n8329_ & new_n6009_;
  assign new_n6013_ = new_n6016_ & new_n8275_ & new_n8278_ & new_n8281_ & new_n6015_;
  assign new_n6014_ = new_n8365_ & new_n8368_ & new_n8356_ & new_n8359_ & new_n8362_;
  assign new_n6015_ = new_n8290_ & new_n8284_ & new_n8287_ & new_n8293_;
  assign new_n6016_ = new_n8299_ & new_n8296_;
  assign new_n6017_ = new_n7860_ & new_n7851_;
  assign new_n6018_ = new_n5648_ & new_n5649_;
  assign new_n6019_ = new_n5559_ & new_n6148_;
  assign new_n6020_ = new_n6019_ & new_n5562_;
  assign new_n6021_ = new_n5615_ & new_n5630_;
  assign new_n6022_ = new_n5619_ & new_n7878_ & new_n6155_;
  assign new_n6023_ = new_n5243_ & new_n7391_;
  assign new_n6024_ = new_n7418_ & new_n7416_;
  assign new_n6025_ = new_n7436_ & new_n7434_;
  assign new_n6026_ = new_n6189_ & new_n5300_;
  assign new_n6027_ = new_n7479_ & new_n7478_;
  assign new_n6028_ = new_n7482_ & new_n7481_;
  assign new_n6029_ = new_n7498_ & new_n7496_;
  assign new_n6030_ = new_n7525_ & new_n7523_;
  assign new_n6031_ = new_n7570_ & new_n7568_;
  assign new_n6032_ = new_n7579_ & new_n7577_;
  assign new_n6033_ = new_n7606_ & new_n7604_;
  assign new_n6034_ = new_n7651_ & new_n7649_;
  assign new_n6035_ = new_n7655_ & pi520;
  assign new_n6036_ = new_n6140_ & new_n6139_ & new_n6156_;
  assign new_n6037_ = new_n7891_ & new_n5639_;
  assign new_n6038_ = new_n5614_ & new_n5559_;
  assign new_n6039_ = new_n6038_ & new_n5562_ & new_n5610_;
  assign new_n6040_ = new_n5554_ & new_n6148_;
  assign new_n6041_ = new_n5635_ & new_n7664_;
  assign new_n6042_ = new_n5635_ & new_n7667_;
  assign new_n6043_ = new_n5635_ & new_n7670_;
  assign new_n6044_ = new_n5635_ & new_n7673_;
  assign new_n6045_ = new_n5635_ & new_n7676_;
  assign new_n6046_ = new_n6047_ & new_n7677_;
  assign new_n6047_ = new_n5635_ & new_n7679_;
  assign new_n6048_ = new_n7680_ & new_n5630_;
  assign new_n6049_ = new_n6050_ & new_n7685_;
  assign new_n6050_ = new_n5635_ & new_n7687_;
  assign new_n6051_ = new_n5635_ & new_n7688_;
  assign new_n6052_ = new_n5635_ & new_n7691_;
  assign new_n6053_ = new_n5635_ & new_n7694_;
  assign new_n6054_ = new_n5635_ & new_n7697_;
  assign new_n6055_ = new_n5635_ & new_n7700_;
  assign new_n6056_ = new_n5635_ & new_n7703_;
  assign new_n6057_ = new_n5635_ & new_n7706_;
  assign new_n6058_ = new_n5635_ & new_n7709_;
  assign new_n6059_ = new_n5635_ & new_n7712_;
  assign new_n6060_ = new_n5635_ & new_n7715_;
  assign new_n6061_ = new_n6062_ & new_n7718_;
  assign new_n6062_ = new_n5635_ & new_n7720_;
  assign new_n6063_ = new_n5635_ & new_n7721_;
  assign new_n6064_ = new_n5635_ & new_n7724_;
  assign new_n6065_ = new_n5635_ & new_n7727_;
  assign new_n6066_ = new_n5635_ & new_n7730_;
  assign new_n6067_ = new_n5635_ & new_n7733_;
  assign new_n6068_ = new_n5635_ & new_n7736_;
  assign new_n6069_ = new_n5635_ & new_n7739_;
  assign new_n6070_ = new_n5635_ & new_n7742_;
  assign new_n6071_ = new_n5635_ & new_n7747_;
  assign new_n6072_ = new_n5635_ & new_n7750_;
  assign new_n6073_ = new_n6074_ & new_n7751_;
  assign new_n6074_ = new_n5635_ & new_n7753_;
  assign new_n6075_ = new_n6076_ & new_n7754_;
  assign new_n6076_ = new_n5635_ & new_n7756_;
  assign new_n6077_ = new_n7759_ & new_n7760_;
  assign new_n6078_ = new_n7762_ & new_n7763_;
  assign new_n6079_ = new_n7784_ & new_n7785_;
  assign new_n6080_ = new_n7787_ & new_n7788_;
  assign new_n6081_ = new_n7790_ & new_n7791_;
  assign new_n6082_ = new_n7793_ & new_n7794_;
  assign new_n6083_ = new_n7796_ & new_n7797_;
  assign new_n6084_ = new_n7799_ & new_n7800_;
  assign new_n6085_ = new_n7802_ & new_n7803_;
  assign new_n6086_ = new_n7805_ & new_n7806_;
  assign new_n6087_ = new_n7808_ & new_n7809_;
  assign new_n6088_ = new_n7811_ & new_n7812_;
  assign new_n6089_ = new_n7817_ & new_n7818_;
  assign new_n6090_ = new_n7820_ & new_n7821_;
  assign new_n6091_ = new_n7823_ & new_n7824_;
  assign new_n6092_ = new_n7826_ & new_n7827_;
  assign new_n6093_ = new_n7829_ & new_n7830_;
  assign new_n6094_ = new_n7832_ & new_n7833_;
  assign new_n6095_ = new_n7835_ & new_n7836_;
  assign new_n6096_ = new_n7838_ & new_n7839_;
  assign new_n6097_ = new_n7841_ & new_n7842_;
  assign new_n6098_ = new_n7844_ & new_n7845_;
  assign new_n6099_ = ~pi309;
  assign new_n6100_ = ~new_n5243_ | ~new_n5553_;
  assign new_n6101_ = ~new_n5797_ | ~new_n5270_;
  assign new_n6102_ = ~new_n5915_ | ~new_n5270_;
  assign new_n6103_ = new_n8142_ & new_n8141_;
  assign new_n6104_ = new_n8144_ & new_n8143_;
  assign new_n6105_ = new_n8146_ & new_n8145_;
  assign new_n6106_ = new_n8148_ & new_n8147_;
  assign new_n6107_ = new_n8150_ & new_n8149_;
  assign new_n6108_ = new_n8152_ & new_n8151_;
  assign new_n6109_ = new_n8154_ & new_n8153_;
  assign new_n6110_ = new_n8156_ & new_n8155_;
  assign new_n6111_ = new_n8158_ & new_n8157_;
  assign new_n6112_ = new_n8160_ & new_n8159_;
  assign new_n6113_ = new_n8162_ & new_n8161_;
  assign new_n6114_ = new_n8164_ & new_n8163_;
  assign new_n6115_ = new_n8166_ & new_n8165_;
  assign new_n6116_ = new_n8168_ & new_n8167_;
  assign new_n6117_ = new_n8170_ & new_n8169_;
  assign new_n6118_ = new_n8172_ & new_n8171_;
  assign new_n6119_ = new_n8174_ & new_n8173_;
  assign new_n6120_ = new_n8176_ & new_n8175_;
  assign new_n6121_ = new_n8178_ & new_n8177_;
  assign new_n6122_ = new_n8180_ & new_n8179_;
  assign new_n6123_ = new_n8182_ & new_n8181_;
  assign new_n6124_ = new_n8184_ & new_n8183_;
  assign new_n6125_ = new_n8186_ & new_n8185_;
  assign new_n6126_ = new_n8188_ & new_n8187_;
  assign new_n6127_ = new_n8190_ & new_n8189_;
  assign new_n6128_ = new_n8192_ & new_n8191_;
  assign new_n6129_ = new_n8194_ & new_n8193_;
  assign new_n6130_ = new_n8196_ & new_n8195_;
  assign new_n6131_ = new_n8198_ & new_n8197_;
  assign new_n6132_ = new_n8200_ & new_n8199_;
  assign new_n6133_ = ~new_n5914_ | ~new_n5278_;
  assign new_n6134_ = new_n8202_ & new_n8201_;
  assign new_n6135_ = new_n8204_ & new_n8203_;
  assign new_n6136_ = ~new_n19224_;
  assign new_n6137_ = new_n8270_ & new_n8269_;
  assign new_n6138_ = ~new_n6014_ | ~new_n6013_ | ~new_n8302_ | ~new_n8305_ | ~new_n6012_;
  assign new_n6139_ = ~new_n5269_ | ~new_n7894_;
  assign new_n6140_ = ~new_n6193_ | ~new_n5638_;
  assign new_n6141_ = ~new_n5610_;
  assign new_n6142_ = ~new_n5562_;
  assign new_n6143_ = ~new_n6196_ | ~new_n5638_;
  assign new_n6144_ = ~new_n5559_;
  assign new_n6145_ = ~new_n5566_;
  assign new_n6146_ = ~new_n5556_;
  assign new_n6147_ = ~new_n5614_;
  assign new_n6148_ = ~new_n6193_ | ~new_n5640_;
  assign new_n6149_ = ~new_n5630_;
  assign new_n6150_ = ~new_n5555_;
  assign new_n6151_ = ~new_n5554_;
  assign new_n6152_ = ~new_n5615_;
  assign new_n6153_ = ~new_n5613_;
  assign new_n6154_ = ~new_n6145_ | ~new_n7894_;
  assign new_n6155_ = ~new_n6183_ | ~new_n5560_;
  assign new_n6156_ = ~new_n6193_ | ~new_n7891_;
  assign new_n6157_ = ~new_n5622_;
  assign new_n6158_ = ~new_n5612_;
  assign new_n6159_ = ~new_n5561_;
  assign new_n6160_ = ~new_n6139_;
  assign new_n6161_ = ~new_n5557_;
  assign new_n6162_ = ~new_n6140_;
  assign new_n6163_ = ~new_n5558_;
  assign new_n6164_ = ~new_n5563_;
  assign new_n6165_ = ~new_n5567_;
  assign new_n6166_ = ~new_n5626_;
  assign po511 = ~new_n5620_;
  assign new_n6168_ = ~new_n5617_;
  assign new_n6169_ = ~new_n5604_;
  assign new_n6170_ = ~new_n5602_;
  assign new_n6171_ = ~new_n5600_;
  assign new_n6172_ = ~new_n5598_;
  assign new_n6173_ = ~new_n5596_;
  assign new_n6174_ = ~new_n5594_;
  assign new_n6175_ = ~new_n5592_;
  assign new_n6176_ = ~new_n5590_;
  assign new_n6177_ = ~new_n5588_;
  assign new_n6178_ = ~new_n5609_;
  assign new_n6179_ = ~new_n5608_;
  assign new_n6180_ = ~new_n5606_;
  assign new_n6181_ = ~new_n5623_;
  assign new_n6182_ = ~new_n5616_;
  assign new_n6183_ = ~new_n5564_;
  assign new_n6184_ = ~new_n5611_;
  assign new_n6185_ = ~new_n6102_;
  assign new_n6186_ = ~new_n6101_;
  assign new_n6187_ = ~new_n6100_;
  assign new_n6188_ = ~new_n6133_;
  assign new_n6189_ = ~new_n5627_;
  assign new_n6190_ = ~new_n5628_ | ~pi520;
  assign new_n6191_ = ~new_n6153_ | ~new_n5243_;
  assign new_n6192_ = ~new_n5625_;
  assign new_n6193_ = ~new_n5624_;
  assign new_n6194_ = ~new_n5560_;
  assign new_n6195_ = ~new_n5552_;
  assign new_n6196_ = ~new_n5565_;
  assign new_n6197_ = ~new_n5619_;
  assign new_n6198_ = ~new_n5549_;
  assign new_n6199_ = ~new_n1594_ | ~po509;
  assign new_n6200_ = ~pi278 | ~new_n5250_;
  assign new_n6201_ = ~pi278 | ~new_n6198_;
  assign new_n6202_ = ~new_n1583_ | ~po509;
  assign new_n6203_ = ~new_n19049_ | ~new_n5250_;
  assign new_n6204_ = ~pi279 | ~new_n6198_;
  assign new_n6205_ = ~new_n1572_ | ~po509;
  assign new_n6206_ = ~new_n19024_ | ~new_n5250_;
  assign new_n6207_ = ~pi280 | ~new_n6198_;
  assign new_n6208_ = ~new_n1569_ | ~po509;
  assign new_n6209_ = ~new_n19025_ | ~new_n5250_;
  assign new_n6210_ = ~pi281 | ~new_n6198_;
  assign new_n6211_ = ~new_n1568_ | ~po509;
  assign new_n6212_ = ~new_n19026_ | ~new_n5250_;
  assign new_n6213_ = ~pi282 | ~new_n6198_;
  assign new_n6214_ = ~new_n1567_ | ~po509;
  assign new_n6215_ = ~new_n19108_ | ~new_n5250_;
  assign new_n6216_ = ~pi283 | ~new_n6198_;
  assign new_n6217_ = ~new_n1566_ | ~po509;
  assign new_n6218_ = ~new_n19027_ | ~new_n5250_;
  assign new_n6219_ = ~pi284 | ~new_n6198_;
  assign new_n6220_ = ~new_n1565_ | ~po509;
  assign new_n6221_ = ~new_n19028_ | ~new_n5250_;
  assign new_n6222_ = ~pi285 | ~new_n6198_;
  assign new_n6223_ = ~new_n1564_ | ~po509;
  assign new_n6224_ = ~new_n19029_ | ~new_n5250_;
  assign new_n6225_ = ~pi286 | ~new_n6198_;
  assign new_n6226_ = ~new_n1563_ | ~po509;
  assign new_n6227_ = ~new_n19106_ | ~new_n5250_;
  assign new_n6228_ = ~pi287 | ~new_n6198_;
  assign new_n6229_ = ~new_n1593_ | ~po509;
  assign new_n6230_ = ~new_n19013_ | ~new_n5250_;
  assign new_n6231_ = ~pi288 | ~new_n6198_;
  assign new_n6232_ = ~new_n1592_ | ~po509;
  assign new_n6233_ = ~new_n19014_ | ~new_n5250_;
  assign new_n6234_ = ~pi289 | ~new_n6198_;
  assign new_n6235_ = ~new_n1591_ | ~po509;
  assign new_n6236_ = ~new_n19015_ | ~new_n5250_;
  assign new_n6237_ = ~pi290 | ~new_n6198_;
  assign new_n6238_ = ~new_n1590_ | ~po509;
  assign new_n6239_ = ~new_n19134_ | ~new_n5250_;
  assign new_n6240_ = ~pi291 | ~new_n6198_;
  assign new_n6241_ = ~new_n1589_ | ~po509;
  assign new_n6242_ = ~new_n19016_ | ~new_n5250_;
  assign new_n6243_ = ~pi292 | ~new_n6198_;
  assign new_n6244_ = ~new_n1588_ | ~po509;
  assign new_n6245_ = ~new_n19017_ | ~new_n5250_;
  assign new_n6246_ = ~pi293 | ~new_n6198_;
  assign new_n6247_ = ~new_n1587_ | ~po509;
  assign new_n6248_ = ~new_n19018_ | ~new_n5250_;
  assign new_n6249_ = ~pi294 | ~new_n6198_;
  assign new_n6250_ = ~new_n1586_ | ~po509;
  assign new_n6251_ = ~new_n19132_ | ~new_n5250_;
  assign new_n6252_ = ~pi295 | ~new_n6198_;
  assign new_n6253_ = ~new_n1585_ | ~po509;
  assign new_n6254_ = ~new_n19019_ | ~new_n5250_;
  assign new_n6255_ = ~pi296 | ~new_n6198_;
  assign new_n6256_ = ~new_n1584_ | ~po509;
  assign new_n6257_ = ~new_n19130_ | ~new_n5250_;
  assign new_n6258_ = ~pi297 | ~new_n6198_;
  assign new_n6259_ = ~new_n1582_ | ~po509;
  assign new_n6260_ = ~new_n19126_ | ~new_n5250_;
  assign new_n6261_ = ~pi298 | ~new_n6198_;
  assign new_n6262_ = ~new_n1581_ | ~po509;
  assign new_n6263_ = ~new_n19123_ | ~new_n5250_;
  assign new_n6264_ = ~pi299 | ~new_n6198_;
  assign new_n6265_ = ~new_n1580_ | ~po509;
  assign new_n6266_ = ~new_n19121_ | ~new_n5250_;
  assign new_n6267_ = ~pi300 | ~new_n6198_;
  assign new_n6268_ = ~new_n1579_ | ~po509;
  assign new_n6269_ = ~new_n19020_ | ~new_n5250_;
  assign new_n6270_ = ~pi301 | ~new_n6198_;
  assign new_n6271_ = ~new_n1578_ | ~po509;
  assign new_n6272_ = ~new_n19021_ | ~new_n5250_;
  assign new_n6273_ = ~pi302 | ~new_n6198_;
  assign new_n6274_ = ~new_n1577_ | ~po509;
  assign new_n6275_ = ~new_n19119_ | ~new_n5250_;
  assign new_n6276_ = ~pi303 | ~new_n6198_;
  assign new_n6277_ = ~new_n1576_ | ~po509;
  assign new_n6278_ = ~new_n19022_ | ~new_n5250_;
  assign new_n6279_ = ~pi304 | ~new_n6198_;
  assign new_n6280_ = ~new_n1575_ | ~po509;
  assign new_n6281_ = ~new_n19117_ | ~new_n5250_;
  assign new_n6282_ = ~pi305 | ~new_n6198_;
  assign new_n6283_ = ~new_n1574_ | ~po509;
  assign new_n6284_ = ~new_n19114_ | ~new_n5250_;
  assign new_n6285_ = ~pi306 | ~new_n6198_;
  assign new_n6286_ = ~new_n1573_ | ~po509;
  assign new_n6287_ = ~new_n19023_ | ~new_n5250_;
  assign new_n6288_ = ~pi307 | ~new_n6198_;
  assign new_n6289_ = ~new_n1571_ | ~po509;
  assign new_n6290_ = ~new_n19111_ | ~new_n5250_;
  assign new_n6291_ = ~pi308 | ~new_n6198_;
  assign new_n6292_ = ~new_n1570_ | ~po509;
  assign new_n6293_ = ~new_n19050_ | ~new_n5250_;
  assign new_n6294_ = ~pi309 | ~new_n6198_;
  assign new_n6295_ = ~new_n6195_ | ~new_n7875_;
  assign new_n6296_ = ~new_n5553_;
  assign new_n6297_ = ~new_n5552_ | ~new_n7866_;
  assign new_n6298_ = ~new_n5552_ | ~new_n7869_;
  assign new_n6299_ = ~new_n6296_ | ~pi320;
  assign new_n6300_ = ~new_n6296_ | ~pi321;
  assign new_n6301_ = ~new_n6296_ | ~pi322;
  assign new_n6302_ = ~new_n6296_ | ~pi323;
  assign new_n6303_ = ~new_n6296_ | ~pi324;
  assign new_n6304_ = ~new_n6296_ | ~pi325;
  assign new_n6305_ = ~new_n6296_ | ~pi326;
  assign new_n6306_ = ~new_n6296_ | ~pi327;
  assign new_n6307_ = ~new_n6296_ | ~pi328;
  assign new_n6308_ = ~new_n6296_ | ~pi329;
  assign new_n6309_ = ~new_n6296_ | ~pi330;
  assign new_n6310_ = ~new_n6296_ | ~pi331;
  assign new_n6311_ = ~new_n6296_ | ~pi332;
  assign new_n6312_ = ~new_n6296_ | ~pi333;
  assign new_n6313_ = ~new_n6296_ | ~pi334;
  assign new_n6314_ = ~new_n6296_ | ~pi335;
  assign new_n6315_ = ~new_n6296_ | ~pi336;
  assign new_n6316_ = ~new_n6296_ | ~pi337;
  assign new_n6317_ = ~new_n6296_ | ~pi338;
  assign new_n6318_ = ~new_n6296_ | ~pi339;
  assign new_n6319_ = ~new_n6296_ | ~pi312;
  assign new_n6320_ = ~new_n6296_ | ~pi340;
  assign new_n6321_ = ~new_n6296_ | ~pi341;
  assign new_n6322_ = ~new_n6296_ | ~pi313;
  assign new_n6323_ = ~new_n6296_ | ~pi314;
  assign new_n6324_ = ~new_n6296_ | ~pi315;
  assign new_n6325_ = ~new_n6296_ | ~pi316;
  assign new_n6326_ = ~new_n6296_ | ~pi317;
  assign new_n6327_ = ~new_n6296_ | ~pi318;
  assign new_n6328_ = ~new_n6296_ | ~pi319;
  assign new_n6329_ = ~new_n7894_ | ~new_n7891_;
  assign new_n6330_ = ~new_n5560_ | ~new_n7913_ | ~new_n7912_;
  assign new_n6331_ = ~new_n5240_ | ~pi407;
  assign new_n6332_ = ~new_n5241_ | ~pi375;
  assign new_n6333_ = ~new_n5242_ | ~pi343;
  assign new_n6334_ = ~pi510 | ~new_n5239_;
  assign new_n6335_ = ~new_n5300_;
  assign new_n6336_ = ~new_n5610_ | ~new_n6154_;
  assign new_n6337_ = ~new_n6151_ | ~new_n23314_;
  assign new_n6338_ = ~new_n6150_ | ~new_n24260_;
  assign new_n6339_ = ~new_n6146_ | ~new_n22890_;
  assign new_n6340_ = ~new_n6161_ | ~new_n20217_;
  assign new_n6341_ = ~new_n6163_ | ~new_n23787_;
  assign new_n6342_ = ~new_n5234_ | ~new_n21268_;
  assign new_n6343_ = ~new_n6142_ | ~new_n21769_;
  assign new_n6344_ = ~new_n5568_;
  assign new_n6345_ = ~new_n5647_ | ~new_n5247_;
  assign new_n6346_ = ~new_n5246_ | ~new_n5300_;
  assign new_n6347_ = ~new_n20768_ | ~new_n5245_;
  assign new_n6348_ = ~new_n5647_ | ~new_n6336_;
  assign new_n6349_ = ~new_n6346_ | ~new_n6344_ | ~new_n5785_ | ~new_n6348_;
  assign new_n6350_ = ~pi408 | ~new_n5240_;
  assign new_n6351_ = ~pi376 | ~new_n5241_;
  assign new_n6352_ = ~pi344 | ~new_n5242_;
  assign new_n6353_ = ~pi495 | ~new_n5239_;
  assign new_n6354_ = ~new_n5290_;
  assign new_n6355_ = ~pi406 | ~new_n5240_;
  assign new_n6356_ = ~pi374 | ~new_n5241_;
  assign new_n6357_ = ~pi342 | ~new_n5242_;
  assign new_n6358_ = ~pi500 | ~new_n5239_;
  assign new_n6359_ = ~new_n5299_;
  assign new_n6360_ = ~new_n5255_ | ~new_n5299_;
  assign new_n6361_ = ~new_n23391_ | ~new_n6151_;
  assign new_n6362_ = ~new_n24337_ | ~new_n6150_;
  assign new_n6363_ = ~new_n22889_ | ~new_n6146_;
  assign new_n6364_ = ~new_n20294_ | ~new_n6161_;
  assign new_n6365_ = ~new_n23864_ | ~new_n6163_;
  assign new_n6366_ = ~new_n21267_ | ~new_n5234_;
  assign new_n6367_ = ~new_n21768_ | ~new_n6142_;
  assign new_n6368_ = ~new_n5569_;
  assign new_n6369_ = ~new_n20098_ | ~new_n5247_;
  assign new_n6370_ = ~new_n5246_ | ~new_n5290_;
  assign new_n6371_ = ~new_n20767_ | ~new_n5245_;
  assign new_n6372_ = ~new_n5652_ | ~new_n6336_;
  assign new_n6373_ = ~new_n5801_ | ~new_n6368_;
  assign new_n6374_ = ~pi409 | ~new_n5240_;
  assign new_n6375_ = ~pi377 | ~new_n5241_;
  assign new_n6376_ = ~pi345 | ~new_n5242_;
  assign new_n6377_ = ~new_n18859_ | ~new_n5239_;
  assign new_n6378_ = ~new_n5286_;
  assign new_n6379_ = ~new_n5255_ | ~new_n5300_;
  assign new_n6380_ = ~new_n23401_ | ~new_n6151_;
  assign new_n6381_ = ~new_n24347_ | ~new_n6150_;
  assign new_n6382_ = ~new_n22811_ | ~new_n6146_;
  assign new_n6383_ = ~new_n20304_ | ~new_n6161_;
  assign new_n6384_ = ~new_n23874_ | ~new_n6163_;
  assign new_n6385_ = ~new_n21189_ | ~new_n5234_;
  assign new_n6386_ = ~new_n21690_ | ~new_n6142_;
  assign new_n6387_ = ~new_n5570_;
  assign new_n6388_ = ~new_n20061_ | ~new_n5247_;
  assign new_n6389_ = ~new_n5246_ | ~new_n5286_;
  assign new_n6390_ = ~new_n20689_ | ~new_n5245_;
  assign new_n6391_ = ~new_n5655_ | ~new_n6336_;
  assign new_n6392_ = ~new_n5805_ | ~new_n6387_;
  assign new_n6393_ = ~pi410 | ~new_n5240_;
  assign new_n6394_ = ~pi378 | ~new_n5241_;
  assign new_n6395_ = ~pi346 | ~new_n5242_;
  assign new_n6396_ = ~new_n18910_ | ~new_n5239_;
  assign new_n6397_ = ~new_n5282_;
  assign new_n6398_ = ~new_n5255_ | ~new_n5290_;
  assign new_n6399_ = ~new_n23311_ | ~new_n6151_;
  assign new_n6400_ = ~new_n24257_ | ~new_n6150_;
  assign new_n6401_ = ~new_n22895_ | ~new_n6146_;
  assign new_n6402_ = ~new_n20214_ | ~new_n6161_;
  assign new_n6403_ = ~new_n23784_ | ~new_n6163_;
  assign new_n6404_ = ~new_n21273_ | ~new_n5234_;
  assign new_n6405_ = ~new_n21774_ | ~new_n6142_;
  assign new_n6406_ = ~new_n5571_;
  assign new_n6407_ = ~new_n20063_ | ~new_n5247_;
  assign new_n6408_ = ~new_n5246_ | ~new_n5282_;
  assign new_n6409_ = ~new_n20773_ | ~new_n5245_;
  assign new_n6410_ = ~new_n5658_ | ~new_n6336_;
  assign new_n6411_ = ~new_n5809_ | ~new_n6406_;
  assign new_n6412_ = ~pi411 | ~new_n5240_;
  assign new_n6413_ = ~pi379 | ~new_n5241_;
  assign new_n6414_ = ~pi347 | ~new_n5242_;
  assign new_n6415_ = ~new_n18909_ | ~new_n5239_;
  assign new_n6416_ = ~new_n5289_;
  assign new_n6417_ = ~new_n5255_ | ~new_n5286_;
  assign new_n6418_ = ~new_n23400_ | ~new_n6151_;
  assign new_n6419_ = ~new_n24346_ | ~new_n6150_;
  assign new_n6420_ = ~new_n22894_ | ~new_n6146_;
  assign new_n6421_ = ~new_n20303_ | ~new_n6161_;
  assign new_n6422_ = ~new_n23873_ | ~new_n6163_;
  assign new_n6423_ = ~new_n21272_ | ~new_n5234_;
  assign new_n6424_ = ~new_n21773_ | ~new_n6142_;
  assign new_n6425_ = ~new_n5572_;
  assign new_n6426_ = ~new_n20064_ | ~new_n5247_;
  assign new_n6427_ = ~new_n5246_ | ~new_n5289_;
  assign new_n6428_ = ~new_n20772_ | ~new_n5245_;
  assign new_n6429_ = ~new_n5661_ | ~new_n6336_;
  assign new_n6430_ = ~new_n5813_ | ~new_n6425_;
  assign new_n6431_ = ~pi412 | ~new_n5240_;
  assign new_n6432_ = ~pi380 | ~new_n5241_;
  assign new_n6433_ = ~pi348 | ~new_n5242_;
  assign new_n6434_ = ~new_n18908_ | ~new_n5239_;
  assign new_n6435_ = ~new_n5293_;
  assign new_n6436_ = ~new_n5255_ | ~new_n5282_;
  assign new_n6437_ = ~new_n23399_ | ~new_n6151_;
  assign new_n6438_ = ~new_n24345_ | ~new_n6150_;
  assign new_n6439_ = ~new_n22812_ | ~new_n6146_;
  assign new_n6440_ = ~new_n20302_ | ~new_n6161_;
  assign new_n6441_ = ~new_n23872_ | ~new_n6163_;
  assign new_n6442_ = ~new_n21190_ | ~new_n5234_;
  assign new_n6443_ = ~new_n21691_ | ~new_n6142_;
  assign new_n6444_ = ~new_n5573_;
  assign new_n6445_ = ~new_n20108_ | ~new_n5247_;
  assign new_n6446_ = ~new_n5246_ | ~new_n5293_;
  assign new_n6447_ = ~new_n20690_ | ~new_n5245_;
  assign new_n6448_ = ~new_n5664_ | ~new_n6336_;
  assign new_n6449_ = ~new_n5817_ | ~new_n6444_;
  assign new_n6450_ = ~pi413 | ~new_n5240_;
  assign new_n6451_ = ~pi381 | ~new_n5241_;
  assign new_n6452_ = ~pi349 | ~new_n5242_;
  assign new_n6453_ = ~new_n18907_ | ~new_n5239_;
  assign new_n6454_ = ~new_n5292_;
  assign new_n6455_ = ~new_n5255_ | ~new_n5289_;
  assign new_n6456_ = ~new_n23312_ | ~new_n6151_;
  assign new_n6457_ = ~new_n24258_ | ~new_n6150_;
  assign new_n6458_ = ~new_n22893_ | ~new_n6146_;
  assign new_n6459_ = ~new_n20215_ | ~new_n6161_;
  assign new_n6460_ = ~new_n23785_ | ~new_n6163_;
  assign new_n6461_ = ~new_n21271_ | ~new_n5234_;
  assign new_n6462_ = ~new_n21772_ | ~new_n6142_;
  assign new_n6463_ = ~new_n5574_;
  assign new_n6464_ = ~new_n20065_ | ~new_n5247_;
  assign new_n6465_ = ~new_n5246_ | ~new_n5292_;
  assign new_n6466_ = ~new_n20771_ | ~new_n5245_;
  assign new_n6467_ = ~new_n5667_ | ~new_n6336_;
  assign new_n6468_ = ~new_n5821_ | ~new_n6463_;
  assign new_n6469_ = ~pi414 | ~new_n5240_;
  assign new_n6470_ = ~pi382 | ~new_n5241_;
  assign new_n6471_ = ~pi350 | ~new_n5242_;
  assign new_n6472_ = ~new_n18906_ | ~new_n5239_;
  assign new_n6473_ = ~new_n5306_;
  assign new_n6474_ = ~new_n5255_ | ~new_n5293_;
  assign new_n6475_ = ~new_n23398_ | ~new_n6151_;
  assign new_n6476_ = ~new_n24344_ | ~new_n6150_;
  assign new_n6477_ = ~new_n22813_ | ~new_n6146_;
  assign new_n6478_ = ~new_n20301_ | ~new_n6161_;
  assign new_n6479_ = ~new_n23871_ | ~new_n6163_;
  assign new_n6480_ = ~new_n21191_ | ~new_n5234_;
  assign new_n6481_ = ~new_n21692_ | ~new_n6142_;
  assign new_n6482_ = ~new_n5575_;
  assign new_n6483_ = ~new_n20066_ | ~new_n5247_;
  assign new_n6484_ = ~new_n5246_ | ~new_n5306_;
  assign new_n6485_ = ~new_n20691_ | ~new_n5245_;
  assign new_n6486_ = ~new_n5670_ | ~new_n6336_;
  assign new_n6487_ = ~new_n5825_ | ~new_n6482_;
  assign new_n6488_ = ~pi415 | ~new_n5240_;
  assign new_n6489_ = ~pi383 | ~new_n5241_;
  assign new_n6490_ = ~pi351 | ~new_n5242_;
  assign new_n6491_ = ~new_n18905_ | ~new_n5239_;
  assign new_n6492_ = ~new_n5305_;
  assign new_n6493_ = ~new_n5255_ | ~new_n5292_;
  assign new_n6494_ = ~new_n23313_ | ~new_n6151_;
  assign new_n6495_ = ~new_n24259_ | ~new_n6150_;
  assign new_n6496_ = ~new_n22892_ | ~new_n6146_;
  assign new_n6497_ = ~new_n20216_ | ~new_n6161_;
  assign new_n6498_ = ~new_n23786_ | ~new_n6163_;
  assign new_n6499_ = ~new_n21270_ | ~new_n5234_;
  assign new_n6500_ = ~new_n21771_ | ~new_n6142_;
  assign new_n6501_ = ~new_n5576_;
  assign new_n6502_ = ~new_n20067_ | ~new_n5247_;
  assign new_n6503_ = ~new_n5246_ | ~new_n5305_;
  assign new_n6504_ = ~new_n20770_ | ~new_n5245_;
  assign new_n6505_ = ~new_n5673_ | ~new_n6336_;
  assign new_n6506_ = ~new_n5829_ | ~new_n6501_;
  assign new_n6507_ = ~pi416 | ~new_n5240_;
  assign new_n6508_ = ~pi384 | ~new_n5241_;
  assign new_n6509_ = ~pi352 | ~new_n5242_;
  assign new_n6510_ = ~new_n18929_ | ~new_n5239_;
  assign new_n6511_ = ~new_n5284_;
  assign new_n6512_ = ~new_n5255_ | ~new_n5306_;
  assign new_n6513_ = ~new_n23397_ | ~new_n6151_;
  assign new_n6514_ = ~new_n24343_ | ~new_n6150_;
  assign new_n6515_ = ~new_n22891_ | ~new_n6146_;
  assign new_n6516_ = ~new_n20300_ | ~new_n6161_;
  assign new_n6517_ = ~new_n23870_ | ~new_n6163_;
  assign new_n6518_ = ~new_n21269_ | ~new_n5234_;
  assign new_n6519_ = ~new_n21770_ | ~new_n6142_;
  assign new_n6520_ = ~new_n5577_;
  assign new_n6521_ = ~new_n20106_ | ~new_n5247_;
  assign new_n6522_ = ~new_n5246_ | ~new_n5284_;
  assign new_n6523_ = ~new_n20769_ | ~new_n5245_;
  assign new_n6524_ = ~new_n5676_ | ~new_n6336_;
  assign new_n6525_ = ~new_n5833_ | ~new_n6520_;
  assign new_n6526_ = ~pi417 | ~new_n5240_;
  assign new_n6527_ = ~pi385 | ~new_n5241_;
  assign new_n6528_ = ~pi353 | ~new_n5242_;
  assign new_n6529_ = ~new_n18928_ | ~new_n5239_;
  assign new_n6530_ = ~new_n5285_;
  assign new_n6531_ = ~new_n5255_ | ~new_n5305_;
  assign new_n6532_ = ~new_n23407_ | ~new_n6151_;
  assign new_n6533_ = ~new_n24353_ | ~new_n6150_;
  assign new_n6534_ = ~new_n22805_ | ~new_n6146_;
  assign new_n6535_ = ~new_n20310_ | ~new_n6161_;
  assign new_n6536_ = ~new_n23880_ | ~new_n6163_;
  assign new_n6537_ = ~new_n21183_ | ~new_n5234_;
  assign new_n6538_ = ~new_n21684_ | ~new_n6142_;
  assign new_n6539_ = ~new_n5578_;
  assign new_n6540_ = ~new_n20049_ | ~new_n5247_;
  assign new_n6541_ = ~new_n5246_ | ~new_n5285_;
  assign new_n6542_ = ~new_n20683_ | ~new_n5245_;
  assign new_n6543_ = ~new_n5679_ | ~new_n6336_;
  assign new_n6544_ = ~new_n5837_ | ~new_n6539_;
  assign new_n6545_ = ~pi418 | ~new_n5240_;
  assign new_n6546_ = ~pi386 | ~new_n5241_;
  assign new_n6547_ = ~pi354 | ~new_n5242_;
  assign new_n6548_ = ~new_n18927_ | ~new_n5239_;
  assign new_n6549_ = ~new_n5294_;
  assign new_n6550_ = ~new_n5255_ | ~new_n5284_;
  assign new_n6551_ = ~new_n23306_ | ~new_n6151_;
  assign new_n6552_ = ~new_n24252_ | ~new_n6150_;
  assign new_n6553_ = ~new_n22909_ | ~new_n6146_;
  assign new_n6554_ = ~new_n20209_ | ~new_n6161_;
  assign new_n6555_ = ~new_n23779_ | ~new_n6163_;
  assign new_n6556_ = ~new_n21287_ | ~new_n5234_;
  assign new_n6557_ = ~new_n21788_ | ~new_n6142_;
  assign new_n6558_ = ~new_n5579_;
  assign new_n6559_ = ~new_n20050_ | ~new_n5247_;
  assign new_n6560_ = ~new_n5246_ | ~new_n5294_;
  assign new_n6561_ = ~new_n20787_ | ~new_n5245_;
  assign new_n6562_ = ~new_n5682_ | ~new_n6336_;
  assign new_n6563_ = ~new_n5841_ | ~new_n6558_;
  assign new_n6564_ = ~pi419 | ~new_n5240_;
  assign new_n6565_ = ~pi387 | ~new_n5241_;
  assign new_n6566_ = ~pi355 | ~new_n5242_;
  assign new_n6567_ = ~new_n18926_ | ~new_n5239_;
  assign new_n6568_ = ~new_n5302_;
  assign new_n6569_ = ~new_n5255_ | ~new_n5285_;
  assign new_n6570_ = ~new_n23396_ | ~new_n6151_;
  assign new_n6571_ = ~new_n24342_ | ~new_n6150_;
  assign new_n6572_ = ~new_n22908_ | ~new_n6146_;
  assign new_n6573_ = ~new_n20299_ | ~new_n6161_;
  assign new_n6574_ = ~new_n23869_ | ~new_n6163_;
  assign new_n6575_ = ~new_n21286_ | ~new_n5234_;
  assign new_n6576_ = ~new_n21787_ | ~new_n6142_;
  assign new_n6577_ = ~new_n5580_;
  assign new_n6578_ = ~new_n20051_ | ~new_n5247_;
  assign new_n6579_ = ~new_n5246_ | ~new_n5302_;
  assign new_n6580_ = ~new_n20786_ | ~new_n5245_;
  assign new_n6581_ = ~new_n5685_ | ~new_n6336_;
  assign new_n6582_ = ~new_n5845_ | ~new_n6577_;
  assign new_n6583_ = ~pi420 | ~new_n5240_;
  assign new_n6584_ = ~pi388 | ~new_n5241_;
  assign new_n6585_ = ~pi356 | ~new_n5242_;
  assign new_n6586_ = ~new_n18925_ | ~new_n5239_;
  assign new_n6587_ = ~new_n5301_;
  assign new_n6588_ = ~new_n5255_ | ~new_n5294_;
  assign new_n6589_ = ~new_n23395_ | ~new_n6151_;
  assign new_n6590_ = ~new_n24341_ | ~new_n6150_;
  assign new_n6591_ = ~new_n22806_ | ~new_n6146_;
  assign new_n6592_ = ~new_n20298_ | ~new_n6161_;
  assign new_n6593_ = ~new_n23868_ | ~new_n6163_;
  assign new_n6594_ = ~new_n21184_ | ~new_n5234_;
  assign new_n6595_ = ~new_n21685_ | ~new_n6142_;
  assign new_n6596_ = ~new_n5581_;
  assign new_n6597_ = ~new_n20129_ | ~new_n5247_;
  assign new_n6598_ = ~new_n5246_ | ~new_n5301_;
  assign new_n6599_ = ~new_n20684_ | ~new_n5245_;
  assign new_n6600_ = ~new_n5688_ | ~new_n6336_;
  assign new_n6601_ = ~new_n5849_ | ~new_n6596_;
  assign new_n6602_ = ~pi421 | ~new_n5240_;
  assign new_n6603_ = ~pi389 | ~new_n5241_;
  assign new_n6604_ = ~pi357 | ~new_n5242_;
  assign new_n6605_ = ~new_n18924_ | ~new_n5239_;
  assign new_n6606_ = ~new_n5296_;
  assign new_n6607_ = ~new_n5255_ | ~new_n5302_;
  assign new_n6608_ = ~new_n23406_ | ~new_n6151_;
  assign new_n6609_ = ~new_n24352_ | ~new_n6150_;
  assign new_n6610_ = ~new_n22907_ | ~new_n6146_;
  assign new_n6611_ = ~new_n20309_ | ~new_n6161_;
  assign new_n6612_ = ~new_n23879_ | ~new_n6163_;
  assign new_n6613_ = ~new_n21285_ | ~new_n5234_;
  assign new_n6614_ = ~new_n21786_ | ~new_n6142_;
  assign new_n6615_ = ~new_n5582_;
  assign new_n6616_ = ~new_n20052_ | ~new_n5247_;
  assign new_n6617_ = ~new_n5246_ | ~new_n5296_;
  assign new_n6618_ = ~new_n20785_ | ~new_n5245_;
  assign new_n6619_ = ~new_n5691_ | ~new_n6336_;
  assign new_n6620_ = ~new_n5853_ | ~new_n6615_;
  assign new_n6621_ = ~pi422 | ~new_n5240_;
  assign new_n6622_ = ~pi390 | ~new_n5241_;
  assign new_n6623_ = ~pi358 | ~new_n5242_;
  assign new_n6624_ = ~new_n18923_ | ~new_n5239_;
  assign new_n6625_ = ~new_n5295_;
  assign new_n6626_ = ~new_n5255_ | ~new_n5301_;
  assign new_n6627_ = ~new_n23405_ | ~new_n6151_;
  assign new_n6628_ = ~new_n24351_ | ~new_n6150_;
  assign new_n6629_ = ~new_n22906_ | ~new_n6146_;
  assign new_n6630_ = ~new_n20308_ | ~new_n6161_;
  assign new_n6631_ = ~new_n23878_ | ~new_n6163_;
  assign new_n6632_ = ~new_n21284_ | ~new_n5234_;
  assign new_n6633_ = ~new_n21785_ | ~new_n6142_;
  assign new_n6634_ = ~new_n5583_;
  assign new_n6635_ = ~new_n20053_ | ~new_n5247_;
  assign new_n6636_ = ~new_n5246_ | ~new_n5295_;
  assign new_n6637_ = ~new_n20784_ | ~new_n5245_;
  assign new_n6638_ = ~new_n5694_ | ~new_n6336_;
  assign new_n6639_ = ~new_n5857_ | ~new_n6634_;
  assign new_n6640_ = ~pi423 | ~new_n5240_;
  assign new_n6641_ = ~pi391 | ~new_n5241_;
  assign new_n6642_ = ~pi359 | ~new_n5242_;
  assign new_n6643_ = ~new_n18922_ | ~new_n5239_;
  assign new_n6644_ = ~new_n5291_;
  assign new_n6645_ = ~new_n5255_ | ~new_n5296_;
  assign new_n6646_ = ~new_n23307_ | ~new_n6151_;
  assign new_n6647_ = ~new_n24253_ | ~new_n6150_;
  assign new_n6648_ = ~new_n22905_ | ~new_n6146_;
  assign new_n6649_ = ~new_n20210_ | ~new_n6161_;
  assign new_n6650_ = ~new_n23780_ | ~new_n6163_;
  assign new_n6651_ = ~new_n21283_ | ~new_n5234_;
  assign new_n6652_ = ~new_n21784_ | ~new_n6142_;
  assign new_n6653_ = ~new_n5584_;
  assign new_n6654_ = ~new_n20054_ | ~new_n5247_;
  assign new_n6655_ = ~new_n5246_ | ~new_n5291_;
  assign new_n6656_ = ~new_n20783_ | ~new_n5245_;
  assign new_n6657_ = ~new_n5697_ | ~new_n6336_;
  assign new_n6658_ = ~new_n5861_ | ~new_n6653_;
  assign new_n6659_ = ~pi424 | ~new_n5240_;
  assign new_n6660_ = ~pi392 | ~new_n5241_;
  assign new_n6661_ = ~pi360 | ~new_n5242_;
  assign new_n6662_ = ~new_n18921_ | ~new_n5239_;
  assign new_n6663_ = ~new_n5304_;
  assign new_n6664_ = ~new_n5255_ | ~new_n5295_;
  assign new_n6665_ = ~new_n23394_ | ~new_n6151_;
  assign new_n6666_ = ~new_n24340_ | ~new_n6150_;
  assign new_n6667_ = ~new_n22807_ | ~new_n6146_;
  assign new_n6668_ = ~new_n20297_ | ~new_n6161_;
  assign new_n6669_ = ~new_n23867_ | ~new_n6163_;
  assign new_n6670_ = ~new_n21185_ | ~new_n5234_;
  assign new_n6671_ = ~new_n21686_ | ~new_n6142_;
  assign new_n6672_ = ~new_n5585_;
  assign new_n6673_ = ~new_n20127_ | ~new_n5247_;
  assign new_n6674_ = ~new_n5246_ | ~new_n5304_;
  assign new_n6675_ = ~new_n20685_ | ~new_n5245_;
  assign new_n6676_ = ~new_n5700_ | ~new_n6336_;
  assign new_n6677_ = ~new_n5865_ | ~new_n6672_;
  assign new_n6678_ = ~pi425 | ~new_n5240_;
  assign new_n6679_ = ~pi393 | ~new_n5241_;
  assign new_n6680_ = ~pi361 | ~new_n5242_;
  assign new_n6681_ = ~new_n18920_ | ~new_n5239_;
  assign new_n6682_ = ~new_n5303_;
  assign new_n6683_ = ~new_n5255_ | ~new_n5291_;
  assign new_n6684_ = ~new_n23393_ | ~new_n6151_;
  assign new_n6685_ = ~new_n24339_ | ~new_n6150_;
  assign new_n6686_ = ~new_n22904_ | ~new_n6146_;
  assign new_n6687_ = ~new_n20296_ | ~new_n6161_;
  assign new_n6688_ = ~new_n23866_ | ~new_n6163_;
  assign new_n6689_ = ~new_n21282_ | ~new_n5234_;
  assign new_n6690_ = ~new_n21783_ | ~new_n6142_;
  assign new_n6691_ = ~new_n5586_;
  assign new_n6692_ = ~new_n20055_ | ~new_n5247_;
  assign new_n6693_ = ~new_n5246_ | ~new_n5303_;
  assign new_n6694_ = ~new_n20782_ | ~new_n5245_;
  assign new_n6695_ = ~new_n5703_ | ~new_n6336_;
  assign new_n6696_ = ~new_n5869_ | ~new_n6691_;
  assign new_n6697_ = ~pi426 | ~new_n5240_;
  assign new_n6698_ = ~pi394 | ~new_n5241_;
  assign new_n6699_ = ~pi362 | ~new_n5242_;
  assign new_n6700_ = ~new_n18919_ | ~new_n5239_;
  assign new_n6701_ = ~new_n5298_;
  assign new_n6702_ = ~new_n5255_ | ~new_n5304_;
  assign new_n6703_ = ~new_n23392_ | ~new_n6151_;
  assign new_n6704_ = ~new_n24338_ | ~new_n6150_;
  assign new_n6705_ = ~new_n22903_ | ~new_n6146_;
  assign new_n6706_ = ~new_n20295_ | ~new_n6161_;
  assign new_n6707_ = ~new_n23865_ | ~new_n6163_;
  assign new_n6708_ = ~new_n21281_ | ~new_n5234_;
  assign new_n6709_ = ~new_n21782_ | ~new_n6142_;
  assign new_n6710_ = ~new_n5587_;
  assign new_n6711_ = ~new_n20125_ | ~new_n5247_;
  assign new_n6712_ = ~new_n5246_ | ~new_n5298_;
  assign new_n6713_ = ~new_n20781_ | ~new_n5245_;
  assign new_n6714_ = ~new_n5705_ | ~new_n6336_;
  assign new_n6715_ = ~new_n5873_ | ~new_n6710_;
  assign new_n6716_ = ~pi427 | ~new_n5240_;
  assign new_n6717_ = ~pi395 | ~new_n5241_;
  assign new_n6718_ = ~pi363 | ~new_n5242_;
  assign new_n6719_ = ~new_n18918_ | ~new_n5239_;
  assign new_n6720_ = ~new_n5297_;
  assign new_n6721_ = ~new_n5255_ | ~new_n5303_;
  assign new_n6722_ = ~new_n23390_ | ~new_n6151_;
  assign new_n6723_ = ~new_n24336_ | ~new_n6150_;
  assign new_n6724_ = ~new_n22808_ | ~new_n6146_;
  assign new_n6725_ = ~new_n20293_ | ~new_n6161_;
  assign new_n6726_ = ~new_n23863_ | ~new_n6163_;
  assign new_n6727_ = ~new_n21186_ | ~new_n5234_;
  assign new_n6728_ = ~new_n21687_ | ~new_n6142_;
  assign new_n6729_ = ~new_n5589_;
  assign new_n6730_ = ~new_n20056_ | ~new_n5247_;
  assign new_n6731_ = ~new_n5246_ | ~new_n5297_;
  assign new_n6732_ = ~new_n20686_ | ~new_n5245_;
  assign new_n6733_ = ~new_n6177_ | ~new_n6336_;
  assign new_n6734_ = ~new_n5877_ | ~new_n6729_;
  assign new_n6735_ = ~pi428 | ~new_n5240_;
  assign new_n6736_ = ~pi396 | ~new_n5241_;
  assign new_n6737_ = ~pi364 | ~new_n5242_;
  assign new_n6738_ = ~new_n18917_ | ~new_n5239_;
  assign new_n6739_ = ~new_n5283_;
  assign new_n6740_ = ~new_n5255_ | ~new_n5298_;
  assign new_n6741_ = ~new_n23404_ | ~new_n6151_;
  assign new_n6742_ = ~new_n24350_ | ~new_n6150_;
  assign new_n6743_ = ~new_n22809_ | ~new_n6146_;
  assign new_n6744_ = ~new_n20307_ | ~new_n6161_;
  assign new_n6745_ = ~new_n23877_ | ~new_n6163_;
  assign new_n6746_ = ~new_n21187_ | ~new_n5234_;
  assign new_n6747_ = ~new_n21688_ | ~new_n6142_;
  assign new_n6748_ = ~new_n5591_;
  assign new_n6749_ = ~new_n20121_ | ~new_n5247_;
  assign new_n6750_ = ~new_n5246_ | ~new_n5283_;
  assign new_n6751_ = ~new_n20687_ | ~new_n5245_;
  assign new_n6752_ = ~new_n6176_ | ~new_n6336_;
  assign new_n6753_ = ~new_n5881_ | ~new_n6748_;
  assign new_n6754_ = ~pi429 | ~new_n5240_;
  assign new_n6755_ = ~pi397 | ~new_n5241_;
  assign new_n6756_ = ~pi365 | ~new_n5242_;
  assign new_n6757_ = ~new_n18916_ | ~new_n5239_;
  assign new_n6758_ = ~new_n5288_;
  assign new_n6759_ = ~new_n5255_ | ~new_n5297_;
  assign new_n6760_ = ~new_n23403_ | ~new_n6151_;
  assign new_n6761_ = ~new_n24349_ | ~new_n6150_;
  assign new_n6762_ = ~new_n22902_ | ~new_n6146_;
  assign new_n6763_ = ~new_n20306_ | ~new_n6161_;
  assign new_n6764_ = ~new_n23876_ | ~new_n6163_;
  assign new_n6765_ = ~new_n21280_ | ~new_n5234_;
  assign new_n6766_ = ~new_n21781_ | ~new_n6142_;
  assign new_n6767_ = ~new_n5593_;
  assign new_n6768_ = ~new_n20057_ | ~new_n5247_;
  assign new_n6769_ = ~new_n5246_ | ~new_n5288_;
  assign new_n6770_ = ~new_n20780_ | ~new_n5245_;
  assign new_n6771_ = ~new_n6175_ | ~new_n6336_;
  assign new_n6772_ = ~new_n5885_ | ~new_n6767_;
  assign new_n6773_ = ~pi430 | ~new_n5240_;
  assign new_n6774_ = ~pi398 | ~new_n5241_;
  assign new_n6775_ = ~pi366 | ~new_n5242_;
  assign new_n6776_ = ~new_n18915_ | ~new_n5239_;
  assign new_n6777_ = ~new_n5287_;
  assign new_n6778_ = ~new_n5255_ | ~new_n5283_;
  assign new_n6779_ = ~new_n23308_ | ~new_n6151_;
  assign new_n6780_ = ~new_n24254_ | ~new_n6150_;
  assign new_n6781_ = ~new_n22901_ | ~new_n6146_;
  assign new_n6782_ = ~new_n20211_ | ~new_n6161_;
  assign new_n6783_ = ~new_n23781_ | ~new_n6163_;
  assign new_n6784_ = ~new_n21279_ | ~new_n5234_;
  assign new_n6785_ = ~new_n21780_ | ~new_n6142_;
  assign new_n6786_ = ~new_n5595_;
  assign new_n6787_ = ~new_n20119_ | ~new_n5247_;
  assign new_n6788_ = ~new_n5246_ | ~new_n5287_;
  assign new_n6789_ = ~new_n20779_ | ~new_n5245_;
  assign new_n6790_ = ~new_n6174_ | ~new_n6336_;
  assign new_n6791_ = ~new_n5889_ | ~new_n6786_;
  assign new_n6792_ = ~pi431 | ~new_n5240_;
  assign new_n6793_ = ~pi399 | ~new_n5241_;
  assign new_n6794_ = ~pi367 | ~new_n5242_;
  assign new_n6795_ = ~new_n18914_ | ~new_n5239_;
  assign new_n6796_ = ~new_n5280_;
  assign new_n6797_ = ~new_n5255_ | ~new_n5288_;
  assign new_n6798_ = ~new_n23389_ | ~new_n6151_;
  assign new_n6799_ = ~new_n24335_ | ~new_n6150_;
  assign new_n6800_ = ~new_n22900_ | ~new_n6146_;
  assign new_n6801_ = ~new_n20292_ | ~new_n6161_;
  assign new_n6802_ = ~new_n23862_ | ~new_n6163_;
  assign new_n6803_ = ~new_n21278_ | ~new_n5234_;
  assign new_n6804_ = ~new_n21779_ | ~new_n6142_;
  assign new_n6805_ = ~new_n5597_;
  assign new_n6806_ = ~new_n20058_ | ~new_n5247_;
  assign new_n6807_ = ~new_n5246_ | ~new_n5280_;
  assign new_n6808_ = ~new_n20778_ | ~new_n5245_;
  assign new_n6809_ = ~new_n6173_ | ~new_n6336_;
  assign new_n6810_ = ~new_n5893_ | ~new_n6805_;
  assign new_n6811_ = ~pi432 | ~new_n5240_;
  assign new_n6812_ = ~pi400 | ~new_n5241_;
  assign new_n6813_ = ~pi368 | ~new_n5242_;
  assign new_n6814_ = ~new_n18913_ | ~new_n5239_;
  assign new_n6815_ = ~new_n5279_;
  assign new_n6816_ = ~new_n5255_ | ~new_n5287_;
  assign new_n6817_ = ~new_n23388_ | ~new_n6151_;
  assign new_n6818_ = ~new_n24334_ | ~new_n6150_;
  assign new_n6819_ = ~new_n22899_ | ~new_n6146_;
  assign new_n6820_ = ~new_n20291_ | ~new_n6161_;
  assign new_n6821_ = ~new_n23861_ | ~new_n6163_;
  assign new_n6822_ = ~new_n21277_ | ~new_n5234_;
  assign new_n6823_ = ~new_n21778_ | ~new_n6142_;
  assign new_n6824_ = ~new_n5599_;
  assign new_n6825_ = ~new_n20117_ | ~new_n5247_;
  assign new_n6826_ = ~new_n5246_ | ~new_n5279_;
  assign new_n6827_ = ~new_n20777_ | ~new_n5245_;
  assign new_n6828_ = ~new_n6172_ | ~new_n6336_;
  assign new_n6829_ = ~new_n5897_ | ~new_n6824_;
  assign new_n6830_ = ~pi433 | ~new_n5240_;
  assign new_n6831_ = ~pi401 | ~new_n5241_;
  assign new_n6832_ = ~pi369 | ~new_n5242_;
  assign new_n6833_ = ~new_n18912_ | ~new_n5239_;
  assign new_n6834_ = ~new_n5275_;
  assign new_n6835_ = ~new_n5255_ | ~new_n5280_;
  assign new_n6836_ = ~new_n23402_ | ~new_n6151_;
  assign new_n6837_ = ~new_n24348_ | ~new_n6150_;
  assign new_n6838_ = ~new_n22810_ | ~new_n6146_;
  assign new_n6839_ = ~new_n20305_ | ~new_n6161_;
  assign new_n6840_ = ~new_n23875_ | ~new_n6163_;
  assign new_n6841_ = ~new_n21188_ | ~new_n5234_;
  assign new_n6842_ = ~new_n21689_ | ~new_n6142_;
  assign new_n6843_ = ~new_n5601_;
  assign new_n6844_ = ~new_n20059_ | ~new_n5247_;
  assign new_n6845_ = ~new_n5246_ | ~new_n5275_;
  assign new_n6846_ = ~new_n20688_ | ~new_n5245_;
  assign new_n6847_ = ~new_n6171_ | ~new_n6336_;
  assign new_n6848_ = ~new_n5901_ | ~new_n6843_;
  assign new_n6849_ = ~pi434 | ~new_n5240_;
  assign new_n6850_ = ~pi402 | ~new_n5241_;
  assign new_n6851_ = ~pi370 | ~new_n5242_;
  assign new_n6852_ = ~new_n18911_ | ~new_n5239_;
  assign new_n6853_ = ~new_n5276_;
  assign new_n6854_ = ~new_n5255_ | ~new_n5279_;
  assign new_n6855_ = ~new_n23309_ | ~new_n6151_;
  assign new_n6856_ = ~new_n24255_ | ~new_n6150_;
  assign new_n6857_ = ~new_n22898_ | ~new_n6146_;
  assign new_n6858_ = ~new_n20212_ | ~new_n6161_;
  assign new_n6859_ = ~new_n23782_ | ~new_n6163_;
  assign new_n6860_ = ~new_n21276_ | ~new_n5234_;
  assign new_n6861_ = ~new_n21777_ | ~new_n6142_;
  assign new_n6862_ = ~new_n5603_;
  assign new_n6863_ = ~new_n20115_ | ~new_n5247_;
  assign new_n6864_ = ~new_n5246_ | ~new_n5276_;
  assign new_n6865_ = ~new_n20776_ | ~new_n5245_;
  assign new_n6866_ = ~new_n6170_ | ~new_n6336_;
  assign new_n6867_ = ~new_n5905_ | ~new_n6862_;
  assign new_n6868_ = ~new_n18860_ | ~new_n5239_;
  assign new_n6869_ = ~pi435 | ~new_n5240_;
  assign new_n6870_ = ~pi403 | ~new_n5241_;
  assign new_n6871_ = ~pi371 | ~new_n5242_;
  assign new_n6872_ = ~new_n5277_;
  assign new_n6873_ = ~new_n5255_ | ~new_n5275_;
  assign new_n6874_ = ~new_n23387_ | ~new_n6151_;
  assign new_n6875_ = ~new_n24333_ | ~new_n6150_;
  assign new_n6876_ = ~new_n22897_ | ~new_n6146_;
  assign new_n6877_ = ~new_n20290_ | ~new_n6161_;
  assign new_n6878_ = ~new_n23860_ | ~new_n6163_;
  assign new_n6879_ = ~new_n21275_ | ~new_n5234_;
  assign new_n6880_ = ~new_n21776_ | ~new_n6142_;
  assign new_n6881_ = ~new_n5605_;
  assign new_n6882_ = ~new_n20060_ | ~new_n5247_;
  assign new_n6883_ = ~new_n5246_ | ~new_n5277_;
  assign new_n6884_ = ~new_n20775_ | ~new_n5245_;
  assign new_n6885_ = ~new_n6169_ | ~new_n6336_;
  assign new_n6886_ = ~new_n5908_ | ~new_n6881_;
  assign new_n6887_ = ~pi436 | ~new_n5240_;
  assign new_n6888_ = ~pi404 | ~new_n5241_;
  assign new_n6889_ = ~pi372 | ~new_n5242_;
  assign new_n6890_ = ~new_n5281_;
  assign new_n6891_ = ~new_n7903_ | ~new_n5551_;
  assign new_n6892_ = ~new_n5567_ | ~new_n6891_;
  assign new_n6893_ = ~new_n5909_ | ~new_n5281_;
  assign new_n6894_ = ~new_n5255_ | ~new_n5276_;
  assign new_n6895_ = ~new_n23310_ | ~new_n6151_;
  assign new_n6896_ = ~new_n24256_ | ~new_n6150_;
  assign new_n6897_ = ~new_n22896_ | ~new_n6146_;
  assign new_n6898_ = ~new_n20213_ | ~new_n6161_;
  assign new_n6899_ = ~new_n23783_ | ~new_n6163_;
  assign new_n6900_ = ~new_n21274_ | ~new_n5234_;
  assign new_n6901_ = ~new_n21775_ | ~new_n6142_;
  assign new_n6902_ = ~new_n5607_;
  assign new_n6903_ = ~new_n20113_ | ~new_n5247_;
  assign new_n6904_ = ~new_n20774_ | ~new_n5245_;
  assign new_n6905_ = ~new_n6180_ | ~new_n6336_;
  assign new_n6906_ = ~new_n5913_ | ~new_n6902_;
  assign new_n6907_ = ~pi437 | ~new_n5240_;
  assign new_n6908_ = ~pi405 | ~new_n5241_;
  assign new_n6909_ = ~pi373 | ~new_n5242_;
  assign new_n6910_ = ~new_n5278_;
  assign new_n6911_ = ~new_n20062_ | ~new_n5247_;
  assign new_n6912_ = ~new_n6179_ | ~new_n6336_;
  assign new_n6913_ = ~new_n6911_ | ~new_n6912_ | ~new_n6133_;
  assign new_n6914_ = ~new_n20111_ | ~new_n5247_;
  assign new_n6915_ = ~new_n6178_ | ~new_n6336_;
  assign new_n6916_ = ~new_n6914_ | ~new_n6915_ | ~new_n6133_;
  assign new_n6917_ = ~new_n5916_ | ~new_n5236_;
  assign new_n6918_ = ~new_n5613_ | ~new_n6917_;
  assign new_n6919_ = ~new_n6141_ | ~new_n5638_;
  assign new_n6920_ = ~new_n5618_;
  assign new_n6921_ = ~new_n5257_ | ~new_n5300_;
  assign new_n6922_ = ~new_n5254_ | ~new_n20768_;
  assign new_n6923_ = ~new_n5253_ | ~pi500;
  assign new_n6924_ = ~new_n5252_ | ~new_n5647_;
  assign new_n6925_ = ~new_n5251_ | ~new_n5647_;
  assign new_n6926_ = ~new_n5257_ | ~new_n5290_;
  assign new_n6927_ = ~new_n5254_ | ~new_n20767_;
  assign new_n6928_ = ~new_n5253_ | ~pi510;
  assign new_n6929_ = ~new_n5252_ | ~new_n5652_;
  assign new_n6930_ = ~new_n5251_ | ~new_n20098_;
  assign new_n6931_ = ~new_n5257_ | ~new_n5286_;
  assign new_n6932_ = ~new_n5254_ | ~new_n20689_;
  assign new_n6933_ = ~new_n5253_ | ~pi495;
  assign new_n6934_ = ~new_n5252_ | ~new_n5655_;
  assign new_n6935_ = ~new_n5251_ | ~new_n20061_;
  assign new_n6936_ = ~new_n5257_ | ~new_n5282_;
  assign new_n6937_ = ~new_n5254_ | ~new_n20773_;
  assign new_n6938_ = ~new_n5253_ | ~new_n18859_;
  assign new_n6939_ = ~new_n5252_ | ~new_n5658_;
  assign new_n6940_ = ~new_n5251_ | ~new_n20063_;
  assign new_n6941_ = ~new_n5257_ | ~new_n5289_;
  assign new_n6942_ = ~new_n5254_ | ~new_n20772_;
  assign new_n6943_ = ~new_n5253_ | ~new_n18910_;
  assign new_n6944_ = ~new_n5252_ | ~new_n5661_;
  assign new_n6945_ = ~new_n5251_ | ~new_n20064_;
  assign new_n6946_ = ~new_n5257_ | ~new_n5293_;
  assign new_n6947_ = ~new_n5254_ | ~new_n20690_;
  assign new_n6948_ = ~new_n5253_ | ~new_n18909_;
  assign new_n6949_ = ~new_n5252_ | ~new_n5664_;
  assign new_n6950_ = ~new_n5251_ | ~new_n20108_;
  assign new_n6951_ = ~new_n5257_ | ~new_n5292_;
  assign new_n6952_ = ~new_n5254_ | ~new_n20771_;
  assign new_n6953_ = ~new_n5253_ | ~new_n18908_;
  assign new_n6954_ = ~new_n5252_ | ~new_n5667_;
  assign new_n6955_ = ~new_n5251_ | ~new_n20065_;
  assign new_n6956_ = ~new_n5257_ | ~new_n5306_;
  assign new_n6957_ = ~new_n5254_ | ~new_n20691_;
  assign new_n6958_ = ~new_n5253_ | ~new_n18907_;
  assign new_n6959_ = ~new_n5252_ | ~new_n5670_;
  assign new_n6960_ = ~new_n5251_ | ~new_n20066_;
  assign new_n6961_ = ~new_n5257_ | ~new_n5305_;
  assign new_n6962_ = ~new_n5254_ | ~new_n20770_;
  assign new_n6963_ = ~new_n5253_ | ~new_n18906_;
  assign new_n6964_ = ~new_n5252_ | ~new_n5673_;
  assign new_n6965_ = ~new_n5251_ | ~new_n20067_;
  assign new_n6966_ = ~new_n5257_ | ~new_n5284_;
  assign new_n6967_ = ~new_n5254_ | ~new_n20769_;
  assign new_n6968_ = ~new_n5253_ | ~new_n18905_;
  assign new_n6969_ = ~new_n5252_ | ~new_n5676_;
  assign new_n6970_ = ~new_n5251_ | ~new_n20106_;
  assign new_n6971_ = ~new_n5257_ | ~new_n5285_;
  assign new_n6972_ = ~new_n5254_ | ~new_n20683_;
  assign new_n6973_ = ~new_n5253_ | ~new_n18929_;
  assign new_n6974_ = ~new_n5252_ | ~new_n5679_;
  assign new_n6975_ = ~new_n5251_ | ~new_n20049_;
  assign new_n6976_ = ~new_n5257_ | ~new_n5294_;
  assign new_n6977_ = ~new_n5254_ | ~new_n20787_;
  assign new_n6978_ = ~new_n5253_ | ~new_n18928_;
  assign new_n6979_ = ~new_n5252_ | ~new_n5682_;
  assign new_n6980_ = ~new_n5251_ | ~new_n20050_;
  assign new_n6981_ = ~new_n5257_ | ~new_n5302_;
  assign new_n6982_ = ~new_n5254_ | ~new_n20786_;
  assign new_n6983_ = ~new_n5253_ | ~new_n18927_;
  assign new_n6984_ = ~new_n5252_ | ~new_n5685_;
  assign new_n6985_ = ~new_n5251_ | ~new_n20051_;
  assign new_n6986_ = ~new_n5257_ | ~new_n5301_;
  assign new_n6987_ = ~new_n5254_ | ~new_n20684_;
  assign new_n6988_ = ~new_n5253_ | ~new_n18926_;
  assign new_n6989_ = ~new_n5252_ | ~new_n5688_;
  assign new_n6990_ = ~new_n5251_ | ~new_n20129_;
  assign new_n6991_ = ~new_n5257_ | ~new_n5296_;
  assign new_n6992_ = ~new_n5254_ | ~new_n20785_;
  assign new_n6993_ = ~new_n5253_ | ~new_n18925_;
  assign new_n6994_ = ~new_n5252_ | ~new_n5691_;
  assign new_n6995_ = ~new_n5251_ | ~new_n20052_;
  assign new_n6996_ = ~new_n5257_ | ~new_n5295_;
  assign new_n6997_ = ~new_n5254_ | ~new_n20784_;
  assign new_n6998_ = ~new_n5253_ | ~new_n18924_;
  assign new_n6999_ = ~new_n5252_ | ~new_n5694_;
  assign new_n7000_ = ~new_n5251_ | ~new_n20053_;
  assign new_n7001_ = ~new_n5257_ | ~new_n5291_;
  assign new_n7002_ = ~new_n5254_ | ~new_n20783_;
  assign new_n7003_ = ~new_n5253_ | ~new_n18923_;
  assign new_n7004_ = ~new_n5252_ | ~new_n5697_;
  assign new_n7005_ = ~new_n5251_ | ~new_n20054_;
  assign new_n7006_ = ~new_n5257_ | ~new_n5304_;
  assign new_n7007_ = ~new_n5254_ | ~new_n20685_;
  assign new_n7008_ = ~new_n5253_ | ~new_n18922_;
  assign new_n7009_ = ~new_n5252_ | ~new_n5700_;
  assign new_n7010_ = ~new_n5251_ | ~new_n20127_;
  assign new_n7011_ = ~new_n5257_ | ~new_n5303_;
  assign new_n7012_ = ~new_n5254_ | ~new_n20782_;
  assign new_n7013_ = ~new_n5253_ | ~new_n18921_;
  assign new_n7014_ = ~new_n5252_ | ~new_n5703_;
  assign new_n7015_ = ~new_n5251_ | ~new_n20055_;
  assign new_n7016_ = ~new_n5257_ | ~new_n5298_;
  assign new_n7017_ = ~new_n5254_ | ~new_n20781_;
  assign new_n7018_ = ~new_n5253_ | ~new_n18920_;
  assign new_n7019_ = ~new_n5252_ | ~new_n5705_;
  assign new_n7020_ = ~new_n5251_ | ~new_n20125_;
  assign new_n7021_ = ~new_n5257_ | ~new_n5297_;
  assign new_n7022_ = ~new_n5254_ | ~new_n20686_;
  assign new_n7023_ = ~new_n5253_ | ~new_n18919_;
  assign new_n7024_ = ~new_n5252_ | ~new_n6177_;
  assign new_n7025_ = ~new_n5251_ | ~new_n20056_;
  assign new_n7026_ = ~new_n5257_ | ~new_n5283_;
  assign new_n7027_ = ~new_n5254_ | ~new_n20687_;
  assign new_n7028_ = ~new_n5253_ | ~new_n18918_;
  assign new_n7029_ = ~new_n5252_ | ~new_n6176_;
  assign new_n7030_ = ~new_n5251_ | ~new_n20121_;
  assign new_n7031_ = ~new_n5257_ | ~new_n5288_;
  assign new_n7032_ = ~new_n5254_ | ~new_n20780_;
  assign new_n7033_ = ~new_n5253_ | ~new_n18917_;
  assign new_n7034_ = ~new_n5252_ | ~new_n6175_;
  assign new_n7035_ = ~new_n5251_ | ~new_n20057_;
  assign new_n7036_ = ~new_n5257_ | ~new_n5287_;
  assign new_n7037_ = ~new_n5254_ | ~new_n20779_;
  assign new_n7038_ = ~new_n5253_ | ~new_n18916_;
  assign new_n7039_ = ~new_n5252_ | ~new_n6174_;
  assign new_n7040_ = ~new_n5251_ | ~new_n20119_;
  assign new_n7041_ = ~new_n5257_ | ~new_n5280_;
  assign new_n7042_ = ~new_n5254_ | ~new_n20778_;
  assign new_n7043_ = ~new_n5253_ | ~new_n18915_;
  assign new_n7044_ = ~new_n5252_ | ~new_n6173_;
  assign new_n7045_ = ~new_n5251_ | ~new_n20058_;
  assign new_n7046_ = ~new_n5257_ | ~new_n5279_;
  assign new_n7047_ = ~new_n5254_ | ~new_n20777_;
  assign new_n7048_ = ~new_n5253_ | ~new_n18914_;
  assign new_n7049_ = ~new_n5252_ | ~new_n6172_;
  assign new_n7050_ = ~new_n5251_ | ~new_n20117_;
  assign new_n7051_ = ~new_n5257_ | ~new_n5275_;
  assign new_n7052_ = ~new_n5254_ | ~new_n20688_;
  assign new_n7053_ = ~new_n5253_ | ~new_n18913_;
  assign new_n7054_ = ~new_n5252_ | ~new_n6171_;
  assign new_n7055_ = ~new_n5251_ | ~new_n20059_;
  assign new_n7056_ = ~new_n5257_ | ~new_n5276_;
  assign new_n7057_ = ~new_n5254_ | ~new_n20776_;
  assign new_n7058_ = ~new_n5253_ | ~new_n18912_;
  assign new_n7059_ = ~new_n5252_ | ~new_n6170_;
  assign new_n7060_ = ~new_n5251_ | ~new_n20115_;
  assign new_n7061_ = ~new_n5257_ | ~new_n5277_;
  assign new_n7062_ = ~new_n5254_ | ~new_n20775_;
  assign new_n7063_ = ~new_n5253_ | ~new_n18911_;
  assign new_n7064_ = ~new_n5252_ | ~new_n6169_;
  assign new_n7065_ = ~new_n5251_ | ~new_n20060_;
  assign new_n7066_ = ~new_n5254_ | ~new_n20774_;
  assign new_n7067_ = ~new_n5253_ | ~new_n18860_;
  assign new_n7068_ = ~new_n5252_ | ~new_n6180_;
  assign new_n7069_ = ~new_n5251_ | ~new_n20113_;
  assign new_n7070_ = ~new_n5252_ | ~new_n6179_;
  assign new_n7071_ = ~new_n5251_ | ~new_n20062_;
  assign new_n7072_ = ~new_n5252_ | ~new_n6178_;
  assign new_n7073_ = ~new_n5251_ | ~new_n20111_;
  assign new_n7074_ = ~new_n5975_ | ~new_n5613_ | ~new_n6920_ | ~new_n5271_ | ~new_n5615_;
  assign new_n7075_ = ~new_n19753_ | ~new_n5263_;
  assign new_n7076_ = ~new_n5261_ | ~new_n5644_;
  assign new_n7077_ = ~new_n19448_ | ~new_n5259_;
  assign new_n7078_ = ~new_n7077_ | ~new_n7076_ | ~new_n7075_;
  assign new_n7079_ = ~new_n19753_ | ~new_n5238_;
  assign new_n7080_ = ~new_n5237_ | ~new_n19448_;
  assign new_n7081_ = ~new_n7903_ | ~new_n5644_;
  assign new_n7082_ = ~new_n7081_ | ~new_n7080_ | ~new_n7079_;
  assign new_n7083_ = ~new_n5621_;
  assign new_n7084_ = ~new_n5265_ | ~new_n7078_;
  assign new_n7085_ = ~po511 | ~new_n7082_;
  assign new_n7086_ = ~new_n5264_ | ~new_n19753_;
  assign new_n7087_ = ~pi513 | ~po509;
  assign new_n7088_ = ~new_n5262_ | ~new_n5644_;
  assign new_n7089_ = ~new_n5260_ | ~new_n19448_;
  assign new_n7090_ = ~pi438 | ~new_n7083_;
  assign new_n7091_ = ~new_n19815_ | ~new_n5263_;
  assign new_n7092_ = ~new_n5261_ | ~new_n5702_;
  assign new_n7093_ = ~new_n19510_ | ~new_n5259_;
  assign new_n7094_ = ~new_n7093_ | ~new_n7092_ | ~new_n7091_;
  assign new_n7095_ = ~new_n19815_ | ~new_n5238_;
  assign new_n7096_ = ~new_n19510_ | ~new_n5237_;
  assign new_n7097_ = ~new_n7903_ | ~new_n5702_;
  assign new_n7098_ = ~new_n7097_ | ~new_n7096_ | ~new_n7095_;
  assign new_n7099_ = ~new_n5265_ | ~new_n7094_;
  assign new_n7100_ = ~po511 | ~new_n7098_;
  assign new_n7101_ = ~new_n19815_ | ~new_n5264_;
  assign new_n7102_ = ~pi494 | ~po509;
  assign new_n7103_ = ~new_n5262_ | ~new_n5702_;
  assign new_n7104_ = ~new_n19510_ | ~new_n5260_;
  assign new_n7105_ = ~pi439 | ~new_n7083_;
  assign new_n7106_ = ~new_n19752_ | ~new_n5263_;
  assign new_n7107_ = ~new_n5261_ | ~new_n5699_;
  assign new_n7108_ = ~new_n19447_ | ~new_n5259_;
  assign new_n7109_ = ~new_n7108_ | ~new_n7107_ | ~new_n7106_;
  assign new_n7110_ = ~new_n19752_ | ~new_n5238_;
  assign new_n7111_ = ~new_n19447_ | ~new_n5237_;
  assign new_n7112_ = ~new_n7903_ | ~new_n5699_;
  assign new_n7113_ = ~new_n7112_ | ~new_n7111_ | ~new_n7110_;
  assign new_n7114_ = ~new_n5265_ | ~new_n7109_;
  assign new_n7115_ = ~po511 | ~new_n7113_;
  assign new_n7116_ = ~new_n19752_ | ~new_n5264_;
  assign new_n7117_ = ~pi504 | ~po509;
  assign new_n7118_ = ~new_n5262_ | ~new_n5699_;
  assign new_n7119_ = ~new_n19447_ | ~new_n5260_;
  assign new_n7120_ = ~pi440 | ~new_n7083_;
  assign new_n7121_ = ~new_n19816_ | ~new_n5263_;
  assign new_n7122_ = ~new_n5261_ | ~new_n5696_;
  assign new_n7123_ = ~new_n19511_ | ~new_n5259_;
  assign new_n7124_ = ~new_n7123_ | ~new_n7122_ | ~new_n7121_;
  assign new_n7125_ = ~new_n19816_ | ~new_n5238_;
  assign new_n7126_ = ~new_n19511_ | ~new_n5237_;
  assign new_n7127_ = ~new_n7903_ | ~new_n5696_;
  assign new_n7128_ = ~new_n7127_ | ~new_n7126_ | ~new_n7125_;
  assign new_n7129_ = ~new_n5265_ | ~new_n7124_;
  assign new_n7130_ = ~po511 | ~new_n7128_;
  assign new_n7131_ = ~new_n19816_ | ~new_n5264_;
  assign new_n7132_ = ~pi506 | ~po509;
  assign new_n7133_ = ~new_n5262_ | ~new_n5696_;
  assign new_n7134_ = ~new_n19511_ | ~new_n5260_;
  assign new_n7135_ = ~pi441 | ~new_n7083_;
  assign new_n7136_ = ~new_n19817_ | ~new_n5263_;
  assign new_n7137_ = ~new_n5261_ | ~new_n5693_;
  assign new_n7138_ = ~new_n19512_ | ~new_n5259_;
  assign new_n7139_ = ~new_n7138_ | ~new_n7137_ | ~new_n7136_;
  assign new_n7140_ = ~new_n19817_ | ~new_n5238_;
  assign new_n7141_ = ~new_n19512_ | ~new_n5237_;
  assign new_n7142_ = ~new_n7903_ | ~new_n5693_;
  assign new_n7143_ = ~new_n7142_ | ~new_n7141_ | ~new_n7140_;
  assign new_n7144_ = ~new_n5265_ | ~new_n7139_;
  assign new_n7145_ = ~po511 | ~new_n7143_;
  assign new_n7146_ = ~new_n19817_ | ~new_n5264_;
  assign new_n7147_ = ~pi491 | ~po509;
  assign new_n7148_ = ~new_n5262_ | ~new_n5693_;
  assign new_n7149_ = ~new_n19512_ | ~new_n5260_;
  assign new_n7150_ = ~pi442 | ~new_n7083_;
  assign new_n7151_ = ~new_n19818_ | ~new_n5263_;
  assign new_n7152_ = ~new_n5261_ | ~new_n5690_;
  assign new_n7153_ = ~new_n19513_ | ~new_n5259_;
  assign new_n7154_ = ~new_n7153_ | ~new_n7152_ | ~new_n7151_;
  assign new_n7155_ = ~new_n19818_ | ~new_n5238_;
  assign new_n7156_ = ~new_n19513_ | ~new_n5237_;
  assign new_n7157_ = ~new_n7903_ | ~new_n5690_;
  assign new_n7158_ = ~new_n7157_ | ~new_n7156_ | ~new_n7155_;
  assign new_n7159_ = ~new_n5265_ | ~new_n7154_;
  assign new_n7160_ = ~po511 | ~new_n7158_;
  assign new_n7161_ = ~new_n19818_ | ~new_n5264_;
  assign new_n7162_ = ~pi517 | ~po509;
  assign new_n7163_ = ~new_n5262_ | ~new_n5690_;
  assign new_n7164_ = ~new_n19513_ | ~new_n5260_;
  assign new_n7165_ = ~pi443 | ~new_n7083_;
  assign new_n7166_ = ~new_n19751_ | ~new_n5263_;
  assign new_n7167_ = ~new_n5261_ | ~new_n5687_;
  assign new_n7168_ = ~new_n19446_ | ~new_n5259_;
  assign new_n7169_ = ~new_n7168_ | ~new_n7167_ | ~new_n7166_;
  assign new_n7170_ = ~new_n19751_ | ~new_n5238_;
  assign new_n7171_ = ~new_n19446_ | ~new_n5237_;
  assign new_n7172_ = ~new_n7903_ | ~new_n5687_;
  assign new_n7173_ = ~new_n7172_ | ~new_n7171_ | ~new_n7170_;
  assign new_n7174_ = ~new_n5265_ | ~new_n7169_;
  assign new_n7175_ = ~po511 | ~new_n7173_;
  assign new_n7176_ = ~new_n19751_ | ~new_n5264_;
  assign new_n7177_ = ~pi498 | ~po509;
  assign new_n7178_ = ~new_n5262_ | ~new_n5687_;
  assign new_n7179_ = ~new_n19446_ | ~new_n5260_;
  assign new_n7180_ = ~pi444 | ~new_n7083_;
  assign new_n7181_ = ~new_n19819_ | ~new_n5263_;
  assign new_n7182_ = ~new_n5261_ | ~new_n5684_;
  assign new_n7183_ = ~new_n19514_ | ~new_n5259_;
  assign new_n7184_ = ~new_n7183_ | ~new_n7182_ | ~new_n7181_;
  assign new_n7185_ = ~new_n19819_ | ~new_n5238_;
  assign new_n7186_ = ~new_n19514_ | ~new_n5237_;
  assign new_n7187_ = ~new_n7903_ | ~new_n5684_;
  assign new_n7188_ = ~new_n7187_ | ~new_n7186_ | ~new_n7185_;
  assign new_n7189_ = ~new_n5265_ | ~new_n7184_;
  assign new_n7190_ = ~po511 | ~new_n7188_;
  assign new_n7191_ = ~new_n19819_ | ~new_n5264_;
  assign new_n7192_ = ~pi508 | ~po509;
  assign new_n7193_ = ~new_n5262_ | ~new_n5684_;
  assign new_n7194_ = ~new_n19514_ | ~new_n5260_;
  assign new_n7195_ = ~pi445 | ~new_n7083_;
  assign new_n7196_ = ~new_n19820_ | ~new_n5263_;
  assign new_n7197_ = ~new_n5261_ | ~new_n5681_;
  assign new_n7198_ = ~new_n19515_ | ~new_n5259_;
  assign new_n7199_ = ~new_n7198_ | ~new_n7197_ | ~new_n7196_;
  assign new_n7200_ = ~new_n19820_ | ~new_n5238_;
  assign new_n7201_ = ~new_n19515_ | ~new_n5237_;
  assign new_n7202_ = ~new_n7903_ | ~new_n5681_;
  assign new_n7203_ = ~new_n7202_ | ~new_n7201_ | ~new_n7200_;
  assign new_n7204_ = ~new_n5265_ | ~new_n7199_;
  assign new_n7205_ = ~po511 | ~new_n7203_;
  assign new_n7206_ = ~new_n19820_ | ~new_n5264_;
  assign new_n7207_ = ~pi496 | ~po509;
  assign new_n7208_ = ~new_n5262_ | ~new_n5681_;
  assign new_n7209_ = ~new_n19515_ | ~new_n5260_;
  assign new_n7210_ = ~pi446 | ~new_n7083_;
  assign new_n7211_ = ~new_n19750_ | ~new_n5263_;
  assign new_n7212_ = ~new_n5261_ | ~new_n5678_;
  assign new_n7213_ = ~new_n19445_ | ~new_n5259_;
  assign new_n7214_ = ~new_n7213_ | ~new_n7212_ | ~new_n7211_;
  assign new_n7215_ = ~new_n19750_ | ~new_n5238_;
  assign new_n7216_ = ~new_n19445_ | ~new_n5237_;
  assign new_n7217_ = ~new_n7903_ | ~new_n5678_;
  assign new_n7218_ = ~new_n7217_ | ~new_n7216_ | ~new_n7215_;
  assign new_n7219_ = ~new_n5265_ | ~new_n7214_;
  assign new_n7220_ = ~po511 | ~new_n7218_;
  assign new_n7221_ = ~new_n19750_ | ~new_n5264_;
  assign new_n7222_ = ~pi515 | ~po509;
  assign new_n7223_ = ~new_n5262_ | ~new_n5678_;
  assign new_n7224_ = ~new_n19445_ | ~new_n5260_;
  assign new_n7225_ = ~pi447 | ~new_n7083_;
  assign new_n7226_ = ~new_n19810_ | ~new_n5263_;
  assign new_n7227_ = ~new_n5261_ | ~new_n5675_;
  assign new_n7228_ = ~new_n19505_ | ~new_n5259_;
  assign new_n7229_ = ~new_n7228_ | ~new_n7227_ | ~new_n7226_;
  assign new_n7230_ = ~new_n19810_ | ~new_n5238_;
  assign new_n7231_ = ~new_n19505_ | ~new_n5237_;
  assign new_n7232_ = ~new_n7903_ | ~new_n5675_;
  assign new_n7233_ = ~new_n7232_ | ~new_n7231_ | ~new_n7230_;
  assign new_n7234_ = ~new_n5265_ | ~new_n7229_;
  assign new_n7235_ = ~po511 | ~new_n7233_;
  assign new_n7236_ = ~new_n19810_ | ~new_n5264_;
  assign new_n7237_ = ~pi501 | ~po509;
  assign new_n7238_ = ~new_n5262_ | ~new_n5675_;
  assign new_n7239_ = ~new_n19505_ | ~new_n5260_;
  assign new_n7240_ = ~pi448 | ~new_n7083_;
  assign new_n7241_ = ~new_n19811_ | ~new_n5263_;
  assign new_n7242_ = ~new_n5261_ | ~new_n5672_;
  assign new_n7243_ = ~new_n19506_ | ~new_n5259_;
  assign new_n7244_ = ~new_n7243_ | ~new_n7242_ | ~new_n7241_;
  assign new_n7245_ = ~new_n19811_ | ~new_n5238_;
  assign new_n7246_ = ~new_n19506_ | ~new_n5237_;
  assign new_n7247_ = ~new_n7903_ | ~new_n5672_;
  assign new_n7248_ = ~new_n7247_ | ~new_n7246_ | ~new_n7245_;
  assign new_n7249_ = ~new_n5265_ | ~new_n7244_;
  assign new_n7250_ = ~po511 | ~new_n7248_;
  assign new_n7251_ = ~new_n19811_ | ~new_n5264_;
  assign new_n7252_ = ~pi511 | ~po509;
  assign new_n7253_ = ~new_n5262_ | ~new_n5672_;
  assign new_n7254_ = ~new_n19506_ | ~new_n5260_;
  assign new_n7255_ = ~pi449 | ~new_n7083_;
  assign new_n7256_ = ~new_n19756_ | ~new_n5263_;
  assign new_n7257_ = ~new_n5261_ | ~new_n5669_;
  assign new_n7258_ = ~new_n19451_ | ~new_n5259_;
  assign new_n7259_ = ~new_n7258_ | ~new_n7257_ | ~new_n7256_;
  assign new_n7260_ = ~new_n19756_ | ~new_n5238_;
  assign new_n7261_ = ~new_n19451_ | ~new_n5237_;
  assign new_n7262_ = ~new_n7903_ | ~new_n5669_;
  assign new_n7263_ = ~new_n7262_ | ~new_n7261_ | ~new_n7260_;
  assign new_n7264_ = ~new_n5265_ | ~new_n7259_;
  assign new_n7265_ = ~po511 | ~new_n7263_;
  assign new_n7266_ = ~new_n19756_ | ~new_n5264_;
  assign new_n7267_ = ~pi519 | ~po509;
  assign new_n7268_ = ~new_n5262_ | ~new_n5669_;
  assign new_n7269_ = ~new_n19451_ | ~new_n5260_;
  assign new_n7270_ = ~pi450 | ~new_n7083_;
  assign new_n7271_ = ~new_n19812_ | ~new_n5263_;
  assign new_n7272_ = ~new_n5261_ | ~new_n5666_;
  assign new_n7273_ = ~new_n19507_ | ~new_n5259_;
  assign new_n7274_ = ~new_n7273_ | ~new_n7272_ | ~new_n7271_;
  assign new_n7275_ = ~new_n19812_ | ~new_n5238_;
  assign new_n7276_ = ~new_n19507_ | ~new_n5237_;
  assign new_n7277_ = ~new_n7903_ | ~new_n5666_;
  assign new_n7278_ = ~new_n7277_ | ~new_n7276_ | ~new_n7275_;
  assign new_n7279_ = ~new_n5265_ | ~new_n7274_;
  assign new_n7280_ = ~po511 | ~new_n7278_;
  assign new_n7281_ = ~new_n19812_ | ~new_n5264_;
  assign new_n7282_ = ~pi493 | ~po509;
  assign new_n7283_ = ~new_n5262_ | ~new_n5666_;
  assign new_n7284_ = ~new_n19507_ | ~new_n5260_;
  assign new_n7285_ = ~pi451 | ~new_n7083_;
  assign new_n7286_ = ~new_n19755_ | ~new_n5263_;
  assign new_n7287_ = ~new_n5261_ | ~new_n5663_;
  assign new_n7288_ = ~new_n19450_ | ~new_n5259_;
  assign new_n7289_ = ~new_n7288_ | ~new_n7287_ | ~new_n7286_;
  assign new_n7290_ = ~new_n19755_ | ~new_n5238_;
  assign new_n7291_ = ~new_n19450_ | ~new_n5237_;
  assign new_n7292_ = ~new_n7903_ | ~new_n5663_;
  assign new_n7293_ = ~new_n7292_ | ~new_n7291_ | ~new_n7290_;
  assign new_n7294_ = ~new_n5265_ | ~new_n7289_;
  assign new_n7295_ = ~po511 | ~new_n7293_;
  assign new_n7296_ = ~new_n19755_ | ~new_n5264_;
  assign new_n7297_ = ~pi505 | ~po509;
  assign new_n7298_ = ~new_n5262_ | ~new_n5663_;
  assign new_n7299_ = ~new_n19450_ | ~new_n5260_;
  assign new_n7300_ = ~pi452 | ~new_n7083_;
  assign new_n7301_ = ~new_n19813_ | ~new_n5263_;
  assign new_n7302_ = ~new_n5261_ | ~new_n5660_;
  assign new_n7303_ = ~new_n19508_ | ~new_n5259_;
  assign new_n7304_ = ~new_n7303_ | ~new_n7302_ | ~new_n7301_;
  assign new_n7305_ = ~new_n19813_ | ~new_n5238_;
  assign new_n7306_ = ~new_n19508_ | ~new_n5237_;
  assign new_n7307_ = ~new_n7903_ | ~new_n5660_;
  assign new_n7308_ = ~new_n7307_ | ~new_n7306_ | ~new_n7305_;
  assign new_n7309_ = ~new_n5265_ | ~new_n7304_;
  assign new_n7310_ = ~po511 | ~new_n7308_;
  assign new_n7311_ = ~new_n19813_ | ~new_n5264_;
  assign new_n7312_ = ~pi502 | ~po509;
  assign new_n7313_ = ~new_n5262_ | ~new_n5660_;
  assign new_n7314_ = ~new_n19508_ | ~new_n5260_;
  assign new_n7315_ = ~pi453 | ~new_n7083_;
  assign new_n7316_ = ~new_n19814_ | ~new_n5263_;
  assign new_n7317_ = ~new_n5261_ | ~new_n5657_;
  assign new_n7318_ = ~new_n19509_ | ~new_n5259_;
  assign new_n7319_ = ~new_n7318_ | ~new_n7317_ | ~new_n7316_;
  assign new_n7320_ = ~new_n19814_ | ~new_n5238_;
  assign new_n7321_ = ~new_n19509_ | ~new_n5237_;
  assign new_n7322_ = ~new_n7903_ | ~new_n5657_;
  assign new_n7323_ = ~new_n7322_ | ~new_n7321_ | ~new_n7320_;
  assign new_n7324_ = ~new_n5265_ | ~new_n7319_;
  assign new_n7325_ = ~po511 | ~new_n7323_;
  assign new_n7326_ = ~new_n19814_ | ~new_n5264_;
  assign new_n7327_ = ~pi514 | ~po509;
  assign new_n7328_ = ~new_n5262_ | ~new_n5657_;
  assign new_n7329_ = ~new_n19509_ | ~new_n5260_;
  assign new_n7330_ = ~pi454 | ~new_n7083_;
  assign new_n7331_ = ~new_n19754_ | ~new_n5263_;
  assign new_n7332_ = ~new_n5261_ | ~new_n5654_;
  assign new_n7333_ = ~new_n19449_ | ~new_n5259_;
  assign new_n7334_ = ~new_n7333_ | ~new_n7332_ | ~new_n7331_;
  assign new_n7335_ = ~new_n19754_ | ~new_n5238_;
  assign new_n7336_ = ~new_n19449_ | ~new_n5237_;
  assign new_n7337_ = ~new_n7903_ | ~new_n5654_;
  assign new_n7338_ = ~new_n7337_ | ~new_n7336_ | ~new_n7335_;
  assign new_n7339_ = ~new_n5265_ | ~new_n7334_;
  assign new_n7340_ = ~po511 | ~new_n7338_;
  assign new_n7341_ = ~new_n19754_ | ~new_n5264_;
  assign new_n7342_ = ~pi495 | ~po509;
  assign new_n7343_ = ~new_n5262_ | ~new_n5654_;
  assign new_n7344_ = ~new_n19449_ | ~new_n5260_;
  assign new_n7345_ = ~pi455 | ~new_n7083_;
  assign new_n7346_ = ~new_n19808_ | ~new_n5263_;
  assign new_n7347_ = ~new_n5261_ | ~new_n5651_;
  assign new_n7348_ = ~new_n19503_ | ~new_n5259_;
  assign new_n7349_ = ~new_n7348_ | ~new_n7347_ | ~new_n7346_;
  assign new_n7350_ = ~new_n19808_ | ~new_n5238_;
  assign new_n7351_ = ~new_n19503_ | ~new_n5237_;
  assign new_n7352_ = ~new_n7903_ | ~new_n5651_;
  assign new_n7353_ = ~new_n7352_ | ~new_n7351_ | ~new_n7350_;
  assign new_n7354_ = ~new_n5265_ | ~new_n7349_;
  assign new_n7355_ = ~po511 | ~new_n7353_;
  assign new_n7356_ = ~new_n19808_ | ~new_n5264_;
  assign new_n7357_ = ~pi510 | ~po509;
  assign new_n7358_ = ~new_n5262_ | ~new_n5651_;
  assign new_n7359_ = ~new_n19503_ | ~new_n5260_;
  assign new_n7360_ = ~pi456 | ~new_n7083_;
  assign new_n7361_ = ~new_n19809_ | ~new_n5263_;
  assign new_n7362_ = ~new_n5261_ | ~new_n5645_;
  assign new_n7363_ = ~new_n19504_ | ~new_n5259_;
  assign new_n7364_ = ~new_n7363_ | ~new_n7362_ | ~new_n7361_;
  assign new_n7365_ = ~new_n19809_ | ~new_n5238_;
  assign new_n7366_ = ~new_n19504_ | ~new_n5237_;
  assign new_n7367_ = ~new_n7903_ | ~new_n5645_;
  assign new_n7368_ = ~new_n7367_ | ~new_n7366_ | ~new_n7365_;
  assign new_n7369_ = ~new_n5265_ | ~new_n7364_;
  assign new_n7370_ = ~po511 | ~new_n7368_;
  assign new_n7371_ = ~new_n19809_ | ~new_n5264_;
  assign new_n7372_ = ~pi500 | ~po509;
  assign new_n7373_ = ~new_n5262_ | ~new_n5645_;
  assign new_n7374_ = ~new_n19504_ | ~new_n5260_;
  assign new_n7375_ = ~pi457 | ~new_n7083_;
  assign new_n7376_ = ~new_n6138_;
  assign new_n7377_ = ~new_n5557_ | ~new_n6156_ | ~new_n5554_;
  assign new_n7378_ = ~new_n7885_ | ~new_n7891_;
  assign new_n7379_ = ~new_n5644_ | ~new_n7378_;
  assign new_n7380_ = ~new_n5639_ | ~new_n7379_;
  assign new_n7381_ = ~new_n5560_ | ~new_n7380_;
  assign new_n7382_ = ~new_n5272_ | ~new_n8272_ | ~new_n8271_;
  assign new_n7383_ = ~pi490 | ~new_n7382_;
  assign new_n7384_ = ~new_n5258_ | ~new_n5301_;
  assign new_n7385_ = ~new_n5256_ | ~new_n5295_;
  assign new_n7386_ = ~new_n18924_ | ~new_n5626_;
  assign new_n7387_ = ~new_n7386_ | ~new_n7385_ | ~new_n7384_;
  assign new_n7388_ = ~new_n5374_;
  assign new_n7389_ = ~new_n6143_ | ~new_n5566_;
  assign new_n7390_ = ~new_n5639_ | ~new_n7389_;
  assign new_n7391_ = ~new_n6021_ | ~new_n6020_ | ~new_n7390_;
  assign new_n7392_ = ~new_n7391_ | ~new_n5626_;
  assign new_n7393_ = ~new_n5628_;
  assign new_n7394_ = ~new_n5694_ | ~new_n7856_;
  assign new_n7395_ = ~new_n18924_ | ~new_n7855_;
  assign new_n7396_ = ~new_n22286_ | ~new_n5248_;
  assign new_n7397_ = ~new_n6189_ | ~new_n7387_;
  assign new_n7398_ = ~pi491 | ~po509;
  assign new_n7399_ = ~new_n5258_ | ~new_n5280_;
  assign new_n7400_ = ~new_n5256_ | ~new_n5275_;
  assign new_n7401_ = ~new_n18913_ | ~new_n5626_;
  assign new_n7402_ = ~new_n7400_ | ~new_n7401_ | ~new_n7399_;
  assign new_n7403_ = ~new_n5618_ | ~new_n5626_;
  assign new_n7404_ = ~new_n7393_ | ~new_n7403_;
  assign new_n7405_ = ~new_n6166_ | ~new_n5618_;
  assign new_n7406_ = ~new_n5613_ | ~new_n7405_;
  assign new_n7407_ = ~new_n5267_ | ~new_n6171_;
  assign new_n7408_ = ~new_n5266_ | ~new_n18913_;
  assign new_n7409_ = ~new_n22191_ | ~new_n5248_;
  assign new_n7410_ = ~new_n6189_ | ~new_n7402_;
  assign new_n7411_ = ~pi492 | ~po509;
  assign new_n7412_ = ~new_n5258_ | ~new_n5289_;
  assign new_n7413_ = ~new_n5256_ | ~new_n5292_;
  assign new_n7414_ = ~new_n18908_ | ~new_n5626_;
  assign new_n7415_ = ~new_n7414_ | ~new_n7413_ | ~new_n7412_;
  assign new_n7416_ = ~new_n5667_ | ~new_n7856_;
  assign new_n7417_ = ~new_n18908_ | ~new_n7855_;
  assign new_n7418_ = ~new_n22271_ | ~new_n5248_;
  assign new_n7419_ = ~new_n6189_ | ~new_n7415_;
  assign new_n7420_ = ~pi493 | ~po509;
  assign new_n7421_ = ~new_n5258_ | ~new_n5291_;
  assign new_n7422_ = ~new_n5256_ | ~new_n5303_;
  assign new_n7423_ = ~new_n18921_ | ~new_n5626_;
  assign new_n7424_ = ~new_n7423_ | ~new_n7422_ | ~new_n7421_;
  assign new_n7425_ = ~new_n5703_ | ~new_n7856_;
  assign new_n7426_ = ~new_n18921_ | ~new_n7855_;
  assign new_n7427_ = ~new_n22284_ | ~new_n5248_;
  assign new_n7428_ = ~new_n6189_ | ~new_n7424_;
  assign new_n7429_ = ~pi494 | ~po509;
  assign new_n7430_ = ~new_n5258_ | ~new_n5300_;
  assign new_n7431_ = ~new_n5256_ | ~new_n5286_;
  assign new_n7432_ = ~pi495 | ~new_n5626_;
  assign new_n7433_ = ~new_n7432_ | ~new_n7431_ | ~new_n7430_;
  assign new_n7434_ = ~new_n5655_ | ~new_n7856_;
  assign new_n7435_ = ~pi495 | ~new_n7855_;
  assign new_n7436_ = ~new_n22274_ | ~new_n5248_;
  assign new_n7437_ = ~new_n6189_ | ~new_n7433_;
  assign new_n7438_ = ~pi495 | ~po509;
  assign new_n7439_ = ~new_n5258_ | ~new_n5284_;
  assign new_n7440_ = ~new_n5256_ | ~new_n5294_;
  assign new_n7441_ = ~new_n18928_ | ~new_n5626_;
  assign new_n7442_ = ~new_n7441_ | ~new_n7440_ | ~new_n7439_;
  assign new_n7443_ = ~new_n5682_ | ~new_n7856_;
  assign new_n7444_ = ~new_n18928_ | ~new_n7855_;
  assign new_n7445_ = ~new_n22289_ | ~new_n5248_;
  assign new_n7446_ = ~new_n6189_ | ~new_n7442_;
  assign new_n7447_ = ~pi496 | ~po509;
  assign new_n7448_ = ~new_n5258_ | ~new_n5297_;
  assign new_n7449_ = ~new_n5256_ | ~new_n5288_;
  assign new_n7450_ = ~new_n18917_ | ~new_n5626_;
  assign new_n7451_ = ~new_n7450_ | ~new_n7449_ | ~new_n7448_;
  assign new_n7452_ = ~new_n5267_ | ~new_n6175_;
  assign new_n7453_ = ~new_n5266_ | ~new_n18917_;
  assign new_n7454_ = ~new_n22280_ | ~new_n5248_;
  assign new_n7455_ = ~new_n6189_ | ~new_n7451_;
  assign new_n7456_ = ~pi497 | ~po509;
  assign new_n7457_ = ~new_n5258_ | ~new_n5294_;
  assign new_n7458_ = ~new_n5256_ | ~new_n5301_;
  assign new_n7459_ = ~new_n18926_ | ~new_n5626_;
  assign new_n7460_ = ~new_n7459_ | ~new_n7458_ | ~new_n7457_;
  assign new_n7461_ = ~new_n5688_ | ~new_n7856_;
  assign new_n7462_ = ~new_n18926_ | ~new_n7855_;
  assign new_n7463_ = ~new_n22188_ | ~new_n5248_;
  assign new_n7464_ = ~new_n6189_ | ~new_n7460_;
  assign new_n7465_ = ~pi498 | ~po509;
  assign new_n7466_ = ~new_n5258_ | ~new_n5303_;
  assign new_n7467_ = ~new_n5256_ | ~new_n5297_;
  assign new_n7468_ = ~new_n18919_ | ~new_n5626_;
  assign new_n7469_ = ~new_n7468_ | ~new_n7467_ | ~new_n7466_;
  assign new_n7470_ = ~new_n5267_ | ~new_n6177_;
  assign new_n7471_ = ~new_n5266_ | ~new_n18919_;
  assign new_n7472_ = ~new_n22281_ | ~new_n5248_;
  assign new_n7473_ = ~new_n6189_ | ~new_n7469_;
  assign new_n7474_ = ~pi499 | ~po509;
  assign new_n7475_ = ~new_n5627_ | ~new_n5625_;
  assign new_n7476_ = ~new_n7475_ | ~new_n5626_;
  assign new_n7477_ = ~new_n6190_ | ~new_n7476_;
  assign new_n7478_ = ~new_n6026_ | ~new_n5256_;
  assign new_n7479_ = ~new_n5647_ | ~new_n7856_;
  assign new_n7480_ = ~pi500 | ~new_n7477_;
  assign new_n7481_ = ~new_n22268_ | ~new_n5248_;
  assign new_n7482_ = ~pi500 | ~po509;
  assign new_n7483_ = ~new_n5258_ | ~new_n5306_;
  assign new_n7484_ = ~new_n5256_ | ~new_n5284_;
  assign new_n7485_ = ~new_n18905_ | ~new_n5626_;
  assign new_n7486_ = ~new_n7485_ | ~new_n7484_ | ~new_n7483_;
  assign new_n7487_ = ~new_n5676_ | ~new_n7856_;
  assign new_n7488_ = ~new_n18905_ | ~new_n7855_;
  assign new_n7489_ = ~new_n22269_ | ~new_n5248_;
  assign new_n7490_ = ~new_n6189_ | ~new_n7486_;
  assign new_n7491_ = ~pi501 | ~po509;
  assign new_n7492_ = ~new_n5258_ | ~new_n5286_;
  assign new_n7493_ = ~new_n5256_ | ~new_n5289_;
  assign new_n7494_ = ~new_n18910_ | ~new_n5626_;
  assign new_n7495_ = ~new_n7494_ | ~new_n7493_ | ~new_n7492_;
  assign new_n7496_ = ~new_n5661_ | ~new_n7856_;
  assign new_n7497_ = ~new_n18910_ | ~new_n7855_;
  assign new_n7498_ = ~new_n22273_ | ~new_n5248_;
  assign new_n7499_ = ~new_n6189_ | ~new_n7495_;
  assign new_n7500_ = ~pi502 | ~po509;
  assign new_n7501_ = ~new_n5258_ | ~new_n5288_;
  assign new_n7502_ = ~new_n5256_ | ~new_n5280_;
  assign new_n7503_ = ~new_n18915_ | ~new_n5626_;
  assign new_n7504_ = ~new_n7503_ | ~new_n7502_ | ~new_n7501_;
  assign new_n7505_ = ~new_n5267_ | ~new_n6173_;
  assign new_n7506_ = ~new_n5266_ | ~new_n18915_;
  assign new_n7507_ = ~new_n22278_ | ~new_n5248_;
  assign new_n7508_ = ~new_n6189_ | ~new_n7504_;
  assign new_n7509_ = ~pi503 | ~po509;
  assign new_n7510_ = ~new_n5258_ | ~new_n5295_;
  assign new_n7511_ = ~new_n5256_ | ~new_n5304_;
  assign new_n7512_ = ~new_n18922_ | ~new_n5626_;
  assign new_n7513_ = ~new_n7512_ | ~new_n7511_ | ~new_n7510_;
  assign new_n7514_ = ~new_n5700_ | ~new_n7856_;
  assign new_n7515_ = ~new_n18922_ | ~new_n7855_;
  assign new_n7516_ = ~new_n22189_ | ~new_n5248_;
  assign new_n7517_ = ~new_n6189_ | ~new_n7513_;
  assign new_n7518_ = ~pi504 | ~po509;
  assign new_n7519_ = ~new_n5258_ | ~new_n5282_;
  assign new_n7520_ = ~new_n5256_ | ~new_n5293_;
  assign new_n7521_ = ~new_n18909_ | ~new_n5626_;
  assign new_n7522_ = ~new_n7521_ | ~new_n7520_ | ~new_n7519_;
  assign new_n7523_ = ~new_n5664_ | ~new_n7856_;
  assign new_n7524_ = ~new_n18909_ | ~new_n7855_;
  assign new_n7525_ = ~new_n22272_ | ~new_n5248_;
  assign new_n7526_ = ~new_n6189_ | ~new_n7522_;
  assign new_n7527_ = ~pi505 | ~po509;
  assign new_n7528_ = ~new_n5258_ | ~new_n5296_;
  assign new_n7529_ = ~new_n5256_ | ~new_n5291_;
  assign new_n7530_ = ~new_n18923_ | ~new_n5626_;
  assign new_n7531_ = ~new_n7530_ | ~new_n7529_ | ~new_n7528_;
  assign new_n7532_ = ~new_n5697_ | ~new_n7856_;
  assign new_n7533_ = ~new_n18923_ | ~new_n7855_;
  assign new_n7534_ = ~new_n22285_ | ~new_n5248_;
  assign new_n7535_ = ~new_n6189_ | ~new_n7531_;
  assign new_n7536_ = ~pi506 | ~po509;
  assign new_n7537_ = ~new_n5258_ | ~new_n5287_;
  assign new_n7538_ = ~new_n5256_ | ~new_n5279_;
  assign new_n7539_ = ~new_n18914_ | ~new_n5626_;
  assign new_n7540_ = ~new_n7539_ | ~new_n7538_ | ~new_n7537_;
  assign new_n7541_ = ~new_n5267_ | ~new_n6172_;
  assign new_n7542_ = ~new_n5266_ | ~new_n18914_;
  assign new_n7543_ = ~new_n22277_ | ~new_n5248_;
  assign new_n7544_ = ~new_n6189_ | ~new_n7540_;
  assign new_n7545_ = ~pi507 | ~po509;
  assign new_n7546_ = ~new_n5258_ | ~new_n5285_;
  assign new_n7547_ = ~new_n5256_ | ~new_n5302_;
  assign new_n7548_ = ~new_n18927_ | ~new_n5626_;
  assign new_n7549_ = ~new_n7548_ | ~new_n7547_ | ~new_n7546_;
  assign new_n7550_ = ~new_n5685_ | ~new_n7856_;
  assign new_n7551_ = ~new_n18927_ | ~new_n7855_;
  assign new_n7552_ = ~new_n22288_ | ~new_n5248_;
  assign new_n7553_ = ~new_n6189_ | ~new_n7549_;
  assign new_n7554_ = ~pi508 | ~po509;
  assign new_n7555_ = ~new_n5258_ | ~new_n5298_;
  assign new_n7556_ = ~new_n5256_ | ~new_n5283_;
  assign new_n7557_ = ~new_n18918_ | ~new_n5626_;
  assign new_n7558_ = ~new_n7557_ | ~new_n7556_ | ~new_n7555_;
  assign new_n7559_ = ~new_n5267_ | ~new_n6176_;
  assign new_n7560_ = ~new_n5266_ | ~new_n18918_;
  assign new_n7561_ = ~new_n22190_ | ~new_n5248_;
  assign new_n7562_ = ~new_n6189_ | ~new_n7558_;
  assign new_n7563_ = ~pi509 | ~po509;
  assign new_n7564_ = ~new_n5258_ | ~new_n5299_;
  assign new_n7565_ = ~new_n5256_ | ~new_n5290_;
  assign new_n7566_ = ~pi510 | ~new_n5626_;
  assign new_n7567_ = ~new_n7566_ | ~new_n7565_ | ~new_n7564_;
  assign new_n7568_ = ~new_n5652_ | ~new_n7856_;
  assign new_n7569_ = ~pi510 | ~new_n7855_;
  assign new_n7570_ = ~new_n22282_ | ~new_n5248_;
  assign new_n7571_ = ~new_n6189_ | ~new_n7567_;
  assign new_n7572_ = ~pi510 | ~po509;
  assign new_n7573_ = ~new_n5258_ | ~new_n5292_;
  assign new_n7574_ = ~new_n5256_ | ~new_n5305_;
  assign new_n7575_ = ~new_n18906_ | ~new_n5626_;
  assign new_n7576_ = ~new_n7575_ | ~new_n7574_ | ~new_n7573_;
  assign new_n7577_ = ~new_n5673_ | ~new_n7856_;
  assign new_n7578_ = ~new_n18906_ | ~new_n7855_;
  assign new_n7579_ = ~new_n22270_ | ~new_n5248_;
  assign new_n7580_ = ~new_n6189_ | ~new_n7576_;
  assign new_n7581_ = ~pi511 | ~po509;
  assign new_n7582_ = ~new_n5258_ | ~new_n5275_;
  assign new_n7583_ = ~new_n5256_ | ~new_n5277_;
  assign new_n7584_ = ~new_n18911_ | ~new_n5626_;
  assign new_n7585_ = ~new_n7582_ | ~new_n7583_ | ~new_n7584_;
  assign new_n7586_ = ~new_n5267_ | ~new_n6169_;
  assign new_n7587_ = ~new_n5266_ | ~new_n18911_;
  assign new_n7588_ = ~new_n22275_ | ~new_n5248_;
  assign new_n7589_ = ~new_n6189_ | ~new_n7585_;
  assign new_n7590_ = ~pi512 | ~po509;
  assign new_n7591_ = ~new_n5258_ | ~new_n5304_;
  assign new_n7592_ = ~new_n5256_ | ~new_n5298_;
  assign new_n7593_ = ~new_n18920_ | ~new_n5626_;
  assign new_n7594_ = ~new_n7593_ | ~new_n7592_ | ~new_n7591_;
  assign new_n7595_ = ~new_n5705_ | ~new_n7856_;
  assign new_n7596_ = ~new_n18920_ | ~new_n7855_;
  assign new_n7597_ = ~new_n22283_ | ~new_n5248_;
  assign new_n7598_ = ~new_n6189_ | ~new_n7594_;
  assign new_n7599_ = ~pi513 | ~po509;
  assign new_n7600_ = ~new_n5258_ | ~new_n5290_;
  assign new_n7601_ = ~new_n5256_ | ~new_n5282_;
  assign new_n7602_ = ~new_n18859_ | ~new_n5626_;
  assign new_n7603_ = ~new_n7602_ | ~new_n7601_ | ~new_n7600_;
  assign new_n7604_ = ~new_n5658_ | ~new_n7856_;
  assign new_n7605_ = ~new_n18859_ | ~new_n7855_;
  assign new_n7606_ = ~new_n22192_ | ~new_n5248_;
  assign new_n7607_ = ~new_n6189_ | ~new_n7603_;
  assign new_n7608_ = ~pi514 | ~po509;
  assign new_n7609_ = ~new_n5258_ | ~new_n5305_;
  assign new_n7610_ = ~new_n5256_ | ~new_n5285_;
  assign new_n7611_ = ~new_n18929_ | ~new_n5626_;
  assign new_n7612_ = ~new_n7611_ | ~new_n7610_ | ~new_n7609_;
  assign new_n7613_ = ~new_n5679_ | ~new_n7856_;
  assign new_n7614_ = ~new_n18929_ | ~new_n7855_;
  assign new_n7615_ = ~new_n22290_ | ~new_n5248_;
  assign new_n7616_ = ~new_n6189_ | ~new_n7612_;
  assign new_n7617_ = ~pi515 | ~po509;
  assign new_n7618_ = ~new_n5258_ | ~new_n5283_;
  assign new_n7619_ = ~new_n5256_ | ~new_n5287_;
  assign new_n7620_ = ~new_n18916_ | ~new_n5626_;
  assign new_n7621_ = ~new_n7620_ | ~new_n7619_ | ~new_n7618_;
  assign new_n7622_ = ~new_n5267_ | ~new_n6174_;
  assign new_n7623_ = ~new_n5266_ | ~new_n18916_;
  assign new_n7624_ = ~new_n22279_ | ~new_n5248_;
  assign new_n7625_ = ~new_n6189_ | ~new_n7621_;
  assign new_n7626_ = ~pi516 | ~po509;
  assign new_n7627_ = ~new_n5258_ | ~new_n5302_;
  assign new_n7628_ = ~new_n5256_ | ~new_n5296_;
  assign new_n7629_ = ~new_n18925_ | ~new_n5626_;
  assign new_n7630_ = ~new_n7629_ | ~new_n7628_ | ~new_n7627_;
  assign new_n7631_ = ~new_n5691_ | ~new_n7856_;
  assign new_n7632_ = ~new_n18925_ | ~new_n7855_;
  assign new_n7633_ = ~new_n22287_ | ~new_n5248_;
  assign new_n7634_ = ~new_n6189_ | ~new_n7630_;
  assign new_n7635_ = ~pi517 | ~po509;
  assign new_n7636_ = ~new_n5258_ | ~new_n5279_;
  assign new_n7637_ = ~new_n5256_ | ~new_n5276_;
  assign new_n7638_ = ~new_n18912_ | ~new_n5626_;
  assign new_n7639_ = ~new_n7637_ | ~new_n7638_ | ~new_n7636_;
  assign new_n7640_ = ~new_n5267_ | ~new_n6170_;
  assign new_n7641_ = ~new_n5266_ | ~new_n18912_;
  assign new_n7642_ = ~new_n22276_ | ~new_n5248_;
  assign new_n7643_ = ~new_n6189_ | ~new_n7639_;
  assign new_n7644_ = ~pi518 | ~po509;
  assign new_n7645_ = ~new_n5258_ | ~new_n5293_;
  assign new_n7646_ = ~new_n5256_ | ~new_n5306_;
  assign new_n7647_ = ~new_n18907_ | ~new_n5626_;
  assign new_n7648_ = ~new_n7647_ | ~new_n7646_ | ~new_n7645_;
  assign new_n7649_ = ~new_n5670_ | ~new_n7856_;
  assign new_n7650_ = ~new_n18907_ | ~new_n7855_;
  assign new_n7651_ = ~new_n22193_ | ~new_n5248_;
  assign new_n7652_ = ~new_n6189_ | ~new_n7648_;
  assign new_n7653_ = ~pi519 | ~po509;
  assign new_n7654_ = ~new_n6168_ | ~new_n5268_;
  assign new_n7655_ = ~new_n5635_ | ~new_n5567_;
  assign new_n7656_ = ~new_n5639_ | ~new_n5638_;
  assign new_n7657_ = ~new_n6036_ | ~new_n5271_;
  assign new_n7658_ = ~new_n5631_;
  assign new_n7659_ = ~new_n5235_ | ~new_n5635_;
  assign new_n7660_ = ~new_n5631_ | ~new_n5629_;
  assign new_n7661_ = ~new_n5273_ | ~new_n7660_;
  assign new_n7662_ = ~new_n5305_ | ~new_n5249_;
  assign new_n7663_ = ~new_n7661_ | ~new_n5305_;
  assign new_n7664_ = ~new_n6149_ | ~new_n5676_;
  assign new_n7665_ = ~new_n5306_ | ~new_n5249_;
  assign new_n7666_ = ~new_n7661_ | ~new_n5306_;
  assign new_n7667_ = ~new_n6149_ | ~new_n5673_;
  assign new_n7668_ = ~new_n5292_ | ~new_n5249_;
  assign new_n7669_ = ~new_n7661_ | ~new_n5292_;
  assign new_n7670_ = ~new_n6149_ | ~new_n5670_;
  assign new_n7671_ = ~new_n5293_ | ~new_n5249_;
  assign new_n7672_ = ~new_n7661_ | ~new_n5293_;
  assign new_n7673_ = ~new_n6149_ | ~new_n5667_;
  assign new_n7674_ = ~new_n5289_ | ~new_n5249_;
  assign new_n7675_ = ~new_n7661_ | ~new_n5289_;
  assign new_n7676_ = ~new_n6149_ | ~new_n5664_;
  assign new_n7677_ = ~new_n5282_ | ~new_n5249_;
  assign new_n7678_ = ~new_n7661_ | ~new_n5282_;
  assign new_n7679_ = ~new_n6149_ | ~new_n5661_;
  assign new_n7680_ = ~new_n19436_ | ~new_n5249_;
  assign new_n7681_ = ~new_n7661_ | ~new_n5278_;
  assign new_n7682_ = ~new_n19434_ | ~new_n5249_;
  assign new_n7683_ = ~new_n7661_ | ~new_n5281_;
  assign new_n7684_ = ~new_n1571_ | ~new_n6149_ | ~new_n5567_;
  assign new_n7685_ = ~new_n5286_ | ~new_n5249_;
  assign new_n7686_ = ~new_n7661_ | ~new_n5286_;
  assign new_n7687_ = ~new_n6149_ | ~new_n5658_;
  assign new_n7688_ = ~new_n5277_ | ~new_n5249_;
  assign new_n7689_ = ~new_n7661_ | ~new_n5277_;
  assign new_n7690_ = ~new_n6149_ | ~new_n6180_;
  assign new_n7691_ = ~new_n5276_ | ~new_n5249_;
  assign new_n7692_ = ~new_n7661_ | ~new_n5276_;
  assign new_n7693_ = ~new_n6149_ | ~new_n6169_;
  assign new_n7694_ = ~new_n5275_ | ~new_n5249_;
  assign new_n7695_ = ~new_n7661_ | ~new_n5275_;
  assign new_n7696_ = ~new_n6149_ | ~new_n6170_;
  assign new_n7697_ = ~new_n5279_ | ~new_n5249_;
  assign new_n7698_ = ~new_n7661_ | ~new_n5279_;
  assign new_n7699_ = ~new_n6149_ | ~new_n6171_;
  assign new_n7700_ = ~new_n5280_ | ~new_n5249_;
  assign new_n7701_ = ~new_n7661_ | ~new_n5280_;
  assign new_n7702_ = ~new_n6149_ | ~new_n6172_;
  assign new_n7703_ = ~new_n5287_ | ~new_n5249_;
  assign new_n7704_ = ~new_n7661_ | ~new_n5287_;
  assign new_n7705_ = ~new_n6149_ | ~new_n6173_;
  assign new_n7706_ = ~new_n5288_ | ~new_n5249_;
  assign new_n7707_ = ~new_n7661_ | ~new_n5288_;
  assign new_n7708_ = ~new_n6149_ | ~new_n6174_;
  assign new_n7709_ = ~new_n5283_ | ~new_n5249_;
  assign new_n7710_ = ~new_n7661_ | ~new_n5283_;
  assign new_n7711_ = ~new_n6149_ | ~new_n6175_;
  assign new_n7712_ = ~new_n5297_ | ~new_n5249_;
  assign new_n7713_ = ~new_n7661_ | ~new_n5297_;
  assign new_n7714_ = ~new_n6149_ | ~new_n6176_;
  assign new_n7715_ = ~new_n5298_ | ~new_n5249_;
  assign new_n7716_ = ~new_n7661_ | ~new_n5298_;
  assign new_n7717_ = ~new_n6149_ | ~new_n6177_;
  assign new_n7718_ = ~new_n5290_ | ~new_n5249_;
  assign new_n7719_ = ~new_n7661_ | ~new_n5290_;
  assign new_n7720_ = ~new_n6149_ | ~new_n5655_;
  assign new_n7721_ = ~new_n5303_ | ~new_n5249_;
  assign new_n7722_ = ~new_n7661_ | ~new_n5303_;
  assign new_n7723_ = ~new_n6149_ | ~new_n5705_;
  assign new_n7724_ = ~new_n5304_ | ~new_n5249_;
  assign new_n7725_ = ~new_n7661_ | ~new_n5304_;
  assign new_n7726_ = ~new_n6149_ | ~new_n5703_;
  assign new_n7727_ = ~new_n5291_ | ~new_n5249_;
  assign new_n7728_ = ~new_n7661_ | ~new_n5291_;
  assign new_n7729_ = ~new_n6149_ | ~new_n5700_;
  assign new_n7730_ = ~new_n5295_ | ~new_n5249_;
  assign new_n7731_ = ~new_n7661_ | ~new_n5295_;
  assign new_n7732_ = ~new_n6149_ | ~new_n5697_;
  assign new_n7733_ = ~new_n5296_ | ~new_n5249_;
  assign new_n7734_ = ~new_n7661_ | ~new_n5296_;
  assign new_n7735_ = ~new_n6149_ | ~new_n5694_;
  assign new_n7736_ = ~new_n5301_ | ~new_n5249_;
  assign new_n7737_ = ~new_n7661_ | ~new_n5301_;
  assign new_n7738_ = ~new_n6149_ | ~new_n5691_;
  assign new_n7739_ = ~new_n5302_ | ~new_n5249_;
  assign new_n7740_ = ~new_n7661_ | ~new_n5302_;
  assign new_n7741_ = ~new_n6149_ | ~new_n5688_;
  assign new_n7742_ = ~new_n5294_ | ~new_n5249_;
  assign new_n7743_ = ~new_n7661_ | ~new_n5294_;
  assign new_n7744_ = ~new_n6149_ | ~new_n5685_;
  assign new_n7745_ = ~new_n5285_ | ~new_n5249_;
  assign new_n7746_ = ~new_n7661_ | ~new_n5285_;
  assign new_n7747_ = ~new_n6149_ | ~new_n5682_;
  assign new_n7748_ = ~new_n5284_ | ~new_n5249_;
  assign new_n7749_ = ~new_n7661_ | ~new_n5284_;
  assign new_n7750_ = ~new_n6149_ | ~new_n5679_;
  assign new_n7751_ = ~new_n5300_ | ~new_n5249_;
  assign new_n7752_ = ~new_n7661_ | ~new_n5300_;
  assign new_n7753_ = ~new_n6149_ | ~new_n5652_;
  assign new_n7754_ = ~new_n5299_ | ~new_n5249_;
  assign new_n7755_ = ~new_n7661_ | ~new_n5299_;
  assign new_n7756_ = ~new_n6149_ | ~new_n5647_;
  assign new_n7757_ = ~new_n7658_ | ~new_n5273_;
  assign new_n7758_ = ~new_n5676_ | ~new_n7757_;
  assign new_n7759_ = ~new_n6149_ | ~new_n5305_;
  assign new_n7760_ = ~new_n7878_ | ~new_n5306_;
  assign new_n7761_ = ~new_n5673_ | ~new_n7757_;
  assign new_n7762_ = ~new_n6149_ | ~new_n5306_;
  assign new_n7763_ = ~new_n7878_ | ~new_n5292_;
  assign new_n7764_ = ~new_n5670_ | ~new_n7757_;
  assign new_n7765_ = ~new_n6149_ | ~new_n5292_;
  assign new_n7766_ = ~new_n7878_ | ~new_n5293_;
  assign new_n7767_ = ~new_n5667_ | ~new_n7757_;
  assign new_n7768_ = ~new_n6149_ | ~new_n5293_;
  assign new_n7769_ = ~new_n7878_ | ~new_n5289_;
  assign new_n7770_ = ~new_n5664_ | ~new_n7757_;
  assign new_n7771_ = ~new_n6149_ | ~new_n5289_;
  assign new_n7772_ = ~new_n7878_ | ~new_n5282_;
  assign new_n7773_ = ~new_n5661_ | ~new_n7757_;
  assign new_n7774_ = ~new_n6149_ | ~new_n5282_;
  assign new_n7775_ = ~new_n7878_ | ~new_n5286_;
  assign new_n7776_ = ~new_n1570_ | ~new_n7757_ | ~new_n5567_;
  assign new_n7777_ = ~new_n6149_ | ~new_n5278_;
  assign new_n7778_ = ~new_n6179_ | ~new_n7757_;
  assign new_n7779_ = ~new_n6149_ | ~new_n5281_;
  assign new_n7780_ = ~new_n5658_ | ~new_n7757_;
  assign new_n7781_ = ~new_n6149_ | ~new_n5286_;
  assign new_n7782_ = ~new_n7878_ | ~new_n5290_;
  assign new_n7783_ = ~new_n6180_ | ~new_n7757_;
  assign new_n7784_ = ~new_n6149_ | ~new_n5277_;
  assign new_n7785_ = ~new_n7878_ | ~new_n5276_;
  assign new_n7786_ = ~new_n6169_ | ~new_n7757_;
  assign new_n7787_ = ~new_n6149_ | ~new_n5276_;
  assign new_n7788_ = ~new_n7878_ | ~new_n5275_;
  assign new_n7789_ = ~new_n6170_ | ~new_n7757_;
  assign new_n7790_ = ~new_n6149_ | ~new_n5275_;
  assign new_n7791_ = ~new_n7878_ | ~new_n5279_;
  assign new_n7792_ = ~new_n6171_ | ~new_n7757_;
  assign new_n7793_ = ~new_n6149_ | ~new_n5279_;
  assign new_n7794_ = ~new_n7878_ | ~new_n5280_;
  assign new_n7795_ = ~new_n6172_ | ~new_n7757_;
  assign new_n7796_ = ~new_n6149_ | ~new_n5280_;
  assign new_n7797_ = ~new_n7878_ | ~new_n5287_;
  assign new_n7798_ = ~new_n6173_ | ~new_n7757_;
  assign new_n7799_ = ~new_n6149_ | ~new_n5287_;
  assign new_n7800_ = ~new_n7878_ | ~new_n5288_;
  assign new_n7801_ = ~new_n6174_ | ~new_n7757_;
  assign new_n7802_ = ~new_n6149_ | ~new_n5288_;
  assign new_n7803_ = ~new_n7878_ | ~new_n5283_;
  assign new_n7804_ = ~new_n6175_ | ~new_n7757_;
  assign new_n7805_ = ~new_n6149_ | ~new_n5283_;
  assign new_n7806_ = ~new_n7878_ | ~new_n5297_;
  assign new_n7807_ = ~new_n6176_ | ~new_n7757_;
  assign new_n7808_ = ~new_n6149_ | ~new_n5297_;
  assign new_n7809_ = ~new_n7878_ | ~new_n5298_;
  assign new_n7810_ = ~new_n6177_ | ~new_n7757_;
  assign new_n7811_ = ~new_n6149_ | ~new_n5298_;
  assign new_n7812_ = ~new_n7878_ | ~new_n5303_;
  assign new_n7813_ = ~new_n5655_ | ~new_n7757_;
  assign new_n7814_ = ~new_n6149_ | ~new_n5290_;
  assign new_n7815_ = ~new_n7878_ | ~new_n5300_;
  assign new_n7816_ = ~new_n5705_ | ~new_n7757_;
  assign new_n7817_ = ~new_n6149_ | ~new_n5303_;
  assign new_n7818_ = ~new_n7878_ | ~new_n5304_;
  assign new_n7819_ = ~new_n5703_ | ~new_n7757_;
  assign new_n7820_ = ~new_n6149_ | ~new_n5304_;
  assign new_n7821_ = ~new_n7878_ | ~new_n5291_;
  assign new_n7822_ = ~new_n5700_ | ~new_n7757_;
  assign new_n7823_ = ~new_n6149_ | ~new_n5291_;
  assign new_n7824_ = ~new_n7878_ | ~new_n5295_;
  assign new_n7825_ = ~new_n5697_ | ~new_n7757_;
  assign new_n7826_ = ~new_n6149_ | ~new_n5295_;
  assign new_n7827_ = ~new_n7878_ | ~new_n5296_;
  assign new_n7828_ = ~new_n5694_ | ~new_n7757_;
  assign new_n7829_ = ~new_n6149_ | ~new_n5296_;
  assign new_n7830_ = ~new_n7878_ | ~new_n5301_;
  assign new_n7831_ = ~new_n5691_ | ~new_n7757_;
  assign new_n7832_ = ~new_n6149_ | ~new_n5301_;
  assign new_n7833_ = ~new_n7878_ | ~new_n5302_;
  assign new_n7834_ = ~new_n5688_ | ~new_n7757_;
  assign new_n7835_ = ~new_n6149_ | ~new_n5302_;
  assign new_n7836_ = ~new_n7878_ | ~new_n5294_;
  assign new_n7837_ = ~new_n5685_ | ~new_n7757_;
  assign new_n7838_ = ~new_n6149_ | ~new_n5294_;
  assign new_n7839_ = ~new_n7878_ | ~new_n5285_;
  assign new_n7840_ = ~new_n5682_ | ~new_n7757_;
  assign new_n7841_ = ~new_n6149_ | ~new_n5285_;
  assign new_n7842_ = ~new_n7878_ | ~new_n5284_;
  assign new_n7843_ = ~new_n5679_ | ~new_n7757_;
  assign new_n7844_ = ~new_n6149_ | ~new_n5284_;
  assign new_n7845_ = ~new_n7878_ | ~new_n5305_;
  assign new_n7846_ = ~new_n5652_ | ~new_n7757_;
  assign new_n7847_ = ~new_n6149_ | ~new_n5300_;
  assign new_n7848_ = ~new_n7878_ | ~new_n5299_;
  assign new_n7849_ = ~new_n5647_ | ~new_n7757_;
  assign new_n7850_ = ~new_n6149_ | ~new_n5299_;
  assign new_n7851_ = ~new_n7383_ | ~po509;
  assign new_n7852_ = ~new_n6048_ | ~new_n7681_;
  assign new_n7853_ = ~new_n6192_ | ~new_n5626_;
  assign new_n7854_ = ~new_n6166_ | ~new_n6192_;
  assign new_n7855_ = ~new_n7853_ | ~new_n6190_;
  assign new_n7856_ = ~new_n7854_ | ~new_n6191_;
  assign new_n7857_ = ~new_n5274_ | ~new_n6165_;
  assign new_n7858_ = ~new_n5274_ | ~new_n5550_;
  assign new_n7859_ = ~new_n6181_ | ~new_n5243_;
  assign new_n7860_ = ~new_n6007_ | ~new_n7383_;
  assign new_n7861_ = ~new_n8369_ | ~new_n6137_ | ~new_n7383_ | ~new_n8370_;
  assign new_n7862_ = ~new_n7872_ | ~new_n7866_;
  assign new_n7863_ = ~new_n5635_ | ~new_n5567_;
  assign new_n7864_ = ~pi302 | ~new_n6099_;
  assign new_n7865_ = ~pi309 | ~new_n19021_;
  assign new_n7866_ = ~new_n5632_;
  assign new_n7867_ = ~pi303 | ~new_n6099_;
  assign new_n7868_ = ~pi309 | ~new_n19119_;
  assign new_n7869_ = ~new_n5633_;
  assign new_n7870_ = ~pi304 | ~new_n6099_;
  assign new_n7871_ = ~pi309 | ~new_n19022_;
  assign new_n7872_ = ~new_n5634_;
  assign new_n7873_ = ~new_n7866_ | ~pi490;
  assign new_n7874_ = ~new_n5632_ | ~new_n5551_;
  assign new_n7875_ = ~new_n7874_ | ~new_n7873_;
  assign new_n7876_ = ~pi301 | ~new_n6099_;
  assign new_n7877_ = ~pi309 | ~new_n19020_;
  assign new_n7878_ = ~new_n5635_;
  assign new_n7879_ = ~pi310 | ~new_n6100_;
  assign new_n7880_ = ~new_n6187_ | ~new_n6297_;
  assign new_n7881_ = ~pi311 | ~new_n6100_;
  assign new_n7882_ = ~new_n6187_ | ~new_n6298_;
  assign new_n7883_ = ~pi300 | ~new_n6099_;
  assign new_n7884_ = ~pi309 | ~new_n19121_;
  assign new_n7885_ = ~new_n5640_;
  assign new_n7886_ = ~pi297 | ~new_n6099_;
  assign new_n7887_ = ~pi309 | ~new_n19130_;
  assign new_n7888_ = ~new_n5644_;
  assign new_n7889_ = ~pi298 | ~new_n6099_;
  assign new_n7890_ = ~pi309 | ~new_n19126_;
  assign new_n7891_ = ~new_n5638_;
  assign new_n7892_ = ~pi299 | ~new_n6099_;
  assign new_n7893_ = ~pi309 | ~new_n19123_;
  assign new_n7894_ = ~new_n5639_;
  assign new_n7895_ = ~pi308 | ~new_n6099_;
  assign new_n7896_ = ~pi309 | ~new_n19111_;
  assign new_n7897_ = ~new_n5641_;
  assign new_n7898_ = ~pi307 | ~new_n6099_;
  assign new_n7899_ = ~pi309 | ~new_n19023_;
  assign new_n7900_ = ~new_n5642_;
  assign new_n7901_ = ~pi306 | ~new_n6099_;
  assign new_n7902_ = ~pi309 | ~new_n19114_;
  assign new_n7903_ = ~new_n5643_;
  assign new_n7904_ = ~pi278 | ~new_n6099_;
  assign new_n7905_ = ~pi309 | ~pi278;
  assign new_n7906_ = ~pi305 | ~new_n6099_;
  assign new_n7907_ = ~pi309 | ~new_n19117_;
  assign new_n7908_ = ~new_n5646_;
  assign new_n7909_ = ~new_n1594_ | ~new_n5567_;
  assign new_n7910_ = ~new_n5645_ | ~new_n6165_;
  assign new_n7911_ = ~new_n5647_;
  assign new_n7912_ = ~new_n5640_ | ~new_n7894_;
  assign new_n7913_ = ~new_n7885_ | ~new_n6329_;
  assign new_n7914_ = ~pi311 | ~new_n6296_;
  assign new_n7915_ = ~new_n6298_ | ~new_n5553_;
  assign new_n7916_ = ~new_n5649_;
  assign new_n7917_ = ~new_n7862_ | ~new_n5553_;
  assign new_n7918_ = ~pi310 | ~new_n6296_;
  assign new_n7919_ = ~new_n5648_;
  assign new_n7920_ = ~pi342 | ~new_n6101_;
  assign new_n7921_ = ~new_n6186_ | ~new_n6349_;
  assign new_n7922_ = ~pi279 | ~new_n6099_;
  assign new_n7923_ = ~pi309 | ~new_n19049_;
  assign new_n7924_ = ~new_n1583_ | ~new_n5567_;
  assign new_n7925_ = ~new_n5651_ | ~new_n6165_;
  assign new_n7926_ = ~new_n5652_;
  assign new_n7927_ = ~pi343 | ~new_n6101_;
  assign new_n7928_ = ~new_n6186_ | ~new_n6373_;
  assign new_n7929_ = ~pi280 | ~new_n6099_;
  assign new_n7930_ = ~pi309 | ~new_n19024_;
  assign new_n7931_ = ~new_n1572_ | ~new_n5567_;
  assign new_n7932_ = ~new_n5654_ | ~new_n6165_;
  assign new_n7933_ = ~new_n5655_;
  assign new_n7934_ = ~pi344 | ~new_n6101_;
  assign new_n7935_ = ~new_n6186_ | ~new_n6392_;
  assign new_n7936_ = ~pi281 | ~new_n6099_;
  assign new_n7937_ = ~pi309 | ~new_n19025_;
  assign new_n7938_ = ~new_n1569_ | ~new_n5567_;
  assign new_n7939_ = ~new_n5657_ | ~new_n6165_;
  assign new_n7940_ = ~new_n5658_;
  assign new_n7941_ = ~pi345 | ~new_n6101_;
  assign new_n7942_ = ~new_n6186_ | ~new_n6411_;
  assign new_n7943_ = ~pi282 | ~new_n6099_;
  assign new_n7944_ = ~pi309 | ~new_n19026_;
  assign new_n7945_ = ~new_n1568_ | ~new_n5567_;
  assign new_n7946_ = ~new_n5660_ | ~new_n6165_;
  assign new_n7947_ = ~new_n5661_;
  assign new_n7948_ = ~pi346 | ~new_n6101_;
  assign new_n7949_ = ~new_n6186_ | ~new_n6430_;
  assign new_n7950_ = ~pi283 | ~new_n6099_;
  assign new_n7951_ = ~pi309 | ~new_n19108_;
  assign new_n7952_ = ~new_n1567_ | ~new_n5567_;
  assign new_n7953_ = ~new_n5663_ | ~new_n6165_;
  assign new_n7954_ = ~new_n5664_;
  assign new_n7955_ = ~pi347 | ~new_n6101_;
  assign new_n7956_ = ~new_n6186_ | ~new_n6449_;
  assign new_n7957_ = ~pi284 | ~new_n6099_;
  assign new_n7958_ = ~pi309 | ~new_n19027_;
  assign new_n7959_ = ~new_n1566_ | ~new_n5567_;
  assign new_n7960_ = ~new_n5666_ | ~new_n6165_;
  assign new_n7961_ = ~new_n5667_;
  assign new_n7962_ = ~pi348 | ~new_n6101_;
  assign new_n7963_ = ~new_n6186_ | ~new_n6468_;
  assign new_n7964_ = ~pi285 | ~new_n6099_;
  assign new_n7965_ = ~pi309 | ~new_n19028_;
  assign new_n7966_ = ~new_n1565_ | ~new_n5567_;
  assign new_n7967_ = ~new_n5669_ | ~new_n6165_;
  assign new_n7968_ = ~new_n5670_;
  assign new_n7969_ = ~pi349 | ~new_n6101_;
  assign new_n7970_ = ~new_n6186_ | ~new_n6487_;
  assign new_n7971_ = ~pi286 | ~new_n6099_;
  assign new_n7972_ = ~pi309 | ~new_n19029_;
  assign new_n7973_ = ~new_n1564_ | ~new_n5567_;
  assign new_n7974_ = ~new_n5672_ | ~new_n6165_;
  assign new_n7975_ = ~new_n5673_;
  assign new_n7976_ = ~pi350 | ~new_n6101_;
  assign new_n7977_ = ~new_n6186_ | ~new_n6506_;
  assign new_n7978_ = ~pi287 | ~new_n6099_;
  assign new_n7979_ = ~pi309 | ~new_n19106_;
  assign new_n7980_ = ~new_n1563_ | ~new_n5567_;
  assign new_n7981_ = ~new_n5675_ | ~new_n6165_;
  assign new_n7982_ = ~new_n5676_;
  assign new_n7983_ = ~pi351 | ~new_n6101_;
  assign new_n7984_ = ~new_n6186_ | ~new_n6525_;
  assign new_n7985_ = ~pi288 | ~new_n6099_;
  assign new_n7986_ = ~pi309 | ~new_n19013_;
  assign new_n7987_ = ~new_n1593_ | ~new_n5567_;
  assign new_n7988_ = ~new_n5678_ | ~new_n6165_;
  assign new_n7989_ = ~new_n5679_;
  assign new_n7990_ = ~pi352 | ~new_n6101_;
  assign new_n7991_ = ~new_n6186_ | ~new_n6544_;
  assign new_n7992_ = ~pi289 | ~new_n6099_;
  assign new_n7993_ = ~pi309 | ~new_n19014_;
  assign new_n7994_ = ~new_n1592_ | ~new_n5567_;
  assign new_n7995_ = ~new_n5681_ | ~new_n6165_;
  assign new_n7996_ = ~new_n5682_;
  assign new_n7997_ = ~pi353 | ~new_n6101_;
  assign new_n7998_ = ~new_n6186_ | ~new_n6563_;
  assign new_n7999_ = ~pi290 | ~new_n6099_;
  assign new_n8000_ = ~pi309 | ~new_n19015_;
  assign new_n8001_ = ~new_n1591_ | ~new_n5567_;
  assign new_n8002_ = ~new_n5684_ | ~new_n6165_;
  assign new_n8003_ = ~new_n5685_;
  assign new_n8004_ = ~pi354 | ~new_n6101_;
  assign new_n8005_ = ~new_n6186_ | ~new_n6582_;
  assign new_n8006_ = ~pi291 | ~new_n6099_;
  assign new_n8007_ = ~pi309 | ~new_n19134_;
  assign new_n8008_ = ~new_n1590_ | ~new_n5567_;
  assign new_n8009_ = ~new_n5687_ | ~new_n6165_;
  assign new_n8010_ = ~new_n5688_;
  assign new_n8011_ = ~pi355 | ~new_n6101_;
  assign new_n8012_ = ~new_n6186_ | ~new_n6601_;
  assign new_n8013_ = ~pi292 | ~new_n6099_;
  assign new_n8014_ = ~pi309 | ~new_n19016_;
  assign new_n8015_ = ~new_n1589_ | ~new_n5567_;
  assign new_n8016_ = ~new_n5690_ | ~new_n6165_;
  assign new_n8017_ = ~new_n5691_;
  assign new_n8018_ = ~pi356 | ~new_n6101_;
  assign new_n8019_ = ~new_n6186_ | ~new_n6620_;
  assign new_n8020_ = ~pi293 | ~new_n6099_;
  assign new_n8021_ = ~pi309 | ~new_n19017_;
  assign new_n8022_ = ~new_n1588_ | ~new_n5567_;
  assign new_n8023_ = ~new_n5693_ | ~new_n6165_;
  assign new_n8024_ = ~new_n5694_;
  assign new_n8025_ = ~pi357 | ~new_n6101_;
  assign new_n8026_ = ~new_n6186_ | ~new_n6639_;
  assign new_n8027_ = ~pi294 | ~new_n6099_;
  assign new_n8028_ = ~pi309 | ~new_n19018_;
  assign new_n8029_ = ~new_n1587_ | ~new_n5567_;
  assign new_n8030_ = ~new_n5696_ | ~new_n6165_;
  assign new_n8031_ = ~new_n5697_;
  assign new_n8032_ = ~pi358 | ~new_n6101_;
  assign new_n8033_ = ~new_n6186_ | ~new_n6658_;
  assign new_n8034_ = ~pi295 | ~new_n6099_;
  assign new_n8035_ = ~pi309 | ~new_n19132_;
  assign new_n8036_ = ~new_n1586_ | ~new_n5567_;
  assign new_n8037_ = ~new_n5699_ | ~new_n6165_;
  assign new_n8038_ = ~new_n5700_;
  assign new_n8039_ = ~pi359 | ~new_n6101_;
  assign new_n8040_ = ~new_n6186_ | ~new_n6677_;
  assign new_n8041_ = ~pi296 | ~new_n6099_;
  assign new_n8042_ = ~pi309 | ~new_n19019_;
  assign new_n8043_ = ~new_n1585_ | ~new_n5567_;
  assign new_n8044_ = ~new_n5702_ | ~new_n6165_;
  assign new_n8045_ = ~new_n5703_;
  assign new_n8046_ = ~pi360 | ~new_n6101_;
  assign new_n8047_ = ~new_n6186_ | ~new_n6696_;
  assign new_n8048_ = ~new_n1584_ | ~new_n5567_;
  assign new_n8049_ = ~new_n5644_ | ~new_n6165_;
  assign new_n8050_ = ~new_n5705_;
  assign new_n8051_ = ~pi361 | ~new_n6101_;
  assign new_n8052_ = ~new_n6186_ | ~new_n6715_;
  assign new_n8053_ = ~pi362 | ~new_n6101_;
  assign new_n8054_ = ~new_n6186_ | ~new_n6734_;
  assign new_n8055_ = ~pi363 | ~new_n6101_;
  assign new_n8056_ = ~new_n6186_ | ~new_n6753_;
  assign new_n8057_ = ~pi364 | ~new_n6101_;
  assign new_n8058_ = ~new_n6186_ | ~new_n6772_;
  assign new_n8059_ = ~pi365 | ~new_n6101_;
  assign new_n8060_ = ~new_n6186_ | ~new_n6791_;
  assign new_n8061_ = ~pi366 | ~new_n6101_;
  assign new_n8062_ = ~new_n6186_ | ~new_n6810_;
  assign new_n8063_ = ~pi367 | ~new_n6101_;
  assign new_n8064_ = ~new_n6186_ | ~new_n6829_;
  assign new_n8065_ = ~pi368 | ~new_n6101_;
  assign new_n8066_ = ~new_n6186_ | ~new_n6848_;
  assign new_n8067_ = ~pi369 | ~new_n6101_;
  assign new_n8068_ = ~new_n6186_ | ~new_n6867_;
  assign new_n8069_ = ~pi370 | ~new_n6101_;
  assign new_n8070_ = ~new_n6186_ | ~new_n6886_;
  assign new_n8071_ = ~pi371 | ~new_n6101_;
  assign new_n8072_ = ~new_n6186_ | ~new_n6906_;
  assign new_n8073_ = ~pi372 | ~new_n6101_;
  assign new_n8074_ = ~new_n6186_ | ~new_n6913_;
  assign new_n8075_ = ~pi373 | ~new_n6101_;
  assign new_n8076_ = ~new_n6186_ | ~new_n6916_;
  assign new_n8077_ = ~pi374 | ~new_n6102_;
  assign new_n8078_ = ~new_n6185_ | ~new_n6349_;
  assign new_n8079_ = ~pi375 | ~new_n6102_;
  assign new_n8080_ = ~new_n6185_ | ~new_n6373_;
  assign new_n8081_ = ~pi376 | ~new_n6102_;
  assign new_n8082_ = ~new_n6185_ | ~new_n6392_;
  assign new_n8083_ = ~pi377 | ~new_n6102_;
  assign new_n8084_ = ~new_n6185_ | ~new_n6411_;
  assign new_n8085_ = ~pi378 | ~new_n6102_;
  assign new_n8086_ = ~new_n6185_ | ~new_n6430_;
  assign new_n8087_ = ~pi379 | ~new_n6102_;
  assign new_n8088_ = ~new_n6185_ | ~new_n6449_;
  assign new_n8089_ = ~pi380 | ~new_n6102_;
  assign new_n8090_ = ~new_n6185_ | ~new_n6468_;
  assign new_n8091_ = ~pi381 | ~new_n6102_;
  assign new_n8092_ = ~new_n6185_ | ~new_n6487_;
  assign new_n8093_ = ~pi382 | ~new_n6102_;
  assign new_n8094_ = ~new_n6185_ | ~new_n6506_;
  assign new_n8095_ = ~pi383 | ~new_n6102_;
  assign new_n8096_ = ~new_n6185_ | ~new_n6525_;
  assign new_n8097_ = ~pi384 | ~new_n6102_;
  assign new_n8098_ = ~new_n6185_ | ~new_n6544_;
  assign new_n8099_ = ~pi385 | ~new_n6102_;
  assign new_n8100_ = ~new_n6185_ | ~new_n6563_;
  assign new_n8101_ = ~pi386 | ~new_n6102_;
  assign new_n8102_ = ~new_n6185_ | ~new_n6582_;
  assign new_n8103_ = ~pi387 | ~new_n6102_;
  assign new_n8104_ = ~new_n6185_ | ~new_n6601_;
  assign new_n8105_ = ~pi388 | ~new_n6102_;
  assign new_n8106_ = ~new_n6185_ | ~new_n6620_;
  assign new_n8107_ = ~pi389 | ~new_n6102_;
  assign new_n8108_ = ~new_n6185_ | ~new_n6639_;
  assign new_n8109_ = ~pi390 | ~new_n6102_;
  assign new_n8110_ = ~new_n6185_ | ~new_n6658_;
  assign new_n8111_ = ~pi391 | ~new_n6102_;
  assign new_n8112_ = ~new_n6185_ | ~new_n6677_;
  assign new_n8113_ = ~pi392 | ~new_n6102_;
  assign new_n8114_ = ~new_n6185_ | ~new_n6696_;
  assign new_n8115_ = ~pi393 | ~new_n6102_;
  assign new_n8116_ = ~new_n6185_ | ~new_n6715_;
  assign new_n8117_ = ~pi394 | ~new_n6102_;
  assign new_n8118_ = ~new_n6185_ | ~new_n6734_;
  assign new_n8119_ = ~pi395 | ~new_n6102_;
  assign new_n8120_ = ~new_n6185_ | ~new_n6753_;
  assign new_n8121_ = ~pi396 | ~new_n6102_;
  assign new_n8122_ = ~new_n6185_ | ~new_n6772_;
  assign new_n8123_ = ~pi397 | ~new_n6102_;
  assign new_n8124_ = ~new_n6185_ | ~new_n6791_;
  assign new_n8125_ = ~pi398 | ~new_n6102_;
  assign new_n8126_ = ~new_n6185_ | ~new_n6810_;
  assign new_n8127_ = ~pi399 | ~new_n6102_;
  assign new_n8128_ = ~new_n6185_ | ~new_n6829_;
  assign new_n8129_ = ~pi400 | ~new_n6102_;
  assign new_n8130_ = ~new_n6185_ | ~new_n6848_;
  assign new_n8131_ = ~pi401 | ~new_n6102_;
  assign new_n8132_ = ~new_n6185_ | ~new_n6867_;
  assign new_n8133_ = ~pi402 | ~new_n6102_;
  assign new_n8134_ = ~new_n6185_ | ~new_n6886_;
  assign new_n8135_ = ~pi403 | ~new_n6102_;
  assign new_n8136_ = ~new_n6185_ | ~new_n6906_;
  assign new_n8137_ = ~pi404 | ~new_n6102_;
  assign new_n8138_ = ~new_n6185_ | ~new_n6913_;
  assign new_n8139_ = ~pi405 | ~new_n6102_;
  assign new_n8140_ = ~new_n6185_ | ~new_n6916_;
  assign new_n8141_ = ~pi406 | ~new_n5611_;
  assign new_n8142_ = ~new_n6184_ | ~new_n5568_;
  assign new_n8143_ = ~pi407 | ~new_n5611_;
  assign new_n8144_ = ~new_n6184_ | ~new_n5569_;
  assign new_n8145_ = ~pi408 | ~new_n5611_;
  assign new_n8146_ = ~new_n6184_ | ~new_n5570_;
  assign new_n8147_ = ~pi409 | ~new_n5611_;
  assign new_n8148_ = ~new_n6184_ | ~new_n5571_;
  assign new_n8149_ = ~pi410 | ~new_n5611_;
  assign new_n8150_ = ~new_n6184_ | ~new_n5572_;
  assign new_n8151_ = ~pi411 | ~new_n5611_;
  assign new_n8152_ = ~new_n6184_ | ~new_n5573_;
  assign new_n8153_ = ~pi412 | ~new_n5611_;
  assign new_n8154_ = ~new_n6184_ | ~new_n5574_;
  assign new_n8155_ = ~pi413 | ~new_n5611_;
  assign new_n8156_ = ~new_n6184_ | ~new_n5575_;
  assign new_n8157_ = ~pi414 | ~new_n5611_;
  assign new_n8158_ = ~new_n6184_ | ~new_n5576_;
  assign new_n8159_ = ~pi415 | ~new_n5611_;
  assign new_n8160_ = ~new_n6184_ | ~new_n5577_;
  assign new_n8161_ = ~pi416 | ~new_n5611_;
  assign new_n8162_ = ~new_n6184_ | ~new_n5578_;
  assign new_n8163_ = ~pi417 | ~new_n5611_;
  assign new_n8164_ = ~new_n6184_ | ~new_n5579_;
  assign new_n8165_ = ~pi418 | ~new_n5611_;
  assign new_n8166_ = ~new_n6184_ | ~new_n5580_;
  assign new_n8167_ = ~pi419 | ~new_n5611_;
  assign new_n8168_ = ~new_n6184_ | ~new_n5581_;
  assign new_n8169_ = ~pi420 | ~new_n5611_;
  assign new_n8170_ = ~new_n6184_ | ~new_n5582_;
  assign new_n8171_ = ~pi421 | ~new_n5611_;
  assign new_n8172_ = ~new_n6184_ | ~new_n5583_;
  assign new_n8173_ = ~pi422 | ~new_n5611_;
  assign new_n8174_ = ~new_n6184_ | ~new_n5584_;
  assign new_n8175_ = ~pi423 | ~new_n5611_;
  assign new_n8176_ = ~new_n6184_ | ~new_n5585_;
  assign new_n8177_ = ~pi424 | ~new_n5611_;
  assign new_n8178_ = ~new_n6184_ | ~new_n5586_;
  assign new_n8179_ = ~pi425 | ~new_n5611_;
  assign new_n8180_ = ~new_n6184_ | ~new_n5587_;
  assign new_n8181_ = ~pi426 | ~new_n5611_;
  assign new_n8182_ = ~new_n6184_ | ~new_n5589_;
  assign new_n8183_ = ~pi427 | ~new_n5611_;
  assign new_n8184_ = ~new_n6184_ | ~new_n5591_;
  assign new_n8185_ = ~pi428 | ~new_n5611_;
  assign new_n8186_ = ~new_n6184_ | ~new_n5593_;
  assign new_n8187_ = ~pi429 | ~new_n5611_;
  assign new_n8188_ = ~new_n6184_ | ~new_n5595_;
  assign new_n8189_ = ~pi430 | ~new_n5611_;
  assign new_n8190_ = ~new_n6184_ | ~new_n5597_;
  assign new_n8191_ = ~pi431 | ~new_n5611_;
  assign new_n8192_ = ~new_n6184_ | ~new_n5599_;
  assign new_n8193_ = ~pi432 | ~new_n5611_;
  assign new_n8194_ = ~new_n6184_ | ~new_n5601_;
  assign new_n8195_ = ~pi433 | ~new_n5611_;
  assign new_n8196_ = ~new_n6184_ | ~new_n5603_;
  assign new_n8197_ = ~pi434 | ~new_n5611_;
  assign new_n8198_ = ~new_n6184_ | ~new_n5605_;
  assign new_n8199_ = ~pi435 | ~new_n5611_;
  assign new_n8200_ = ~new_n6184_ | ~new_n5607_;
  assign new_n8201_ = ~pi436 | ~new_n5611_;
  assign new_n8202_ = ~new_n6188_ | ~new_n6184_;
  assign new_n8203_ = ~pi437 | ~new_n5611_;
  assign new_n8204_ = ~new_n6188_ | ~new_n6184_;
  assign new_n8205_ = ~pi458 | ~new_n5620_;
  assign new_n8206_ = ~po511 | ~new_n5299_;
  assign new_n8207_ = ~pi459 | ~new_n5620_;
  assign new_n8208_ = ~po511 | ~new_n5300_;
  assign new_n8209_ = ~pi460 | ~new_n5620_;
  assign new_n8210_ = ~po511 | ~new_n5290_;
  assign new_n8211_ = ~pi461 | ~new_n5620_;
  assign new_n8212_ = ~po511 | ~new_n5286_;
  assign new_n8213_ = ~pi462 | ~new_n5620_;
  assign new_n8214_ = ~po511 | ~new_n5282_;
  assign new_n8215_ = ~pi463 | ~new_n5620_;
  assign new_n8216_ = ~po511 | ~new_n5289_;
  assign new_n8217_ = ~pi464 | ~new_n5620_;
  assign new_n8218_ = ~po511 | ~new_n5293_;
  assign new_n8219_ = ~pi465 | ~new_n5620_;
  assign new_n8220_ = ~po511 | ~new_n5292_;
  assign new_n8221_ = ~pi466 | ~new_n5620_;
  assign new_n8222_ = ~po511 | ~new_n5306_;
  assign new_n8223_ = ~pi467 | ~new_n5620_;
  assign new_n8224_ = ~po511 | ~new_n5305_;
  assign new_n8225_ = ~pi468 | ~new_n5620_;
  assign new_n8226_ = ~po511 | ~new_n5284_;
  assign new_n8227_ = ~pi469 | ~new_n5620_;
  assign new_n8228_ = ~po511 | ~new_n5285_;
  assign new_n8229_ = ~pi470 | ~new_n5620_;
  assign new_n8230_ = ~po511 | ~new_n5294_;
  assign new_n8231_ = ~pi471 | ~new_n5620_;
  assign new_n8232_ = ~po511 | ~new_n5302_;
  assign new_n8233_ = ~pi472 | ~new_n5620_;
  assign new_n8234_ = ~po511 | ~new_n5301_;
  assign new_n8235_ = ~pi473 | ~new_n5620_;
  assign new_n8236_ = ~po511 | ~new_n5296_;
  assign new_n8237_ = ~pi474 | ~new_n5620_;
  assign new_n8238_ = ~po511 | ~new_n5295_;
  assign new_n8239_ = ~pi475 | ~new_n5620_;
  assign new_n8240_ = ~po511 | ~new_n5291_;
  assign new_n8241_ = ~pi476 | ~new_n5620_;
  assign new_n8242_ = ~po511 | ~new_n5304_;
  assign new_n8243_ = ~pi477 | ~new_n5620_;
  assign new_n8244_ = ~po511 | ~new_n5303_;
  assign new_n8245_ = ~pi478 | ~new_n5620_;
  assign new_n8246_ = ~po511 | ~new_n5298_;
  assign new_n8247_ = ~pi479 | ~new_n5620_;
  assign new_n8248_ = ~po511 | ~new_n5297_;
  assign new_n8249_ = ~pi480 | ~new_n5620_;
  assign new_n8250_ = ~po511 | ~new_n5283_;
  assign new_n8251_ = ~pi481 | ~new_n5620_;
  assign new_n8252_ = ~po511 | ~new_n5288_;
  assign new_n8253_ = ~pi482 | ~new_n5620_;
  assign new_n8254_ = ~po511 | ~new_n5287_;
  assign new_n8255_ = ~pi483 | ~new_n5620_;
  assign new_n8256_ = ~po511 | ~new_n5280_;
  assign new_n8257_ = ~pi484 | ~new_n5620_;
  assign new_n8258_ = ~po511 | ~new_n5279_;
  assign new_n8259_ = ~pi485 | ~new_n5620_;
  assign new_n8260_ = ~po511 | ~new_n5275_;
  assign new_n8261_ = ~pi486 | ~new_n5620_;
  assign new_n8262_ = ~po511 | ~new_n5276_;
  assign new_n8263_ = ~pi487 | ~new_n5620_;
  assign new_n8264_ = ~po511 | ~new_n5277_;
  assign new_n8265_ = ~pi488 | ~new_n5620_;
  assign new_n8266_ = ~po511 | ~new_n5281_;
  assign new_n8267_ = ~pi489 | ~new_n5620_;
  assign new_n8268_ = ~po511 | ~new_n5278_;
  assign new_n8269_ = ~new_n19224_ | ~new_n7377_;
  assign new_n8270_ = ~new_n7381_ | ~new_n6136_;
  assign new_n8271_ = ~new_n7878_ | ~new_n5623_;
  assign new_n8272_ = ~new_n5640_ | ~new_n5635_;
  assign new_n8273_ = ~new_n6180_ | ~new_n5277_;
  assign new_n8274_ = ~new_n5606_ | ~new_n6872_;
  assign new_n8275_ = ~new_n8274_ | ~new_n8273_;
  assign new_n8276_ = ~new_n6169_ | ~new_n5276_;
  assign new_n8277_ = ~new_n5604_ | ~new_n6853_;
  assign new_n8278_ = ~new_n8277_ | ~new_n8276_;
  assign new_n8279_ = ~new_n6170_ | ~new_n5275_;
  assign new_n8280_ = ~new_n5602_ | ~new_n6834_;
  assign new_n8281_ = ~new_n8280_ | ~new_n8279_;
  assign new_n8282_ = ~new_n6173_ | ~new_n5287_;
  assign new_n8283_ = ~new_n5596_ | ~new_n6777_;
  assign new_n8284_ = ~new_n8283_ | ~new_n8282_;
  assign new_n8285_ = ~new_n6174_ | ~new_n5288_;
  assign new_n8286_ = ~new_n5594_ | ~new_n6758_;
  assign new_n8287_ = ~new_n8286_ | ~new_n8285_;
  assign new_n8288_ = ~new_n6176_ | ~new_n5297_;
  assign new_n8289_ = ~new_n5590_ | ~new_n6720_;
  assign new_n8290_ = ~new_n8289_ | ~new_n8288_;
  assign new_n8291_ = ~new_n6175_ | ~new_n5283_;
  assign new_n8292_ = ~new_n5592_ | ~new_n6739_;
  assign new_n8293_ = ~new_n8292_ | ~new_n8291_;
  assign new_n8294_ = ~new_n6172_ | ~new_n5280_;
  assign new_n8295_ = ~new_n5598_ | ~new_n6796_;
  assign new_n8296_ = ~new_n8295_ | ~new_n8294_;
  assign new_n8297_ = ~new_n6171_ | ~new_n5279_;
  assign new_n8298_ = ~new_n5600_ | ~new_n6815_;
  assign new_n8299_ = ~new_n8298_ | ~new_n8297_;
  assign new_n8300_ = ~new_n6179_ | ~new_n5281_;
  assign new_n8301_ = ~new_n5608_ | ~new_n6890_;
  assign new_n8302_ = ~new_n8301_ | ~new_n8300_;
  assign new_n8303_ = ~new_n6178_ | ~new_n5278_;
  assign new_n8304_ = ~new_n5609_ | ~new_n6910_;
  assign new_n8305_ = ~new_n8304_ | ~new_n8303_;
  assign new_n8306_ = ~new_n8017_ | ~new_n6587_;
  assign new_n8307_ = ~new_n5691_ | ~new_n5301_;
  assign new_n8308_ = ~new_n8307_ | ~new_n8306_;
  assign new_n8309_ = ~new_n7926_ | ~new_n6335_;
  assign new_n8310_ = ~new_n5652_ | ~new_n5300_;
  assign new_n8311_ = ~new_n8310_ | ~new_n8309_;
  assign new_n8312_ = ~new_n7911_ | ~new_n6359_;
  assign new_n8313_ = ~new_n5647_ | ~new_n5299_;
  assign new_n8314_ = ~new_n8313_ | ~new_n8312_;
  assign new_n8315_ = ~new_n8024_ | ~new_n6606_;
  assign new_n8316_ = ~new_n5694_ | ~new_n5296_;
  assign new_n8317_ = ~new_n8316_ | ~new_n8315_;
  assign new_n8318_ = ~new_n7975_ | ~new_n6473_;
  assign new_n8319_ = ~new_n5673_ | ~new_n5306_;
  assign new_n8320_ = ~new_n8319_ | ~new_n8318_;
  assign new_n8321_ = ~new_n7982_ | ~new_n6492_;
  assign new_n8322_ = ~new_n5676_ | ~new_n5305_;
  assign new_n8323_ = ~new_n8322_ | ~new_n8321_;
  assign new_n8324_ = ~new_n8010_ | ~new_n6568_;
  assign new_n8325_ = ~new_n5688_ | ~new_n5302_;
  assign new_n8326_ = ~new_n8325_ | ~new_n8324_;
  assign new_n8327_ = ~new_n8045_ | ~new_n6663_;
  assign new_n8328_ = ~new_n5703_ | ~new_n5304_;
  assign new_n8329_ = ~new_n8328_ | ~new_n8327_;
  assign new_n8330_ = ~new_n8031_ | ~new_n6625_;
  assign new_n8331_ = ~new_n5697_ | ~new_n5295_;
  assign new_n8332_ = ~new_n8331_ | ~new_n8330_;
  assign new_n8333_ = ~new_n8003_ | ~new_n6549_;
  assign new_n8334_ = ~new_n5685_ | ~new_n5294_;
  assign new_n8335_ = ~new_n8334_ | ~new_n8333_;
  assign new_n8336_ = ~new_n7961_ | ~new_n6435_;
  assign new_n8337_ = ~new_n5667_ | ~new_n5293_;
  assign new_n8338_ = ~new_n8337_ | ~new_n8336_;
  assign new_n8339_ = ~new_n7968_ | ~new_n6454_;
  assign new_n8340_ = ~new_n5670_ | ~new_n5292_;
  assign new_n8341_ = ~new_n8340_ | ~new_n8339_;
  assign new_n8342_ = ~new_n7954_ | ~new_n6416_;
  assign new_n8343_ = ~new_n5664_ | ~new_n5289_;
  assign new_n8344_ = ~new_n8343_ | ~new_n8342_;
  assign new_n8345_ = ~new_n7940_ | ~new_n6378_;
  assign new_n8346_ = ~new_n5658_ | ~new_n5286_;
  assign new_n8347_ = ~new_n8346_ | ~new_n8345_;
  assign new_n8348_ = ~new_n7933_ | ~new_n6354_;
  assign new_n8349_ = ~new_n5655_ | ~new_n5290_;
  assign new_n8350_ = ~new_n8349_ | ~new_n8348_;
  assign new_n8351_ = ~new_n8038_ | ~new_n6644_;
  assign new_n8352_ = ~new_n5700_ | ~new_n5291_;
  assign new_n8353_ = ~new_n8352_ | ~new_n8351_;
  assign new_n8354_ = ~new_n8050_ | ~new_n6682_;
  assign new_n8355_ = ~new_n5705_ | ~new_n5303_;
  assign new_n8356_ = ~new_n8355_ | ~new_n8354_;
  assign new_n8357_ = ~new_n7947_ | ~new_n6397_;
  assign new_n8358_ = ~new_n5661_ | ~new_n5282_;
  assign new_n8359_ = ~new_n8358_ | ~new_n8357_;
  assign new_n8360_ = ~new_n7996_ | ~new_n6530_;
  assign new_n8361_ = ~new_n5682_ | ~new_n5285_;
  assign new_n8362_ = ~new_n8361_ | ~new_n8360_;
  assign new_n8363_ = ~new_n7989_ | ~new_n6511_;
  assign new_n8364_ = ~new_n5679_ | ~new_n5284_;
  assign new_n8365_ = ~new_n8364_ | ~new_n8363_;
  assign new_n8366_ = ~new_n6177_ | ~new_n5298_;
  assign new_n8367_ = ~new_n5588_ | ~new_n6701_;
  assign new_n8368_ = ~new_n8367_ | ~new_n8366_;
  assign new_n8369_ = ~new_n6160_ | ~new_n7376_;
  assign new_n8370_ = ~new_n6162_ | ~new_n6138_;
  assign new_n8371_ = ~new_n8446_ | ~new_n30318_;
  assign new_n8372_ = ~new_n30528_ | ~new_n8374_;
  assign new_n8373_ = ~new_n30618_ | ~new_n30420_;
  assign new_n8374_ = ~new_n8375_ | ~new_n8376_;
  assign new_n8375_ = ~new_n8821_ | ~new_n30334_;
  assign new_n8376_ = ~new_n8459_ | ~new_n30333_;
  assign new_n8377_ = ~new_n8379_ | ~new_n30574_;
  assign new_n8378_ = ~new_n30617_ | ~new_n30349_;
  assign new_n8379_ = ~new_n8380_ | ~new_n8381_;
  assign new_n8380_ = ~new_n8823_ | ~new_n30337_;
  assign new_n8381_ = ~new_n8458_ | ~new_n30336_;
  assign new_n8382_ = ~new_n30586_ | ~new_n30289_;
  assign new_n8383_ = ~new_n30440_ | ~new_n30419_;
  assign new_n8384_ = ~new_n9285_ | ~new_n30348_;
  assign new_n8385_ = ~new_n8453_ | ~new_n30339_;
  assign new_n8386_ = ~new_n8387_ | ~new_n8388_;
  assign new_n8387_ = ~new_n9284_ | ~new_n30313_;
  assign new_n8388_ = ~new_n8452_ | ~new_n30312_;
  assign new_n8389_ = ~new_n9284_ | ~new_n30313_;
  assign new_n8390_ = ~new_n8452_ | ~new_n30312_;
  assign new_n8391_ = new_n8758_ & new_n10828_;
  assign new_n8392_ = new_n8758_ & new_n8757_;
  assign new_n8393_ = new_n10831_ & new_n8757_;
  assign new_n8394_ = new_n10831_ & new_n10828_;
  assign new_n8395_ = new_n9252_ & new_n10825_;
  assign new_n8396_ = new_n8965_ & new_n8960_;
  assign new_n8397_ = new_n8759_ & new_n8760_;
  assign new_n8398_ = new_n10840_ & new_n8759_;
  assign new_n8399_ = new_n10837_ & new_n8760_;
  assign new_n8400_ = new_n10840_ & new_n10837_;
  assign new_n8401_ = new_n8424_ & pi765;
  assign new_n8402_ = new_n9074_ & new_n8744_;
  assign new_n8403_ = new_n9289_ & new_n9451_;
  assign new_n8404_ = new_n8393_ & new_n10825_;
  assign new_n8405_ = new_n8675_ & pi765;
  assign new_n8406_ = new_n9264_ & new_n9290_;
  assign new_n8407_ = new_n9290_ & new_n8743_;
  assign new_n8408_ = new_n9071_ & new_n9290_;
  assign new_n8409_ = new_n9268_ & new_n8401_;
  assign new_n8410_ = new_n9273_ & new_n9451_;
  assign new_n8411_ = new_n9289_ & new_n9467_;
  assign new_n8412_ = new_n9290_ & new_n8403_;
  assign new_n8413_ = new_n8401_ & new_n10367_;
  assign new_n8414_ = new_n9273_ & new_n9467_;
  assign new_n8415_ = new_n10846_ & new_n10132_;
  assign new_n8416_ = new_n8402_ & new_n10846_;
  assign new_n8417_ = new_n10843_ & new_n10132_;
  assign new_n8418_ = new_n9270_ & new_n10132_;
  assign new_n8419_ = new_n8402_ & new_n9270_;
  assign new_n8420_ = new_n8401_ & new_n8744_;
  assign new_n8421_ = new_n8401_ & new_n8743_;
  assign new_n8422_ = new_n10382_ & pi765;
  assign new_n8423_ = new_n8401_ & new_n10384_;
  assign new_n8424_ = new_n10818_ & new_n8740_;
  assign new_n8425_ = new_n9070_ & new_n8396_;
  assign new_n8426_ = new_n9069_ & new_n8396_;
  assign new_n8427_ = new_n10127_ & new_n10126_;
  assign new_n8428_ = new_n10137_ & pi765;
  assign new_n8429_ = po756 & new_n10139_;
  assign new_n8430_ = ~new_n9915_ | ~new_n9916_ | ~new_n9913_ | ~new_n9914_;
  assign new_n8431_ = ~new_n9933_ | ~new_n9931_ | ~new_n9932_ | ~new_n9934_;
  assign new_n8432_ = ~new_n9951_ | ~new_n9949_ | ~new_n9950_ | ~new_n9952_;
  assign new_n8433_ = ~new_n9989_ | ~new_n9987_ | ~new_n9988_ | ~new_n9990_;
  assign new_n8434_ = ~new_n9897_ | ~new_n9895_ | ~new_n9896_ | ~new_n9898_;
  assign new_n8435_ = ~new_n9879_ | ~new_n9877_ | ~new_n9878_ | ~new_n9880_;
  assign new_n8436_ = ~new_n9969_ | ~new_n9967_ | ~new_n9968_ | ~new_n9970_;
  assign new_n8437_ = ~new_n9501_ | ~new_n9499_ | ~new_n9500_ | ~new_n9502_;
  assign new_n8438_ = ~new_n9825_ | ~new_n9823_ | ~new_n9824_ | ~new_n9826_;
  assign new_n8439_ = ~new_n9609_ | ~new_n9607_ | ~new_n9608_ | ~new_n9610_;
  assign new_n8440_ = ~new_n9627_ | ~new_n9625_ | ~new_n9626_ | ~new_n9628_;
  assign new_n8441_ = ~new_n9483_ | ~new_n9481_ | ~new_n9482_ | ~new_n9484_;
  assign new_n8442_ = ~new_n9861_ | ~new_n9859_ | ~new_n9860_ | ~new_n9862_;
  assign new_n8443_ = ~new_n9843_ | ~new_n9841_ | ~new_n9842_ | ~new_n9844_;
  assign new_n8444_ = ~new_n9519_ | ~new_n9517_ | ~new_n9518_ | ~new_n9520_;
  assign new_n8445_ = ~new_n9458_ | ~new_n9456_ | ~new_n9457_ | ~new_n9459_;
  assign new_n8446_ = ~new_n9735_ | ~new_n9733_ | ~new_n9734_ | ~new_n9736_;
  assign new_n8447_ = ~new_n9555_ | ~new_n9553_ | ~new_n9554_ | ~new_n9556_;
  assign new_n8448_ = ~new_n9537_ | ~new_n9535_ | ~new_n9536_ | ~new_n9538_;
  assign new_n8449_ = ~new_n9645_ | ~new_n9643_ | ~new_n9644_ | ~new_n9646_;
  assign new_n8450_ = ~new_n9717_ | ~new_n9715_ | ~new_n9716_ | ~new_n9718_;
  assign new_n8451_ = ~new_n9699_ | ~new_n9697_ | ~new_n9698_ | ~new_n9700_;
  assign new_n8452_ = ~new_n9807_ | ~new_n9805_ | ~new_n9806_ | ~new_n9808_;
  assign new_n8453_ = ~new_n9789_ | ~new_n9787_ | ~new_n9788_ | ~new_n9790_;
  assign new_n8454_ = ~new_n9463_ | ~new_n9461_ | ~new_n9462_ | ~new_n9464_;
  assign new_n8455_ = ~new_n9439_ | ~new_n9437_ | ~new_n9438_ | ~new_n9440_;
  assign new_n8456_ = ~new_n9681_ | ~new_n9679_ | ~new_n9680_ | ~new_n9682_;
  assign new_n8457_ = ~new_n9663_ | ~new_n9661_ | ~new_n9662_ | ~new_n9664_;
  assign new_n8458_ = ~new_n9771_ | ~new_n9769_ | ~new_n9770_ | ~new_n9772_;
  assign new_n8459_ = ~new_n9753_ | ~new_n9751_ | ~new_n9752_ | ~new_n9754_;
  assign new_n8460_ = ~new_n9591_ | ~new_n9589_ | ~new_n9590_ | ~new_n9592_;
  assign new_n8461_ = ~new_n9573_ | ~new_n9571_ | ~new_n9572_ | ~new_n9574_;
  assign new_n8462_ = ~new_n10719_ | ~new_n10718_;
  assign new_n8463_ = ~new_n10721_ | ~new_n10720_;
  assign new_n8464_ = ~new_n10726_ | ~new_n10727_ | ~new_n10725_;
  assign new_n8465_ = ~new_n10729_ | ~new_n10730_ | ~new_n10728_;
  assign new_n8466_ = ~new_n10732_ | ~new_n10733_ | ~new_n10731_;
  assign new_n8467_ = ~new_n10735_ | ~new_n10736_ | ~new_n10734_;
  assign new_n8468_ = ~new_n10738_ | ~new_n10739_ | ~new_n10737_;
  assign new_n8469_ = ~new_n10741_ | ~new_n10742_ | ~new_n10740_;
  assign new_n8470_ = ~new_n10744_ | ~new_n10745_ | ~new_n10743_;
  assign new_n8471_ = ~new_n10747_ | ~new_n10748_ | ~new_n10746_;
  assign new_n8472_ = ~new_n10750_ | ~new_n10751_ | ~new_n10749_;
  assign new_n8473_ = ~new_n10753_ | ~new_n10754_ | ~new_n10752_;
  assign new_n8474_ = ~new_n10758_ | ~new_n10759_ | ~new_n10760_;
  assign new_n8475_ = ~new_n10761_ | ~new_n10762_ | ~new_n10763_;
  assign new_n8476_ = ~new_n10764_ | ~new_n10765_ | ~new_n10766_;
  assign new_n8477_ = ~new_n10767_ | ~new_n10768_ | ~new_n10769_;
  assign new_n8478_ = ~new_n10770_ | ~new_n10771_ | ~new_n10772_;
  assign new_n8479_ = ~new_n10773_ | ~new_n10774_ | ~new_n10775_;
  assign new_n8480_ = ~new_n10778_ | ~new_n10777_ | ~new_n10776_;
  assign new_n8481_ = ~new_n10781_ | ~new_n10780_ | ~new_n10779_;
  assign new_n8482_ = ~new_n10784_ | ~new_n10783_ | ~new_n10782_;
  assign new_n8483_ = ~new_n10787_ | ~new_n10786_ | ~new_n10785_;
  assign new_n8484_ = ~new_n10702_ | ~new_n10701_ | ~new_n10700_;
  assign new_n8485_ = ~new_n10705_ | ~new_n10704_ | ~new_n10703_;
  assign new_n8486_ = ~new_n10708_ | ~new_n10707_ | ~new_n10706_;
  assign new_n8487_ = ~new_n10711_ | ~new_n10710_ | ~new_n10709_;
  assign new_n8488_ = ~new_n10714_ | ~new_n10713_ | ~new_n10712_;
  assign new_n8489_ = ~new_n10717_ | ~new_n10716_ | ~new_n10715_;
  assign new_n8490_ = ~new_n10724_ | ~new_n10723_ | ~new_n10722_;
  assign new_n8491_ = ~new_n10757_ | ~new_n10756_ | ~new_n10755_;
  assign new_n8492_ = ~new_n10790_ | ~new_n10789_ | ~new_n10788_;
  assign new_n8493_ = ~new_n10792_ | ~new_n10791_;
  assign new_n8494_ = ~new_n10649_ | ~new_n10648_;
  assign new_n8495_ = ~new_n10651_ | ~new_n10650_;
  assign new_n8496_ = ~new_n10654_ | ~new_n10655_ | ~new_n8753_;
  assign new_n8497_ = ~new_n10656_ | ~new_n10657_ | ~new_n8753_;
  assign new_n8498_ = ~new_n10658_ | ~new_n10659_ | ~new_n8753_;
  assign new_n8499_ = ~new_n10660_ | ~new_n10661_ | ~new_n8753_;
  assign new_n8500_ = ~new_n10662_ | ~new_n10663_ | ~new_n8753_;
  assign new_n8501_ = ~new_n10664_ | ~new_n10665_ | ~new_n8753_;
  assign new_n8502_ = ~new_n10666_ | ~new_n10667_ | ~new_n8753_;
  assign new_n8503_ = ~new_n10668_ | ~new_n10669_ | ~new_n8753_;
  assign new_n8504_ = ~new_n10670_ | ~new_n10671_ | ~new_n8753_;
  assign new_n8505_ = ~new_n10672_ | ~new_n10673_ | ~new_n8753_;
  assign new_n8506_ = ~new_n10676_ | ~new_n10677_ | ~new_n8753_;
  assign new_n8507_ = ~new_n10678_ | ~new_n10679_ | ~new_n8753_;
  assign new_n8508_ = ~new_n10680_ | ~new_n10681_ | ~new_n8753_;
  assign new_n8509_ = ~new_n10682_ | ~new_n10683_ | ~new_n8753_;
  assign new_n8510_ = ~new_n10684_ | ~new_n10685_ | ~new_n8753_;
  assign new_n8511_ = ~new_n10686_ | ~new_n10687_ | ~new_n8753_;
  assign new_n8512_ = ~new_n9203_ | ~new_n10689_;
  assign new_n8513_ = ~new_n9204_ | ~new_n10691_;
  assign new_n8514_ = ~new_n9205_ | ~new_n10693_;
  assign new_n8515_ = ~new_n9206_ | ~new_n10695_;
  assign new_n8516_ = ~new_n9195_ | ~new_n10637_;
  assign new_n8517_ = ~new_n9196_ | ~new_n10639_;
  assign new_n8518_ = ~new_n9197_ | ~new_n10641_;
  assign new_n8519_ = ~new_n9198_ | ~new_n10643_;
  assign new_n8520_ = ~new_n9199_ | ~new_n10645_;
  assign new_n8521_ = ~new_n9200_ | ~new_n10647_;
  assign new_n8522_ = ~new_n9201_ | ~new_n10653_;
  assign new_n8523_ = ~new_n9202_ | ~new_n10675_;
  assign new_n8524_ = ~new_n9207_ | ~new_n10697_;
  assign new_n8525_ = ~new_n9208_ | ~new_n10699_;
  assign new_n8526_ = ~new_n8753_ | ~new_n8763_ | ~new_n10831_;
  assign new_n8527_ = ~new_n9191_ | ~new_n8391_;
  assign po755 = ~new_n9190_ | ~new_n10631_;
  assign po754 = ~pi765;
  assign new_n8530_ = ~new_n8737_ | ~new_n11322_ | ~new_n11321_;
  assign po753 = ~new_n10626_ | ~new_n10628_ | ~new_n9189_ | ~new_n10627_;
  assign po752 = ~new_n9188_ | ~new_n10619_ | ~new_n10617_ | ~new_n10618_;
  assign po751 = ~new_n10608_ | ~new_n10610_ | ~new_n9187_ | ~new_n10609_;
  assign po750 = ~new_n9186_ | ~new_n10601_ | ~new_n10599_ | ~new_n10600_;
  assign po749 = ~new_n10590_ | ~new_n10592_ | ~new_n9185_ | ~new_n10591_;
  assign po748 = ~new_n9184_ | ~new_n9183_ | ~new_n10582_;
  assign po747 = ~new_n9182_ | ~new_n10574_ | ~new_n10572_ | ~new_n10573_;
  assign po746 = ~new_n9181_ | ~new_n10565_ | ~new_n10563_ | ~new_n10564_;
  assign po745 = ~new_n10554_ | ~new_n10556_ | ~new_n9180_ | ~new_n10555_;
  assign po744 = ~new_n9179_ | ~new_n9178_ | ~new_n10546_;
  assign po743 = ~new_n9177_ | ~new_n10538_ | ~new_n10536_ | ~new_n10537_;
  assign po742 = ~new_n10527_ | ~new_n10529_ | ~new_n9176_ | ~new_n10528_;
  assign po741 = ~new_n9175_ | ~new_n10520_ | ~new_n10518_ | ~new_n10519_;
  assign po740 = ~new_n10509_ | ~new_n10511_ | ~new_n9174_ | ~new_n10510_;
  assign po739 = ~new_n10500_ | ~new_n10502_ | ~new_n9173_ | ~new_n10501_;
  assign po738 = ~new_n10491_ | ~new_n10493_ | ~new_n9172_ | ~new_n10492_;
  assign po737 = ~new_n9171_ | ~new_n10484_ | ~new_n10482_ | ~new_n10483_;
  assign po736 = ~new_n9170_ | ~new_n9169_ | ~new_n10474_;
  assign po735 = ~new_n10464_ | ~new_n10466_ | ~new_n9168_ | ~new_n10465_;
  assign po734 = ~new_n10457_ | ~new_n9167_;
  assign po733 = ~new_n9164_ | ~new_n10450_ | ~new_n10448_ | ~new_n10449_;
  assign po732 = ~new_n10439_ | ~new_n10441_ | ~new_n9163_ | ~new_n10440_;
  assign po731 = ~new_n9162_ | ~new_n10432_ | ~new_n10430_ | ~new_n10431_;
  assign po730 = ~new_n10421_ | ~new_n10423_ | ~new_n9161_ | ~new_n10422_;
  assign po729 = ~new_n9160_ | ~new_n9159_ | ~new_n10413_;
  assign po728 = ~new_n10403_ | ~new_n10405_ | ~new_n9158_ | ~new_n10404_;
  assign po727 = ~new_n10394_ | ~new_n10396_ | ~new_n9157_ | ~new_n10395_;
  assign po726 = ~new_n9156_ | ~new_n10387_ | ~new_n10385_ | ~new_n10386_;
  assign po725 = ~new_n10372_ | ~new_n10374_ | ~new_n9155_ | ~new_n10373_;
  assign po691 = ~new_n10351_ | ~new_n9134_;
  assign po690 = ~new_n10340_ | ~new_n9131_;
  assign po689 = ~new_n10329_ | ~new_n9128_;
  assign po688 = ~new_n9125_ | ~new_n10319_ | ~new_n10318_;
  assign po687 = ~new_n9122_ | ~new_n10308_ | ~new_n10307_;
  assign po686 = ~new_n9119_ | ~new_n10294_ | ~new_n9121_ | ~new_n10296_;
  assign po685 = ~new_n10283_ | ~new_n10285_ | ~new_n9116_;
  assign po684 = ~new_n10274_ | ~new_n9113_;
  assign po683 = ~new_n10263_ | ~new_n9110_;
  assign po682 = ~new_n10252_ | ~new_n9107_;
  assign po681 = ~new_n10241_ | ~new_n9104_;
  assign po680 = ~new_n10230_ | ~new_n9101_;
  assign po679 = ~new_n10219_ | ~new_n9098_;
  assign po678 = ~new_n10208_ | ~new_n9095_;
  assign po677 = ~new_n10197_ | ~new_n9092_;
  assign po676 = ~new_n10186_ | ~new_n9089_;
  assign po675 = ~new_n10175_ | ~new_n9086_;
  assign po674 = ~new_n10164_ | ~new_n9083_;
  assign po673 = ~new_n10153_ | ~new_n9080_;
  assign po672 = ~new_n10142_ | ~new_n9077_;
  assign po671 = ~new_n10130_ | ~new_n10131_ | ~new_n8427_;
  assign po670 = ~new_n10128_ | ~new_n10129_ | ~new_n8427_;
  assign po669 = ~new_n10125_ | ~new_n9244_ | ~new_n10123_ | ~new_n10124_;
  assign po668 = ~new_n10121_ | ~new_n9243_ | ~new_n10120_ | ~new_n10122_ | ~new_n10119_;
  assign po667 = ~new_n10117_ | ~new_n9242_ | ~new_n10116_ | ~new_n10118_ | ~new_n10115_;
  assign po666 = ~new_n10113_ | ~new_n9241_ | ~new_n10112_ | ~new_n10114_ | ~new_n10111_;
  assign po665 = ~new_n10109_ | ~new_n9240_ | ~new_n10108_ | ~new_n10110_ | ~new_n10107_;
  assign po664 = ~new_n10105_ | ~new_n9239_ | ~new_n10104_ | ~new_n10106_ | ~new_n10103_;
  assign po663 = ~new_n10101_ | ~new_n9238_ | ~new_n10100_ | ~new_n10102_ | ~new_n10099_;
  assign po662 = ~new_n10097_ | ~new_n9237_ | ~new_n10096_ | ~new_n10098_ | ~new_n10095_;
  assign po661 = ~new_n10093_ | ~new_n9236_ | ~new_n10092_ | ~new_n10094_ | ~new_n10091_;
  assign po660 = ~new_n10089_ | ~new_n9235_ | ~new_n10088_ | ~new_n10090_ | ~new_n10087_;
  assign po659 = ~new_n10085_ | ~new_n9234_ | ~new_n10084_ | ~new_n10086_ | ~new_n10083_;
  assign po658 = ~new_n10081_ | ~new_n9233_ | ~new_n10080_ | ~new_n10082_ | ~new_n10079_;
  assign po657 = ~new_n10077_ | ~new_n9232_ | ~new_n10076_ | ~new_n10078_ | ~new_n10075_;
  assign po656 = ~new_n10073_ | ~new_n9231_ | ~new_n10072_ | ~new_n10074_ | ~new_n10071_;
  assign po655 = ~new_n10069_ | ~new_n9230_ | ~new_n10068_ | ~new_n10070_ | ~new_n10067_;
  assign po654 = ~new_n10065_ | ~new_n9229_ | ~new_n10064_ | ~new_n10066_ | ~new_n10063_;
  assign po653 = ~new_n10062_ | ~new_n9228_ | ~new_n10059_ | ~new_n10061_ | ~new_n10060_;
  assign po652 = ~new_n10058_ | ~new_n9227_ | ~new_n10055_ | ~new_n10056_ | ~new_n10057_;
  assign po651 = ~new_n10054_ | ~new_n9226_ | ~new_n10051_ | ~new_n10053_ | ~new_n10052_;
  assign po650 = ~new_n10050_ | ~new_n9225_ | ~new_n10047_ | ~new_n10048_ | ~new_n10049_;
  assign po649 = ~new_n10044_ | ~new_n10046_ | ~new_n9224_ | ~new_n10045_ | ~new_n10043_;
  assign po648 = ~new_n10040_ | ~new_n10042_ | ~new_n9223_ | ~new_n10041_ | ~new_n10039_;
  assign po647 = ~new_n10036_ | ~new_n10038_ | ~new_n9222_ | ~new_n10037_ | ~new_n10035_;
  assign po646 = ~new_n10032_ | ~new_n10034_ | ~new_n9221_ | ~new_n10033_ | ~new_n10031_;
  assign po645 = ~new_n10028_ | ~new_n10030_ | ~new_n9220_ | ~new_n10029_ | ~new_n10027_;
  assign po644 = ~new_n10024_ | ~new_n10026_ | ~new_n9219_ | ~new_n10025_ | ~new_n10023_;
  assign po643 = ~new_n10020_ | ~new_n10022_ | ~new_n9218_ | ~new_n10021_ | ~new_n10019_;
  assign po642 = ~new_n10016_ | ~new_n10018_ | ~new_n9217_ | ~new_n10017_ | ~new_n10015_;
  assign po641 = ~new_n10012_ | ~new_n10014_ | ~new_n9216_ | ~new_n10013_ | ~new_n10011_;
  assign po640 = ~new_n10008_ | ~new_n10010_ | ~new_n9215_ | ~new_n10009_ | ~new_n10007_;
  assign po575 = pi586 & new_n9210_;
  assign po574 = pi585 & new_n9210_;
  assign po573 = pi584 & new_n9210_;
  assign po572 = pi583 & new_n9210_;
  assign po571 = pi582 & new_n9210_;
  assign po570 = pi581 & new_n9210_;
  assign po569 = pi580 & new_n9210_;
  assign po568 = pi579 & new_n9210_;
  assign po567 = pi578 & new_n9210_;
  assign po566 = pi577 & new_n9210_;
  assign po565 = pi576 & new_n9210_;
  assign po564 = pi575 & new_n9210_;
  assign po563 = pi574 & new_n9210_;
  assign po562 = pi573 & new_n9210_;
  assign po561 = pi572 & new_n9210_;
  assign po560 = pi571 & new_n9210_;
  assign po559 = pi570 & new_n9210_;
  assign po558 = pi569 & new_n9210_;
  assign po557 = pi568 & new_n9210_;
  assign po556 = pi567 & new_n9210_;
  assign po555 = pi566 & new_n9210_;
  assign po554 = pi565 & new_n9210_;
  assign po553 = pi564 & new_n9210_;
  assign po552 = pi563 & new_n9210_;
  assign po551 = pi562 & new_n9210_;
  assign po550 = pi561 & new_n9210_;
  assign po549 = pi560 & new_n9210_;
  assign po548 = pi559 & new_n9210_;
  assign po547 = pi558 & new_n9210_;
  assign po546 = pi557 & new_n9210_;
  assign po543 = ~new_n9393_ | ~new_n9394_ | ~new_n9395_;
  assign po542 = ~new_n9390_ | ~new_n9391_ | ~new_n9392_;
  assign po541 = ~new_n9387_ | ~new_n9388_ | ~new_n9389_;
  assign po540 = ~new_n9384_ | ~new_n9385_ | ~new_n9386_;
  assign po539 = ~new_n9381_ | ~new_n9382_ | ~new_n9383_;
  assign po538 = ~new_n9378_ | ~new_n9379_ | ~new_n9380_;
  assign po537 = ~new_n9375_ | ~new_n9376_ | ~new_n9377_;
  assign po536 = ~new_n9372_ | ~new_n9373_ | ~new_n9374_;
  assign po535 = ~new_n9369_ | ~new_n9370_ | ~new_n9371_;
  assign po534 = ~new_n9366_ | ~new_n9367_ | ~new_n9368_;
  assign po533 = ~new_n9363_ | ~new_n9364_ | ~new_n9365_;
  assign po532 = ~new_n9360_ | ~new_n9361_ | ~new_n9362_;
  assign po531 = ~new_n9357_ | ~new_n9358_ | ~new_n9359_;
  assign po530 = ~new_n9354_ | ~new_n9355_ | ~new_n9356_;
  assign po529 = ~new_n9351_ | ~new_n9352_ | ~new_n9353_;
  assign po528 = ~new_n9348_ | ~new_n9349_ | ~new_n9350_;
  assign po527 = ~new_n9345_ | ~new_n9346_ | ~new_n9347_;
  assign po526 = ~new_n9342_ | ~new_n9343_ | ~new_n9344_;
  assign po525 = ~new_n9339_ | ~new_n9340_ | ~new_n9341_;
  assign po524 = ~new_n9336_ | ~new_n9337_ | ~new_n9338_;
  assign po523 = ~new_n9333_ | ~new_n9334_ | ~new_n9335_;
  assign po522 = ~new_n9330_ | ~new_n9331_ | ~new_n9332_;
  assign po521 = ~new_n9327_ | ~new_n9328_ | ~new_n9329_;
  assign po520 = ~new_n9324_ | ~new_n9325_ | ~new_n9326_;
  assign po519 = ~new_n9321_ | ~new_n9322_ | ~new_n9323_;
  assign po518 = ~new_n9318_ | ~new_n9319_ | ~new_n9320_;
  assign po517 = ~new_n9315_ | ~new_n9316_ | ~new_n9317_;
  assign po516 = ~new_n9312_ | ~new_n9313_ | ~new_n9314_;
  assign po515 = ~new_n9309_ | ~new_n9310_ | ~new_n9311_;
  assign po514 = ~new_n9306_ | ~new_n9307_ | ~new_n9308_;
  assign po513 = ~new_n9303_ | ~new_n9304_ | ~new_n9305_;
  assign po512 = ~new_n9300_ | ~new_n9301_ | ~new_n9302_;
  assign po724 = new_n9153_ & new_n10799_;
  assign new_n8675_ = ~pi765 | ~new_n9209_;
  assign new_n8676_ = ~pi735;
  assign new_n8677_ = ~new_n8752_ | ~new_n10809_;
  assign new_n8678_ = ~new_n8752_ | ~new_n9396_;
  assign new_n8679_ = ~new_n8391_ | ~new_n10825_;
  assign new_n8680_ = ~new_n8392_ | ~new_n10834_;
  assign new_n8681_ = ~new_n8966_ | ~new_n8396_;
  assign new_n8682_ = ~new_n8967_ | ~new_n8396_;
  assign new_n8683_ = ~new_n8392_ | ~new_n10825_;
  assign new_n8684_ = ~new_n8392_ | ~new_n8756_;
  assign new_n8685_ = ~new_n8391_ | ~new_n8756_;
  assign new_n8686_ = ~new_n8756_ | ~new_n8763_ | ~new_n8757_;
  assign new_n8687_ = ~new_n8756_ | ~new_n10828_ | ~new_n8763_;
  assign new_n8688_ = ~new_n10834_ | ~new_n8391_;
  assign new_n8689_ = ~new_n9256_ | ~new_n10825_;
  assign new_n8690_ = ~new_n8394_ | ~new_n8763_;
  assign new_n8691_ = ~new_n8763_ | ~new_n8758_;
  assign new_n8692_ = ~new_n9448_ | ~new_n8953_ | ~new_n8954_ | ~new_n9449_ | ~new_n9447_;
  assign new_n8693_ = ~new_n9468_ | ~new_n8970_ | ~new_n8968_ | ~new_n9469_;
  assign new_n8694_ = ~new_n9486_ | ~new_n8974_ | ~new_n8972_ | ~new_n9487_;
  assign new_n8695_ = ~new_n9504_ | ~new_n8978_ | ~new_n8976_ | ~new_n9505_;
  assign new_n8696_ = ~new_n9523_ | ~new_n8981_ | ~new_n9525_ | ~new_n9524_ | ~new_n9522_;
  assign new_n8697_ = ~new_n9541_ | ~new_n8984_ | ~new_n9543_ | ~new_n9542_ | ~new_n9540_;
  assign new_n8698_ = ~new_n9559_ | ~new_n8987_ | ~new_n9561_ | ~new_n9560_ | ~new_n9558_;
  assign new_n8699_ = ~new_n9577_ | ~new_n8990_ | ~new_n9579_ | ~new_n9578_ | ~new_n9576_;
  assign new_n8700_ = ~new_n9595_ | ~new_n8993_ | ~new_n9597_ | ~new_n9596_ | ~new_n9594_;
  assign new_n8701_ = ~new_n9612_ | ~new_n8997_ | ~new_n8995_ | ~new_n9613_;
  assign new_n8702_ = ~new_n9630_ | ~new_n9001_ | ~new_n8999_ | ~new_n9631_;
  assign new_n8703_ = ~new_n9649_ | ~new_n9004_ | ~new_n9651_ | ~new_n9650_ | ~new_n9648_;
  assign new_n8704_ = ~new_n9666_ | ~new_n9008_ | ~new_n9006_ | ~new_n9667_;
  assign new_n8705_ = ~new_n9684_ | ~new_n9012_ | ~new_n9010_ | ~new_n9685_;
  assign new_n8706_ = ~new_n9703_ | ~new_n9015_ | ~new_n9705_ | ~new_n9704_ | ~new_n9702_;
  assign new_n8707_ = ~new_n9721_ | ~new_n9018_ | ~new_n9723_ | ~new_n9722_ | ~new_n9720_;
  assign new_n8708_ = ~new_n9739_ | ~new_n9021_ | ~new_n9741_ | ~new_n9740_ | ~new_n9738_;
  assign new_n8709_ = ~new_n9756_ | ~new_n9025_ | ~new_n9023_ | ~new_n9757_;
  assign new_n8710_ = ~new_n9775_ | ~new_n9028_ | ~new_n9777_ | ~new_n9776_ | ~new_n9774_;
  assign new_n8711_ = ~new_n9793_ | ~new_n9031_ | ~new_n9795_ | ~new_n9794_ | ~new_n9792_;
  assign new_n8712_ = ~new_n1550_ | ~new_n9211_;
  assign new_n8713_ = ~new_n9811_ | ~new_n9034_ | ~new_n9813_ | ~new_n9812_ | ~new_n9810_;
  assign new_n8714_ = ~new_n1549_ | ~new_n9211_;
  assign new_n8715_ = ~new_n9829_ | ~new_n9037_ | ~new_n9831_ | ~new_n9830_ | ~new_n9828_;
  assign new_n8716_ = ~new_n1548_ | ~new_n9211_;
  assign new_n8717_ = ~new_n9847_ | ~new_n9040_ | ~new_n9849_ | ~new_n9848_ | ~new_n9846_;
  assign new_n8718_ = ~new_n1547_ | ~new_n9211_;
  assign new_n8719_ = ~new_n9865_ | ~new_n9043_ | ~new_n9867_ | ~new_n9866_ | ~new_n9864_;
  assign new_n8720_ = ~new_n1546_ | ~new_n9211_;
  assign new_n8721_ = ~new_n9882_ | ~new_n9047_ | ~new_n9045_ | ~new_n9883_;
  assign new_n8722_ = ~new_n1545_ | ~new_n9211_;
  assign new_n8723_ = ~new_n9900_ | ~new_n9051_ | ~new_n9049_ | ~new_n9901_;
  assign new_n8724_ = ~new_n1544_ | ~new_n9211_;
  assign new_n8725_ = ~new_n9918_ | ~new_n9055_ | ~new_n9053_ | ~new_n9919_;
  assign new_n8726_ = ~new_n1543_ | ~new_n9211_;
  assign new_n8727_ = ~new_n9936_ | ~new_n9059_ | ~new_n9057_ | ~new_n9937_;
  assign new_n8728_ = ~new_n1542_ | ~new_n9211_;
  assign new_n8729_ = ~new_n9954_ | ~new_n9063_ | ~new_n9061_ | ~new_n9955_;
  assign new_n8730_ = ~new_n8761_ | ~new_n8762_;
  assign new_n8731_ = ~new_n1541_ | ~new_n9211_;
  assign new_n8732_ = ~new_n9975_ | ~new_n9067_ | ~new_n9065_ | ~new_n9976_ | ~new_n9974_;
  assign new_n8733_ = ~new_n1539_ | ~new_n9211_;
  assign new_n8734_ = ~new_n1538_ | ~new_n9211_;
  assign new_n8735_ = ~new_n8393_ | ~new_n10834_;
  assign new_n8736_ = ~new_n8401_ | ~new_n10005_;
  assign new_n8737_ = ~new_n10825_ | ~new_n8763_;
  assign new_n8738_ = ~new_n9257_ | ~new_n10825_;
  assign new_n8739_ = ~new_n8433_ | ~new_n9289_ | ~new_n9973_;
  assign new_n8740_ = ~new_n8750_ | ~new_n8751_ | ~new_n8752_;
  assign new_n8741_ = ~new_n9072_ | ~new_n9288_;
  assign new_n8742_ = ~new_n8691_ | ~new_n9211_;
  assign new_n8743_ = ~new_n9255_ | ~new_n10801_;
  assign new_n8744_ = ~new_n9073_ | ~new_n8428_;
  assign new_n8745_ = ~new_n9260_ | ~new_n8763_;
  assign new_n8746_ = ~new_n9137_ | ~new_n9268_;
  assign new_n8747_ = ~new_n9254_ | ~new_n8756_;
  assign new_n8748_ = ~new_n9154_ | ~new_n10370_ | ~new_n10369_;
  assign new_n8749_ = ~new_n10795_ | ~new_n9295_;
  assign new_n8750_ = ~new_n10805_ | ~new_n10804_;
  assign new_n8751_ = ~new_n10808_ | ~new_n10807_;
  assign new_n8752_ = ~new_n10811_ | ~new_n10810_;
  assign new_n8753_ = ~new_n10817_ | ~new_n10816_;
  assign po544 = ~new_n10820_ | ~new_n10819_;
  assign po545 = ~new_n10822_ | ~new_n10821_;
  assign new_n8756_ = ~new_n10824_ | ~new_n10823_;
  assign new_n8757_ = ~new_n10827_ | ~new_n10826_;
  assign new_n8758_ = ~new_n10830_ | ~new_n10829_;
  assign new_n8759_ = ~new_n10836_ | ~new_n10835_;
  assign new_n8760_ = ~new_n10839_ | ~new_n10838_;
  assign new_n8761_ = ~new_n10842_ | ~new_n10841_;
  assign new_n8762_ = ~new_n10845_ | ~new_n10844_;
  assign new_n8763_ = ~new_n10833_ | ~new_n10832_;
  assign new_n8764_ = ~new_n10848_ | ~new_n10847_;
  assign new_n8765_ = ~new_n10850_ | ~new_n10849_;
  assign new_n8766_ = ~new_n10853_ | ~new_n10852_;
  assign new_n8767_ = ~new_n10856_ | ~new_n10855_;
  assign po576 = ~new_n10862_ | ~new_n10861_;
  assign new_n8769_ = ~new_n10864_ | ~new_n10863_;
  assign new_n8770_ = ~new_n10866_ | ~new_n10865_;
  assign po577 = ~new_n10869_ | ~new_n10868_;
  assign new_n8772_ = ~new_n10871_ | ~new_n10870_;
  assign new_n8773_ = ~new_n10873_ | ~new_n10872_;
  assign po578 = ~new_n10876_ | ~new_n10875_;
  assign new_n8775_ = ~new_n10878_ | ~new_n10877_;
  assign new_n8776_ = ~new_n10880_ | ~new_n10879_;
  assign po579 = ~new_n10883_ | ~new_n10882_;
  assign new_n8778_ = ~new_n10885_ | ~new_n10884_;
  assign new_n8779_ = ~new_n10887_ | ~new_n10886_;
  assign po580 = ~new_n10890_ | ~new_n10889_;
  assign new_n8781_ = ~new_n10892_ | ~new_n10891_;
  assign new_n8782_ = ~new_n10894_ | ~new_n10893_;
  assign po581 = ~new_n10897_ | ~new_n10896_;
  assign new_n8784_ = ~new_n10899_ | ~new_n10898_;
  assign new_n8785_ = ~new_n10901_ | ~new_n10900_;
  assign po582 = ~new_n10904_ | ~new_n10903_;
  assign new_n8787_ = ~new_n10906_ | ~new_n10905_;
  assign new_n8788_ = ~new_n10908_ | ~new_n10907_;
  assign po583 = ~new_n10911_ | ~new_n10910_;
  assign new_n8790_ = ~new_n10913_ | ~new_n10912_;
  assign new_n8791_ = ~new_n10915_ | ~new_n10914_;
  assign po584 = ~new_n10918_ | ~new_n10917_;
  assign new_n8793_ = ~new_n10920_ | ~new_n10919_;
  assign new_n8794_ = ~new_n10922_ | ~new_n10921_;
  assign po585 = ~new_n10925_ | ~new_n10924_;
  assign new_n8796_ = ~new_n10927_ | ~new_n10926_;
  assign new_n8797_ = ~new_n10929_ | ~new_n10928_;
  assign po586 = ~new_n10932_ | ~new_n10931_;
  assign new_n8799_ = ~new_n10934_ | ~new_n10933_;
  assign new_n8800_ = ~new_n10936_ | ~new_n10935_;
  assign po587 = ~new_n10939_ | ~new_n10938_;
  assign new_n8802_ = ~new_n10941_ | ~new_n10940_;
  assign new_n8803_ = ~new_n10943_ | ~new_n10942_;
  assign po588 = ~new_n10946_ | ~new_n10945_;
  assign new_n8805_ = ~new_n10948_ | ~new_n10947_;
  assign new_n8806_ = ~new_n10950_ | ~new_n10949_;
  assign po589 = ~new_n10953_ | ~new_n10952_;
  assign new_n8808_ = ~new_n10955_ | ~new_n10954_;
  assign new_n8809_ = ~new_n10957_ | ~new_n10956_;
  assign po590 = ~new_n10960_ | ~new_n10959_;
  assign new_n8811_ = ~new_n10962_ | ~new_n10961_;
  assign new_n8812_ = ~new_n10964_ | ~new_n10963_;
  assign po591 = ~new_n10967_ | ~new_n10966_;
  assign new_n8814_ = ~new_n10969_ | ~new_n10968_;
  assign new_n8815_ = ~new_n10971_ | ~new_n10970_;
  assign po592 = ~new_n10974_ | ~new_n10973_;
  assign new_n8817_ = ~new_n10976_ | ~new_n10975_;
  assign new_n8818_ = ~new_n10978_ | ~new_n10977_;
  assign po593 = ~new_n10981_ | ~new_n10980_;
  assign new_n8820_ = ~new_n10983_ | ~new_n10982_;
  assign new_n8821_ = ~new_n10985_ | ~new_n10984_;
  assign po594 = ~new_n10988_ | ~new_n10987_;
  assign new_n8823_ = ~new_n10990_ | ~new_n10989_;
  assign po595 = ~new_n10993_ | ~new_n10992_;
  assign po596 = ~new_n10995_ | ~new_n10994_;
  assign po597 = ~new_n10997_ | ~new_n10996_;
  assign po598 = ~new_n10999_ | ~new_n10998_;
  assign po599 = ~new_n11001_ | ~new_n11000_;
  assign po600 = ~new_n11003_ | ~new_n11002_;
  assign po601 = ~new_n11005_ | ~new_n11004_;
  assign po602 = ~new_n11007_ | ~new_n11006_;
  assign po603 = ~new_n11009_ | ~new_n11008_;
  assign po604 = ~new_n11011_ | ~new_n11010_;
  assign po605 = ~new_n11013_ | ~new_n11012_;
  assign po606 = ~new_n11015_ | ~new_n11014_;
  assign po607 = ~new_n11017_ | ~new_n11016_;
  assign po608 = ~new_n11021_ | ~new_n11020_;
  assign po609 = ~new_n11023_ | ~new_n11022_;
  assign po610 = ~new_n11025_ | ~new_n11024_;
  assign po611 = ~new_n11027_ | ~new_n11026_;
  assign po612 = ~new_n11029_ | ~new_n11028_;
  assign po613 = ~new_n11031_ | ~new_n11030_;
  assign po614 = ~new_n11033_ | ~new_n11032_;
  assign po615 = ~new_n11035_ | ~new_n11034_;
  assign po616 = ~new_n11037_ | ~new_n11036_;
  assign po617 = ~new_n11039_ | ~new_n11038_;
  assign po618 = ~new_n11041_ | ~new_n11040_;
  assign po619 = ~new_n11043_ | ~new_n11042_;
  assign po620 = ~new_n11045_ | ~new_n11044_;
  assign po621 = ~new_n11047_ | ~new_n11046_;
  assign po622 = ~new_n11049_ | ~new_n11048_;
  assign po623 = ~new_n11051_ | ~new_n11050_;
  assign po624 = ~new_n11053_ | ~new_n11052_;
  assign po625 = ~new_n11055_ | ~new_n11054_;
  assign po626 = ~new_n11057_ | ~new_n11056_;
  assign po627 = ~new_n11059_ | ~new_n11058_;
  assign po628 = ~new_n11061_ | ~new_n11060_;
  assign po629 = ~new_n11063_ | ~new_n11062_;
  assign po630 = ~new_n11065_ | ~new_n11064_;
  assign po631 = ~new_n11067_ | ~new_n11066_;
  assign po632 = ~new_n11069_ | ~new_n11068_;
  assign po633 = ~new_n11071_ | ~new_n11070_;
  assign po634 = ~new_n11073_ | ~new_n11072_;
  assign po635 = ~new_n11075_ | ~new_n11074_;
  assign po636 = ~new_n11077_ | ~new_n11076_;
  assign po637 = ~new_n11079_ | ~new_n11078_;
  assign po638 = ~new_n11081_ | ~new_n11080_;
  assign po639 = ~new_n11083_ | ~new_n11082_;
  assign po692 = ~new_n11148_ | ~new_n11147_;
  assign po693 = ~new_n11150_ | ~new_n11149_;
  assign po694 = ~new_n11152_ | ~new_n11151_;
  assign po695 = ~new_n11154_ | ~new_n11153_;
  assign po696 = ~new_n11156_ | ~new_n11155_;
  assign po697 = ~new_n11158_ | ~new_n11157_;
  assign po698 = ~new_n11160_ | ~new_n11159_;
  assign po699 = ~new_n11162_ | ~new_n11161_;
  assign po700 = ~new_n11164_ | ~new_n11163_;
  assign po701 = ~new_n11166_ | ~new_n11165_;
  assign po702 = ~new_n11168_ | ~new_n11167_;
  assign po703 = ~new_n11170_ | ~new_n11169_;
  assign po704 = ~new_n11172_ | ~new_n11171_;
  assign po705 = ~new_n11174_ | ~new_n11173_;
  assign po706 = ~new_n11176_ | ~new_n11175_;
  assign po707 = ~new_n11178_ | ~new_n11177_;
  assign po708 = ~new_n11180_ | ~new_n11179_;
  assign po709 = ~new_n11182_ | ~new_n11181_;
  assign po710 = ~new_n11184_ | ~new_n11183_;
  assign po711 = ~new_n11186_ | ~new_n11185_;
  assign po712 = ~new_n11188_ | ~new_n11187_;
  assign po713 = ~new_n11190_ | ~new_n11189_;
  assign po714 = ~new_n11192_ | ~new_n11191_;
  assign po715 = ~new_n11194_ | ~new_n11193_;
  assign po716 = ~new_n11196_ | ~new_n11195_;
  assign po717 = ~new_n11198_ | ~new_n11197_;
  assign po718 = ~new_n11200_ | ~new_n11199_;
  assign po719 = ~new_n11202_ | ~new_n11201_;
  assign po720 = ~new_n11204_ | ~new_n11203_;
  assign po721 = ~new_n11206_ | ~new_n11205_;
  assign po722 = ~new_n11208_ | ~new_n11207_;
  assign po723 = ~new_n11210_ | ~new_n11209_;
  assign new_n8901_ = ~new_n11324_ | ~new_n11323_;
  assign new_n8902_ = ~new_n11326_ | ~new_n11325_;
  assign new_n8903_ = ~new_n11328_ | ~new_n11327_;
  assign new_n8904_ = ~new_n11330_ | ~new_n11329_;
  assign new_n8905_ = ~new_n11332_ | ~new_n11331_;
  assign new_n8906_ = ~new_n11334_ | ~new_n11333_;
  assign new_n8907_ = ~new_n11336_ | ~new_n11335_;
  assign new_n8908_ = ~new_n11338_ | ~new_n11337_;
  assign new_n8909_ = ~new_n11340_ | ~new_n11339_;
  assign new_n8910_ = ~new_n11342_ | ~new_n11341_;
  assign new_n8911_ = ~new_n11344_ | ~new_n11343_;
  assign new_n8912_ = ~new_n11346_ | ~new_n11345_;
  assign new_n8913_ = ~new_n11348_ | ~new_n11347_;
  assign new_n8914_ = ~new_n11350_ | ~new_n11349_;
  assign new_n8915_ = ~new_n11352_ | ~new_n11351_;
  assign new_n8916_ = ~new_n11354_ | ~new_n11353_;
  assign new_n8917_ = ~new_n11356_ | ~new_n11355_;
  assign new_n8918_ = ~new_n11358_ | ~new_n11357_;
  assign new_n8919_ = ~new_n11360_ | ~new_n11359_;
  assign new_n8920_ = ~new_n11362_ | ~new_n11361_;
  assign new_n8921_ = ~new_n11364_ | ~new_n11363_;
  assign new_n8922_ = ~new_n11366_ | ~new_n11365_;
  assign new_n8923_ = ~new_n11368_ | ~new_n11367_;
  assign new_n8924_ = ~new_n11370_ | ~new_n11369_;
  assign new_n8925_ = ~new_n11372_ | ~new_n11371_;
  assign new_n8926_ = ~new_n11374_ | ~new_n11373_;
  assign new_n8927_ = ~new_n11376_ | ~new_n11375_;
  assign new_n8928_ = ~new_n11378_ | ~new_n11377_;
  assign new_n8929_ = ~new_n11380_ | ~new_n11379_;
  assign new_n8930_ = ~new_n11382_ | ~new_n11381_;
  assign new_n8931_ = ~new_n11384_ | ~new_n11383_;
  assign new_n8932_ = ~new_n11386_ | ~new_n11385_;
  assign new_n8933_ = ~new_n11388_ | ~new_n11387_;
  assign new_n8934_ = ~new_n11390_ | ~new_n11389_;
  assign new_n8935_ = ~new_n11392_ | ~new_n11391_;
  assign new_n8936_ = ~new_n11394_ | ~new_n11393_;
  assign new_n8937_ = ~new_n11396_ | ~new_n11395_;
  assign new_n8938_ = ~new_n11398_ | ~new_n11397_;
  assign new_n8939_ = ~new_n11400_ | ~new_n11399_;
  assign new_n8940_ = ~new_n11402_ | ~new_n11401_;
  assign new_n8941_ = ~new_n11404_ | ~new_n11403_;
  assign new_n8942_ = ~new_n11406_ | ~new_n11405_;
  assign new_n8943_ = ~new_n11408_ | ~new_n11407_;
  assign new_n8944_ = ~new_n11410_ | ~new_n11409_;
  assign new_n8945_ = ~new_n11412_ | ~new_n11411_;
  assign new_n8946_ = ~new_n11414_ | ~new_n11413_;
  assign new_n8947_ = ~new_n11416_ | ~new_n11415_;
  assign new_n8948_ = ~new_n11418_ | ~new_n11417_;
  assign new_n8949_ = ~new_n11420_ | ~new_n11419_;
  assign new_n8950_ = ~new_n11422_ | ~new_n11421_;
  assign new_n8951_ = ~new_n11424_ | ~new_n11423_;
  assign new_n8952_ = ~new_n11426_ | ~new_n11425_;
  assign new_n8953_ = new_n9444_ & new_n9443_;
  assign new_n8954_ = new_n9446_ & new_n9445_;
  assign new_n8955_ = new_n9453_ & new_n9454_ & new_n9452_;
  assign new_n8956_ = new_n9402_ & new_n9400_ & new_n9401_ & new_n9403_;
  assign new_n8957_ = new_n9406_ & new_n9404_ & new_n9405_ & new_n9407_;
  assign new_n8958_ = new_n9410_ & new_n9408_ & new_n9409_ & new_n9411_;
  assign new_n8959_ = new_n9414_ & new_n9413_ & new_n9412_;
  assign new_n8960_ = new_n8958_ & new_n8956_ & new_n8957_ & new_n8959_;
  assign new_n8961_ = new_n9417_ & new_n9415_ & new_n9416_ & new_n9418_;
  assign new_n8962_ = new_n9421_ & new_n9419_ & new_n9420_ & new_n9422_;
  assign new_n8963_ = new_n9425_ & new_n9423_ & new_n9424_ & new_n9426_;
  assign new_n8964_ = new_n9429_ & new_n9428_ & new_n9427_;
  assign new_n8965_ = new_n8963_ & new_n8961_ & new_n8962_ & new_n8964_;
  assign new_n8966_ = new_n8767_ & new_n8766_;
  assign new_n8967_ = new_n10857_ & new_n10854_;
  assign new_n8968_ = new_n9471_ & new_n9470_;
  assign new_n8969_ = new_n9473_ & new_n9472_;
  assign new_n8970_ = new_n8969_ & new_n9475_ & new_n9474_;
  assign new_n8971_ = new_n9477_ & new_n9478_ & new_n9479_;
  assign new_n8972_ = new_n9489_ & new_n9488_;
  assign new_n8973_ = new_n9491_ & new_n9490_;
  assign new_n8974_ = new_n8973_ & new_n9493_ & new_n9492_;
  assign new_n8975_ = new_n9495_ & new_n9496_ & new_n9497_;
  assign new_n8976_ = new_n9507_ & new_n9506_;
  assign new_n8977_ = new_n9509_ & new_n9508_;
  assign new_n8978_ = new_n8977_ & new_n9511_ & new_n9510_;
  assign new_n8979_ = new_n9513_ & new_n9514_ & new_n9515_;
  assign new_n8980_ = new_n9527_ & new_n9526_;
  assign new_n8981_ = new_n8980_ & new_n9529_ & new_n9528_;
  assign new_n8982_ = new_n9531_ & new_n9532_ & new_n9533_;
  assign new_n8983_ = new_n9545_ & new_n9544_;
  assign new_n8984_ = new_n8983_ & new_n9547_ & new_n9546_;
  assign new_n8985_ = new_n9549_ & new_n9550_ & new_n9551_;
  assign new_n8986_ = new_n9563_ & new_n9562_;
  assign new_n8987_ = new_n8986_ & new_n9565_ & new_n9564_;
  assign new_n8988_ = new_n9567_ & new_n9568_ & new_n9569_;
  assign new_n8989_ = new_n9581_ & new_n9580_;
  assign new_n8990_ = new_n8989_ & new_n9583_ & new_n9582_;
  assign new_n8991_ = new_n9585_ & new_n9586_ & new_n9587_;
  assign new_n8992_ = new_n9599_ & new_n9598_;
  assign new_n8993_ = new_n8992_ & new_n9601_ & new_n9600_;
  assign new_n8994_ = new_n9603_ & new_n9604_ & new_n9605_;
  assign new_n8995_ = new_n9615_ & new_n9614_;
  assign new_n8996_ = new_n9617_ & new_n9616_;
  assign new_n8997_ = new_n8996_ & new_n9619_ & new_n9618_;
  assign new_n8998_ = new_n9621_ & new_n9622_ & new_n9623_;
  assign new_n8999_ = new_n9633_ & new_n9632_;
  assign new_n9000_ = new_n9635_ & new_n9634_;
  assign new_n9001_ = new_n9000_ & new_n9637_ & new_n9636_;
  assign new_n9002_ = new_n9639_ & new_n9640_ & new_n9641_;
  assign new_n9003_ = new_n9653_ & new_n9652_;
  assign new_n9004_ = new_n9003_ & new_n9655_ & new_n9654_;
  assign new_n9005_ = new_n9657_ & new_n9658_ & new_n9659_;
  assign new_n9006_ = new_n9669_ & new_n9668_;
  assign new_n9007_ = new_n9671_ & new_n9670_;
  assign new_n9008_ = new_n9007_ & new_n9673_ & new_n9672_;
  assign new_n9009_ = new_n9675_ & new_n9676_ & new_n9677_;
  assign new_n9010_ = new_n9687_ & new_n9686_;
  assign new_n9011_ = new_n9689_ & new_n9688_;
  assign new_n9012_ = new_n9011_ & new_n9691_ & new_n9690_;
  assign new_n9013_ = new_n9693_ & new_n9694_ & new_n9695_;
  assign new_n9014_ = new_n9707_ & new_n9706_;
  assign new_n9015_ = new_n9014_ & new_n9709_ & new_n9708_;
  assign new_n9016_ = new_n9711_ & new_n9712_ & new_n9713_;
  assign new_n9017_ = new_n9725_ & new_n9724_;
  assign new_n9018_ = new_n9017_ & new_n9727_ & new_n9726_;
  assign new_n9019_ = new_n9729_ & new_n9730_ & new_n9731_;
  assign new_n9020_ = new_n9743_ & new_n9742_;
  assign new_n9021_ = new_n9020_ & new_n9745_ & new_n9744_;
  assign new_n9022_ = new_n9747_ & new_n9748_ & new_n9749_;
  assign new_n9023_ = new_n9759_ & new_n9758_;
  assign new_n9024_ = new_n9761_ & new_n9760_;
  assign new_n9025_ = new_n9024_ & new_n9763_ & new_n9762_;
  assign new_n9026_ = new_n9765_ & new_n9766_ & new_n9767_;
  assign new_n9027_ = new_n9779_ & new_n9778_;
  assign new_n9028_ = new_n9027_ & new_n9781_ & new_n9780_;
  assign new_n9029_ = new_n9783_ & new_n9784_ & new_n9785_;
  assign new_n9030_ = new_n9797_ & new_n9796_;
  assign new_n9031_ = new_n9030_ & new_n9799_ & new_n9798_;
  assign new_n9032_ = new_n9801_ & new_n9802_ & new_n9803_;
  assign new_n9033_ = new_n9815_ & new_n9814_;
  assign new_n9034_ = new_n9033_ & new_n9817_ & new_n9816_;
  assign new_n9035_ = new_n9819_ & new_n9820_ & new_n9821_;
  assign new_n9036_ = new_n9833_ & new_n9832_;
  assign new_n9037_ = new_n9036_ & new_n9835_ & new_n9834_;
  assign new_n9038_ = new_n9837_ & new_n9838_ & new_n9839_;
  assign new_n9039_ = new_n9851_ & new_n9850_;
  assign new_n9040_ = new_n9039_ & new_n9853_ & new_n9852_;
  assign new_n9041_ = new_n9855_ & new_n9856_ & new_n9857_;
  assign new_n9042_ = new_n9869_ & new_n9868_;
  assign new_n9043_ = new_n9042_ & new_n9871_ & new_n9870_;
  assign new_n9044_ = new_n9873_ & new_n9874_ & new_n9875_;
  assign new_n9045_ = new_n9885_ & new_n9884_;
  assign new_n9046_ = new_n9887_ & new_n9886_;
  assign new_n9047_ = new_n9046_ & new_n9889_ & new_n9888_;
  assign new_n9048_ = new_n9891_ & new_n9892_ & new_n9893_;
  assign new_n9049_ = new_n9903_ & new_n9902_;
  assign new_n9050_ = new_n9905_ & new_n9904_;
  assign new_n9051_ = new_n9050_ & new_n9907_ & new_n9906_;
  assign new_n9052_ = new_n9909_ & new_n9910_ & new_n9911_;
  assign new_n9053_ = new_n9921_ & new_n9920_;
  assign new_n9054_ = new_n9923_ & new_n9922_;
  assign new_n9055_ = new_n9054_ & new_n9925_ & new_n9924_;
  assign new_n9056_ = new_n9927_ & new_n9928_ & new_n9929_;
  assign new_n9057_ = new_n9939_ & new_n9938_;
  assign new_n9058_ = new_n9941_ & new_n9940_;
  assign new_n9059_ = new_n9058_ & new_n9943_ & new_n9942_;
  assign new_n9060_ = new_n9945_ & new_n9946_ & new_n9947_;
  assign new_n9061_ = new_n9957_ & new_n9956_;
  assign new_n9062_ = new_n9959_ & new_n9958_;
  assign new_n9063_ = new_n9062_ & new_n9961_ & new_n9960_;
  assign new_n9064_ = new_n9963_ & new_n9964_ & new_n9965_;
  assign new_n9065_ = new_n9978_ & new_n9977_;
  assign new_n9066_ = new_n9980_ & new_n9979_;
  assign new_n9067_ = new_n9066_ & new_n9982_ & new_n9981_;
  assign new_n9068_ = new_n9985_ & new_n9984_;
  assign new_n9069_ = new_n10854_ & new_n8767_;
  assign new_n9070_ = new_n10857_ & new_n8766_;
  assign new_n9071_ = new_n9298_ & new_n8757_;
  assign new_n9072_ = new_n10818_ & pi765;
  assign new_n9073_ = new_n10802_ & new_n8742_;
  assign new_n9074_ = new_n8753_ & pi765;
  assign new_n9075_ = new_n8679_ & new_n8685_ & new_n8684_ & new_n8683_ & new_n8686_;
  assign new_n9076_ = new_n8687_ & new_n8738_;
  assign new_n9077_ = new_n10140_ & new_n9079_ & new_n10143_ & new_n10141_;
  assign new_n9078_ = new_n10146_ & new_n10144_;
  assign new_n9079_ = new_n9078_ & new_n10145_;
  assign new_n9080_ = new_n10151_ & new_n9082_ & new_n10154_ & new_n10152_;
  assign new_n9081_ = new_n10157_ & new_n10155_;
  assign new_n9082_ = new_n9081_ & new_n10156_;
  assign new_n9083_ = new_n10162_ & new_n9085_ & new_n10165_ & new_n10163_;
  assign new_n9084_ = new_n10168_ & new_n10166_;
  assign new_n9085_ = new_n9084_ & new_n10167_;
  assign new_n9086_ = new_n10173_ & new_n9088_ & new_n10176_ & new_n10174_;
  assign new_n9087_ = new_n10179_ & new_n10177_;
  assign new_n9088_ = new_n9087_ & new_n10178_;
  assign new_n9089_ = new_n10184_ & new_n9091_ & new_n10187_ & new_n10185_;
  assign new_n9090_ = new_n10190_ & new_n10188_;
  assign new_n9091_ = new_n9090_ & new_n10189_;
  assign new_n9092_ = new_n10195_ & new_n9094_ & new_n10198_ & new_n10196_;
  assign new_n9093_ = new_n10201_ & new_n10199_;
  assign new_n9094_ = new_n9093_ & new_n10200_;
  assign new_n9095_ = new_n10206_ & new_n9097_ & new_n10209_ & new_n10207_;
  assign new_n9096_ = new_n10212_ & new_n10210_;
  assign new_n9097_ = new_n9096_ & new_n10211_;
  assign new_n9098_ = new_n10217_ & new_n9100_ & new_n10220_ & new_n10218_;
  assign new_n9099_ = new_n10223_ & new_n10221_;
  assign new_n9100_ = new_n9099_ & new_n10222_;
  assign new_n9101_ = new_n10228_ & new_n9103_ & new_n10231_ & new_n10229_;
  assign new_n9102_ = new_n10234_ & new_n10232_;
  assign new_n9103_ = new_n9102_ & new_n10233_;
  assign new_n9104_ = new_n10239_ & new_n9106_ & new_n10242_ & new_n10240_;
  assign new_n9105_ = new_n10245_ & new_n10243_;
  assign new_n9106_ = new_n9105_ & new_n10244_;
  assign new_n9107_ = new_n10250_ & new_n9109_ & new_n10253_ & new_n10251_;
  assign new_n9108_ = new_n10256_ & new_n10254_;
  assign new_n9109_ = new_n9108_ & new_n10255_;
  assign new_n9110_ = new_n10264_ & new_n9112_ & new_n10261_ & new_n10262_;
  assign new_n9111_ = new_n10267_ & new_n10265_;
  assign new_n9112_ = new_n9111_ & new_n10266_;
  assign new_n9113_ = new_n10275_ & new_n9115_ & new_n10272_ & new_n10273_;
  assign new_n9114_ = new_n10278_ & new_n10276_;
  assign new_n9115_ = new_n9114_ & new_n10277_;
  assign new_n9116_ = new_n9118_ & new_n10286_ & new_n10284_;
  assign new_n9117_ = new_n10289_ & new_n10287_;
  assign new_n9118_ = new_n9117_ & new_n10288_;
  assign new_n9119_ = new_n10297_ & new_n10295_;
  assign new_n9120_ = new_n10300_ & new_n10298_;
  assign new_n9121_ = new_n9120_ & new_n10299_;
  assign new_n9122_ = new_n10305_ & new_n10306_ & new_n9124_;
  assign new_n9123_ = new_n10311_ & new_n10309_;
  assign new_n9124_ = new_n9123_ & new_n10310_;
  assign new_n9125_ = new_n10316_ & new_n10317_ & new_n9127_;
  assign new_n9126_ = new_n10322_ & new_n10320_;
  assign new_n9127_ = new_n9126_ & new_n10321_;
  assign new_n9128_ = new_n10330_ & new_n9130_ & new_n10327_ & new_n10328_;
  assign new_n9129_ = new_n10333_ & new_n10331_;
  assign new_n9130_ = new_n9129_ & new_n10332_;
  assign new_n9131_ = new_n10338_ & new_n9133_ & new_n10341_ & new_n10339_;
  assign new_n9132_ = new_n10344_ & new_n10342_;
  assign new_n9133_ = new_n9132_ & new_n10343_;
  assign new_n9134_ = new_n10349_ & new_n9136_ & new_n10352_ & new_n10350_;
  assign new_n9135_ = new_n10355_ & new_n10353_;
  assign new_n9136_ = new_n9135_ & new_n10354_;
  assign new_n9137_ = new_n10846_ & new_n8761_;
  assign new_n9138_ = ~new_n11212_ | ~new_n11211_;
  assign new_n9139_ = new_n11293_ & new_n11290_;
  assign new_n9140_ = new_n9141_ & new_n11275_ & new_n9139_ & new_n9142_;
  assign new_n9141_ = new_n11281_ & new_n11278_;
  assign new_n9142_ = new_n11287_ & new_n11284_;
  assign new_n9143_ = new_n11257_ & new_n11263_ & new_n11260_;
  assign new_n9144_ = new_n11266_ & new_n11272_ & new_n11269_;
  assign new_n9145_ = new_n9143_ & new_n11251_ & new_n11254_ & new_n9144_;
  assign new_n9146_ = new_n11242_ & new_n11236_ & new_n11239_ & new_n11245_;
  assign new_n9147_ = new_n11233_ & new_n11230_;
  assign new_n9148_ = new_n11305_ & new_n11299_ & new_n11302_ & new_n11308_;
  assign new_n9149_ = new_n11224_ & new_n11221_ & new_n11218_;
  assign new_n9150_ = new_n9146_ & new_n9149_ & new_n11227_ & new_n11248_ & new_n9147_;
  assign new_n9151_ = new_n9140_ & new_n11311_ & new_n9148_ & new_n11296_ & new_n9145_;
  assign new_n9152_ = new_n10358_ & new_n10359_ & new_n9248_;
  assign new_n9153_ = new_n10794_ & new_n10793_;
  assign new_n9154_ = new_n8740_ & new_n9258_ & new_n10368_ & new_n10818_;
  assign new_n9155_ = new_n10376_ & new_n10375_;
  assign new_n9156_ = new_n10389_ & new_n10388_;
  assign new_n9157_ = new_n10398_ & new_n10397_;
  assign new_n9158_ = new_n10407_ & new_n10406_;
  assign new_n9159_ = new_n10414_ & new_n10412_;
  assign new_n9160_ = new_n10416_ & new_n10415_;
  assign new_n9161_ = new_n10425_ & new_n10424_;
  assign new_n9162_ = new_n10434_ & new_n10433_;
  assign new_n9163_ = new_n10443_ & new_n10442_;
  assign new_n9164_ = new_n10452_ & new_n10451_;
  assign new_n9165_ = new_n8409_ & new_n8455_;
  assign new_n9166_ = new_n10456_ & new_n10455_;
  assign new_n9167_ = new_n9166_ & new_n10459_ & new_n10458_;
  assign new_n9168_ = new_n10468_ & new_n10467_;
  assign new_n9169_ = new_n10475_ & new_n10473_;
  assign new_n9170_ = new_n10477_ & new_n10476_;
  assign new_n9171_ = new_n10486_ & new_n10485_;
  assign new_n9172_ = new_n10495_ & new_n10494_;
  assign new_n9173_ = new_n10504_ & new_n10503_;
  assign new_n9174_ = new_n10513_ & new_n10512_;
  assign new_n9175_ = new_n10522_ & new_n10521_;
  assign new_n9176_ = new_n10531_ & new_n10530_;
  assign new_n9177_ = new_n10540_ & new_n10539_;
  assign new_n9178_ = new_n10547_ & new_n10545_;
  assign new_n9179_ = new_n10549_ & new_n10548_;
  assign new_n9180_ = new_n10558_ & new_n10557_;
  assign new_n9181_ = new_n10567_ & new_n10566_;
  assign new_n9182_ = new_n10576_ & new_n10575_;
  assign new_n9183_ = new_n10583_ & new_n10581_;
  assign new_n9184_ = new_n10585_ & new_n10584_;
  assign new_n9185_ = new_n10594_ & new_n10593_;
  assign new_n9186_ = new_n10603_ & new_n10602_;
  assign new_n9187_ = new_n10612_ & new_n10611_;
  assign new_n9188_ = new_n10621_ & new_n10620_;
  assign new_n9189_ = new_n10630_ & new_n10629_;
  assign new_n9190_ = new_n10632_ & pi765;
  assign new_n9191_ = new_n10818_ & new_n8763_;
  assign new_n9192_ = new_n8763_ & new_n8753_;
  assign new_n9193_ = new_n8680_ & new_n9253_ & new_n8690_;
  assign new_n9194_ = new_n8688_ & new_n8735_ & new_n9255_;
  assign new_n9195_ = new_n8753_ & new_n10636_;
  assign new_n9196_ = new_n8753_ & new_n10638_;
  assign new_n9197_ = new_n8753_ & new_n10640_;
  assign new_n9198_ = new_n8753_ & new_n10642_;
  assign new_n9199_ = new_n8753_ & new_n10644_;
  assign new_n9200_ = new_n8753_ & new_n10646_;
  assign new_n9201_ = new_n8753_ & new_n10652_;
  assign new_n9202_ = new_n8753_ & new_n10674_;
  assign new_n9203_ = new_n8753_ & new_n10688_;
  assign new_n9204_ = new_n8753_ & new_n10690_;
  assign new_n9205_ = new_n8753_ & new_n10692_;
  assign new_n9206_ = new_n8753_ & new_n10694_;
  assign new_n9207_ = new_n8753_ & new_n10696_;
  assign new_n9208_ = new_n8753_ & new_n10698_;
  assign new_n9209_ = ~pi554;
  assign new_n9210_ = ~new_n8401_ | ~new_n8678_;
  assign new_n9211_ = ~new_n10846_ | ~new_n10843_;
  assign new_n9212_ = ~new_n10834_ | ~new_n10825_;
  assign new_n9213_ = ~new_n8401_ | ~new_n9436_;
  assign new_n9214_ = ~new_n8401_ | ~new_n10000_;
  assign new_n9215_ = new_n11085_ & new_n11084_;
  assign new_n9216_ = new_n11087_ & new_n11086_;
  assign new_n9217_ = new_n11089_ & new_n11088_;
  assign new_n9218_ = new_n11091_ & new_n11090_;
  assign new_n9219_ = new_n11093_ & new_n11092_;
  assign new_n9220_ = new_n11095_ & new_n11094_;
  assign new_n9221_ = new_n11097_ & new_n11096_;
  assign new_n9222_ = new_n11099_ & new_n11098_;
  assign new_n9223_ = new_n11101_ & new_n11100_;
  assign new_n9224_ = new_n11103_ & new_n11102_;
  assign new_n9225_ = new_n11105_ & new_n11104_;
  assign new_n9226_ = new_n11107_ & new_n11106_;
  assign new_n9227_ = new_n11109_ & new_n11108_;
  assign new_n9228_ = new_n11111_ & new_n11110_;
  assign new_n9229_ = new_n11113_ & new_n11112_;
  assign new_n9230_ = new_n11115_ & new_n11114_;
  assign new_n9231_ = new_n11117_ & new_n11116_;
  assign new_n9232_ = new_n11119_ & new_n11118_;
  assign new_n9233_ = new_n11121_ & new_n11120_;
  assign new_n9234_ = new_n11123_ & new_n11122_;
  assign new_n9235_ = new_n11125_ & new_n11124_;
  assign new_n9236_ = new_n11127_ & new_n11126_;
  assign new_n9237_ = new_n11129_ & new_n11128_;
  assign new_n9238_ = new_n11131_ & new_n11130_;
  assign new_n9239_ = new_n11133_ & new_n11132_;
  assign new_n9240_ = new_n11135_ & new_n11134_;
  assign new_n9241_ = new_n11137_ & new_n11136_;
  assign new_n9242_ = new_n11139_ & new_n11138_;
  assign new_n9243_ = new_n11141_ & new_n11140_;
  assign new_n9244_ = new_n11143_ & new_n11142_;
  assign new_n9245_ = ~new_n27167_;
  assign new_n9246_ = ~new_n9151_ | ~new_n9150_;
  assign new_n9247_ = ~new_n24882_;
  assign new_n9248_ = new_n11318_ & new_n11317_;
  assign new_n9249_ = ~new_n27860_;
  assign new_n9250_ = ~new_n8734_;
  assign new_n9251_ = ~new_n8733_;
  assign new_n9252_ = ~new_n8690_;
  assign new_n9253_ = ~new_n8393_ | ~new_n8763_;
  assign new_n9254_ = ~new_n8680_;
  assign new_n9255_ = ~new_n8394_ | ~new_n10834_;
  assign new_n9256_ = ~new_n8688_;
  assign new_n9257_ = ~new_n8735_;
  assign new_n9258_ = ~new_n8392_ | ~new_n8763_;
  assign new_n9259_ = ~new_n8686_;
  assign new_n9260_ = ~new_n8679_;
  assign new_n9261_ = ~new_n8683_;
  assign new_n9262_ = ~new_n8685_;
  assign new_n9263_ = ~new_n8684_;
  assign new_n9264_ = ~new_n8738_;
  assign new_n9265_ = ~new_n8689_;
  assign new_n9266_ = ~new_n9256_ | ~new_n8756_;
  assign new_n9267_ = ~new_n8747_;
  assign new_n9268_ = ~new_n8745_;
  assign new_n9269_ = ~new_n8687_;
  assign new_n9270_ = ~new_n8730_;
  assign new_n9271_ = ~new_n9211_;
  assign new_n9272_ = ~new_n8681_;
  assign new_n9273_ = ~new_n8682_;
  assign new_n9274_ = ~new_n10843_ | ~new_n8762_;
  assign po756 = ~new_n8741_;
  assign new_n9276_ = ~new_n8742_;
  assign new_n9277_ = ~new_n8728_;
  assign new_n9278_ = ~new_n8726_;
  assign new_n9279_ = ~new_n8724_;
  assign new_n9280_ = ~new_n8722_;
  assign new_n9281_ = ~new_n8720_;
  assign new_n9282_ = ~new_n8718_;
  assign new_n9283_ = ~new_n8716_;
  assign new_n9284_ = ~new_n8714_;
  assign new_n9285_ = ~new_n8712_;
  assign new_n9286_ = ~new_n8731_;
  assign new_n9287_ = ~new_n8746_;
  assign new_n9288_ = ~new_n8740_;
  assign new_n9289_ = ~new_n8691_;
  assign new_n9290_ = ~new_n8736_;
  assign new_n9291_ = ~new_n9214_;
  assign new_n9292_ = ~new_n9213_;
  assign new_n9293_ = ~new_n9210_;
  assign new_n9294_ = ~new_n8739_;
  assign new_n9295_ = ~new_n8748_ | ~pi765;
  assign new_n9296_ = ~new_n9264_ | ~new_n8401_;
  assign new_n9297_ = ~new_n8677_;
  assign new_n9298_ = ~new_n8737_;
  assign new_n9299_ = ~new_n8675_;
  assign new_n9300_ = ~new_n1562_ | ~po754;
  assign new_n9301_ = ~pi523 | ~new_n8405_;
  assign new_n9302_ = ~pi523 | ~new_n9299_;
  assign new_n9303_ = ~new_n1551_ | ~po754;
  assign new_n9304_ = ~new_n24764_ | ~new_n8405_;
  assign new_n9305_ = ~pi524 | ~new_n9299_;
  assign new_n9306_ = ~new_n1540_ | ~po754;
  assign new_n9307_ = ~new_n24735_ | ~new_n8405_;
  assign new_n9308_ = ~pi525 | ~new_n9299_;
  assign new_n9309_ = ~new_n1537_ | ~po754;
  assign new_n9310_ = ~new_n24736_ | ~new_n8405_;
  assign new_n9311_ = ~pi526 | ~new_n9299_;
  assign new_n9312_ = ~new_n1536_ | ~po754;
  assign new_n9313_ = ~new_n24737_ | ~new_n8405_;
  assign new_n9314_ = ~pi527 | ~new_n9299_;
  assign new_n9315_ = ~new_n1535_ | ~po754;
  assign new_n9316_ = ~new_n24787_ | ~new_n8405_;
  assign new_n9317_ = ~pi528 | ~new_n9299_;
  assign new_n9318_ = ~new_n1534_ | ~po754;
  assign new_n9319_ = ~new_n24738_ | ~new_n8405_;
  assign new_n9320_ = ~pi529 | ~new_n9299_;
  assign new_n9321_ = ~new_n1533_ | ~po754;
  assign new_n9322_ = ~new_n24739_ | ~new_n8405_;
  assign new_n9323_ = ~pi530 | ~new_n9299_;
  assign new_n9324_ = ~new_n1532_ | ~po754;
  assign new_n9325_ = ~new_n24740_ | ~new_n8405_;
  assign new_n9326_ = ~pi531 | ~new_n9299_;
  assign new_n9327_ = ~new_n1531_ | ~po754;
  assign new_n9328_ = ~new_n24785_ | ~new_n8405_;
  assign new_n9329_ = ~pi532 | ~new_n9299_;
  assign new_n9330_ = ~new_n1561_ | ~po754;
  assign new_n9331_ = ~new_n24720_ | ~new_n8405_;
  assign new_n9332_ = ~pi533 | ~new_n9299_;
  assign new_n9333_ = ~new_n1560_ | ~po754;
  assign new_n9334_ = ~new_n24721_ | ~new_n8405_;
  assign new_n9335_ = ~pi534 | ~new_n9299_;
  assign new_n9336_ = ~new_n1559_ | ~po754;
  assign new_n9337_ = ~new_n24722_ | ~new_n8405_;
  assign new_n9338_ = ~pi535 | ~new_n9299_;
  assign new_n9339_ = ~new_n1558_ | ~po754;
  assign new_n9340_ = ~new_n24802_ | ~new_n8405_;
  assign new_n9341_ = ~pi536 | ~new_n9299_;
  assign new_n9342_ = ~new_n1557_ | ~po754;
  assign new_n9343_ = ~new_n24723_ | ~new_n8405_;
  assign new_n9344_ = ~pi537 | ~new_n9299_;
  assign new_n9345_ = ~new_n1556_ | ~po754;
  assign new_n9346_ = ~new_n24724_ | ~new_n8405_;
  assign new_n9347_ = ~pi538 | ~new_n9299_;
  assign new_n9348_ = ~new_n1555_ | ~po754;
  assign new_n9349_ = ~new_n24725_ | ~new_n8405_;
  assign new_n9350_ = ~pi539 | ~new_n9299_;
  assign new_n9351_ = ~new_n1554_ | ~po754;
  assign new_n9352_ = ~new_n24800_ | ~new_n8405_;
  assign new_n9353_ = ~pi540 | ~new_n9299_;
  assign new_n9354_ = ~new_n1553_ | ~po754;
  assign new_n9355_ = ~new_n24726_ | ~new_n8405_;
  assign new_n9356_ = ~pi541 | ~new_n9299_;
  assign new_n9357_ = ~new_n1552_ | ~po754;
  assign new_n9358_ = ~new_n24727_ | ~new_n8405_;
  assign new_n9359_ = ~pi542 | ~new_n9299_;
  assign new_n9360_ = ~new_n1550_ | ~po754;
  assign new_n9361_ = ~new_n24728_ | ~new_n8405_;
  assign new_n9362_ = ~pi543 | ~new_n9299_;
  assign new_n9363_ = ~new_n1549_ | ~po754;
  assign new_n9364_ = ~new_n24796_ | ~new_n8405_;
  assign new_n9365_ = ~pi544 | ~new_n9299_;
  assign new_n9366_ = ~new_n1548_ | ~po754;
  assign new_n9367_ = ~new_n24729_ | ~new_n8405_;
  assign new_n9368_ = ~pi545 | ~new_n9299_;
  assign new_n9369_ = ~new_n1547_ | ~po754;
  assign new_n9370_ = ~new_n24730_ | ~new_n8405_;
  assign new_n9371_ = ~pi546 | ~new_n9299_;
  assign new_n9372_ = ~new_n1546_ | ~po754;
  assign new_n9373_ = ~new_n24731_ | ~new_n8405_;
  assign new_n9374_ = ~pi547 | ~new_n9299_;
  assign new_n9375_ = ~new_n1545_ | ~po754;
  assign new_n9376_ = ~new_n24794_ | ~new_n8405_;
  assign new_n9377_ = ~pi548 | ~new_n9299_;
  assign new_n9378_ = ~new_n1544_ | ~po754;
  assign new_n9379_ = ~new_n24732_ | ~new_n8405_;
  assign new_n9380_ = ~pi549 | ~new_n9299_;
  assign new_n9381_ = ~new_n1543_ | ~po754;
  assign new_n9382_ = ~new_n24792_ | ~new_n8405_;
  assign new_n9383_ = ~pi550 | ~new_n9299_;
  assign new_n9384_ = ~new_n1542_ | ~po754;
  assign new_n9385_ = ~new_n24733_ | ~new_n8405_;
  assign new_n9386_ = ~pi551 | ~new_n9299_;
  assign new_n9387_ = ~new_n1541_ | ~po754;
  assign new_n9388_ = ~new_n24734_ | ~new_n8405_;
  assign new_n9389_ = ~pi552 | ~new_n9299_;
  assign new_n9390_ = ~new_n1539_ | ~po754;
  assign new_n9391_ = ~new_n24790_ | ~new_n8405_;
  assign new_n9392_ = ~pi553 | ~new_n9299_;
  assign new_n9393_ = ~new_n1538_ | ~po754;
  assign new_n9394_ = ~new_n24765_ | ~new_n8405_;
  assign new_n9395_ = ~pi554 | ~new_n9299_;
  assign new_n9396_ = ~new_n9297_ | ~new_n10815_;
  assign new_n9397_ = ~new_n8678_;
  assign new_n9398_ = ~new_n8677_ | ~new_n10806_;
  assign new_n9399_ = ~new_n8677_ | ~new_n10809_;
  assign new_n9400_ = ~new_n9397_ | ~pi565;
  assign new_n9401_ = ~new_n9397_ | ~pi566;
  assign new_n9402_ = ~new_n9397_ | ~pi567;
  assign new_n9403_ = ~new_n9397_ | ~pi568;
  assign new_n9404_ = ~new_n9397_ | ~pi569;
  assign new_n9405_ = ~new_n9397_ | ~pi570;
  assign new_n9406_ = ~new_n9397_ | ~pi571;
  assign new_n9407_ = ~new_n9397_ | ~pi572;
  assign new_n9408_ = ~new_n9397_ | ~pi573;
  assign new_n9409_ = ~new_n9397_ | ~pi574;
  assign new_n9410_ = ~new_n9397_ | ~pi575;
  assign new_n9411_ = ~new_n9397_ | ~pi576;
  assign new_n9412_ = ~new_n9397_ | ~pi577;
  assign new_n9413_ = ~new_n9397_ | ~pi578;
  assign new_n9414_ = ~new_n9397_ | ~pi579;
  assign new_n9415_ = ~new_n9397_ | ~pi580;
  assign new_n9416_ = ~new_n9397_ | ~pi581;
  assign new_n9417_ = ~new_n9397_ | ~pi582;
  assign new_n9418_ = ~new_n9397_ | ~pi583;
  assign new_n9419_ = ~new_n9397_ | ~pi584;
  assign new_n9420_ = ~new_n9397_ | ~pi557;
  assign new_n9421_ = ~new_n9397_ | ~pi585;
  assign new_n9422_ = ~new_n9397_ | ~pi586;
  assign new_n9423_ = ~new_n9397_ | ~pi558;
  assign new_n9424_ = ~new_n9397_ | ~pi559;
  assign new_n9425_ = ~new_n9397_ | ~pi560;
  assign new_n9426_ = ~new_n9397_ | ~pi561;
  assign new_n9427_ = ~new_n9397_ | ~pi562;
  assign new_n9428_ = ~new_n9397_ | ~pi563;
  assign new_n9429_ = ~new_n9397_ | ~pi564;
  assign new_n9430_ = ~new_n9212_;
  assign new_n9431_ = ~new_n10834_ | ~new_n10828_;
  assign new_n9432_ = ~new_n10860_ | ~new_n9431_;
  assign new_n9433_ = ~new_n8747_ | ~new_n8745_;
  assign new_n9434_ = ~new_n9272_ | ~new_n9433_;
  assign new_n9435_ = ~new_n9273_ | ~new_n9432_;
  assign new_n9436_ = ~new_n9435_ | ~new_n9434_;
  assign new_n9437_ = ~new_n8400_ | ~pi588;
  assign new_n9438_ = ~pi620 | ~new_n8399_;
  assign new_n9439_ = ~pi652 | ~new_n8398_;
  assign new_n9440_ = ~pi755 | ~new_n8397_;
  assign new_n9441_ = ~new_n8455_;
  assign new_n9442_ = ~new_n9255_ | ~new_n8735_;
  assign new_n9443_ = ~new_n9261_ | ~new_n27450_;
  assign new_n9444_ = ~new_n9263_ | ~new_n27953_;
  assign new_n9445_ = ~new_n9262_ | ~new_n25193_;
  assign new_n9446_ = ~new_n9259_ | ~new_n28454_;
  assign new_n9447_ = ~new_n9269_ | ~new_n30353_;
  assign new_n9448_ = ~new_n9265_ | ~new_n29511_;
  assign new_n9449_ = ~new_n8395_ | ~new_n26220_;
  assign new_n9450_ = ~new_n8692_;
  assign new_n9451_ = ~new_n8730_ | ~new_n9211_;
  assign new_n9452_ = ~new_n26700_ | ~new_n8404_;
  assign new_n9453_ = ~new_n8403_ | ~new_n8455_;
  assign new_n9454_ = ~new_n8765_ | ~new_n9442_;
  assign new_n9455_ = ~new_n8955_ | ~new_n9450_;
  assign new_n9456_ = ~pi589 | ~new_n8400_;
  assign new_n9457_ = ~pi621 | ~new_n8399_;
  assign new_n9458_ = ~pi653 | ~new_n8398_;
  assign new_n9459_ = ~pi740 | ~new_n8397_;
  assign new_n9460_ = ~new_n8445_;
  assign new_n9461_ = ~pi587 | ~new_n8400_;
  assign new_n9462_ = ~pi619 | ~new_n8399_;
  assign new_n9463_ = ~pi651 | ~new_n8398_;
  assign new_n9464_ = ~pi745 | ~new_n8397_;
  assign new_n9465_ = ~new_n8454_;
  assign new_n9466_ = ~new_n10846_ | ~new_n8761_;
  assign new_n9467_ = ~new_n9274_ | ~new_n9466_;
  assign new_n9468_ = ~new_n8411_ | ~new_n8454_;
  assign new_n9469_ = ~new_n27449_ | ~new_n9261_;
  assign new_n9470_ = ~new_n27952_ | ~new_n9263_;
  assign new_n9471_ = ~new_n25269_ | ~new_n9262_;
  assign new_n9472_ = ~new_n28453_ | ~new_n9259_;
  assign new_n9473_ = ~new_n30352_ | ~new_n9269_;
  assign new_n9474_ = ~new_n29587_ | ~new_n9265_;
  assign new_n9475_ = ~new_n26296_ | ~new_n8395_;
  assign new_n9476_ = ~new_n8693_;
  assign new_n9477_ = ~new_n26776_ | ~new_n8404_;
  assign new_n9478_ = ~new_n8403_ | ~new_n8445_;
  assign new_n9479_ = ~new_n8770_ | ~new_n9442_;
  assign new_n9480_ = ~new_n8971_ | ~new_n9476_;
  assign new_n9481_ = ~pi590 | ~new_n8400_;
  assign new_n9482_ = ~pi622 | ~new_n8399_;
  assign new_n9483_ = ~pi654 | ~new_n8398_;
  assign new_n9484_ = ~new_n25084_ | ~new_n8397_;
  assign new_n9485_ = ~new_n8441_;
  assign new_n9486_ = ~new_n8411_ | ~new_n8455_;
  assign new_n9487_ = ~new_n27371_ | ~new_n9261_;
  assign new_n9488_ = ~new_n27874_ | ~new_n9263_;
  assign new_n9489_ = ~new_n25279_ | ~new_n9262_;
  assign new_n9490_ = ~new_n28375_ | ~new_n9259_;
  assign new_n9491_ = ~new_n30274_ | ~new_n9269_;
  assign new_n9492_ = ~new_n29597_ | ~new_n9265_;
  assign new_n9493_ = ~new_n26306_ | ~new_n8395_;
  assign new_n9494_ = ~new_n8694_;
  assign new_n9495_ = ~new_n26786_ | ~new_n8404_;
  assign new_n9496_ = ~new_n8403_ | ~new_n8441_;
  assign new_n9497_ = ~new_n8773_ | ~new_n9442_;
  assign new_n9498_ = ~new_n8975_ | ~new_n9494_;
  assign new_n9499_ = ~pi591 | ~new_n8400_;
  assign new_n9500_ = ~pi623 | ~new_n8399_;
  assign new_n9501_ = ~pi655 | ~new_n8398_;
  assign new_n9502_ = ~new_n25088_ | ~new_n8397_;
  assign new_n9503_ = ~new_n8437_;
  assign new_n9504_ = ~new_n8411_ | ~new_n8445_;
  assign new_n9505_ = ~new_n27455_ | ~new_n9261_;
  assign new_n9506_ = ~new_n27958_ | ~new_n9263_;
  assign new_n9507_ = ~new_n25190_ | ~new_n9262_;
  assign new_n9508_ = ~new_n28459_ | ~new_n9259_;
  assign new_n9509_ = ~new_n30358_ | ~new_n9269_;
  assign new_n9510_ = ~new_n29508_ | ~new_n9265_;
  assign new_n9511_ = ~new_n26217_ | ~new_n8395_;
  assign new_n9512_ = ~new_n8695_;
  assign new_n9513_ = ~new_n26697_ | ~new_n8404_;
  assign new_n9514_ = ~new_n8403_ | ~new_n8437_;
  assign new_n9515_ = ~new_n8776_ | ~new_n9442_;
  assign new_n9516_ = ~new_n8979_ | ~new_n9512_;
  assign new_n9517_ = ~pi592 | ~new_n8400_;
  assign new_n9518_ = ~pi624 | ~new_n8399_;
  assign new_n9519_ = ~pi656 | ~new_n8398_;
  assign new_n9520_ = ~new_n25112_ | ~new_n8397_;
  assign new_n9521_ = ~new_n8444_;
  assign new_n9522_ = ~new_n8411_ | ~new_n8441_;
  assign new_n9523_ = ~new_n27454_ | ~new_n9261_;
  assign new_n9524_ = ~new_n27957_ | ~new_n9263_;
  assign new_n9525_ = ~new_n25278_ | ~new_n9262_;
  assign new_n9526_ = ~new_n28458_ | ~new_n9259_;
  assign new_n9527_ = ~new_n30357_ | ~new_n9269_;
  assign new_n9528_ = ~new_n29596_ | ~new_n9265_;
  assign new_n9529_ = ~new_n26305_ | ~new_n8395_;
  assign new_n9530_ = ~new_n8696_;
  assign new_n9531_ = ~new_n26785_ | ~new_n8404_;
  assign new_n9532_ = ~new_n8403_ | ~new_n8444_;
  assign new_n9533_ = ~new_n8779_ | ~new_n9442_;
  assign new_n9534_ = ~new_n8982_ | ~new_n9530_;
  assign new_n9535_ = ~pi593 | ~new_n8400_;
  assign new_n9536_ = ~pi625 | ~new_n8399_;
  assign new_n9537_ = ~pi657 | ~new_n8398_;
  assign new_n9538_ = ~new_n25067_ | ~new_n8397_;
  assign new_n9539_ = ~new_n8448_;
  assign new_n9540_ = ~new_n8411_ | ~new_n8437_;
  assign new_n9541_ = ~new_n27372_ | ~new_n9261_;
  assign new_n9542_ = ~new_n27875_ | ~new_n9263_;
  assign new_n9543_ = ~new_n25277_ | ~new_n9262_;
  assign new_n9544_ = ~new_n28376_ | ~new_n9259_;
  assign new_n9545_ = ~new_n30275_ | ~new_n9269_;
  assign new_n9546_ = ~new_n29595_ | ~new_n9265_;
  assign new_n9547_ = ~new_n26304_ | ~new_n8395_;
  assign new_n9548_ = ~new_n8697_;
  assign new_n9549_ = ~new_n26784_ | ~new_n8404_;
  assign new_n9550_ = ~new_n8403_ | ~new_n8448_;
  assign new_n9551_ = ~new_n8782_ | ~new_n9442_;
  assign new_n9552_ = ~new_n8985_ | ~new_n9548_;
  assign new_n9553_ = ~pi594 | ~new_n8400_;
  assign new_n9554_ = ~pi626 | ~new_n8399_;
  assign new_n9555_ = ~pi658 | ~new_n8398_;
  assign new_n9556_ = ~new_n25077_ | ~new_n8397_;
  assign new_n9557_ = ~new_n8447_;
  assign new_n9558_ = ~new_n8411_ | ~new_n8444_;
  assign new_n9559_ = ~new_n27453_ | ~new_n9261_;
  assign new_n9560_ = ~new_n27956_ | ~new_n9263_;
  assign new_n9561_ = ~new_n25191_ | ~new_n9262_;
  assign new_n9562_ = ~new_n28457_ | ~new_n9259_;
  assign new_n9563_ = ~new_n30356_ | ~new_n9269_;
  assign new_n9564_ = ~new_n29509_ | ~new_n9265_;
  assign new_n9565_ = ~new_n26218_ | ~new_n8395_;
  assign new_n9566_ = ~new_n8698_;
  assign new_n9567_ = ~new_n26698_ | ~new_n8404_;
  assign new_n9568_ = ~new_n8403_ | ~new_n8447_;
  assign new_n9569_ = ~new_n8785_ | ~new_n9442_;
  assign new_n9570_ = ~new_n8988_ | ~new_n9566_;
  assign new_n9571_ = ~pi595 | ~new_n8400_;
  assign new_n9572_ = ~pi627 | ~new_n8399_;
  assign new_n9573_ = ~pi659 | ~new_n8398_;
  assign new_n9574_ = ~new_n25071_ | ~new_n8397_;
  assign new_n9575_ = ~new_n8461_;
  assign new_n9576_ = ~new_n8411_ | ~new_n8448_;
  assign new_n9577_ = ~new_n27373_ | ~new_n9261_;
  assign new_n9578_ = ~new_n27876_ | ~new_n9263_;
  assign new_n9579_ = ~new_n25276_ | ~new_n9262_;
  assign new_n9580_ = ~new_n28377_ | ~new_n9259_;
  assign new_n9581_ = ~new_n30276_ | ~new_n9269_;
  assign new_n9582_ = ~new_n29594_ | ~new_n9265_;
  assign new_n9583_ = ~new_n26303_ | ~new_n8395_;
  assign new_n9584_ = ~new_n8699_;
  assign new_n9585_ = ~new_n26783_ | ~new_n8404_;
  assign new_n9586_ = ~new_n8403_ | ~new_n8461_;
  assign new_n9587_ = ~new_n8788_ | ~new_n9442_;
  assign new_n9588_ = ~new_n8991_ | ~new_n9584_;
  assign new_n9589_ = ~pi596 | ~new_n8400_;
  assign new_n9590_ = ~pi628 | ~new_n8399_;
  assign new_n9591_ = ~pi660 | ~new_n8398_;
  assign new_n9592_ = ~new_n25073_ | ~new_n8397_;
  assign new_n9593_ = ~new_n8460_;
  assign new_n9594_ = ~new_n8411_ | ~new_n8447_;
  assign new_n9595_ = ~new_n27452_ | ~new_n9261_;
  assign new_n9596_ = ~new_n27955_ | ~new_n9263_;
  assign new_n9597_ = ~new_n25192_ | ~new_n9262_;
  assign new_n9598_ = ~new_n28456_ | ~new_n9259_;
  assign new_n9599_ = ~new_n30355_ | ~new_n9269_;
  assign new_n9600_ = ~new_n29510_ | ~new_n9265_;
  assign new_n9601_ = ~new_n26219_ | ~new_n8395_;
  assign new_n9602_ = ~new_n8700_;
  assign new_n9603_ = ~new_n26699_ | ~new_n8404_;
  assign new_n9604_ = ~new_n8403_ | ~new_n8460_;
  assign new_n9605_ = ~new_n8791_ | ~new_n9442_;
  assign new_n9606_ = ~new_n8994_ | ~new_n9602_;
  assign new_n9607_ = ~pi597 | ~new_n8400_;
  assign new_n9608_ = ~pi629 | ~new_n8399_;
  assign new_n9609_ = ~pi661 | ~new_n8398_;
  assign new_n9610_ = ~new_n25072_ | ~new_n8397_;
  assign new_n9611_ = ~new_n8439_;
  assign new_n9612_ = ~new_n8411_ | ~new_n8461_;
  assign new_n9613_ = ~new_n27451_ | ~new_n9261_;
  assign new_n9614_ = ~new_n27954_ | ~new_n9263_;
  assign new_n9615_ = ~new_n25275_ | ~new_n9262_;
  assign new_n9616_ = ~new_n28455_ | ~new_n9259_;
  assign new_n9617_ = ~new_n30354_ | ~new_n9269_;
  assign new_n9618_ = ~new_n29593_ | ~new_n9265_;
  assign new_n9619_ = ~new_n26302_ | ~new_n8395_;
  assign new_n9620_ = ~new_n8701_;
  assign new_n9621_ = ~new_n26782_ | ~new_n8404_;
  assign new_n9622_ = ~new_n8403_ | ~new_n8439_;
  assign new_n9623_ = ~new_n8794_ | ~new_n9442_;
  assign new_n9624_ = ~new_n8998_ | ~new_n9620_;
  assign new_n9625_ = ~pi598 | ~new_n8400_;
  assign new_n9626_ = ~pi630 | ~new_n8399_;
  assign new_n9627_ = ~pi662 | ~new_n8398_;
  assign new_n9628_ = ~new_n25068_ | ~new_n8397_;
  assign new_n9629_ = ~new_n8440_;
  assign new_n9630_ = ~new_n8411_ | ~new_n8460_;
  assign new_n9631_ = ~new_n27365_ | ~new_n9261_;
  assign new_n9632_ = ~new_n27868_ | ~new_n9263_;
  assign new_n9633_ = ~new_n25285_ | ~new_n9262_;
  assign new_n9634_ = ~new_n28369_ | ~new_n9259_;
  assign new_n9635_ = ~new_n30268_ | ~new_n9269_;
  assign new_n9636_ = ~new_n29603_ | ~new_n9265_;
  assign new_n9637_ = ~new_n26312_ | ~new_n8395_;
  assign new_n9638_ = ~new_n8702_;
  assign new_n9639_ = ~new_n26792_ | ~new_n8404_;
  assign new_n9640_ = ~new_n8403_ | ~new_n8440_;
  assign new_n9641_ = ~new_n8797_ | ~new_n9442_;
  assign new_n9642_ = ~new_n9002_ | ~new_n9638_;
  assign new_n9643_ = ~pi599 | ~new_n8400_;
  assign new_n9644_ = ~pi631 | ~new_n8399_;
  assign new_n9645_ = ~pi663 | ~new_n8398_;
  assign new_n9646_ = ~new_n25082_ | ~new_n8397_;
  assign new_n9647_ = ~new_n8449_;
  assign new_n9648_ = ~new_n8411_ | ~new_n8439_;
  assign new_n9649_ = ~new_n27469_ | ~new_n9261_;
  assign new_n9650_ = ~new_n27972_ | ~new_n9263_;
  assign new_n9651_ = ~new_n25185_ | ~new_n9262_;
  assign new_n9652_ = ~new_n28473_ | ~new_n9259_;
  assign new_n9653_ = ~new_n30372_ | ~new_n9269_;
  assign new_n9654_ = ~new_n29503_ | ~new_n9265_;
  assign new_n9655_ = ~new_n26212_ | ~new_n8395_;
  assign new_n9656_ = ~new_n8703_;
  assign new_n9657_ = ~new_n26692_ | ~new_n8404_;
  assign new_n9658_ = ~new_n8403_ | ~new_n8449_;
  assign new_n9659_ = ~new_n8800_ | ~new_n9442_;
  assign new_n9660_ = ~new_n9005_ | ~new_n9656_;
  assign new_n9661_ = ~pi600 | ~new_n8400_;
  assign new_n9662_ = ~pi632 | ~new_n8399_;
  assign new_n9663_ = ~pi664 | ~new_n8398_;
  assign new_n9664_ = ~new_n25083_ | ~new_n8397_;
  assign new_n9665_ = ~new_n8457_;
  assign new_n9666_ = ~new_n8411_ | ~new_n8440_;
  assign new_n9667_ = ~new_n27468_ | ~new_n9261_;
  assign new_n9668_ = ~new_n27971_ | ~new_n9263_;
  assign new_n9669_ = ~new_n25274_ | ~new_n9262_;
  assign new_n9670_ = ~new_n28472_ | ~new_n9259_;
  assign new_n9671_ = ~new_n30371_ | ~new_n9269_;
  assign new_n9672_ = ~new_n29592_ | ~new_n9265_;
  assign new_n9673_ = ~new_n26301_ | ~new_n8395_;
  assign new_n9674_ = ~new_n8704_;
  assign new_n9675_ = ~new_n26781_ | ~new_n8404_;
  assign new_n9676_ = ~new_n8403_ | ~new_n8457_;
  assign new_n9677_ = ~new_n8803_ | ~new_n9442_;
  assign new_n9678_ = ~new_n9009_ | ~new_n9674_;
  assign new_n9679_ = ~pi601 | ~new_n8400_;
  assign new_n9680_ = ~pi633 | ~new_n8399_;
  assign new_n9681_ = ~pi665 | ~new_n8398_;
  assign new_n9682_ = ~new_n25089_ | ~new_n8397_;
  assign new_n9683_ = ~new_n8456_;
  assign new_n9684_ = ~new_n8411_ | ~new_n8449_;
  assign new_n9685_ = ~new_n27366_ | ~new_n9261_;
  assign new_n9686_ = ~new_n27869_ | ~new_n9263_;
  assign new_n9687_ = ~new_n25273_ | ~new_n9262_;
  assign new_n9688_ = ~new_n28370_ | ~new_n9259_;
  assign new_n9689_ = ~new_n30269_ | ~new_n9269_;
  assign new_n9690_ = ~new_n29591_ | ~new_n9265_;
  assign new_n9691_ = ~new_n26300_ | ~new_n8395_;
  assign new_n9692_ = ~new_n8705_;
  assign new_n9693_ = ~new_n26780_ | ~new_n8404_;
  assign new_n9694_ = ~new_n8403_ | ~new_n8456_;
  assign new_n9695_ = ~new_n8806_ | ~new_n9442_;
  assign new_n9696_ = ~new_n9013_ | ~new_n9692_;
  assign new_n9697_ = ~pi602 | ~new_n8400_;
  assign new_n9698_ = ~pi634 | ~new_n8399_;
  assign new_n9699_ = ~pi666 | ~new_n8398_;
  assign new_n9700_ = ~new_n25080_ | ~new_n8397_;
  assign new_n9701_ = ~new_n8451_;
  assign new_n9702_ = ~new_n8411_ | ~new_n8457_;
  assign new_n9703_ = ~new_n27467_ | ~new_n9261_;
  assign new_n9704_ = ~new_n27970_ | ~new_n9263_;
  assign new_n9705_ = ~new_n25284_ | ~new_n9262_;
  assign new_n9706_ = ~new_n28471_ | ~new_n9259_;
  assign new_n9707_ = ~new_n30370_ | ~new_n9269_;
  assign new_n9708_ = ~new_n29602_ | ~new_n9265_;
  assign new_n9709_ = ~new_n26311_ | ~new_n8395_;
  assign new_n9710_ = ~new_n8706_;
  assign new_n9711_ = ~new_n26791_ | ~new_n8404_;
  assign new_n9712_ = ~new_n8403_ | ~new_n8451_;
  assign new_n9713_ = ~new_n8809_ | ~new_n9442_;
  assign new_n9714_ = ~new_n9016_ | ~new_n9710_;
  assign new_n9715_ = ~pi603 | ~new_n8400_;
  assign new_n9716_ = ~pi635 | ~new_n8399_;
  assign new_n9717_ = ~pi667 | ~new_n8398_;
  assign new_n9718_ = ~new_n25066_ | ~new_n8397_;
  assign new_n9719_ = ~new_n8450_;
  assign new_n9720_ = ~new_n8411_ | ~new_n8456_;
  assign new_n9721_ = ~new_n27466_ | ~new_n9261_;
  assign new_n9722_ = ~new_n27969_ | ~new_n9263_;
  assign new_n9723_ = ~new_n25283_ | ~new_n9262_;
  assign new_n9724_ = ~new_n28470_ | ~new_n9259_;
  assign new_n9725_ = ~new_n30369_ | ~new_n9269_;
  assign new_n9726_ = ~new_n29601_ | ~new_n9265_;
  assign new_n9727_ = ~new_n26310_ | ~new_n8395_;
  assign new_n9728_ = ~new_n8707_;
  assign new_n9729_ = ~new_n26790_ | ~new_n8404_;
  assign new_n9730_ = ~new_n8403_ | ~new_n8450_;
  assign new_n9731_ = ~new_n8812_ | ~new_n9442_;
  assign new_n9732_ = ~new_n9019_ | ~new_n9728_;
  assign new_n9733_ = ~pi604 | ~new_n8400_;
  assign new_n9734_ = ~pi636 | ~new_n8399_;
  assign new_n9735_ = ~pi668 | ~new_n8398_;
  assign new_n9736_ = ~new_n25078_ | ~new_n8397_;
  assign new_n9737_ = ~new_n8446_;
  assign new_n9738_ = ~new_n8411_ | ~new_n8451_;
  assign new_n9739_ = ~new_n27465_ | ~new_n9261_;
  assign new_n9740_ = ~new_n27968_ | ~new_n9263_;
  assign new_n9741_ = ~new_n25186_ | ~new_n9262_;
  assign new_n9742_ = ~new_n28469_ | ~new_n9259_;
  assign new_n9743_ = ~new_n30368_ | ~new_n9269_;
  assign new_n9744_ = ~new_n29504_ | ~new_n9265_;
  assign new_n9745_ = ~new_n26213_ | ~new_n8395_;
  assign new_n9746_ = ~new_n8708_;
  assign new_n9747_ = ~new_n26693_ | ~new_n8404_;
  assign new_n9748_ = ~new_n8403_ | ~new_n8446_;
  assign new_n9749_ = ~new_n8815_ | ~new_n9442_;
  assign new_n9750_ = ~new_n9022_ | ~new_n9746_;
  assign new_n9751_ = ~pi605 | ~new_n8400_;
  assign new_n9752_ = ~pi637 | ~new_n8399_;
  assign new_n9753_ = ~pi669 | ~new_n8398_;
  assign new_n9754_ = ~new_n25070_ | ~new_n8397_;
  assign new_n9755_ = ~new_n8459_;
  assign new_n9756_ = ~new_n8411_ | ~new_n8450_;
  assign new_n9757_ = ~new_n27367_ | ~new_n9261_;
  assign new_n9758_ = ~new_n27870_ | ~new_n9263_;
  assign new_n9759_ = ~new_n25272_ | ~new_n9262_;
  assign new_n9760_ = ~new_n28371_ | ~new_n9259_;
  assign new_n9761_ = ~new_n30270_ | ~new_n9269_;
  assign new_n9762_ = ~new_n29590_ | ~new_n9265_;
  assign new_n9763_ = ~new_n26299_ | ~new_n8395_;
  assign new_n9764_ = ~new_n8709_;
  assign new_n9765_ = ~new_n26779_ | ~new_n8404_;
  assign new_n9766_ = ~new_n8403_ | ~new_n8459_;
  assign new_n9767_ = ~new_n8818_ | ~new_n9442_;
  assign new_n9768_ = ~new_n9026_ | ~new_n9764_;
  assign new_n9769_ = ~pi606 | ~new_n8400_;
  assign new_n9770_ = ~pi638 | ~new_n8399_;
  assign new_n9771_ = ~pi670 | ~new_n8398_;
  assign new_n9772_ = ~new_n25074_ | ~new_n8397_;
  assign new_n9773_ = ~new_n8458_;
  assign new_n9774_ = ~new_n8411_ | ~new_n8446_;
  assign new_n9775_ = ~new_n27464_ | ~new_n9261_;
  assign new_n9776_ = ~new_n27967_ | ~new_n9263_;
  assign new_n9777_ = ~new_n25271_ | ~new_n9262_;
  assign new_n9778_ = ~new_n28468_ | ~new_n9259_;
  assign new_n9779_ = ~new_n30367_ | ~new_n9269_;
  assign new_n9780_ = ~new_n29589_ | ~new_n9265_;
  assign new_n9781_ = ~new_n26298_ | ~new_n8395_;
  assign new_n9782_ = ~new_n8710_;
  assign new_n9783_ = ~new_n26778_ | ~new_n8404_;
  assign new_n9784_ = ~new_n8403_ | ~new_n8458_;
  assign new_n9785_ = ~new_n8821_ | ~new_n9442_;
  assign new_n9786_ = ~new_n9029_ | ~new_n9782_;
  assign new_n9787_ = ~pi671 | ~new_n8398_;
  assign new_n9788_ = ~pi639 | ~new_n8399_;
  assign new_n9789_ = ~pi607 | ~new_n8400_;
  assign new_n9790_ = ~new_n25079_ | ~new_n8397_;
  assign new_n9791_ = ~new_n8453_;
  assign new_n9792_ = ~new_n8411_ | ~new_n8459_;
  assign new_n9793_ = ~new_n27463_ | ~new_n9261_;
  assign new_n9794_ = ~new_n27966_ | ~new_n9263_;
  assign new_n9795_ = ~new_n25270_ | ~new_n9262_;
  assign new_n9796_ = ~new_n28467_ | ~new_n9259_;
  assign new_n9797_ = ~new_n30366_ | ~new_n9269_;
  assign new_n9798_ = ~new_n29588_ | ~new_n9265_;
  assign new_n9799_ = ~new_n26297_ | ~new_n8395_;
  assign new_n9800_ = ~new_n8711_;
  assign new_n9801_ = ~new_n26777_ | ~new_n8404_;
  assign new_n9802_ = ~new_n8403_ | ~new_n8453_;
  assign new_n9803_ = ~new_n8823_ | ~new_n9442_;
  assign new_n9804_ = ~new_n9032_ | ~new_n9800_;
  assign new_n9805_ = ~pi672 | ~new_n8398_;
  assign new_n9806_ = ~pi640 | ~new_n8399_;
  assign new_n9807_ = ~pi608 | ~new_n8400_;
  assign new_n9808_ = ~new_n25086_ | ~new_n8397_;
  assign new_n9809_ = ~new_n8452_;
  assign new_n9810_ = ~new_n8411_ | ~new_n8458_;
  assign new_n9811_ = ~new_n27368_ | ~new_n9261_;
  assign new_n9812_ = ~new_n27871_ | ~new_n9263_;
  assign new_n9813_ = ~new_n25268_ | ~new_n9262_;
  assign new_n9814_ = ~new_n28372_ | ~new_n9259_;
  assign new_n9815_ = ~new_n30271_ | ~new_n9269_;
  assign new_n9816_ = ~new_n29586_ | ~new_n9265_;
  assign new_n9817_ = ~new_n26295_ | ~new_n8395_;
  assign new_n9818_ = ~new_n8713_;
  assign new_n9819_ = ~new_n26775_ | ~new_n8404_;
  assign new_n9820_ = ~new_n8403_ | ~new_n8452_;
  assign new_n9821_ = ~new_n9285_ | ~new_n9442_;
  assign new_n9822_ = ~new_n9035_ | ~new_n9818_;
  assign new_n9823_ = ~pi673 | ~new_n8398_;
  assign new_n9824_ = ~pi641 | ~new_n8399_;
  assign new_n9825_ = ~pi609 | ~new_n8400_;
  assign new_n9826_ = ~new_n25076_ | ~new_n8397_;
  assign new_n9827_ = ~new_n8438_;
  assign new_n9828_ = ~new_n8411_ | ~new_n8453_;
  assign new_n9829_ = ~new_n27369_ | ~new_n9261_;
  assign new_n9830_ = ~new_n27872_ | ~new_n9263_;
  assign new_n9831_ = ~new_n25282_ | ~new_n9262_;
  assign new_n9832_ = ~new_n28373_ | ~new_n9259_;
  assign new_n9833_ = ~new_n30272_ | ~new_n9269_;
  assign new_n9834_ = ~new_n29600_ | ~new_n9265_;
  assign new_n9835_ = ~new_n26309_ | ~new_n8395_;
  assign new_n9836_ = ~new_n8715_;
  assign new_n9837_ = ~new_n26789_ | ~new_n8404_;
  assign new_n9838_ = ~new_n8403_ | ~new_n8438_;
  assign new_n9839_ = ~new_n9284_ | ~new_n9442_;
  assign new_n9840_ = ~new_n9038_ | ~new_n9836_;
  assign new_n9841_ = ~pi674 | ~new_n8398_;
  assign new_n9842_ = ~pi642 | ~new_n8399_;
  assign new_n9843_ = ~pi610 | ~new_n8400_;
  assign new_n9844_ = ~new_n25065_ | ~new_n8397_;
  assign new_n9845_ = ~new_n8443_;
  assign new_n9846_ = ~new_n8411_ | ~new_n8452_;
  assign new_n9847_ = ~new_n27462_ | ~new_n9261_;
  assign new_n9848_ = ~new_n27965_ | ~new_n9263_;
  assign new_n9849_ = ~new_n25281_ | ~new_n9262_;
  assign new_n9850_ = ~new_n28466_ | ~new_n9259_;
  assign new_n9851_ = ~new_n30365_ | ~new_n9269_;
  assign new_n9852_ = ~new_n29599_ | ~new_n9265_;
  assign new_n9853_ = ~new_n26308_ | ~new_n8395_;
  assign new_n9854_ = ~new_n8717_;
  assign new_n9855_ = ~new_n26788_ | ~new_n8404_;
  assign new_n9856_ = ~new_n8403_ | ~new_n8443_;
  assign new_n9857_ = ~new_n9283_ | ~new_n9442_;
  assign new_n9858_ = ~new_n9041_ | ~new_n9854_;
  assign new_n9859_ = ~pi675 | ~new_n8398_;
  assign new_n9860_ = ~pi643 | ~new_n8399_;
  assign new_n9861_ = ~pi611 | ~new_n8400_;
  assign new_n9862_ = ~new_n25069_ | ~new_n8397_;
  assign new_n9863_ = ~new_n8442_;
  assign new_n9864_ = ~new_n8411_ | ~new_n8438_;
  assign new_n9865_ = ~new_n27461_ | ~new_n9261_;
  assign new_n9866_ = ~new_n27964_ | ~new_n9263_;
  assign new_n9867_ = ~new_n25187_ | ~new_n9262_;
  assign new_n9868_ = ~new_n28465_ | ~new_n9259_;
  assign new_n9869_ = ~new_n30364_ | ~new_n9269_;
  assign new_n9870_ = ~new_n29505_ | ~new_n9265_;
  assign new_n9871_ = ~new_n26214_ | ~new_n8395_;
  assign new_n9872_ = ~new_n8719_;
  assign new_n9873_ = ~new_n26694_ | ~new_n8404_;
  assign new_n9874_ = ~new_n8403_ | ~new_n8442_;
  assign new_n9875_ = ~new_n9282_ | ~new_n9442_;
  assign new_n9876_ = ~new_n9044_ | ~new_n9872_;
  assign new_n9877_ = ~pi676 | ~new_n8398_;
  assign new_n9878_ = ~pi644 | ~new_n8399_;
  assign new_n9879_ = ~pi612 | ~new_n8400_;
  assign new_n9880_ = ~new_n25075_ | ~new_n8397_;
  assign new_n9881_ = ~new_n8435_;
  assign new_n9882_ = ~new_n8411_ | ~new_n8443_;
  assign new_n9883_ = ~new_n27460_ | ~new_n9261_;
  assign new_n9884_ = ~new_n27963_ | ~new_n9263_;
  assign new_n9885_ = ~new_n25267_ | ~new_n9262_;
  assign new_n9886_ = ~new_n28464_ | ~new_n9259_;
  assign new_n9887_ = ~new_n30363_ | ~new_n9269_;
  assign new_n9888_ = ~new_n29585_ | ~new_n9265_;
  assign new_n9889_ = ~new_n26294_ | ~new_n8395_;
  assign new_n9890_ = ~new_n8721_;
  assign new_n9891_ = ~new_n26774_ | ~new_n8404_;
  assign new_n9892_ = ~new_n8403_ | ~new_n8435_;
  assign new_n9893_ = ~new_n9281_ | ~new_n9442_;
  assign new_n9894_ = ~new_n9048_ | ~new_n9890_;
  assign new_n9895_ = ~pi677 | ~new_n8398_;
  assign new_n9896_ = ~pi645 | ~new_n8399_;
  assign new_n9897_ = ~pi613 | ~new_n8400_;
  assign new_n9898_ = ~new_n25085_ | ~new_n8397_;
  assign new_n9899_ = ~new_n8434_;
  assign new_n9900_ = ~new_n8411_ | ~new_n8442_;
  assign new_n9901_ = ~new_n27459_ | ~new_n9261_;
  assign new_n9902_ = ~new_n27962_ | ~new_n9263_;
  assign new_n9903_ = ~new_n25266_ | ~new_n9262_;
  assign new_n9904_ = ~new_n28463_ | ~new_n9259_;
  assign new_n9905_ = ~new_n30362_ | ~new_n9269_;
  assign new_n9906_ = ~new_n29584_ | ~new_n9265_;
  assign new_n9907_ = ~new_n26293_ | ~new_n8395_;
  assign new_n9908_ = ~new_n8723_;
  assign new_n9909_ = ~new_n26773_ | ~new_n8404_;
  assign new_n9910_ = ~new_n8403_ | ~new_n8434_;
  assign new_n9911_ = ~new_n9280_ | ~new_n9442_;
  assign new_n9912_ = ~new_n9052_ | ~new_n9908_;
  assign new_n9913_ = ~pi678 | ~new_n8398_;
  assign new_n9914_ = ~pi646 | ~new_n8399_;
  assign new_n9915_ = ~pi614 | ~new_n8400_;
  assign new_n9916_ = ~new_n25081_ | ~new_n8397_;
  assign new_n9917_ = ~new_n8430_;
  assign new_n9918_ = ~new_n8411_ | ~new_n8435_;
  assign new_n9919_ = ~new_n27370_ | ~new_n9261_;
  assign new_n9920_ = ~new_n27873_ | ~new_n9263_;
  assign new_n9921_ = ~new_n25280_ | ~new_n9262_;
  assign new_n9922_ = ~new_n28374_ | ~new_n9259_;
  assign new_n9923_ = ~new_n30273_ | ~new_n9269_;
  assign new_n9924_ = ~new_n29598_ | ~new_n9265_;
  assign new_n9925_ = ~new_n26307_ | ~new_n8395_;
  assign new_n9926_ = ~new_n8725_;
  assign new_n9927_ = ~new_n26787_ | ~new_n8404_;
  assign new_n9928_ = ~new_n8403_ | ~new_n8430_;
  assign new_n9929_ = ~new_n9279_ | ~new_n9442_;
  assign new_n9930_ = ~new_n9056_ | ~new_n9926_;
  assign new_n9931_ = ~pi679 | ~new_n8398_;
  assign new_n9932_ = ~pi647 | ~new_n8399_;
  assign new_n9933_ = ~pi615 | ~new_n8400_;
  assign new_n9934_ = ~new_n25087_ | ~new_n8397_;
  assign new_n9935_ = ~new_n8431_;
  assign new_n9936_ = ~new_n8411_ | ~new_n8434_;
  assign new_n9937_ = ~new_n27458_ | ~new_n9261_;
  assign new_n9938_ = ~new_n27961_ | ~new_n9263_;
  assign new_n9939_ = ~new_n25188_ | ~new_n9262_;
  assign new_n9940_ = ~new_n28462_ | ~new_n9259_;
  assign new_n9941_ = ~new_n30361_ | ~new_n9269_;
  assign new_n9942_ = ~new_n29506_ | ~new_n9265_;
  assign new_n9943_ = ~new_n26215_ | ~new_n8395_;
  assign new_n9944_ = ~new_n8727_;
  assign new_n9945_ = ~new_n26695_ | ~new_n8404_;
  assign new_n9946_ = ~new_n8403_ | ~new_n8431_;
  assign new_n9947_ = ~new_n9278_ | ~new_n9442_;
  assign new_n9948_ = ~new_n9060_ | ~new_n9944_;
  assign new_n9949_ = ~new_n25151_ | ~new_n8397_;
  assign new_n9950_ = ~pi680 | ~new_n8398_;
  assign new_n9951_ = ~pi648 | ~new_n8399_;
  assign new_n9952_ = ~pi616 | ~new_n8400_;
  assign new_n9953_ = ~new_n8432_;
  assign new_n9954_ = ~new_n8411_ | ~new_n8430_;
  assign new_n9955_ = ~new_n27457_ | ~new_n9261_;
  assign new_n9956_ = ~new_n27960_ | ~new_n9263_;
  assign new_n9957_ = ~new_n25265_ | ~new_n9262_;
  assign new_n9958_ = ~new_n28461_ | ~new_n9259_;
  assign new_n9959_ = ~new_n30360_ | ~new_n9269_;
  assign new_n9960_ = ~new_n29583_ | ~new_n9265_;
  assign new_n9961_ = ~new_n26292_ | ~new_n8395_;
  assign new_n9962_ = ~new_n8729_;
  assign new_n9963_ = ~new_n26772_ | ~new_n8404_;
  assign new_n9964_ = ~new_n8403_ | ~new_n8432_;
  assign new_n9965_ = ~new_n9277_ | ~new_n9442_;
  assign new_n9966_ = ~new_n9064_ | ~new_n9962_;
  assign new_n9967_ = ~pi681 | ~new_n8398_;
  assign new_n9968_ = ~pi649 | ~new_n8399_;
  assign new_n9969_ = ~pi617 | ~new_n8400_;
  assign new_n9970_ = ~new_n25151_ | ~new_n8397_;
  assign new_n9971_ = ~new_n8436_;
  assign new_n9972_ = ~new_n9270_ | ~new_n8676_;
  assign new_n9973_ = ~new_n9211_ | ~new_n9972_;
  assign new_n9974_ = ~new_n8436_ | ~new_n9973_ | ~new_n9289_;
  assign new_n9975_ = ~new_n8411_ | ~new_n8431_;
  assign new_n9976_ = ~new_n27456_ | ~new_n9261_;
  assign new_n9977_ = ~new_n27959_ | ~new_n9263_;
  assign new_n9978_ = ~new_n25189_ | ~new_n9262_;
  assign new_n9979_ = ~new_n28460_ | ~new_n9259_;
  assign new_n9980_ = ~new_n30359_ | ~new_n9269_;
  assign new_n9981_ = ~new_n29507_ | ~new_n9265_;
  assign new_n9982_ = ~new_n26216_ | ~new_n8395_;
  assign new_n9983_ = ~new_n8732_;
  assign new_n9984_ = ~new_n26696_ | ~new_n8404_;
  assign new_n9985_ = ~new_n9286_ | ~new_n9442_;
  assign new_n9986_ = ~new_n9068_ | ~new_n9983_;
  assign new_n9987_ = ~new_n25151_ | ~new_n8397_;
  assign new_n9988_ = ~pi682 | ~new_n8398_;
  assign new_n9989_ = ~pi650 | ~new_n8399_;
  assign new_n9990_ = ~pi618 | ~new_n8400_;
  assign new_n9991_ = ~new_n8433_;
  assign new_n9992_ = ~new_n9251_ | ~new_n9442_;
  assign new_n9993_ = ~new_n8739_ | ~new_n9992_;
  assign new_n9994_ = ~new_n9250_ | ~new_n9442_;
  assign new_n9995_ = ~new_n8739_ | ~new_n9994_;
  assign new_n9996_ = ~new_n8680_ | ~new_n11019_ | ~new_n11018_;
  assign new_n9997_ = ~new_n9266_ | ~new_n8745_;
  assign new_n9998_ = ~new_n8426_ | ~new_n9997_;
  assign new_n9999_ = ~new_n8425_ | ~new_n9996_;
  assign new_n10000_ = ~new_n9999_ | ~new_n9998_;
  assign new_n10001_ = ~new_n10834_ | ~new_n8757_;
  assign new_n10002_ = ~new_n9212_ | ~new_n10001_ | ~new_n8758_;
  assign new_n10003_ = ~new_n8426_ | ~new_n10002_;
  assign new_n10004_ = ~new_n8425_ | ~new_n9997_;
  assign new_n10005_ = ~new_n10004_ | ~new_n10003_ | ~new_n8738_;
  assign new_n10006_ = ~new_n8743_;
  assign new_n10007_ = ~new_n8412_ | ~new_n8455_;
  assign new_n10008_ = ~new_n8408_ | ~new_n26700_;
  assign new_n10009_ = ~new_n8407_ | ~new_n8765_;
  assign new_n10010_ = ~new_n8406_ | ~pi745;
  assign new_n10011_ = ~new_n8412_ | ~new_n8445_;
  assign new_n10012_ = ~new_n8408_ | ~new_n26776_;
  assign new_n10013_ = ~new_n8407_ | ~new_n8770_;
  assign new_n10014_ = ~new_n8406_ | ~pi755;
  assign new_n10015_ = ~new_n8412_ | ~new_n8441_;
  assign new_n10016_ = ~new_n8408_ | ~new_n26786_;
  assign new_n10017_ = ~new_n8407_ | ~new_n8773_;
  assign new_n10018_ = ~new_n8406_ | ~pi740;
  assign new_n10019_ = ~new_n8412_ | ~new_n8437_;
  assign new_n10020_ = ~new_n8408_ | ~new_n26697_;
  assign new_n10021_ = ~new_n8407_ | ~new_n8776_;
  assign new_n10022_ = ~new_n8406_ | ~new_n25084_;
  assign new_n10023_ = ~new_n8412_ | ~new_n8444_;
  assign new_n10024_ = ~new_n8408_ | ~new_n26785_;
  assign new_n10025_ = ~new_n8407_ | ~new_n8779_;
  assign new_n10026_ = ~new_n8406_ | ~new_n25088_;
  assign new_n10027_ = ~new_n8412_ | ~new_n8448_;
  assign new_n10028_ = ~new_n8408_ | ~new_n26784_;
  assign new_n10029_ = ~new_n8407_ | ~new_n8782_;
  assign new_n10030_ = ~new_n8406_ | ~new_n25112_;
  assign new_n10031_ = ~new_n8412_ | ~new_n8447_;
  assign new_n10032_ = ~new_n8408_ | ~new_n26698_;
  assign new_n10033_ = ~new_n8407_ | ~new_n8785_;
  assign new_n10034_ = ~new_n8406_ | ~new_n25067_;
  assign new_n10035_ = ~new_n8412_ | ~new_n8461_;
  assign new_n10036_ = ~new_n8408_ | ~new_n26783_;
  assign new_n10037_ = ~new_n8407_ | ~new_n8788_;
  assign new_n10038_ = ~new_n8406_ | ~new_n25077_;
  assign new_n10039_ = ~new_n8412_ | ~new_n8460_;
  assign new_n10040_ = ~new_n8408_ | ~new_n26699_;
  assign new_n10041_ = ~new_n8407_ | ~new_n8791_;
  assign new_n10042_ = ~new_n8406_ | ~new_n25071_;
  assign new_n10043_ = ~new_n8412_ | ~new_n8439_;
  assign new_n10044_ = ~new_n8408_ | ~new_n26782_;
  assign new_n10045_ = ~new_n8407_ | ~new_n8794_;
  assign new_n10046_ = ~new_n8406_ | ~new_n25073_;
  assign new_n10047_ = ~new_n8412_ | ~new_n8440_;
  assign new_n10048_ = ~new_n8408_ | ~new_n26792_;
  assign new_n10049_ = ~new_n8407_ | ~new_n8797_;
  assign new_n10050_ = ~new_n8406_ | ~new_n25072_;
  assign new_n10051_ = ~new_n8412_ | ~new_n8449_;
  assign new_n10052_ = ~new_n8408_ | ~new_n26692_;
  assign new_n10053_ = ~new_n8407_ | ~new_n8800_;
  assign new_n10054_ = ~new_n8406_ | ~new_n25068_;
  assign new_n10055_ = ~new_n8412_ | ~new_n8457_;
  assign new_n10056_ = ~new_n8408_ | ~new_n26781_;
  assign new_n10057_ = ~new_n8407_ | ~new_n8803_;
  assign new_n10058_ = ~new_n8406_ | ~new_n25082_;
  assign new_n10059_ = ~new_n8412_ | ~new_n8456_;
  assign new_n10060_ = ~new_n8408_ | ~new_n26780_;
  assign new_n10061_ = ~new_n8407_ | ~new_n8806_;
  assign new_n10062_ = ~new_n8406_ | ~new_n25083_;
  assign new_n10063_ = ~new_n8412_ | ~new_n8451_;
  assign new_n10064_ = ~new_n8408_ | ~new_n26791_;
  assign new_n10065_ = ~new_n8407_ | ~new_n8809_;
  assign new_n10066_ = ~new_n8406_ | ~new_n25089_;
  assign new_n10067_ = ~new_n8412_ | ~new_n8450_;
  assign new_n10068_ = ~new_n8408_ | ~new_n26790_;
  assign new_n10069_ = ~new_n8407_ | ~new_n8812_;
  assign new_n10070_ = ~new_n8406_ | ~new_n25080_;
  assign new_n10071_ = ~new_n8412_ | ~new_n8446_;
  assign new_n10072_ = ~new_n8408_ | ~new_n26693_;
  assign new_n10073_ = ~new_n8407_ | ~new_n8815_;
  assign new_n10074_ = ~new_n8406_ | ~new_n25066_;
  assign new_n10075_ = ~new_n8412_ | ~new_n8459_;
  assign new_n10076_ = ~new_n8408_ | ~new_n26779_;
  assign new_n10077_ = ~new_n8407_ | ~new_n8818_;
  assign new_n10078_ = ~new_n8406_ | ~new_n25078_;
  assign new_n10079_ = ~new_n8412_ | ~new_n8458_;
  assign new_n10080_ = ~new_n8408_ | ~new_n26778_;
  assign new_n10081_ = ~new_n8407_ | ~new_n8821_;
  assign new_n10082_ = ~new_n8406_ | ~new_n25070_;
  assign new_n10083_ = ~new_n8412_ | ~new_n8453_;
  assign new_n10084_ = ~new_n8408_ | ~new_n26777_;
  assign new_n10085_ = ~new_n8407_ | ~new_n8823_;
  assign new_n10086_ = ~new_n8406_ | ~new_n25074_;
  assign new_n10087_ = ~new_n8412_ | ~new_n8452_;
  assign new_n10088_ = ~new_n8408_ | ~new_n26775_;
  assign new_n10089_ = ~new_n8407_ | ~new_n9285_;
  assign new_n10090_ = ~new_n8406_ | ~new_n25079_;
  assign new_n10091_ = ~new_n8412_ | ~new_n8438_;
  assign new_n10092_ = ~new_n8408_ | ~new_n26789_;
  assign new_n10093_ = ~new_n8407_ | ~new_n9284_;
  assign new_n10094_ = ~new_n8406_ | ~new_n25086_;
  assign new_n10095_ = ~new_n8412_ | ~new_n8443_;
  assign new_n10096_ = ~new_n8408_ | ~new_n26788_;
  assign new_n10097_ = ~new_n8407_ | ~new_n9283_;
  assign new_n10098_ = ~new_n8406_ | ~new_n25076_;
  assign new_n10099_ = ~new_n8412_ | ~new_n8442_;
  assign new_n10100_ = ~new_n8408_ | ~new_n26694_;
  assign new_n10101_ = ~new_n8407_ | ~new_n9282_;
  assign new_n10102_ = ~new_n8406_ | ~new_n25065_;
  assign new_n10103_ = ~new_n8412_ | ~new_n8435_;
  assign new_n10104_ = ~new_n8408_ | ~new_n26774_;
  assign new_n10105_ = ~new_n8407_ | ~new_n9281_;
  assign new_n10106_ = ~new_n8406_ | ~new_n25069_;
  assign new_n10107_ = ~new_n8412_ | ~new_n8434_;
  assign new_n10108_ = ~new_n8408_ | ~new_n26773_;
  assign new_n10109_ = ~new_n8407_ | ~new_n9280_;
  assign new_n10110_ = ~new_n8406_ | ~new_n25075_;
  assign new_n10111_ = ~new_n8412_ | ~new_n8430_;
  assign new_n10112_ = ~new_n8408_ | ~new_n26787_;
  assign new_n10113_ = ~new_n8407_ | ~new_n9279_;
  assign new_n10114_ = ~new_n8406_ | ~new_n25085_;
  assign new_n10115_ = ~new_n8412_ | ~new_n8431_;
  assign new_n10116_ = ~new_n8408_ | ~new_n26695_;
  assign new_n10117_ = ~new_n8407_ | ~new_n9278_;
  assign new_n10118_ = ~new_n8406_ | ~new_n25081_;
  assign new_n10119_ = ~new_n8412_ | ~new_n8432_;
  assign new_n10120_ = ~new_n8408_ | ~new_n26772_;
  assign new_n10121_ = ~new_n8407_ | ~new_n9277_;
  assign new_n10122_ = ~new_n8406_ | ~new_n25087_;
  assign new_n10123_ = ~new_n8408_ | ~new_n26696_;
  assign new_n10124_ = ~new_n8407_ | ~new_n9286_;
  assign new_n10125_ = ~new_n8406_ | ~new_n25151_;
  assign new_n10126_ = ~new_n8406_ | ~new_n25151_;
  assign new_n10127_ = ~new_n9294_ | ~new_n9290_;
  assign new_n10128_ = ~new_n8407_ | ~new_n9251_;
  assign new_n10129_ = ~pi681 | ~new_n8736_;
  assign new_n10130_ = ~new_n8407_ | ~new_n9250_;
  assign new_n10131_ = ~pi682 | ~new_n8736_;
  assign new_n10132_ = ~new_n8737_ | ~new_n9075_ | ~new_n9076_ | ~new_n10006_;
  assign new_n10133_ = ~new_n25655_ | ~new_n8418_;
  assign new_n10134_ = ~new_n8417_ | ~new_n8757_;
  assign new_n10135_ = ~new_n25926_ | ~new_n8415_;
  assign new_n10136_ = ~new_n10135_ | ~new_n10134_ | ~new_n10133_;
  assign new_n10137_ = ~new_n9288_ | ~new_n10818_;
  assign new_n10138_ = ~new_n8744_;
  assign new_n10139_ = ~new_n9211_ | ~new_n9274_;
  assign new_n10140_ = ~new_n30034_ | ~new_n8429_;
  assign new_n10141_ = ~new_n11146_ | ~new_n8757_;
  assign new_n10142_ = ~new_n8420_ | ~new_n10136_;
  assign new_n10143_ = ~new_n8419_ | ~new_n25655_;
  assign new_n10144_ = ~pi758 | ~po754;
  assign new_n10145_ = ~new_n8416_ | ~new_n25926_;
  assign new_n10146_ = ~pi683 | ~new_n10138_;
  assign new_n10147_ = ~new_n25707_ | ~new_n8418_;
  assign new_n10148_ = ~new_n8417_ | ~new_n8820_;
  assign new_n10149_ = ~new_n25978_ | ~new_n8415_;
  assign new_n10150_ = ~new_n10149_ | ~new_n10148_ | ~new_n10147_;
  assign new_n10151_ = ~new_n30035_ | ~new_n8429_;
  assign new_n10152_ = ~new_n11146_ | ~new_n8820_;
  assign new_n10153_ = ~new_n8420_ | ~new_n10150_;
  assign new_n10154_ = ~new_n25707_ | ~new_n8419_;
  assign new_n10155_ = ~pi739 | ~po754;
  assign new_n10156_ = ~new_n25978_ | ~new_n8416_;
  assign new_n10157_ = ~pi684 | ~new_n10138_;
  assign new_n10158_ = ~new_n25708_ | ~new_n8418_;
  assign new_n10159_ = ~new_n8417_ | ~new_n8817_;
  assign new_n10160_ = ~new_n25979_ | ~new_n8415_;
  assign new_n10161_ = ~new_n10160_ | ~new_n10159_ | ~new_n10158_;
  assign new_n10162_ = ~new_n30036_ | ~new_n8429_;
  assign new_n10163_ = ~new_n11146_ | ~new_n8817_;
  assign new_n10164_ = ~new_n8420_ | ~new_n10161_;
  assign new_n10165_ = ~new_n25708_ | ~new_n8419_;
  assign new_n10166_ = ~pi749 | ~po754;
  assign new_n10167_ = ~new_n25979_ | ~new_n8416_;
  assign new_n10168_ = ~pi685 | ~new_n10138_;
  assign new_n10169_ = ~new_n25709_ | ~new_n8418_;
  assign new_n10170_ = ~new_n8417_ | ~new_n8814_;
  assign new_n10171_ = ~new_n25980_ | ~new_n8415_;
  assign new_n10172_ = ~new_n10171_ | ~new_n10170_ | ~new_n10169_;
  assign new_n10173_ = ~new_n29980_ | ~new_n8429_;
  assign new_n10174_ = ~new_n11146_ | ~new_n8814_;
  assign new_n10175_ = ~new_n8420_ | ~new_n10172_;
  assign new_n10176_ = ~new_n25709_ | ~new_n8419_;
  assign new_n10177_ = ~pi751 | ~po754;
  assign new_n10178_ = ~new_n25980_ | ~new_n8416_;
  assign new_n10179_ = ~pi686 | ~new_n10138_;
  assign new_n10180_ = ~new_n25710_ | ~new_n8418_;
  assign new_n10181_ = ~new_n8417_ | ~new_n8811_;
  assign new_n10182_ = ~new_n25981_ | ~new_n8415_;
  assign new_n10183_ = ~new_n10182_ | ~new_n10181_ | ~new_n10180_;
  assign new_n10184_ = ~new_n30044_ | ~new_n8429_;
  assign new_n10185_ = ~new_n11146_ | ~new_n8811_;
  assign new_n10186_ = ~new_n8420_ | ~new_n10183_;
  assign new_n10187_ = ~new_n25710_ | ~new_n8419_;
  assign new_n10188_ = ~pi736 | ~po754;
  assign new_n10189_ = ~new_n25981_ | ~new_n8416_;
  assign new_n10190_ = ~pi687 | ~new_n10138_;
  assign new_n10191_ = ~new_n25711_ | ~new_n8418_;
  assign new_n10192_ = ~new_n8417_ | ~new_n8808_;
  assign new_n10193_ = ~new_n25982_ | ~new_n8415_;
  assign new_n10194_ = ~new_n10193_ | ~new_n10192_ | ~new_n10191_;
  assign new_n10195_ = ~new_n30045_ | ~new_n8429_;
  assign new_n10196_ = ~new_n11146_ | ~new_n8808_;
  assign new_n10197_ = ~new_n8420_ | ~new_n10194_;
  assign new_n10198_ = ~new_n25711_ | ~new_n8419_;
  assign new_n10199_ = ~pi762 | ~po754;
  assign new_n10200_ = ~new_n25982_ | ~new_n8416_;
  assign new_n10201_ = ~pi688 | ~new_n10138_;
  assign new_n10202_ = ~new_n25712_ | ~new_n8418_;
  assign new_n10203_ = ~new_n8417_ | ~new_n8805_;
  assign new_n10204_ = ~new_n25983_ | ~new_n8415_;
  assign new_n10205_ = ~new_n10204_ | ~new_n10203_ | ~new_n10202_;
  assign new_n10206_ = ~new_n30037_ | ~new_n8429_;
  assign new_n10207_ = ~new_n11146_ | ~new_n8805_;
  assign new_n10208_ = ~new_n8420_ | ~new_n10205_;
  assign new_n10209_ = ~new_n25712_ | ~new_n8419_;
  assign new_n10210_ = ~pi743 | ~po754;
  assign new_n10211_ = ~new_n25983_ | ~new_n8416_;
  assign new_n10212_ = ~pi689 | ~new_n10138_;
  assign new_n10213_ = ~new_n25713_ | ~new_n8418_;
  assign new_n10214_ = ~new_n8417_ | ~new_n8802_;
  assign new_n10215_ = ~new_n25984_ | ~new_n8415_;
  assign new_n10216_ = ~new_n10215_ | ~new_n10214_ | ~new_n10213_;
  assign new_n10217_ = ~new_n30038_ | ~new_n8429_;
  assign new_n10218_ = ~new_n11146_ | ~new_n8802_;
  assign new_n10219_ = ~new_n8420_ | ~new_n10216_;
  assign new_n10220_ = ~new_n25713_ | ~new_n8419_;
  assign new_n10221_ = ~pi753 | ~po754;
  assign new_n10222_ = ~new_n25984_ | ~new_n8416_;
  assign new_n10223_ = ~pi690 | ~new_n10138_;
  assign new_n10224_ = ~new_n25714_ | ~new_n8418_;
  assign new_n10225_ = ~new_n8417_ | ~new_n8799_;
  assign new_n10226_ = ~new_n25985_ | ~new_n8415_;
  assign new_n10227_ = ~new_n10226_ | ~new_n10225_ | ~new_n10224_;
  assign new_n10228_ = ~new_n29979_ | ~new_n8429_;
  assign new_n10229_ = ~new_n11146_ | ~new_n8799_;
  assign new_n10230_ = ~new_n8420_ | ~new_n10227_;
  assign new_n10231_ = ~new_n25714_ | ~new_n8419_;
  assign new_n10232_ = ~pi741 | ~po754;
  assign new_n10233_ = ~new_n25985_ | ~new_n8416_;
  assign new_n10234_ = ~pi691 | ~new_n10138_;
  assign new_n10235_ = ~new_n25715_ | ~new_n8418_;
  assign new_n10236_ = ~new_n8417_ | ~new_n8796_;
  assign new_n10237_ = ~new_n25986_ | ~new_n8415_;
  assign new_n10238_ = ~new_n10237_ | ~new_n10236_ | ~new_n10235_;
  assign new_n10239_ = ~new_n30046_ | ~new_n8429_;
  assign new_n10240_ = ~new_n11146_ | ~new_n8796_;
  assign new_n10241_ = ~new_n8420_ | ~new_n10238_;
  assign new_n10242_ = ~new_n25715_ | ~new_n8419_;
  assign new_n10243_ = ~pi760 | ~po754;
  assign new_n10244_ = ~new_n25986_ | ~new_n8416_;
  assign new_n10245_ = ~pi692 | ~new_n10138_;
  assign new_n10246_ = ~new_n25698_ | ~new_n8418_;
  assign new_n10247_ = ~new_n8417_ | ~new_n8793_;
  assign new_n10248_ = ~new_n25969_ | ~new_n8415_;
  assign new_n10249_ = ~new_n10248_ | ~new_n10247_ | ~new_n10246_;
  assign new_n10250_ = ~new_n30039_ | ~new_n8429_;
  assign new_n10251_ = ~new_n11146_ | ~new_n8793_;
  assign new_n10252_ = ~new_n8420_ | ~new_n10249_;
  assign new_n10253_ = ~new_n25698_ | ~new_n8419_;
  assign new_n10254_ = ~pi746 | ~po754;
  assign new_n10255_ = ~new_n25969_ | ~new_n8416_;
  assign new_n10256_ = ~pi693 | ~new_n10138_;
  assign new_n10257_ = ~new_n25699_ | ~new_n8418_;
  assign new_n10258_ = ~new_n8417_ | ~new_n8790_;
  assign new_n10259_ = ~new_n25970_ | ~new_n8415_;
  assign new_n10260_ = ~new_n10259_ | ~new_n10258_ | ~new_n10257_;
  assign new_n10261_ = ~new_n29983_ | ~new_n8429_;
  assign new_n10262_ = ~new_n11146_ | ~new_n8790_;
  assign new_n10263_ = ~new_n8420_ | ~new_n10260_;
  assign new_n10264_ = ~new_n25699_ | ~new_n8419_;
  assign new_n10265_ = ~pi756 | ~po754;
  assign new_n10266_ = ~new_n25970_ | ~new_n8416_;
  assign new_n10267_ = ~pi694 | ~new_n10138_;
  assign new_n10268_ = ~new_n25700_ | ~new_n8418_;
  assign new_n10269_ = ~new_n8417_ | ~new_n8787_;
  assign new_n10270_ = ~new_n25971_ | ~new_n8415_;
  assign new_n10271_ = ~new_n10270_ | ~new_n10269_ | ~new_n10268_;
  assign new_n10272_ = ~new_n30040_ | ~new_n8429_;
  assign new_n10273_ = ~new_n11146_ | ~new_n8787_;
  assign new_n10274_ = ~new_n8420_ | ~new_n10271_;
  assign new_n10275_ = ~new_n25700_ | ~new_n8419_;
  assign new_n10276_ = ~pi764 | ~po754;
  assign new_n10277_ = ~new_n25971_ | ~new_n8416_;
  assign new_n10278_ = ~pi695 | ~new_n10138_;
  assign new_n10279_ = ~new_n25701_ | ~new_n8418_;
  assign new_n10280_ = ~new_n8417_ | ~new_n8784_;
  assign new_n10281_ = ~new_n25972_ | ~new_n8415_;
  assign new_n10282_ = ~new_n10281_ | ~new_n10280_ | ~new_n10279_;
  assign new_n10283_ = ~new_n29982_ | ~new_n8429_;
  assign new_n10284_ = ~new_n11146_ | ~new_n8784_;
  assign new_n10285_ = ~new_n8420_ | ~new_n10282_;
  assign new_n10286_ = ~new_n25701_ | ~new_n8419_;
  assign new_n10287_ = ~pi738 | ~po754;
  assign new_n10288_ = ~new_n25972_ | ~new_n8416_;
  assign new_n10289_ = ~pi696 | ~new_n10138_;
  assign new_n10290_ = ~new_n25702_ | ~new_n8418_;
  assign new_n10291_ = ~new_n8417_ | ~new_n8781_;
  assign new_n10292_ = ~new_n25973_ | ~new_n8415_;
  assign new_n10293_ = ~new_n10292_ | ~new_n10291_ | ~new_n10290_;
  assign new_n10294_ = ~new_n30041_ | ~new_n8429_;
  assign new_n10295_ = ~new_n11146_ | ~new_n8781_;
  assign new_n10296_ = ~new_n8420_ | ~new_n10293_;
  assign new_n10297_ = ~new_n25702_ | ~new_n8419_;
  assign new_n10298_ = ~pi750 | ~po754;
  assign new_n10299_ = ~new_n25973_ | ~new_n8416_;
  assign new_n10300_ = ~pi697 | ~new_n10138_;
  assign new_n10301_ = ~new_n25703_ | ~new_n8418_;
  assign new_n10302_ = ~new_n8417_ | ~new_n8778_;
  assign new_n10303_ = ~new_n25974_ | ~new_n8415_;
  assign new_n10304_ = ~new_n10303_ | ~new_n10302_ | ~new_n10301_;
  assign new_n10305_ = ~new_n30042_ | ~new_n8429_;
  assign new_n10306_ = ~new_n11146_ | ~new_n8778_;
  assign new_n10307_ = ~new_n8420_ | ~new_n10304_;
  assign new_n10308_ = ~new_n25703_ | ~new_n8419_;
  assign new_n10309_ = ~pi747 | ~po754;
  assign new_n10310_ = ~new_n25974_ | ~new_n8416_;
  assign new_n10311_ = ~pi698 | ~new_n10138_;
  assign new_n10312_ = ~new_n25704_ | ~new_n8418_;
  assign new_n10313_ = ~new_n8417_ | ~new_n8775_;
  assign new_n10314_ = ~new_n25975_ | ~new_n8415_;
  assign new_n10315_ = ~new_n10314_ | ~new_n10313_ | ~new_n10312_;
  assign new_n10316_ = ~new_n29981_ | ~new_n8429_;
  assign new_n10317_ = ~new_n11146_ | ~new_n8775_;
  assign new_n10318_ = ~new_n8420_ | ~new_n10315_;
  assign new_n10319_ = ~new_n25704_ | ~new_n8419_;
  assign new_n10320_ = ~pi759 | ~po754;
  assign new_n10321_ = ~new_n25975_ | ~new_n8416_;
  assign new_n10322_ = ~pi699 | ~new_n10138_;
  assign new_n10323_ = ~new_n25705_ | ~new_n8418_;
  assign new_n10324_ = ~new_n8417_ | ~new_n8772_;
  assign new_n10325_ = ~new_n25976_ | ~new_n8415_;
  assign new_n10326_ = ~new_n10325_ | ~new_n10324_ | ~new_n10323_;
  assign new_n10327_ = ~new_n30043_ | ~new_n8429_;
  assign new_n10328_ = ~new_n11146_ | ~new_n8772_;
  assign new_n10329_ = ~new_n8420_ | ~new_n10326_;
  assign new_n10330_ = ~new_n25705_ | ~new_n8419_;
  assign new_n10331_ = ~pi740 | ~po754;
  assign new_n10332_ = ~new_n25976_ | ~new_n8416_;
  assign new_n10333_ = ~pi700 | ~new_n10138_;
  assign new_n10334_ = ~new_n25706_ | ~new_n8418_;
  assign new_n10335_ = ~new_n8417_ | ~new_n8769_;
  assign new_n10336_ = ~new_n25977_ | ~new_n8415_;
  assign new_n10337_ = ~new_n10336_ | ~new_n10335_ | ~new_n10334_;
  assign new_n10338_ = ~new_n30033_ | ~new_n8429_;
  assign new_n10339_ = ~new_n11146_ | ~new_n8769_;
  assign new_n10340_ = ~new_n8420_ | ~new_n10337_;
  assign new_n10341_ = ~new_n25706_ | ~new_n8419_;
  assign new_n10342_ = ~pi755 | ~po754;
  assign new_n10343_ = ~new_n25977_ | ~new_n8416_;
  assign new_n10344_ = ~pi701 | ~new_n10138_;
  assign new_n10345_ = ~new_n25656_ | ~new_n8418_;
  assign new_n10346_ = ~new_n8417_ | ~new_n8764_;
  assign new_n10347_ = ~new_n25927_ | ~new_n8415_;
  assign new_n10348_ = ~new_n10347_ | ~new_n10346_ | ~new_n10345_;
  assign new_n10349_ = ~new_n29984_ | ~new_n8429_;
  assign new_n10350_ = ~new_n11146_ | ~new_n8764_;
  assign new_n10351_ = ~new_n8420_ | ~new_n10348_;
  assign new_n10352_ = ~new_n25656_ | ~new_n8419_;
  assign new_n10353_ = ~pi745 | ~po754;
  assign new_n10354_ = ~new_n25927_ | ~new_n8416_;
  assign new_n10355_ = ~pi702 | ~new_n10138_;
  assign new_n10356_ = ~new_n9246_;
  assign new_n10357_ = ~new_n8428_ | ~new_n11320_ | ~new_n11319_;
  assign new_n10358_ = ~new_n9245_ | ~new_n8401_ | ~new_n9287_;
  assign new_n10359_ = ~pi735 | ~new_n10357_;
  assign new_n10360_ = ~new_n8414_ | ~new_n8456_;
  assign new_n10361_ = ~new_n8410_ | ~new_n8450_;
  assign new_n10362_ = ~new_n25080_ | ~new_n8682_;
  assign new_n10363_ = ~new_n10362_ | ~new_n10361_ | ~new_n10360_;
  assign new_n10364_ = ~new_n8689_ | ~new_n8690_ | ~new_n10803_ | ~new_n9266_ | ~new_n9253_;
  assign new_n10365_ = ~new_n9272_ | ~new_n10364_;
  assign new_n10366_ = ~new_n9267_ | ~new_n9273_;
  assign new_n10367_ = ~new_n10366_ | ~new_n10365_;
  assign new_n10368_ = ~new_n9289_ | ~new_n8756_;
  assign new_n10369_ = ~new_n9267_ | ~new_n8682_;
  assign new_n10370_ = ~new_n10364_ | ~new_n8681_;
  assign new_n10371_ = ~new_n8748_;
  assign new_n10372_ = ~new_n8812_ | ~new_n10798_;
  assign new_n10373_ = ~new_n25080_ | ~new_n8749_;
  assign new_n10374_ = ~new_n28974_ | ~new_n8413_;
  assign new_n10375_ = ~new_n8409_ | ~new_n10363_;
  assign new_n10376_ = ~pi736 | ~po754;
  assign new_n10377_ = ~new_n8414_ | ~new_n8435_;
  assign new_n10378_ = ~new_n8410_ | ~new_n8430_;
  assign new_n10379_ = ~new_n25085_ | ~new_n8682_;
  assign new_n10380_ = ~new_n10379_ | ~new_n10378_ | ~new_n10377_;
  assign new_n10381_ = ~new_n8743_ | ~new_n8681_;
  assign new_n10382_ = ~new_n10371_ | ~new_n10381_;
  assign new_n10383_ = ~new_n9272_ | ~new_n8743_;
  assign new_n10384_ = ~new_n8738_ | ~new_n10383_;
  assign new_n10385_ = ~new_n8423_ | ~new_n9279_;
  assign new_n10386_ = ~new_n8422_ | ~new_n25085_;
  assign new_n10387_ = ~new_n28876_ | ~new_n8413_;
  assign new_n10388_ = ~new_n8409_ | ~new_n10380_;
  assign new_n10389_ = ~pi737 | ~po754;
  assign new_n10390_ = ~new_n8414_ | ~new_n8444_;
  assign new_n10391_ = ~new_n8410_ | ~new_n8447_;
  assign new_n10392_ = ~new_n25067_ | ~new_n8682_;
  assign new_n10393_ = ~new_n10392_ | ~new_n10391_ | ~new_n10390_;
  assign new_n10394_ = ~new_n8785_ | ~new_n10798_;
  assign new_n10395_ = ~new_n25067_ | ~new_n8749_;
  assign new_n10396_ = ~new_n28957_ | ~new_n8413_;
  assign new_n10397_ = ~new_n8409_ | ~new_n10393_;
  assign new_n10398_ = ~pi738 | ~po754;
  assign new_n10399_ = ~new_n8414_ | ~new_n8446_;
  assign new_n10400_ = ~new_n8410_ | ~new_n8458_;
  assign new_n10401_ = ~new_n25070_ | ~new_n8682_;
  assign new_n10402_ = ~new_n10401_ | ~new_n10400_ | ~new_n10399_;
  assign new_n10403_ = ~new_n8821_ | ~new_n10798_;
  assign new_n10404_ = ~new_n25070_ | ~new_n8749_;
  assign new_n10405_ = ~new_n28972_ | ~new_n8413_;
  assign new_n10406_ = ~new_n8409_ | ~new_n10402_;
  assign new_n10407_ = ~pi739 | ~po754;
  assign new_n10408_ = ~new_n8414_ | ~new_n8455_;
  assign new_n10409_ = ~new_n8410_ | ~new_n8441_;
  assign new_n10410_ = ~pi740 | ~new_n8682_;
  assign new_n10411_ = ~new_n10410_ | ~new_n10409_ | ~new_n10408_;
  assign new_n10412_ = ~new_n8773_ | ~new_n10798_;
  assign new_n10413_ = ~pi740 | ~new_n8749_;
  assign new_n10414_ = ~new_n28960_ | ~new_n8413_;
  assign new_n10415_ = ~new_n8409_ | ~new_n10411_;
  assign new_n10416_ = ~pi740 | ~po754;
  assign new_n10417_ = ~new_n8414_ | ~new_n8439_;
  assign new_n10418_ = ~new_n8410_ | ~new_n8449_;
  assign new_n10419_ = ~new_n25068_ | ~new_n8682_;
  assign new_n10420_ = ~new_n10419_ | ~new_n10418_ | ~new_n10417_;
  assign new_n10421_ = ~new_n8800_ | ~new_n10798_;
  assign new_n10422_ = ~new_n25068_ | ~new_n8749_;
  assign new_n10423_ = ~new_n28977_ | ~new_n8413_;
  assign new_n10424_ = ~new_n8409_ | ~new_n10420_;
  assign new_n10425_ = ~pi741 | ~po754;
  assign new_n10426_ = ~new_n8414_ | ~new_n8452_;
  assign new_n10427_ = ~new_n8410_ | ~new_n8443_;
  assign new_n10428_ = ~new_n25076_ | ~new_n8682_;
  assign new_n10429_ = ~new_n10428_ | ~new_n10427_ | ~new_n10426_;
  assign new_n10430_ = ~new_n8423_ | ~new_n9283_;
  assign new_n10431_ = ~new_n8422_ | ~new_n25076_;
  assign new_n10432_ = ~new_n28968_ | ~new_n8413_;
  assign new_n10433_ = ~new_n8409_ | ~new_n10429_;
  assign new_n10434_ = ~pi742 | ~po754;
  assign new_n10435_ = ~new_n8414_ | ~new_n8449_;
  assign new_n10436_ = ~new_n8410_ | ~new_n8456_;
  assign new_n10437_ = ~new_n25083_ | ~new_n8682_;
  assign new_n10438_ = ~new_n10437_ | ~new_n10436_ | ~new_n10435_;
  assign new_n10439_ = ~new_n8806_ | ~new_n10798_;
  assign new_n10440_ = ~new_n25083_ | ~new_n8749_;
  assign new_n10441_ = ~new_n28873_ | ~new_n8413_;
  assign new_n10442_ = ~new_n8409_ | ~new_n10438_;
  assign new_n10443_ = ~pi743 | ~po754;
  assign new_n10444_ = ~new_n8414_ | ~new_n8458_;
  assign new_n10445_ = ~new_n8410_ | ~new_n8452_;
  assign new_n10446_ = ~new_n25079_ | ~new_n8682_;
  assign new_n10447_ = ~new_n10446_ | ~new_n10445_ | ~new_n10444_;
  assign new_n10448_ = ~new_n8423_ | ~new_n9285_;
  assign new_n10449_ = ~new_n8422_ | ~new_n25079_;
  assign new_n10450_ = ~new_n28969_ | ~new_n8413_;
  assign new_n10451_ = ~new_n8409_ | ~new_n10447_;
  assign new_n10452_ = ~pi744 | ~po754;
  assign new_n10453_ = ~new_n8409_ | ~new_n8682_;
  assign new_n10454_ = ~new_n10797_ | ~new_n10453_;
  assign new_n10455_ = ~new_n9165_ | ~new_n8410_;
  assign new_n10456_ = ~new_n8765_ | ~new_n10798_;
  assign new_n10457_ = ~pi745 | ~new_n10454_;
  assign new_n10458_ = ~new_n28954_ | ~new_n8413_;
  assign new_n10459_ = ~pi745 | ~po754;
  assign new_n10460_ = ~new_n8414_ | ~new_n8461_;
  assign new_n10461_ = ~new_n8410_ | ~new_n8439_;
  assign new_n10462_ = ~new_n25073_ | ~new_n8682_;
  assign new_n10463_ = ~new_n10462_ | ~new_n10461_ | ~new_n10460_;
  assign new_n10464_ = ~new_n8794_ | ~new_n10798_;
  assign new_n10465_ = ~new_n25073_ | ~new_n8749_;
  assign new_n10466_ = ~new_n28955_ | ~new_n8413_;
  assign new_n10467_ = ~new_n8409_ | ~new_n10463_;
  assign new_n10468_ = ~pi746 | ~po754;
  assign new_n10469_ = ~new_n8414_ | ~new_n8441_;
  assign new_n10470_ = ~new_n8410_ | ~new_n8444_;
  assign new_n10471_ = ~new_n25088_ | ~new_n8682_;
  assign new_n10472_ = ~new_n10471_ | ~new_n10470_ | ~new_n10469_;
  assign new_n10473_ = ~new_n8779_ | ~new_n10798_;
  assign new_n10474_ = ~new_n25088_ | ~new_n8749_;
  assign new_n10475_ = ~new_n28959_ | ~new_n8413_;
  assign new_n10476_ = ~new_n8409_ | ~new_n10472_;
  assign new_n10477_ = ~pi747 | ~po754;
  assign new_n10478_ = ~new_n8414_ | ~new_n8443_;
  assign new_n10479_ = ~new_n8410_ | ~new_n8435_;
  assign new_n10480_ = ~new_n25069_ | ~new_n8682_;
  assign new_n10481_ = ~new_n10480_ | ~new_n10479_ | ~new_n10478_;
  assign new_n10482_ = ~new_n8423_ | ~new_n9281_;
  assign new_n10483_ = ~new_n8422_ | ~new_n25069_;
  assign new_n10484_ = ~new_n28966_ | ~new_n8413_;
  assign new_n10485_ = ~new_n8409_ | ~new_n10481_;
  assign new_n10486_ = ~pi748 | ~po754;
  assign new_n10487_ = ~new_n8414_ | ~new_n8450_;
  assign new_n10488_ = ~new_n8410_ | ~new_n8459_;
  assign new_n10489_ = ~new_n25078_ | ~new_n8682_;
  assign new_n10490_ = ~new_n10489_ | ~new_n10488_ | ~new_n10487_;
  assign new_n10491_ = ~new_n8818_ | ~new_n10798_;
  assign new_n10492_ = ~new_n25078_ | ~new_n8749_;
  assign new_n10493_ = ~new_n28874_ | ~new_n8413_;
  assign new_n10494_ = ~new_n8409_ | ~new_n10490_;
  assign new_n10495_ = ~pi749 | ~po754;
  assign new_n10496_ = ~new_n8414_ | ~new_n8437_;
  assign new_n10497_ = ~new_n8410_ | ~new_n8448_;
  assign new_n10498_ = ~new_n25112_ | ~new_n8682_;
  assign new_n10499_ = ~new_n10498_ | ~new_n10497_ | ~new_n10496_;
  assign new_n10500_ = ~new_n8782_ | ~new_n10798_;
  assign new_n10501_ = ~new_n25112_ | ~new_n8749_;
  assign new_n10502_ = ~new_n28958_ | ~new_n8413_;
  assign new_n10503_ = ~new_n8409_ | ~new_n10499_;
  assign new_n10504_ = ~pi750 | ~po754;
  assign new_n10505_ = ~new_n8414_ | ~new_n8451_;
  assign new_n10506_ = ~new_n8410_ | ~new_n8446_;
  assign new_n10507_ = ~new_n25066_ | ~new_n8682_;
  assign new_n10508_ = ~new_n10507_ | ~new_n10506_ | ~new_n10505_;
  assign new_n10509_ = ~new_n8815_ | ~new_n10798_;
  assign new_n10510_ = ~new_n25066_ | ~new_n8749_;
  assign new_n10511_ = ~new_n28973_ | ~new_n8413_;
  assign new_n10512_ = ~new_n8409_ | ~new_n10508_;
  assign new_n10513_ = ~pi751 | ~po754;
  assign new_n10514_ = ~new_n8414_ | ~new_n8442_;
  assign new_n10515_ = ~new_n8410_ | ~new_n8434_;
  assign new_n10516_ = ~new_n25075_ | ~new_n8682_;
  assign new_n10517_ = ~new_n10516_ | ~new_n10515_ | ~new_n10514_;
  assign new_n10518_ = ~new_n8423_ | ~new_n9280_;
  assign new_n10519_ = ~new_n8422_ | ~new_n25075_;
  assign new_n10520_ = ~new_n28965_ | ~new_n8413_;
  assign new_n10521_ = ~new_n8409_ | ~new_n10517_;
  assign new_n10522_ = ~pi752 | ~po754;
  assign new_n10523_ = ~new_n8414_ | ~new_n8440_;
  assign new_n10524_ = ~new_n8410_ | ~new_n8457_;
  assign new_n10525_ = ~new_n25082_ | ~new_n8682_;
  assign new_n10526_ = ~new_n10525_ | ~new_n10524_ | ~new_n10523_;
  assign new_n10527_ = ~new_n8803_ | ~new_n10798_;
  assign new_n10528_ = ~new_n25082_ | ~new_n8749_;
  assign new_n10529_ = ~new_n28976_ | ~new_n8413_;
  assign new_n10530_ = ~new_n8409_ | ~new_n10526_;
  assign new_n10531_ = ~pi753 | ~po754;
  assign new_n10532_ = ~new_n8414_ | ~new_n8453_;
  assign new_n10533_ = ~new_n8410_ | ~new_n8438_;
  assign new_n10534_ = ~new_n25086_ | ~new_n8682_;
  assign new_n10535_ = ~new_n10534_ | ~new_n10533_ | ~new_n10532_;
  assign new_n10536_ = ~new_n8423_ | ~new_n9284_;
  assign new_n10537_ = ~new_n8422_ | ~new_n25086_;
  assign new_n10538_ = ~new_n28875_ | ~new_n8413_;
  assign new_n10539_ = ~new_n8409_ | ~new_n10535_;
  assign new_n10540_ = ~pi754 | ~po754;
  assign new_n10541_ = ~new_n8414_ | ~new_n8454_;
  assign new_n10542_ = ~new_n8410_ | ~new_n8445_;
  assign new_n10543_ = ~pi755 | ~new_n8682_;
  assign new_n10544_ = ~new_n10543_ | ~new_n10542_ | ~new_n10541_;
  assign new_n10545_ = ~new_n8770_ | ~new_n10798_;
  assign new_n10546_ = ~pi755 | ~new_n8749_;
  assign new_n10547_ = ~new_n28970_ | ~new_n8413_;
  assign new_n10548_ = ~new_n8409_ | ~new_n10544_;
  assign new_n10549_ = ~pi755 | ~po754;
  assign new_n10550_ = ~new_n8414_ | ~new_n8447_;
  assign new_n10551_ = ~new_n8410_ | ~new_n8460_;
  assign new_n10552_ = ~new_n25071_ | ~new_n8682_;
  assign new_n10553_ = ~new_n10552_ | ~new_n10551_ | ~new_n10550_;
  assign new_n10554_ = ~new_n8791_ | ~new_n10798_;
  assign new_n10555_ = ~new_n25071_ | ~new_n8749_;
  assign new_n10556_ = ~new_n28956_ | ~new_n8413_;
  assign new_n10557_ = ~new_n8409_ | ~new_n10553_;
  assign new_n10558_ = ~pi756 | ~po754;
  assign new_n10559_ = ~new_n8414_ | ~new_n8430_;
  assign new_n10560_ = ~new_n8410_ | ~new_n8432_;
  assign new_n10561_ = ~new_n25087_ | ~new_n8682_;
  assign new_n10562_ = ~new_n10561_ | ~new_n10560_ | ~new_n10559_;
  assign new_n10563_ = ~new_n8423_ | ~new_n9277_;
  assign new_n10564_ = ~new_n8422_ | ~new_n25087_;
  assign new_n10565_ = ~new_n28961_ | ~new_n8413_;
  assign new_n10566_ = ~new_n8409_ | ~new_n10562_;
  assign new_n10567_ = ~pi757 | ~po754;
  assign new_n10568_ = ~new_n8414_ | ~new_n8459_;
  assign new_n10569_ = ~new_n8410_ | ~new_n8453_;
  assign new_n10570_ = ~new_n25074_ | ~new_n8682_;
  assign new_n10571_ = ~new_n10570_ | ~new_n10569_ | ~new_n10568_;
  assign new_n10572_ = ~new_n8823_ | ~new_n10798_;
  assign new_n10573_ = ~new_n25074_ | ~new_n8749_;
  assign new_n10574_ = ~new_n28971_ | ~new_n8413_;
  assign new_n10575_ = ~new_n8409_ | ~new_n10571_;
  assign new_n10576_ = ~pi758 | ~po754;
  assign new_n10577_ = ~new_n8414_ | ~new_n8445_;
  assign new_n10578_ = ~new_n8410_ | ~new_n8437_;
  assign new_n10579_ = ~new_n25084_ | ~new_n8682_;
  assign new_n10580_ = ~new_n10579_ | ~new_n10578_ | ~new_n10577_;
  assign new_n10581_ = ~new_n8776_ | ~new_n10798_;
  assign new_n10582_ = ~new_n25084_ | ~new_n8749_;
  assign new_n10583_ = ~new_n28877_ | ~new_n8413_;
  assign new_n10584_ = ~new_n8409_ | ~new_n10580_;
  assign new_n10585_ = ~pi759 | ~po754;
  assign new_n10586_ = ~new_n8414_ | ~new_n8460_;
  assign new_n10587_ = ~new_n8410_ | ~new_n8440_;
  assign new_n10588_ = ~new_n25072_ | ~new_n8682_;
  assign new_n10589_ = ~new_n10588_ | ~new_n10587_ | ~new_n10586_;
  assign new_n10590_ = ~new_n8797_ | ~new_n10798_;
  assign new_n10591_ = ~new_n25072_ | ~new_n8749_;
  assign new_n10592_ = ~new_n28978_ | ~new_n8413_;
  assign new_n10593_ = ~new_n8409_ | ~new_n10589_;
  assign new_n10594_ = ~pi760 | ~po754;
  assign new_n10595_ = ~new_n8414_ | ~new_n8438_;
  assign new_n10596_ = ~new_n8410_ | ~new_n8442_;
  assign new_n10597_ = ~new_n25065_ | ~new_n8682_;
  assign new_n10598_ = ~new_n10597_ | ~new_n10596_ | ~new_n10595_;
  assign new_n10599_ = ~new_n8423_ | ~new_n9282_;
  assign new_n10600_ = ~new_n8422_ | ~new_n25065_;
  assign new_n10601_ = ~new_n28967_ | ~new_n8413_;
  assign new_n10602_ = ~new_n8409_ | ~new_n10598_;
  assign new_n10603_ = ~pi761 | ~po754;
  assign new_n10604_ = ~new_n8414_ | ~new_n8457_;
  assign new_n10605_ = ~new_n8410_ | ~new_n8451_;
  assign new_n10606_ = ~new_n25089_ | ~new_n8682_;
  assign new_n10607_ = ~new_n10606_ | ~new_n10605_ | ~new_n10604_;
  assign new_n10608_ = ~new_n8809_ | ~new_n10798_;
  assign new_n10609_ = ~new_n25089_ | ~new_n8749_;
  assign new_n10610_ = ~new_n28975_ | ~new_n8413_;
  assign new_n10611_ = ~new_n8409_ | ~new_n10607_;
  assign new_n10612_ = ~pi762 | ~po754;
  assign new_n10613_ = ~new_n8414_ | ~new_n8434_;
  assign new_n10614_ = ~new_n8410_ | ~new_n8431_;
  assign new_n10615_ = ~new_n25081_ | ~new_n8682_;
  assign new_n10616_ = ~new_n10615_ | ~new_n10614_ | ~new_n10613_;
  assign new_n10617_ = ~new_n8423_ | ~new_n9278_;
  assign new_n10618_ = ~new_n8422_ | ~new_n25081_;
  assign new_n10619_ = ~new_n28962_ | ~new_n8413_;
  assign new_n10620_ = ~new_n8409_ | ~new_n10616_;
  assign new_n10621_ = ~pi763 | ~po754;
  assign new_n10622_ = ~new_n8414_ | ~new_n8448_;
  assign new_n10623_ = ~new_n8410_ | ~new_n8461_;
  assign new_n10624_ = ~new_n25077_ | ~new_n8682_;
  assign new_n10625_ = ~new_n10624_ | ~new_n10623_ | ~new_n10622_;
  assign new_n10626_ = ~new_n8788_ | ~new_n10798_;
  assign new_n10627_ = ~new_n25077_ | ~new_n8749_;
  assign new_n10628_ = ~new_n28878_ | ~new_n8413_;
  assign new_n10629_ = ~new_n8409_ | ~new_n10625_;
  assign new_n10630_ = ~pi764 | ~po754;
  assign new_n10631_ = ~new_n9276_ | ~new_n8424_;
  assign new_n10632_ = ~new_n8753_ | ~new_n9211_;
  assign new_n10633_ = ~new_n9194_ | ~new_n9193_;
  assign new_n10634_ = ~new_n9192_ | ~new_n8391_;
  assign new_n10635_ = ~new_n9258_ | ~new_n10634_;
  assign new_n10636_ = ~new_n8794_ | ~new_n10635_;
  assign new_n10637_ = ~new_n10633_ | ~new_n8460_;
  assign new_n10638_ = ~new_n8791_ | ~new_n10635_;
  assign new_n10639_ = ~new_n10633_ | ~new_n8461_;
  assign new_n10640_ = ~new_n8788_ | ~new_n10635_;
  assign new_n10641_ = ~new_n10633_ | ~new_n8447_;
  assign new_n10642_ = ~new_n8785_ | ~new_n10635_;
  assign new_n10643_ = ~new_n10633_ | ~new_n8448_;
  assign new_n10644_ = ~new_n8782_ | ~new_n10635_;
  assign new_n10645_ = ~new_n10633_ | ~new_n8444_;
  assign new_n10646_ = ~new_n8779_ | ~new_n10635_;
  assign new_n10647_ = ~new_n10633_ | ~new_n8437_;
  assign new_n10648_ = ~new_n9250_ | ~new_n10635_;
  assign new_n10649_ = ~new_n10633_ | ~new_n8433_;
  assign new_n10650_ = ~new_n9251_ | ~new_n10635_;
  assign new_n10651_ = ~new_n10633_ | ~new_n8436_;
  assign new_n10652_ = ~new_n8776_ | ~new_n10635_;
  assign new_n10653_ = ~new_n10633_ | ~new_n8441_;
  assign new_n10654_ = ~new_n9286_ | ~new_n10635_;
  assign new_n10655_ = ~new_n10633_ | ~new_n8432_;
  assign new_n10656_ = ~new_n9277_ | ~new_n10635_;
  assign new_n10657_ = ~new_n10633_ | ~new_n8431_;
  assign new_n10658_ = ~new_n9278_ | ~new_n10635_;
  assign new_n10659_ = ~new_n10633_ | ~new_n8430_;
  assign new_n10660_ = ~new_n9279_ | ~new_n10635_;
  assign new_n10661_ = ~new_n10633_ | ~new_n8434_;
  assign new_n10662_ = ~new_n9280_ | ~new_n10635_;
  assign new_n10663_ = ~new_n10633_ | ~new_n8435_;
  assign new_n10664_ = ~new_n9281_ | ~new_n10635_;
  assign new_n10665_ = ~new_n10633_ | ~new_n8442_;
  assign new_n10666_ = ~new_n9282_ | ~new_n10635_;
  assign new_n10667_ = ~new_n10633_ | ~new_n8443_;
  assign new_n10668_ = ~new_n9283_ | ~new_n10635_;
  assign new_n10669_ = ~new_n10633_ | ~new_n8438_;
  assign new_n10670_ = ~new_n9284_ | ~new_n10635_;
  assign new_n10671_ = ~new_n10633_ | ~new_n8452_;
  assign new_n10672_ = ~new_n9285_ | ~new_n10635_;
  assign new_n10673_ = ~new_n10633_ | ~new_n8453_;
  assign new_n10674_ = ~new_n8773_ | ~new_n10635_;
  assign new_n10675_ = ~new_n10633_ | ~new_n8445_;
  assign new_n10676_ = ~new_n8823_ | ~new_n10635_;
  assign new_n10677_ = ~new_n10633_ | ~new_n8458_;
  assign new_n10678_ = ~new_n8821_ | ~new_n10635_;
  assign new_n10679_ = ~new_n10633_ | ~new_n8459_;
  assign new_n10680_ = ~new_n8818_ | ~new_n10635_;
  assign new_n10681_ = ~new_n10633_ | ~new_n8446_;
  assign new_n10682_ = ~new_n8815_ | ~new_n10635_;
  assign new_n10683_ = ~new_n10633_ | ~new_n8450_;
  assign new_n10684_ = ~new_n8812_ | ~new_n10635_;
  assign new_n10685_ = ~new_n10633_ | ~new_n8451_;
  assign new_n10686_ = ~new_n8809_ | ~new_n10635_;
  assign new_n10687_ = ~new_n10633_ | ~new_n8456_;
  assign new_n10688_ = ~new_n8806_ | ~new_n10635_;
  assign new_n10689_ = ~new_n10633_ | ~new_n8457_;
  assign new_n10690_ = ~new_n8803_ | ~new_n10635_;
  assign new_n10691_ = ~new_n10633_ | ~new_n8449_;
  assign new_n10692_ = ~new_n8800_ | ~new_n10635_;
  assign new_n10693_ = ~new_n10633_ | ~new_n8440_;
  assign new_n10694_ = ~new_n8797_ | ~new_n10635_;
  assign new_n10695_ = ~new_n10633_ | ~new_n8439_;
  assign new_n10696_ = ~new_n8770_ | ~new_n10635_;
  assign new_n10697_ = ~new_n10633_ | ~new_n8455_;
  assign new_n10698_ = ~new_n8765_ | ~new_n10635_;
  assign new_n10699_ = ~new_n10633_ | ~new_n8454_;
  assign new_n10700_ = ~new_n8794_ | ~new_n10633_;
  assign new_n10701_ = ~new_n10635_ | ~new_n8460_;
  assign new_n10702_ = ~new_n10818_ | ~new_n8461_;
  assign new_n10703_ = ~new_n8791_ | ~new_n10633_;
  assign new_n10704_ = ~new_n10635_ | ~new_n8461_;
  assign new_n10705_ = ~new_n10818_ | ~new_n8447_;
  assign new_n10706_ = ~new_n8788_ | ~new_n10633_;
  assign new_n10707_ = ~new_n10635_ | ~new_n8447_;
  assign new_n10708_ = ~new_n10818_ | ~new_n8448_;
  assign new_n10709_ = ~new_n8785_ | ~new_n10633_;
  assign new_n10710_ = ~new_n10635_ | ~new_n8448_;
  assign new_n10711_ = ~new_n10818_ | ~new_n8444_;
  assign new_n10712_ = ~new_n8782_ | ~new_n10633_;
  assign new_n10713_ = ~new_n10635_ | ~new_n8444_;
  assign new_n10714_ = ~new_n10818_ | ~new_n8437_;
  assign new_n10715_ = ~new_n8779_ | ~new_n10633_;
  assign new_n10716_ = ~new_n10635_ | ~new_n8437_;
  assign new_n10717_ = ~new_n10818_ | ~new_n8441_;
  assign new_n10718_ = ~new_n10635_ | ~new_n8433_;
  assign new_n10719_ = ~new_n9250_ | ~new_n10633_;
  assign new_n10720_ = ~new_n10635_ | ~new_n8436_;
  assign new_n10721_ = ~new_n9251_ | ~new_n10633_;
  assign new_n10722_ = ~new_n8776_ | ~new_n10633_;
  assign new_n10723_ = ~new_n10635_ | ~new_n8441_;
  assign new_n10724_ = ~new_n10818_ | ~new_n8445_;
  assign new_n10725_ = ~new_n10635_ | ~new_n8432_;
  assign new_n10726_ = ~new_n9286_ | ~new_n10633_;
  assign new_n10727_ = ~new_n10818_ | ~new_n8431_;
  assign new_n10728_ = ~new_n10635_ | ~new_n8431_;
  assign new_n10729_ = ~new_n9277_ | ~new_n10633_;
  assign new_n10730_ = ~new_n10818_ | ~new_n8430_;
  assign new_n10731_ = ~new_n10635_ | ~new_n8430_;
  assign new_n10732_ = ~new_n9278_ | ~new_n10633_;
  assign new_n10733_ = ~new_n10818_ | ~new_n8434_;
  assign new_n10734_ = ~new_n10635_ | ~new_n8434_;
  assign new_n10735_ = ~new_n9279_ | ~new_n10633_;
  assign new_n10736_ = ~new_n10818_ | ~new_n8435_;
  assign new_n10737_ = ~new_n10635_ | ~new_n8435_;
  assign new_n10738_ = ~new_n9280_ | ~new_n10633_;
  assign new_n10739_ = ~new_n10818_ | ~new_n8442_;
  assign new_n10740_ = ~new_n10635_ | ~new_n8442_;
  assign new_n10741_ = ~new_n9281_ | ~new_n10633_;
  assign new_n10742_ = ~new_n10818_ | ~new_n8443_;
  assign new_n10743_ = ~new_n10635_ | ~new_n8443_;
  assign new_n10744_ = ~new_n9282_ | ~new_n10633_;
  assign new_n10745_ = ~new_n10818_ | ~new_n8438_;
  assign new_n10746_ = ~new_n10635_ | ~new_n8438_;
  assign new_n10747_ = ~new_n9283_ | ~new_n10633_;
  assign new_n10748_ = ~new_n10818_ | ~new_n8452_;
  assign new_n10749_ = ~new_n10635_ | ~new_n8452_;
  assign new_n10750_ = ~new_n9284_ | ~new_n10633_;
  assign new_n10751_ = ~new_n10818_ | ~new_n8453_;
  assign new_n10752_ = ~new_n10635_ | ~new_n8453_;
  assign new_n10753_ = ~new_n9285_ | ~new_n10633_;
  assign new_n10754_ = ~new_n10818_ | ~new_n8458_;
  assign new_n10755_ = ~new_n8773_ | ~new_n10633_;
  assign new_n10756_ = ~new_n10635_ | ~new_n8445_;
  assign new_n10757_ = ~new_n10818_ | ~new_n8455_;
  assign new_n10758_ = ~new_n8823_ | ~new_n10633_;
  assign new_n10759_ = ~new_n10635_ | ~new_n8458_;
  assign new_n10760_ = ~new_n10818_ | ~new_n8459_;
  assign new_n10761_ = ~new_n8821_ | ~new_n10633_;
  assign new_n10762_ = ~new_n10635_ | ~new_n8459_;
  assign new_n10763_ = ~new_n10818_ | ~new_n8446_;
  assign new_n10764_ = ~new_n8818_ | ~new_n10633_;
  assign new_n10765_ = ~new_n10635_ | ~new_n8446_;
  assign new_n10766_ = ~new_n10818_ | ~new_n8450_;
  assign new_n10767_ = ~new_n8815_ | ~new_n10633_;
  assign new_n10768_ = ~new_n10635_ | ~new_n8450_;
  assign new_n10769_ = ~new_n10818_ | ~new_n8451_;
  assign new_n10770_ = ~new_n8812_ | ~new_n10633_;
  assign new_n10771_ = ~new_n10635_ | ~new_n8451_;
  assign new_n10772_ = ~new_n10818_ | ~new_n8456_;
  assign new_n10773_ = ~new_n8809_ | ~new_n10633_;
  assign new_n10774_ = ~new_n10635_ | ~new_n8456_;
  assign new_n10775_ = ~new_n10818_ | ~new_n8457_;
  assign new_n10776_ = ~new_n8806_ | ~new_n10633_;
  assign new_n10777_ = ~new_n10635_ | ~new_n8457_;
  assign new_n10778_ = ~new_n10818_ | ~new_n8449_;
  assign new_n10779_ = ~new_n8803_ | ~new_n10633_;
  assign new_n10780_ = ~new_n10635_ | ~new_n8449_;
  assign new_n10781_ = ~new_n10818_ | ~new_n8440_;
  assign new_n10782_ = ~new_n8800_ | ~new_n10633_;
  assign new_n10783_ = ~new_n10635_ | ~new_n8440_;
  assign new_n10784_ = ~new_n10818_ | ~new_n8439_;
  assign new_n10785_ = ~new_n8797_ | ~new_n10633_;
  assign new_n10786_ = ~new_n10635_ | ~new_n8439_;
  assign new_n10787_ = ~new_n10818_ | ~new_n8460_;
  assign new_n10788_ = ~new_n8770_ | ~new_n10633_;
  assign new_n10789_ = ~new_n10635_ | ~new_n8455_;
  assign new_n10790_ = ~new_n10818_ | ~new_n8454_;
  assign new_n10791_ = ~new_n8765_ | ~new_n10633_;
  assign new_n10792_ = ~new_n10635_ | ~new_n8454_;
  assign new_n10793_ = ~new_n10359_ | ~po754;
  assign new_n10794_ = ~new_n10358_ | ~new_n10359_ | ~new_n10818_;
  assign new_n10795_ = ~new_n8421_ | ~new_n8681_;
  assign new_n10796_ = ~new_n8421_ | ~new_n9272_;
  assign new_n10797_ = ~new_n8749_;
  assign new_n10798_ = ~new_n10796_ | ~new_n9296_;
  assign new_n10799_ = ~new_n9152_ | ~new_n11316_ | ~new_n11315_;
  assign new_n10800_ = ~new_n10812_ | ~new_n10806_;
  assign new_n10801_ = ~new_n9257_ | ~new_n8756_;
  assign new_n10802_ = ~new_n8753_ | ~new_n9211_;
  assign new_n10803_ = ~new_n9254_ | ~new_n10825_;
  assign new_n10804_ = ~pi547 | ~new_n9209_;
  assign new_n10805_ = ~pi554 | ~new_n24731_;
  assign new_n10806_ = ~new_n8750_;
  assign new_n10807_ = ~pi548 | ~new_n9209_;
  assign new_n10808_ = ~pi554 | ~new_n24794_;
  assign new_n10809_ = ~new_n8751_;
  assign new_n10810_ = ~pi549 | ~new_n9209_;
  assign new_n10811_ = ~pi554 | ~new_n24732_;
  assign new_n10812_ = ~new_n8752_;
  assign new_n10813_ = ~new_n10806_ | ~pi735;
  assign new_n10814_ = ~new_n8750_ | ~new_n8676_;
  assign new_n10815_ = ~new_n10814_ | ~new_n10813_;
  assign new_n10816_ = ~pi546 | ~new_n9209_;
  assign new_n10817_ = ~pi554 | ~new_n24730_;
  assign new_n10818_ = ~new_n8753_;
  assign new_n10819_ = ~pi555 | ~new_n9210_;
  assign new_n10820_ = ~new_n9293_ | ~new_n9398_;
  assign new_n10821_ = ~pi556 | ~new_n9210_;
  assign new_n10822_ = ~new_n9293_ | ~new_n9399_;
  assign new_n10823_ = ~pi543 | ~new_n9209_;
  assign new_n10824_ = ~pi554 | ~new_n24728_;
  assign new_n10825_ = ~new_n8756_;
  assign new_n10826_ = ~pi542 | ~new_n9209_;
  assign new_n10827_ = ~pi554 | ~new_n24727_;
  assign new_n10828_ = ~new_n8757_;
  assign new_n10829_ = ~pi545 | ~new_n9209_;
  assign new_n10830_ = ~pi554 | ~new_n24729_;
  assign new_n10831_ = ~new_n8758_;
  assign new_n10832_ = ~pi544 | ~new_n9209_;
  assign new_n10833_ = ~pi554 | ~new_n24796_;
  assign new_n10834_ = ~new_n8763_;
  assign new_n10835_ = ~pi553 | ~new_n9209_;
  assign new_n10836_ = ~pi554 | ~new_n24790_;
  assign new_n10837_ = ~new_n8759_;
  assign new_n10838_ = ~pi552 | ~new_n9209_;
  assign new_n10839_ = ~pi554 | ~new_n24734_;
  assign new_n10840_ = ~new_n8760_;
  assign new_n10841_ = ~pi551 | ~new_n9209_;
  assign new_n10842_ = ~pi554 | ~new_n24733_;
  assign new_n10843_ = ~new_n8761_;
  assign new_n10844_ = ~pi550 | ~new_n9209_;
  assign new_n10845_ = ~pi554 | ~new_n24792_;
  assign new_n10846_ = ~new_n8762_;
  assign new_n10847_ = ~pi523 | ~new_n9209_;
  assign new_n10848_ = ~pi554 | ~pi523;
  assign new_n10849_ = ~new_n1562_ | ~new_n9211_;
  assign new_n10850_ = ~new_n9271_ | ~new_n8764_;
  assign new_n10851_ = ~new_n8765_;
  assign new_n10852_ = ~new_n10800_ | ~new_n8678_;
  assign new_n10853_ = ~pi555 | ~new_n9397_;
  assign new_n10854_ = ~new_n8766_;
  assign new_n10855_ = ~pi556 | ~new_n9397_;
  assign new_n10856_ = ~new_n9399_ | ~new_n8678_;
  assign new_n10857_ = ~new_n8767_;
  assign new_n10858_ = ~new_n9430_ | ~new_n10831_;
  assign new_n10859_ = ~new_n8758_ | ~new_n9212_;
  assign new_n10860_ = ~new_n10859_ | ~new_n10858_;
  assign new_n10861_ = ~pi587 | ~new_n9213_;
  assign new_n10862_ = ~new_n9292_ | ~new_n9455_;
  assign new_n10863_ = ~pi524 | ~new_n9209_;
  assign new_n10864_ = ~pi554 | ~new_n24764_;
  assign new_n10865_ = ~new_n1551_ | ~new_n9211_;
  assign new_n10866_ = ~new_n8769_ | ~new_n9271_;
  assign new_n10867_ = ~new_n8770_;
  assign new_n10868_ = ~pi588 | ~new_n9213_;
  assign new_n10869_ = ~new_n9292_ | ~new_n9480_;
  assign new_n10870_ = ~pi525 | ~new_n9209_;
  assign new_n10871_ = ~pi554 | ~new_n24735_;
  assign new_n10872_ = ~new_n1540_ | ~new_n9211_;
  assign new_n10873_ = ~new_n8772_ | ~new_n9271_;
  assign new_n10874_ = ~new_n8773_;
  assign new_n10875_ = ~pi589 | ~new_n9213_;
  assign new_n10876_ = ~new_n9292_ | ~new_n9498_;
  assign new_n10877_ = ~pi526 | ~new_n9209_;
  assign new_n10878_ = ~pi554 | ~new_n24736_;
  assign new_n10879_ = ~new_n1537_ | ~new_n9211_;
  assign new_n10880_ = ~new_n8775_ | ~new_n9271_;
  assign new_n10881_ = ~new_n8776_;
  assign new_n10882_ = ~pi590 | ~new_n9213_;
  assign new_n10883_ = ~new_n9292_ | ~new_n9516_;
  assign new_n10884_ = ~pi527 | ~new_n9209_;
  assign new_n10885_ = ~pi554 | ~new_n24737_;
  assign new_n10886_ = ~new_n1536_ | ~new_n9211_;
  assign new_n10887_ = ~new_n8778_ | ~new_n9271_;
  assign new_n10888_ = ~new_n8779_;
  assign new_n10889_ = ~pi591 | ~new_n9213_;
  assign new_n10890_ = ~new_n9292_ | ~new_n9534_;
  assign new_n10891_ = ~pi528 | ~new_n9209_;
  assign new_n10892_ = ~pi554 | ~new_n24787_;
  assign new_n10893_ = ~new_n1535_ | ~new_n9211_;
  assign new_n10894_ = ~new_n8781_ | ~new_n9271_;
  assign new_n10895_ = ~new_n8782_;
  assign new_n10896_ = ~pi592 | ~new_n9213_;
  assign new_n10897_ = ~new_n9292_ | ~new_n9552_;
  assign new_n10898_ = ~pi529 | ~new_n9209_;
  assign new_n10899_ = ~pi554 | ~new_n24738_;
  assign new_n10900_ = ~new_n1534_ | ~new_n9211_;
  assign new_n10901_ = ~new_n8784_ | ~new_n9271_;
  assign new_n10902_ = ~new_n8785_;
  assign new_n10903_ = ~pi593 | ~new_n9213_;
  assign new_n10904_ = ~new_n9292_ | ~new_n9570_;
  assign new_n10905_ = ~pi530 | ~new_n9209_;
  assign new_n10906_ = ~pi554 | ~new_n24739_;
  assign new_n10907_ = ~new_n1533_ | ~new_n9211_;
  assign new_n10908_ = ~new_n8787_ | ~new_n9271_;
  assign new_n10909_ = ~new_n8788_;
  assign new_n10910_ = ~pi594 | ~new_n9213_;
  assign new_n10911_ = ~new_n9292_ | ~new_n9588_;
  assign new_n10912_ = ~pi531 | ~new_n9209_;
  assign new_n10913_ = ~pi554 | ~new_n24740_;
  assign new_n10914_ = ~new_n1532_ | ~new_n9211_;
  assign new_n10915_ = ~new_n8790_ | ~new_n9271_;
  assign new_n10916_ = ~new_n8791_;
  assign new_n10917_ = ~pi595 | ~new_n9213_;
  assign new_n10918_ = ~new_n9292_ | ~new_n9606_;
  assign new_n10919_ = ~pi532 | ~new_n9209_;
  assign new_n10920_ = ~pi554 | ~new_n24785_;
  assign new_n10921_ = ~new_n1531_ | ~new_n9211_;
  assign new_n10922_ = ~new_n8793_ | ~new_n9271_;
  assign new_n10923_ = ~new_n8794_;
  assign new_n10924_ = ~pi596 | ~new_n9213_;
  assign new_n10925_ = ~new_n9292_ | ~new_n9624_;
  assign new_n10926_ = ~pi533 | ~new_n9209_;
  assign new_n10927_ = ~pi554 | ~new_n24720_;
  assign new_n10928_ = ~new_n1561_ | ~new_n9211_;
  assign new_n10929_ = ~new_n8796_ | ~new_n9271_;
  assign new_n10930_ = ~new_n8797_;
  assign new_n10931_ = ~pi597 | ~new_n9213_;
  assign new_n10932_ = ~new_n9292_ | ~new_n9642_;
  assign new_n10933_ = ~pi534 | ~new_n9209_;
  assign new_n10934_ = ~pi554 | ~new_n24721_;
  assign new_n10935_ = ~new_n1560_ | ~new_n9211_;
  assign new_n10936_ = ~new_n8799_ | ~new_n9271_;
  assign new_n10937_ = ~new_n8800_;
  assign new_n10938_ = ~pi598 | ~new_n9213_;
  assign new_n10939_ = ~new_n9292_ | ~new_n9660_;
  assign new_n10940_ = ~pi535 | ~new_n9209_;
  assign new_n10941_ = ~pi554 | ~new_n24722_;
  assign new_n10942_ = ~new_n1559_ | ~new_n9211_;
  assign new_n10943_ = ~new_n8802_ | ~new_n9271_;
  assign new_n10944_ = ~new_n8803_;
  assign new_n10945_ = ~pi599 | ~new_n9213_;
  assign new_n10946_ = ~new_n9292_ | ~new_n9678_;
  assign new_n10947_ = ~pi536 | ~new_n9209_;
  assign new_n10948_ = ~pi554 | ~new_n24802_;
  assign new_n10949_ = ~new_n1558_ | ~new_n9211_;
  assign new_n10950_ = ~new_n8805_ | ~new_n9271_;
  assign new_n10951_ = ~new_n8806_;
  assign new_n10952_ = ~pi600 | ~new_n9213_;
  assign new_n10953_ = ~new_n9292_ | ~new_n9696_;
  assign new_n10954_ = ~pi537 | ~new_n9209_;
  assign new_n10955_ = ~pi554 | ~new_n24723_;
  assign new_n10956_ = ~new_n1557_ | ~new_n9211_;
  assign new_n10957_ = ~new_n8808_ | ~new_n9271_;
  assign new_n10958_ = ~new_n8809_;
  assign new_n10959_ = ~pi601 | ~new_n9213_;
  assign new_n10960_ = ~new_n9292_ | ~new_n9714_;
  assign new_n10961_ = ~pi538 | ~new_n9209_;
  assign new_n10962_ = ~pi554 | ~new_n24724_;
  assign new_n10963_ = ~new_n1556_ | ~new_n9211_;
  assign new_n10964_ = ~new_n8811_ | ~new_n9271_;
  assign new_n10965_ = ~new_n8812_;
  assign new_n10966_ = ~pi602 | ~new_n9213_;
  assign new_n10967_ = ~new_n9292_ | ~new_n9732_;
  assign new_n10968_ = ~pi539 | ~new_n9209_;
  assign new_n10969_ = ~pi554 | ~new_n24725_;
  assign new_n10970_ = ~new_n1555_ | ~new_n9211_;
  assign new_n10971_ = ~new_n8814_ | ~new_n9271_;
  assign new_n10972_ = ~new_n8815_;
  assign new_n10973_ = ~pi603 | ~new_n9213_;
  assign new_n10974_ = ~new_n9292_ | ~new_n9750_;
  assign new_n10975_ = ~pi540 | ~new_n9209_;
  assign new_n10976_ = ~pi554 | ~new_n24800_;
  assign new_n10977_ = ~new_n1554_ | ~new_n9211_;
  assign new_n10978_ = ~new_n8817_ | ~new_n9271_;
  assign new_n10979_ = ~new_n8818_;
  assign new_n10980_ = ~pi604 | ~new_n9213_;
  assign new_n10981_ = ~new_n9292_ | ~new_n9768_;
  assign new_n10982_ = ~pi541 | ~new_n9209_;
  assign new_n10983_ = ~pi554 | ~new_n24726_;
  assign new_n10984_ = ~new_n1553_ | ~new_n9211_;
  assign new_n10985_ = ~new_n8820_ | ~new_n9271_;
  assign new_n10986_ = ~new_n8821_;
  assign new_n10987_ = ~pi605 | ~new_n9213_;
  assign new_n10988_ = ~new_n9292_ | ~new_n9786_;
  assign new_n10989_ = ~new_n1552_ | ~new_n9211_;
  assign new_n10990_ = ~new_n9271_ | ~new_n8757_;
  assign new_n10991_ = ~new_n8823_;
  assign new_n10992_ = ~pi606 | ~new_n9213_;
  assign new_n10993_ = ~new_n9292_ | ~new_n9804_;
  assign new_n10994_ = ~pi607 | ~new_n9213_;
  assign new_n10995_ = ~new_n9292_ | ~new_n9822_;
  assign new_n10996_ = ~pi608 | ~new_n9213_;
  assign new_n10997_ = ~new_n9292_ | ~new_n9840_;
  assign new_n10998_ = ~pi609 | ~new_n9213_;
  assign new_n10999_ = ~new_n9292_ | ~new_n9858_;
  assign new_n11000_ = ~pi610 | ~new_n9213_;
  assign new_n11001_ = ~new_n9292_ | ~new_n9876_;
  assign new_n11002_ = ~pi611 | ~new_n9213_;
  assign new_n11003_ = ~new_n9292_ | ~new_n9894_;
  assign new_n11004_ = ~pi612 | ~new_n9213_;
  assign new_n11005_ = ~new_n9292_ | ~new_n9912_;
  assign new_n11006_ = ~pi613 | ~new_n9213_;
  assign new_n11007_ = ~new_n9292_ | ~new_n9930_;
  assign new_n11008_ = ~pi614 | ~new_n9213_;
  assign new_n11009_ = ~new_n9292_ | ~new_n9948_;
  assign new_n11010_ = ~pi615 | ~new_n9213_;
  assign new_n11011_ = ~new_n9292_ | ~new_n9966_;
  assign new_n11012_ = ~pi616 | ~new_n9213_;
  assign new_n11013_ = ~new_n9292_ | ~new_n9986_;
  assign new_n11014_ = ~pi617 | ~new_n9213_;
  assign new_n11015_ = ~new_n9292_ | ~new_n9993_;
  assign new_n11016_ = ~pi618 | ~new_n9213_;
  assign new_n11017_ = ~new_n9292_ | ~new_n9995_;
  assign new_n11018_ = ~new_n10831_ | ~new_n9212_;
  assign new_n11019_ = ~new_n9430_ | ~new_n10828_;
  assign new_n11020_ = ~pi619 | ~new_n9214_;
  assign new_n11021_ = ~new_n9291_ | ~new_n9455_;
  assign new_n11022_ = ~pi620 | ~new_n9214_;
  assign new_n11023_ = ~new_n9291_ | ~new_n9480_;
  assign new_n11024_ = ~pi621 | ~new_n9214_;
  assign new_n11025_ = ~new_n9291_ | ~new_n9498_;
  assign new_n11026_ = ~pi622 | ~new_n9214_;
  assign new_n11027_ = ~new_n9291_ | ~new_n9516_;
  assign new_n11028_ = ~pi623 | ~new_n9214_;
  assign new_n11029_ = ~new_n9291_ | ~new_n9534_;
  assign new_n11030_ = ~pi624 | ~new_n9214_;
  assign new_n11031_ = ~new_n9291_ | ~new_n9552_;
  assign new_n11032_ = ~pi625 | ~new_n9214_;
  assign new_n11033_ = ~new_n9291_ | ~new_n9570_;
  assign new_n11034_ = ~pi626 | ~new_n9214_;
  assign new_n11035_ = ~new_n9291_ | ~new_n9588_;
  assign new_n11036_ = ~pi627 | ~new_n9214_;
  assign new_n11037_ = ~new_n9291_ | ~new_n9606_;
  assign new_n11038_ = ~pi628 | ~new_n9214_;
  assign new_n11039_ = ~new_n9291_ | ~new_n9624_;
  assign new_n11040_ = ~pi629 | ~new_n9214_;
  assign new_n11041_ = ~new_n9291_ | ~new_n9642_;
  assign new_n11042_ = ~pi630 | ~new_n9214_;
  assign new_n11043_ = ~new_n9291_ | ~new_n9660_;
  assign new_n11044_ = ~pi631 | ~new_n9214_;
  assign new_n11045_ = ~new_n9291_ | ~new_n9678_;
  assign new_n11046_ = ~pi632 | ~new_n9214_;
  assign new_n11047_ = ~new_n9291_ | ~new_n9696_;
  assign new_n11048_ = ~pi633 | ~new_n9214_;
  assign new_n11049_ = ~new_n9291_ | ~new_n9714_;
  assign new_n11050_ = ~pi634 | ~new_n9214_;
  assign new_n11051_ = ~new_n9291_ | ~new_n9732_;
  assign new_n11052_ = ~pi635 | ~new_n9214_;
  assign new_n11053_ = ~new_n9291_ | ~new_n9750_;
  assign new_n11054_ = ~pi636 | ~new_n9214_;
  assign new_n11055_ = ~new_n9291_ | ~new_n9768_;
  assign new_n11056_ = ~pi637 | ~new_n9214_;
  assign new_n11057_ = ~new_n9291_ | ~new_n9786_;
  assign new_n11058_ = ~pi638 | ~new_n9214_;
  assign new_n11059_ = ~new_n9291_ | ~new_n9804_;
  assign new_n11060_ = ~pi639 | ~new_n9214_;
  assign new_n11061_ = ~new_n9291_ | ~new_n9822_;
  assign new_n11062_ = ~pi640 | ~new_n9214_;
  assign new_n11063_ = ~new_n9291_ | ~new_n9840_;
  assign new_n11064_ = ~pi641 | ~new_n9214_;
  assign new_n11065_ = ~new_n9291_ | ~new_n9858_;
  assign new_n11066_ = ~pi642 | ~new_n9214_;
  assign new_n11067_ = ~new_n9291_ | ~new_n9876_;
  assign new_n11068_ = ~pi643 | ~new_n9214_;
  assign new_n11069_ = ~new_n9291_ | ~new_n9894_;
  assign new_n11070_ = ~pi644 | ~new_n9214_;
  assign new_n11071_ = ~new_n9291_ | ~new_n9912_;
  assign new_n11072_ = ~pi645 | ~new_n9214_;
  assign new_n11073_ = ~new_n9291_ | ~new_n9930_;
  assign new_n11074_ = ~pi646 | ~new_n9214_;
  assign new_n11075_ = ~new_n9291_ | ~new_n9948_;
  assign new_n11076_ = ~pi647 | ~new_n9214_;
  assign new_n11077_ = ~new_n9291_ | ~new_n9966_;
  assign new_n11078_ = ~pi648 | ~new_n9214_;
  assign new_n11079_ = ~new_n9291_ | ~new_n9986_;
  assign new_n11080_ = ~pi649 | ~new_n9214_;
  assign new_n11081_ = ~new_n9291_ | ~new_n9993_;
  assign new_n11082_ = ~pi650 | ~new_n9214_;
  assign new_n11083_ = ~new_n9291_ | ~new_n9995_;
  assign new_n11084_ = ~pi651 | ~new_n8736_;
  assign new_n11085_ = ~new_n9290_ | ~new_n8692_;
  assign new_n11086_ = ~pi652 | ~new_n8736_;
  assign new_n11087_ = ~new_n9290_ | ~new_n8693_;
  assign new_n11088_ = ~pi653 | ~new_n8736_;
  assign new_n11089_ = ~new_n9290_ | ~new_n8694_;
  assign new_n11090_ = ~pi654 | ~new_n8736_;
  assign new_n11091_ = ~new_n9290_ | ~new_n8695_;
  assign new_n11092_ = ~pi655 | ~new_n8736_;
  assign new_n11093_ = ~new_n9290_ | ~new_n8696_;
  assign new_n11094_ = ~pi656 | ~new_n8736_;
  assign new_n11095_ = ~new_n9290_ | ~new_n8697_;
  assign new_n11096_ = ~pi657 | ~new_n8736_;
  assign new_n11097_ = ~new_n9290_ | ~new_n8698_;
  assign new_n11098_ = ~pi658 | ~new_n8736_;
  assign new_n11099_ = ~new_n9290_ | ~new_n8699_;
  assign new_n11100_ = ~pi659 | ~new_n8736_;
  assign new_n11101_ = ~new_n9290_ | ~new_n8700_;
  assign new_n11102_ = ~pi660 | ~new_n8736_;
  assign new_n11103_ = ~new_n9290_ | ~new_n8701_;
  assign new_n11104_ = ~pi661 | ~new_n8736_;
  assign new_n11105_ = ~new_n9290_ | ~new_n8702_;
  assign new_n11106_ = ~pi662 | ~new_n8736_;
  assign new_n11107_ = ~new_n9290_ | ~new_n8703_;
  assign new_n11108_ = ~pi663 | ~new_n8736_;
  assign new_n11109_ = ~new_n9290_ | ~new_n8704_;
  assign new_n11110_ = ~pi664 | ~new_n8736_;
  assign new_n11111_ = ~new_n9290_ | ~new_n8705_;
  assign new_n11112_ = ~pi665 | ~new_n8736_;
  assign new_n11113_ = ~new_n9290_ | ~new_n8706_;
  assign new_n11114_ = ~pi666 | ~new_n8736_;
  assign new_n11115_ = ~new_n9290_ | ~new_n8707_;
  assign new_n11116_ = ~pi667 | ~new_n8736_;
  assign new_n11117_ = ~new_n9290_ | ~new_n8708_;
  assign new_n11118_ = ~pi668 | ~new_n8736_;
  assign new_n11119_ = ~new_n9290_ | ~new_n8709_;
  assign new_n11120_ = ~pi669 | ~new_n8736_;
  assign new_n11121_ = ~new_n9290_ | ~new_n8710_;
  assign new_n11122_ = ~pi670 | ~new_n8736_;
  assign new_n11123_ = ~new_n9290_ | ~new_n8711_;
  assign new_n11124_ = ~pi671 | ~new_n8736_;
  assign new_n11125_ = ~new_n9290_ | ~new_n8713_;
  assign new_n11126_ = ~pi672 | ~new_n8736_;
  assign new_n11127_ = ~new_n9290_ | ~new_n8715_;
  assign new_n11128_ = ~pi673 | ~new_n8736_;
  assign new_n11129_ = ~new_n9290_ | ~new_n8717_;
  assign new_n11130_ = ~pi674 | ~new_n8736_;
  assign new_n11131_ = ~new_n9290_ | ~new_n8719_;
  assign new_n11132_ = ~pi675 | ~new_n8736_;
  assign new_n11133_ = ~new_n9290_ | ~new_n8721_;
  assign new_n11134_ = ~pi676 | ~new_n8736_;
  assign new_n11135_ = ~new_n9290_ | ~new_n8723_;
  assign new_n11136_ = ~pi677 | ~new_n8736_;
  assign new_n11137_ = ~new_n9290_ | ~new_n8725_;
  assign new_n11138_ = ~pi678 | ~new_n8736_;
  assign new_n11139_ = ~new_n9290_ | ~new_n8727_;
  assign new_n11140_ = ~pi679 | ~new_n8736_;
  assign new_n11141_ = ~new_n9290_ | ~new_n8729_;
  assign new_n11142_ = ~pi680 | ~new_n8736_;
  assign new_n11143_ = ~new_n9290_ | ~new_n8732_;
  assign new_n11144_ = ~new_n10843_ | ~new_n8402_;
  assign new_n11145_ = ~new_n8761_ | ~po756;
  assign new_n11146_ = ~new_n11145_ | ~new_n11144_;
  assign new_n11147_ = ~pi703 | ~new_n8741_;
  assign new_n11148_ = ~po756 | ~new_n8454_;
  assign new_n11149_ = ~pi704 | ~new_n8741_;
  assign new_n11150_ = ~po756 | ~new_n8455_;
  assign new_n11151_ = ~pi705 | ~new_n8741_;
  assign new_n11152_ = ~po756 | ~new_n8445_;
  assign new_n11153_ = ~pi706 | ~new_n8741_;
  assign new_n11154_ = ~po756 | ~new_n8441_;
  assign new_n11155_ = ~pi707 | ~new_n8741_;
  assign new_n11156_ = ~po756 | ~new_n8437_;
  assign new_n11157_ = ~pi708 | ~new_n8741_;
  assign new_n11158_ = ~po756 | ~new_n8444_;
  assign new_n11159_ = ~pi709 | ~new_n8741_;
  assign new_n11160_ = ~po756 | ~new_n8448_;
  assign new_n11161_ = ~pi710 | ~new_n8741_;
  assign new_n11162_ = ~po756 | ~new_n8447_;
  assign new_n11163_ = ~pi711 | ~new_n8741_;
  assign new_n11164_ = ~po756 | ~new_n8461_;
  assign new_n11165_ = ~pi712 | ~new_n8741_;
  assign new_n11166_ = ~po756 | ~new_n8460_;
  assign new_n11167_ = ~pi713 | ~new_n8741_;
  assign new_n11168_ = ~po756 | ~new_n8439_;
  assign new_n11169_ = ~pi714 | ~new_n8741_;
  assign new_n11170_ = ~po756 | ~new_n8440_;
  assign new_n11171_ = ~pi715 | ~new_n8741_;
  assign new_n11172_ = ~po756 | ~new_n8449_;
  assign new_n11173_ = ~pi716 | ~new_n8741_;
  assign new_n11174_ = ~po756 | ~new_n8457_;
  assign new_n11175_ = ~pi717 | ~new_n8741_;
  assign new_n11176_ = ~po756 | ~new_n8456_;
  assign new_n11177_ = ~pi718 | ~new_n8741_;
  assign new_n11178_ = ~po756 | ~new_n8451_;
  assign new_n11179_ = ~pi719 | ~new_n8741_;
  assign new_n11180_ = ~po756 | ~new_n8450_;
  assign new_n11181_ = ~pi720 | ~new_n8741_;
  assign new_n11182_ = ~po756 | ~new_n8446_;
  assign new_n11183_ = ~pi721 | ~new_n8741_;
  assign new_n11184_ = ~po756 | ~new_n8459_;
  assign new_n11185_ = ~pi722 | ~new_n8741_;
  assign new_n11186_ = ~po756 | ~new_n8458_;
  assign new_n11187_ = ~pi723 | ~new_n8741_;
  assign new_n11188_ = ~po756 | ~new_n8453_;
  assign new_n11189_ = ~pi724 | ~new_n8741_;
  assign new_n11190_ = ~po756 | ~new_n8452_;
  assign new_n11191_ = ~pi725 | ~new_n8741_;
  assign new_n11192_ = ~po756 | ~new_n8438_;
  assign new_n11193_ = ~pi726 | ~new_n8741_;
  assign new_n11194_ = ~po756 | ~new_n8443_;
  assign new_n11195_ = ~pi727 | ~new_n8741_;
  assign new_n11196_ = ~po756 | ~new_n8442_;
  assign new_n11197_ = ~pi728 | ~new_n8741_;
  assign new_n11198_ = ~po756 | ~new_n8435_;
  assign new_n11199_ = ~pi729 | ~new_n8741_;
  assign new_n11200_ = ~po756 | ~new_n8434_;
  assign new_n11201_ = ~pi730 | ~new_n8741_;
  assign new_n11202_ = ~po756 | ~new_n8430_;
  assign new_n11203_ = ~pi731 | ~new_n8741_;
  assign new_n11204_ = ~po756 | ~new_n8431_;
  assign new_n11205_ = ~pi732 | ~new_n8741_;
  assign new_n11206_ = ~po756 | ~new_n8432_;
  assign new_n11207_ = ~pi733 | ~new_n8741_;
  assign new_n11208_ = ~po756 | ~new_n8436_;
  assign new_n11209_ = ~pi734 | ~new_n8741_;
  assign new_n11210_ = ~po756 | ~new_n8433_;
  assign new_n11211_ = ~new_n8757_ | ~new_n8691_;
  assign new_n11212_ = ~new_n10828_ | ~new_n9289_;
  assign new_n11213_ = ~new_n9138_;
  assign new_n11214_ = ~new_n27167_ | ~new_n11213_;
  assign new_n11215_ = ~new_n9138_ | ~new_n9245_;
  assign new_n11216_ = ~new_n9278_ | ~new_n8430_;
  assign new_n11217_ = ~new_n8726_ | ~new_n9917_;
  assign new_n11218_ = ~new_n11217_ | ~new_n11216_;
  assign new_n11219_ = ~new_n9277_ | ~new_n8431_;
  assign new_n11220_ = ~new_n8728_ | ~new_n9935_;
  assign new_n11221_ = ~new_n11220_ | ~new_n11219_;
  assign new_n11222_ = ~new_n9250_ | ~new_n8433_;
  assign new_n11223_ = ~new_n8734_ | ~new_n9991_;
  assign new_n11224_ = ~new_n11223_ | ~new_n11222_;
  assign new_n11225_ = ~new_n9286_ | ~new_n8432_;
  assign new_n11226_ = ~new_n8731_ | ~new_n9953_;
  assign new_n11227_ = ~new_n11226_ | ~new_n11225_;
  assign new_n11228_ = ~new_n9284_ | ~new_n8452_;
  assign new_n11229_ = ~new_n8714_ | ~new_n9809_;
  assign new_n11230_ = ~new_n11229_ | ~new_n11228_;
  assign new_n11231_ = ~new_n9285_ | ~new_n8453_;
  assign new_n11232_ = ~new_n8712_ | ~new_n9791_;
  assign new_n11233_ = ~new_n11232_ | ~new_n11231_;
  assign new_n11234_ = ~new_n10881_ | ~new_n9485_;
  assign new_n11235_ = ~new_n8776_ | ~new_n8441_;
  assign new_n11236_ = ~new_n11235_ | ~new_n11234_;
  assign new_n11237_ = ~new_n10937_ | ~new_n9629_;
  assign new_n11238_ = ~new_n8800_ | ~new_n8440_;
  assign new_n11239_ = ~new_n11238_ | ~new_n11237_;
  assign new_n11240_ = ~new_n10930_ | ~new_n9611_;
  assign new_n11241_ = ~new_n8797_ | ~new_n8439_;
  assign new_n11242_ = ~new_n11241_ | ~new_n11240_;
  assign new_n11243_ = ~new_n10888_ | ~new_n9503_;
  assign new_n11244_ = ~new_n8779_ | ~new_n8437_;
  assign new_n11245_ = ~new_n11244_ | ~new_n11243_;
  assign new_n11246_ = ~new_n9283_ | ~new_n8438_;
  assign new_n11247_ = ~new_n8716_ | ~new_n9827_;
  assign new_n11248_ = ~new_n11247_ | ~new_n11246_;
  assign new_n11249_ = ~new_n10979_ | ~new_n9737_;
  assign new_n11250_ = ~new_n8818_ | ~new_n8446_;
  assign new_n11251_ = ~new_n11250_ | ~new_n11249_;
  assign new_n11252_ = ~new_n10972_ | ~new_n9719_;
  assign new_n11253_ = ~new_n8815_ | ~new_n8450_;
  assign new_n11254_ = ~new_n11253_ | ~new_n11252_;
  assign new_n11255_ = ~new_n10965_ | ~new_n9701_;
  assign new_n11256_ = ~new_n8812_ | ~new_n8451_;
  assign new_n11257_ = ~new_n11256_ | ~new_n11255_;
  assign new_n11258_ = ~new_n10944_ | ~new_n9647_;
  assign new_n11259_ = ~new_n8803_ | ~new_n8449_;
  assign new_n11260_ = ~new_n11259_ | ~new_n11258_;
  assign new_n11261_ = ~new_n10902_ | ~new_n9539_;
  assign new_n11262_ = ~new_n8785_ | ~new_n8448_;
  assign new_n11263_ = ~new_n11262_ | ~new_n11261_;
  assign new_n11264_ = ~new_n10909_ | ~new_n9557_;
  assign new_n11265_ = ~new_n8788_ | ~new_n8447_;
  assign new_n11266_ = ~new_n11265_ | ~new_n11264_;
  assign new_n11267_ = ~new_n10874_ | ~new_n9460_;
  assign new_n11268_ = ~new_n8773_ | ~new_n8445_;
  assign new_n11269_ = ~new_n11268_ | ~new_n11267_;
  assign new_n11270_ = ~new_n10895_ | ~new_n9521_;
  assign new_n11271_ = ~new_n8782_ | ~new_n8444_;
  assign new_n11272_ = ~new_n11271_ | ~new_n11270_;
  assign new_n11273_ = ~new_n10986_ | ~new_n9755_;
  assign new_n11274_ = ~new_n8821_ | ~new_n8459_;
  assign new_n11275_ = ~new_n11274_ | ~new_n11273_;
  assign new_n11276_ = ~new_n10951_ | ~new_n9665_;
  assign new_n11277_ = ~new_n8806_ | ~new_n8457_;
  assign new_n11278_ = ~new_n11277_ | ~new_n11276_;
  assign new_n11279_ = ~new_n10958_ | ~new_n9683_;
  assign new_n11280_ = ~new_n8809_ | ~new_n8456_;
  assign new_n11281_ = ~new_n11280_ | ~new_n11279_;
  assign new_n11282_ = ~new_n10867_ | ~new_n9441_;
  assign new_n11283_ = ~new_n8770_ | ~new_n8455_;
  assign new_n11284_ = ~new_n11283_ | ~new_n11282_;
  assign new_n11285_ = ~new_n10851_ | ~new_n9465_;
  assign new_n11286_ = ~new_n8765_ | ~new_n8454_;
  assign new_n11287_ = ~new_n11286_ | ~new_n11285_;
  assign new_n11288_ = ~new_n10916_ | ~new_n9575_;
  assign new_n11289_ = ~new_n8791_ | ~new_n8461_;
  assign new_n11290_ = ~new_n11289_ | ~new_n11288_;
  assign new_n11291_ = ~new_n10923_ | ~new_n9593_;
  assign new_n11292_ = ~new_n8794_ | ~new_n8460_;
  assign new_n11293_ = ~new_n11292_ | ~new_n11291_;
  assign new_n11294_ = ~new_n10991_ | ~new_n9773_;
  assign new_n11295_ = ~new_n8823_ | ~new_n8458_;
  assign new_n11296_ = ~new_n11295_ | ~new_n11294_;
  assign new_n11297_ = ~new_n9279_ | ~new_n8434_;
  assign new_n11298_ = ~new_n8724_ | ~new_n9899_;
  assign new_n11299_ = ~new_n11298_ | ~new_n11297_;
  assign new_n11300_ = ~new_n9280_ | ~new_n8435_;
  assign new_n11301_ = ~new_n8722_ | ~new_n9881_;
  assign new_n11302_ = ~new_n11301_ | ~new_n11300_;
  assign new_n11303_ = ~new_n9282_ | ~new_n8443_;
  assign new_n11304_ = ~new_n8718_ | ~new_n9845_;
  assign new_n11305_ = ~new_n11304_ | ~new_n11303_;
  assign new_n11306_ = ~new_n9281_ | ~new_n8442_;
  assign new_n11307_ = ~new_n8720_ | ~new_n9863_;
  assign new_n11308_ = ~new_n11307_ | ~new_n11306_;
  assign new_n11309_ = ~new_n9251_ | ~new_n8436_;
  assign new_n11310_ = ~new_n8733_ | ~new_n9971_;
  assign new_n11311_ = ~new_n11310_ | ~new_n11309_;
  assign new_n11312_ = ~new_n10356_ | ~new_n10828_;
  assign new_n11313_ = ~new_n8757_ | ~new_n9246_;
  assign new_n11314_ = ~new_n11313_ | ~new_n11312_;
  assign new_n11315_ = ~new_n10825_ | ~new_n11215_ | ~new_n11214_;
  assign new_n11316_ = ~new_n8756_ | ~new_n10834_ | ~new_n11314_;
  assign new_n11317_ = ~new_n9259_ | ~new_n9247_;
  assign new_n11318_ = ~new_n24882_ | ~new_n9269_;
  assign new_n11319_ = ~new_n10818_ | ~new_n8746_;
  assign new_n11320_ = ~new_n8758_ | ~new_n8753_;
  assign new_n11321_ = ~new_n10828_ | ~new_n10825_;
  assign new_n11322_ = ~new_n8756_ | ~new_n8766_ | ~new_n10834_;
  assign new_n11323_ = ~new_n8460_ | ~new_n27860_;
  assign new_n11324_ = ~new_n8460_ | ~new_n9249_;
  assign new_n11325_ = ~new_n8461_ | ~new_n27860_;
  assign new_n11326_ = ~new_n8461_ | ~new_n9249_;
  assign new_n11327_ = ~new_n8447_ | ~new_n27860_;
  assign new_n11328_ = ~new_n8447_ | ~new_n9249_;
  assign new_n11329_ = ~new_n8448_ | ~new_n27860_;
  assign new_n11330_ = ~new_n8448_ | ~new_n9249_;
  assign new_n11331_ = ~new_n8444_ | ~new_n27860_;
  assign new_n11332_ = ~new_n8444_ | ~new_n9249_;
  assign new_n11333_ = ~new_n8437_ | ~new_n27860_;
  assign new_n11334_ = ~new_n8437_ | ~new_n9249_;
  assign new_n11335_ = ~new_n26199_ | ~new_n27860_;
  assign new_n11336_ = ~new_n8433_ | ~new_n9249_;
  assign new_n11337_ = ~new_n26197_ | ~new_n27860_;
  assign new_n11338_ = ~new_n8436_ | ~new_n9249_;
  assign new_n11339_ = ~new_n8441_ | ~new_n27860_;
  assign new_n11340_ = ~new_n8441_ | ~new_n9249_;
  assign new_n11341_ = ~new_n8432_ | ~new_n27860_;
  assign new_n11342_ = ~new_n8432_ | ~new_n9249_;
  assign new_n11343_ = ~new_n8431_ | ~new_n27860_;
  assign new_n11344_ = ~new_n8431_ | ~new_n9249_;
  assign new_n11345_ = ~new_n8430_ | ~new_n27860_;
  assign new_n11346_ = ~new_n8430_ | ~new_n9249_;
  assign new_n11347_ = ~new_n8434_ | ~new_n27860_;
  assign new_n11348_ = ~new_n8434_ | ~new_n9249_;
  assign new_n11349_ = ~new_n8435_ | ~new_n27860_;
  assign new_n11350_ = ~new_n8435_ | ~new_n9249_;
  assign new_n11351_ = ~new_n8442_ | ~new_n27860_;
  assign new_n11352_ = ~new_n8442_ | ~new_n9249_;
  assign new_n11353_ = ~new_n8443_ | ~new_n27860_;
  assign new_n11354_ = ~new_n8443_ | ~new_n9249_;
  assign new_n11355_ = ~new_n8438_ | ~new_n27860_;
  assign new_n11356_ = ~new_n8438_ | ~new_n9249_;
  assign new_n11357_ = ~new_n8452_ | ~new_n27860_;
  assign new_n11358_ = ~new_n8452_ | ~new_n9249_;
  assign new_n11359_ = ~new_n8453_ | ~new_n27860_;
  assign new_n11360_ = ~new_n8453_ | ~new_n9249_;
  assign new_n11361_ = ~new_n8445_ | ~new_n27860_;
  assign new_n11362_ = ~new_n8445_ | ~new_n9249_;
  assign new_n11363_ = ~new_n8458_ | ~new_n27860_;
  assign new_n11364_ = ~new_n8458_ | ~new_n9249_;
  assign new_n11365_ = ~new_n8459_ | ~new_n27860_;
  assign new_n11366_ = ~new_n8459_ | ~new_n9249_;
  assign new_n11367_ = ~new_n8446_ | ~new_n27860_;
  assign new_n11368_ = ~new_n8446_ | ~new_n9249_;
  assign new_n11369_ = ~new_n8450_ | ~new_n27860_;
  assign new_n11370_ = ~new_n8450_ | ~new_n9249_;
  assign new_n11371_ = ~new_n8451_ | ~new_n27860_;
  assign new_n11372_ = ~new_n8451_ | ~new_n9249_;
  assign new_n11373_ = ~new_n8456_ | ~new_n27860_;
  assign new_n11374_ = ~new_n8456_ | ~new_n9249_;
  assign new_n11375_ = ~new_n8457_ | ~new_n27860_;
  assign new_n11376_ = ~new_n8457_ | ~new_n9249_;
  assign new_n11377_ = ~new_n8449_ | ~new_n27860_;
  assign new_n11378_ = ~new_n8449_ | ~new_n9249_;
  assign new_n11379_ = ~new_n8440_ | ~new_n27860_;
  assign new_n11380_ = ~new_n8440_ | ~new_n9249_;
  assign new_n11381_ = ~new_n8439_ | ~new_n27860_;
  assign new_n11382_ = ~new_n8439_ | ~new_n9249_;
  assign new_n11383_ = ~new_n8455_ | ~new_n27860_;
  assign new_n11384_ = ~new_n8455_ | ~new_n9249_;
  assign new_n11385_ = ~new_n8454_ | ~new_n27860_;
  assign new_n11386_ = ~new_n8454_ | ~new_n9249_;
  assign new_n11387_ = ~new_n10846_ | ~pi628;
  assign new_n11388_ = ~new_n8762_ | ~pi660;
  assign new_n11389_ = ~new_n10846_ | ~pi627;
  assign new_n11390_ = ~new_n8762_ | ~pi659;
  assign new_n11391_ = ~new_n10846_ | ~pi626;
  assign new_n11392_ = ~new_n8762_ | ~pi658;
  assign new_n11393_ = ~new_n10846_ | ~pi625;
  assign new_n11394_ = ~new_n8762_ | ~pi657;
  assign new_n11395_ = ~new_n10846_ | ~pi624;
  assign new_n11396_ = ~new_n8762_ | ~pi656;
  assign new_n11397_ = ~new_n10846_ | ~pi623;
  assign new_n11398_ = ~new_n8762_ | ~pi655;
  assign new_n11399_ = ~new_n10846_ | ~pi622;
  assign new_n11400_ = ~new_n8762_ | ~pi654;
  assign new_n11401_ = ~new_n10846_ | ~pi621;
  assign new_n11402_ = ~new_n8762_ | ~pi653;
  assign new_n11403_ = ~new_n10846_ | ~pi638;
  assign new_n11404_ = ~new_n8762_ | ~pi670;
  assign new_n11405_ = ~new_n10846_ | ~pi637;
  assign new_n11406_ = ~new_n8762_ | ~pi669;
  assign new_n11407_ = ~new_n10846_ | ~pi636;
  assign new_n11408_ = ~new_n8762_ | ~pi668;
  assign new_n11409_ = ~new_n10846_ | ~pi635;
  assign new_n11410_ = ~new_n8762_ | ~pi667;
  assign new_n11411_ = ~new_n10846_ | ~pi634;
  assign new_n11412_ = ~new_n8762_ | ~pi666;
  assign new_n11413_ = ~new_n10846_ | ~pi633;
  assign new_n11414_ = ~new_n8762_ | ~pi665;
  assign new_n11415_ = ~new_n10846_ | ~pi632;
  assign new_n11416_ = ~new_n8762_ | ~pi664;
  assign new_n11417_ = ~new_n10846_ | ~pi631;
  assign new_n11418_ = ~new_n8762_ | ~pi663;
  assign new_n11419_ = ~new_n10846_ | ~pi630;
  assign new_n11420_ = ~new_n8762_ | ~pi662;
  assign new_n11421_ = ~new_n10846_ | ~pi629;
  assign new_n11422_ = ~new_n8762_ | ~pi661;
  assign new_n11423_ = ~new_n10846_ | ~pi620;
  assign new_n11424_ = ~new_n8762_ | ~pi652;
  assign new_n11425_ = ~new_n10846_ | ~pi619;
  assign new_n11426_ = ~new_n8762_ | ~pi651;
  assign new_n11427_ = ~new_n30544_ | ~new_n11429_;
  assign new_n11428_ = ~new_n30416_ | ~new_n30417_;
  assign new_n11429_ = ~new_n11430_ | ~new_n11431_;
  assign new_n11430_ = ~new_n9283_ | ~new_n30341_;
  assign new_n11431_ = ~new_n8438_ | ~new_n30340_;
  assign new_n11432_ = ~new_n9283_ | ~new_n30341_;
  assign new_n11433_ = ~new_n8438_ | ~new_n30340_;
  assign new_n11434_ = ~new_n30548_ | ~new_n11436_;
  assign new_n11435_ = ~new_n30414_ | ~new_n30415_;
  assign new_n11436_ = ~new_n11437_ | ~new_n11438_;
  assign new_n11437_ = ~new_n9282_ | ~new_n30343_;
  assign new_n11438_ = ~new_n8443_ | ~new_n30342_;
  assign new_n11439_ = ~new_n9282_ | ~new_n30343_;
  assign new_n11440_ = ~new_n8443_ | ~new_n30342_;
  assign new_n11441_ = ~new_n30552_ | ~new_n11443_;
  assign new_n11442_ = ~new_n30616_ | ~new_n30413_;
  assign new_n11443_ = ~new_n11444_ | ~new_n11445_;
  assign new_n11444_ = ~new_n9281_ | ~new_n30311_;
  assign new_n11445_ = ~new_n8442_ | ~new_n30310_;
  assign new_n11446_ = new_n11634_ & new_n11630_;
  assign new_n11447_ = new_n11642_ & new_n11640_;
  assign new_n11448_ = new_n11447_ & new_n11644_;
  assign new_n11449_ = new_n11652_ & new_n11648_;
  assign new_n11450_ = new_n11449_ & new_n11655_;
  assign new_n11451_ = new_n11803_ & new_n11802_;
  assign new_n11452_ = ~new_n11568_ | ~new_n11763_;
  assign new_n11453_ = ~new_n11615_ | ~new_n11731_;
  assign new_n11454_ = ~pi221;
  assign new_n11455_ = ~pi466;
  assign new_n11456_ = ~pi465;
  assign new_n11457_ = ~pi219;
  assign new_n11458_ = ~pi220;
  assign new_n11459_ = ~pi464;
  assign new_n11460_ = ~pi218;
  assign new_n11461_ = ~new_n11743_ | ~new_n11644_;
  assign new_n11462_ = ~pi217;
  assign new_n11463_ = ~pi458;
  assign new_n11464_ = ~pi214;
  assign new_n11465_ = ~pi462;
  assign new_n11466_ = ~pi460;
  assign new_n11467_ = ~pi461;
  assign new_n11468_ = ~pi215;
  assign new_n11469_ = ~pi216;
  assign new_n11470_ = ~pi463;
  assign new_n11471_ = ~pi467;
  assign new_n11472_ = ~pi222;
  assign new_n11473_ = ~pi225;
  assign new_n11474_ = ~pi470;
  assign new_n11475_ = ~pi469;
  assign new_n11476_ = ~pi468;
  assign new_n11477_ = ~pi224;
  assign new_n11478_ = ~pi223;
  assign new_n11479_ = ~pi222 | ~new_n11471_;
  assign new_n11480_ = ~pi471;
  assign new_n11481_ = ~pi226;
  assign new_n11482_ = ~pi472;
  assign new_n11483_ = ~pi227;
  assign new_n11484_ = ~pi473;
  assign new_n11485_ = ~pi228;
  assign new_n11486_ = ~pi474;
  assign new_n11487_ = ~pi229;
  assign new_n11488_ = ~pi475;
  assign new_n11489_ = ~pi230;
  assign new_n11490_ = ~pi476;
  assign new_n11491_ = ~pi231;
  assign new_n11492_ = ~pi477;
  assign new_n11493_ = ~pi232;
  assign new_n11494_ = ~pi478;
  assign new_n11495_ = ~pi233;
  assign new_n11496_ = ~pi479;
  assign new_n11497_ = ~pi234;
  assign new_n11498_ = ~pi480;
  assign new_n11499_ = ~pi235;
  assign new_n11500_ = ~pi481;
  assign new_n11501_ = ~pi236;
  assign new_n11502_ = ~pi482;
  assign new_n11503_ = ~pi237;
  assign new_n11504_ = ~pi483;
  assign new_n11505_ = ~pi238;
  assign new_n11506_ = ~pi484;
  assign new_n11507_ = ~pi239;
  assign new_n11508_ = ~pi485;
  assign new_n11509_ = ~pi240;
  assign new_n11510_ = ~pi486;
  assign new_n11511_ = ~pi241;
  assign new_n11512_ = ~pi487;
  assign new_n11513_ = ~pi242;
  assign new_n11514_ = ~pi243;
  assign new_n11515_ = ~pi488;
  assign new_n11516_ = ~new_n11748_ | ~new_n11656_;
  assign new_n11517_ = ~new_n11745_ | ~new_n11653_;
  assign new_n11518_ = ~pi213;
  assign new_n11519_ = ~new_n11768_ | ~new_n11767_;
  assign new_n11520_ = ~new_n11773_ | ~new_n11772_;
  assign new_n11521_ = ~new_n11778_ | ~new_n11777_;
  assign new_n11522_ = ~new_n11783_ | ~new_n11782_;
  assign new_n11523_ = ~new_n11788_ | ~new_n11787_;
  assign new_n11524_ = ~new_n11793_ | ~new_n11792_;
  assign new_n11525_ = ~new_n11798_ | ~new_n11797_;
  assign new_n11526_ = ~new_n11810_ | ~new_n11809_;
  assign new_n11527_ = ~new_n11815_ | ~new_n11814_;
  assign new_n11528_ = ~new_n11820_ | ~new_n11819_;
  assign new_n11529_ = ~new_n11825_ | ~new_n11824_;
  assign new_n11530_ = ~new_n11830_ | ~new_n11829_;
  assign new_n11531_ = ~new_n11835_ | ~new_n11834_;
  assign new_n11532_ = ~new_n11840_ | ~new_n11839_;
  assign new_n11533_ = ~new_n11845_ | ~new_n11844_;
  assign new_n11534_ = ~new_n11850_ | ~new_n11849_;
  assign new_n11535_ = ~new_n11855_ | ~new_n11854_;
  assign new_n11536_ = ~new_n11860_ | ~new_n11859_;
  assign new_n11537_ = ~new_n11865_ | ~new_n11864_;
  assign new_n11538_ = ~new_n11870_ | ~new_n11869_;
  assign new_n11539_ = ~new_n11875_ | ~new_n11874_;
  assign new_n11540_ = ~new_n11880_ | ~new_n11879_;
  assign new_n11541_ = ~new_n11885_ | ~new_n11884_;
  assign new_n11542_ = ~new_n11890_ | ~new_n11889_;
  assign new_n11543_ = ~new_n11895_ | ~new_n11894_;
  assign new_n11544_ = ~new_n11900_ | ~new_n11899_;
  assign new_n11545_ = ~new_n11905_ | ~new_n11904_;
  assign new_n11546_ = ~new_n11910_ | ~new_n11909_;
  assign new_n11547_ = ~new_n11915_ | ~new_n11914_;
  assign new_n11548_ = ~new_n11920_ | ~new_n11919_;
  assign new_n11549_ = pi218 & new_n11470_;
  assign new_n11550_ = new_n11645_ & new_n11643_;
  assign new_n11551_ = new_n11637_ & new_n11446_;
  assign new_n11552_ = new_n11739_ & new_n11637_;
  assign new_n11553_ = new_n11738_ & new_n11638_;
  assign new_n11554_ = new_n11646_ & new_n11448_;
  assign new_n11555_ = new_n11742_ & new_n11647_;
  assign new_n11556_ = ~new_n11765_ | ~new_n11764_;
  assign new_n11557_ = ~new_n11770_ | ~new_n11769_;
  assign new_n11558_ = new_n11740_ & new_n11643_;
  assign new_n11559_ = ~new_n11775_ | ~new_n11774_;
  assign new_n11560_ = ~new_n11780_ | ~new_n11779_;
  assign new_n11561_ = ~new_n11785_ | ~new_n11784_;
  assign new_n11562_ = ~new_n11790_ | ~new_n11789_;
  assign new_n11563_ = ~new_n11795_ | ~new_n11794_;
  assign new_n11564_ = new_n11450_ & new_n11658_;
  assign new_n11565_ = new_n11751_ & new_n11659_;
  assign new_n11566_ = new_n11727_ & new_n11451_ & new_n11730_;
  assign new_n11567_ = new_n11729_ & new_n11801_;
  assign new_n11568_ = new_n11601_ & new_n11733_;
  assign new_n11569_ = ~new_n11807_ | ~new_n11806_;
  assign new_n11570_ = ~new_n11812_ | ~new_n11811_;
  assign new_n11571_ = ~new_n11817_ | ~new_n11816_;
  assign new_n11572_ = ~new_n11822_ | ~new_n11821_;
  assign new_n11573_ = ~new_n11827_ | ~new_n11826_;
  assign new_n11574_ = ~new_n11832_ | ~new_n11831_;
  assign new_n11575_ = ~new_n11837_ | ~new_n11836_;
  assign new_n11576_ = ~new_n11842_ | ~new_n11841_;
  assign new_n11577_ = ~new_n11847_ | ~new_n11846_;
  assign new_n11578_ = ~new_n11852_ | ~new_n11851_;
  assign new_n11579_ = ~new_n11857_ | ~new_n11856_;
  assign new_n11580_ = ~new_n11862_ | ~new_n11861_;
  assign new_n11581_ = ~new_n11867_ | ~new_n11866_;
  assign new_n11582_ = ~new_n11872_ | ~new_n11871_;
  assign new_n11583_ = ~new_n11877_ | ~new_n11876_;
  assign new_n11584_ = ~new_n11882_ | ~new_n11881_;
  assign new_n11585_ = ~new_n11887_ | ~new_n11886_;
  assign new_n11586_ = ~new_n11892_ | ~new_n11891_;
  assign new_n11587_ = ~new_n11897_ | ~new_n11896_;
  assign new_n11588_ = ~new_n11902_ | ~new_n11901_;
  assign new_n11589_ = ~new_n11907_ | ~new_n11906_;
  assign new_n11590_ = ~new_n11912_ | ~new_n11911_;
  assign new_n11591_ = ~new_n11917_ | ~new_n11916_;
  assign new_n11592_ = ~new_n11555_ | ~new_n11761_;
  assign new_n11593_ = ~new_n11759_ | ~new_n11461_;
  assign new_n11594_ = ~new_n11558_ | ~new_n11757_;
  assign new_n11595_ = ~new_n11755_ | ~new_n11641_;
  assign new_n11596_ = ~new_n11553_ | ~new_n11737_;
  assign new_n11597_ = ~new_n11736_ | ~new_n11734_;
  assign new_n11598_ = ~new_n11632_ | ~new_n11631_;
  assign new_n11599_ = ~pi489;
  assign new_n11600_ = ~pi244;
  assign new_n11601_ = new_n11805_ & new_n11804_;
  assign new_n11602_ = ~new_n11727_ | ~new_n11726_;
  assign new_n11603_ = ~new_n11732_ | ~new_n11628_ | ~new_n11626_;
  assign new_n11604_ = ~new_n11723_ | ~new_n11722_;
  assign new_n11605_ = ~new_n11719_ | ~new_n11718_;
  assign new_n11606_ = ~new_n11715_ | ~new_n11714_;
  assign new_n11607_ = ~new_n11711_ | ~new_n11710_;
  assign new_n11608_ = ~new_n11707_ | ~new_n11706_;
  assign new_n11609_ = ~new_n11703_ | ~new_n11702_;
  assign new_n11610_ = ~new_n11699_ | ~new_n11698_;
  assign new_n11611_ = ~new_n11695_ | ~new_n11694_;
  assign new_n11612_ = ~new_n11691_ | ~new_n11690_;
  assign new_n11613_ = ~new_n11687_ | ~new_n11686_;
  assign new_n11614_ = ~pi459;
  assign new_n11615_ = ~pi458 | ~new_n11518_;
  assign new_n11616_ = ~new_n11683_ | ~new_n11682_;
  assign new_n11617_ = ~new_n11679_ | ~new_n11678_;
  assign new_n11618_ = ~new_n11675_ | ~new_n11674_;
  assign new_n11619_ = ~new_n11671_ | ~new_n11670_;
  assign new_n11620_ = ~new_n11667_ | ~new_n11666_;
  assign new_n11621_ = ~new_n11663_ | ~new_n11662_;
  assign new_n11622_ = ~new_n11565_ | ~new_n11750_;
  assign new_n11623_ = ~new_n11749_ | ~new_n11747_;
  assign new_n11624_ = ~new_n11746_ | ~new_n11744_;
  assign new_n11625_ = ~new_n11479_ | ~new_n11649_;
  assign new_n11626_ = ~new_n11615_ | ~new_n11614_;
  assign new_n11627_ = ~new_n11615_;
  assign new_n11628_ = ~pi214 | ~new_n11615_;
  assign new_n11629_ = ~new_n11603_;
  assign new_n11630_ = ~pi460 | ~new_n11468_;
  assign new_n11631_ = ~new_n11630_ | ~new_n11752_;
  assign new_n11632_ = ~pi215 | ~new_n11466_;
  assign new_n11633_ = ~new_n11598_;
  assign new_n11634_ = ~pi461 | ~new_n11469_;
  assign new_n11635_ = ~pi216 | ~new_n11467_;
  assign new_n11636_ = ~new_n11597_;
  assign new_n11637_ = ~pi462 | ~new_n11462_;
  assign new_n11638_ = ~pi217 | ~new_n11465_;
  assign new_n11639_ = ~new_n11596_;
  assign new_n11640_ = ~pi463 | ~new_n11460_;
  assign new_n11641_ = ~pi218 | ~new_n11470_;
  assign new_n11642_ = ~pi464 | ~new_n11457_;
  assign new_n11643_ = ~pi219 | ~new_n11459_;
  assign new_n11644_ = ~pi465 | ~new_n11458_;
  assign new_n11645_ = ~pi220 | ~new_n11456_;
  assign new_n11646_ = ~pi466 | ~new_n11454_;
  assign new_n11647_ = ~pi221 | ~new_n11455_;
  assign new_n11648_ = ~pi467 | ~new_n11472_;
  assign new_n11649_ = ~new_n11648_ | ~new_n11592_;
  assign new_n11650_ = ~new_n11479_;
  assign new_n11651_ = ~new_n11625_;
  assign new_n11652_ = ~pi468 | ~new_n11478_;
  assign new_n11653_ = ~pi223 | ~new_n11476_;
  assign new_n11654_ = ~new_n11624_;
  assign new_n11655_ = ~pi469 | ~new_n11477_;
  assign new_n11656_ = ~pi224 | ~new_n11475_;
  assign new_n11657_ = ~new_n11623_;
  assign new_n11658_ = ~pi470 | ~new_n11473_;
  assign new_n11659_ = ~pi225 | ~new_n11474_;
  assign new_n11660_ = ~new_n11622_;
  assign new_n11661_ = ~pi471 | ~new_n11481_;
  assign new_n11662_ = ~new_n11661_ | ~new_n11622_;
  assign new_n11663_ = ~pi226 | ~new_n11480_;
  assign new_n11664_ = ~new_n11621_;
  assign new_n11665_ = ~pi472 | ~new_n11483_;
  assign new_n11666_ = ~new_n11665_ | ~new_n11621_;
  assign new_n11667_ = ~pi227 | ~new_n11482_;
  assign new_n11668_ = ~new_n11620_;
  assign new_n11669_ = ~pi473 | ~new_n11485_;
  assign new_n11670_ = ~new_n11669_ | ~new_n11620_;
  assign new_n11671_ = ~pi228 | ~new_n11484_;
  assign new_n11672_ = ~new_n11619_;
  assign new_n11673_ = ~pi474 | ~new_n11487_;
  assign new_n11674_ = ~new_n11673_ | ~new_n11619_;
  assign new_n11675_ = ~pi229 | ~new_n11486_;
  assign new_n11676_ = ~new_n11618_;
  assign new_n11677_ = ~pi475 | ~new_n11489_;
  assign new_n11678_ = ~new_n11677_ | ~new_n11618_;
  assign new_n11679_ = ~pi230 | ~new_n11488_;
  assign new_n11680_ = ~new_n11617_;
  assign new_n11681_ = ~pi476 | ~new_n11491_;
  assign new_n11682_ = ~new_n11681_ | ~new_n11617_;
  assign new_n11683_ = ~pi231 | ~new_n11490_;
  assign new_n11684_ = ~new_n11616_;
  assign new_n11685_ = ~pi477 | ~new_n11493_;
  assign new_n11686_ = ~new_n11685_ | ~new_n11616_;
  assign new_n11687_ = ~pi232 | ~new_n11492_;
  assign new_n11688_ = ~new_n11613_;
  assign new_n11689_ = ~pi478 | ~new_n11495_;
  assign new_n11690_ = ~new_n11689_ | ~new_n11613_;
  assign new_n11691_ = ~pi233 | ~new_n11494_;
  assign new_n11692_ = ~new_n11612_;
  assign new_n11693_ = ~pi479 | ~new_n11497_;
  assign new_n11694_ = ~new_n11693_ | ~new_n11612_;
  assign new_n11695_ = ~pi234 | ~new_n11496_;
  assign new_n11696_ = ~new_n11611_;
  assign new_n11697_ = ~pi480 | ~new_n11499_;
  assign new_n11698_ = ~new_n11697_ | ~new_n11611_;
  assign new_n11699_ = ~pi235 | ~new_n11498_;
  assign new_n11700_ = ~new_n11610_;
  assign new_n11701_ = ~pi481 | ~new_n11501_;
  assign new_n11702_ = ~new_n11701_ | ~new_n11610_;
  assign new_n11703_ = ~pi236 | ~new_n11500_;
  assign new_n11704_ = ~new_n11609_;
  assign new_n11705_ = ~pi482 | ~new_n11503_;
  assign new_n11706_ = ~new_n11705_ | ~new_n11609_;
  assign new_n11707_ = ~pi237 | ~new_n11502_;
  assign new_n11708_ = ~new_n11608_;
  assign new_n11709_ = ~pi483 | ~new_n11505_;
  assign new_n11710_ = ~new_n11709_ | ~new_n11608_;
  assign new_n11711_ = ~pi238 | ~new_n11504_;
  assign new_n11712_ = ~new_n11607_;
  assign new_n11713_ = ~pi484 | ~new_n11507_;
  assign new_n11714_ = ~new_n11713_ | ~new_n11607_;
  assign new_n11715_ = ~pi239 | ~new_n11506_;
  assign new_n11716_ = ~new_n11606_;
  assign new_n11717_ = ~pi485 | ~new_n11509_;
  assign new_n11718_ = ~new_n11717_ | ~new_n11606_;
  assign new_n11719_ = ~pi240 | ~new_n11508_;
  assign new_n11720_ = ~new_n11605_;
  assign new_n11721_ = ~pi486 | ~new_n11511_;
  assign new_n11722_ = ~new_n11721_ | ~new_n11605_;
  assign new_n11723_ = ~pi241 | ~new_n11510_;
  assign new_n11724_ = ~new_n11604_;
  assign new_n11725_ = ~pi487 | ~new_n11513_;
  assign new_n11726_ = ~new_n11725_ | ~new_n11604_;
  assign new_n11727_ = ~pi242 | ~new_n11512_;
  assign new_n11728_ = ~new_n11602_;
  assign new_n11729_ = ~pi488 | ~new_n11514_;
  assign new_n11730_ = ~pi243 | ~new_n11515_;
  assign new_n11731_ = ~pi213 | ~new_n11463_;
  assign new_n11732_ = ~pi214 | ~new_n11614_;
  assign new_n11733_ = ~new_n11726_ | ~new_n11566_;
  assign new_n11734_ = ~new_n11446_ | ~new_n11603_;
  assign new_n11735_ = ~new_n11635_ | ~new_n11632_;
  assign new_n11736_ = ~new_n11735_ | ~new_n11739_;
  assign new_n11737_ = ~new_n11551_ | ~new_n11603_;
  assign new_n11738_ = ~new_n11552_ | ~new_n11735_;
  assign new_n11739_ = ~pi461 | ~new_n11469_;
  assign new_n11740_ = ~new_n11549_ | ~new_n11642_;
  assign new_n11741_ = ~new_n11461_;
  assign new_n11742_ = ~new_n11741_ | ~new_n11646_;
  assign new_n11743_ = ~new_n11550_ | ~new_n11740_;
  assign new_n11744_ = ~new_n11449_ | ~new_n11592_;
  assign new_n11745_ = ~new_n11650_ | ~new_n11652_;
  assign new_n11746_ = ~new_n11517_;
  assign new_n11747_ = ~new_n11450_ | ~new_n11592_;
  assign new_n11748_ = ~new_n11517_ | ~new_n11655_;
  assign new_n11749_ = ~new_n11516_;
  assign new_n11750_ = ~new_n11564_ | ~new_n11592_;
  assign new_n11751_ = ~new_n11516_ | ~new_n11658_;
  assign new_n11752_ = ~new_n11754_ | ~new_n11753_ | ~new_n11732_;
  assign new_n11753_ = ~pi214 | ~new_n11615_;
  assign new_n11754_ = ~new_n11615_ | ~new_n11614_;
  assign new_n11755_ = ~new_n11640_ | ~new_n11596_;
  assign new_n11756_ = ~new_n11595_;
  assign new_n11757_ = ~new_n11447_ | ~new_n11596_;
  assign new_n11758_ = ~new_n11594_;
  assign new_n11759_ = ~new_n11448_ | ~new_n11596_;
  assign new_n11760_ = ~new_n11593_;
  assign new_n11761_ = ~new_n11554_ | ~new_n11596_;
  assign new_n11762_ = ~new_n11592_;
  assign new_n11763_ = ~new_n11567_ | ~new_n11602_;
  assign new_n11764_ = ~pi467 | ~new_n11472_;
  assign new_n11765_ = ~pi222 | ~new_n11471_;
  assign new_n11766_ = ~new_n11556_;
  assign new_n11767_ = ~new_n11762_ | ~new_n11766_;
  assign new_n11768_ = ~new_n11556_ | ~new_n11592_;
  assign new_n11769_ = ~pi466 | ~new_n11454_;
  assign new_n11770_ = ~pi221 | ~new_n11455_;
  assign new_n11771_ = ~new_n11557_;
  assign new_n11772_ = ~new_n11760_ | ~new_n11771_;
  assign new_n11773_ = ~new_n11557_ | ~new_n11593_;
  assign new_n11774_ = ~pi465 | ~new_n11458_;
  assign new_n11775_ = ~pi220 | ~new_n11456_;
  assign new_n11776_ = ~new_n11559_;
  assign new_n11777_ = ~new_n11758_ | ~new_n11776_;
  assign new_n11778_ = ~new_n11559_ | ~new_n11594_;
  assign new_n11779_ = ~pi464 | ~new_n11457_;
  assign new_n11780_ = ~pi219 | ~new_n11459_;
  assign new_n11781_ = ~new_n11560_;
  assign new_n11782_ = ~new_n11756_ | ~new_n11781_;
  assign new_n11783_ = ~new_n11560_ | ~new_n11595_;
  assign new_n11784_ = ~pi463 | ~new_n11460_;
  assign new_n11785_ = ~pi218 | ~new_n11470_;
  assign new_n11786_ = ~new_n11561_;
  assign new_n11787_ = ~new_n11639_ | ~new_n11786_;
  assign new_n11788_ = ~new_n11561_ | ~new_n11596_;
  assign new_n11789_ = ~pi462 | ~new_n11462_;
  assign new_n11790_ = ~pi217 | ~new_n11465_;
  assign new_n11791_ = ~new_n11562_;
  assign new_n11792_ = ~new_n11636_ | ~new_n11791_;
  assign new_n11793_ = ~new_n11562_ | ~new_n11597_;
  assign new_n11794_ = ~pi461 | ~new_n11469_;
  assign new_n11795_ = ~pi216 | ~new_n11467_;
  assign new_n11796_ = ~new_n11563_;
  assign new_n11797_ = ~new_n11633_ | ~new_n11796_;
  assign new_n11798_ = ~new_n11563_ | ~new_n11598_;
  assign new_n11799_ = ~pi489 | ~new_n11600_;
  assign new_n11800_ = ~pi244 | ~new_n11599_;
  assign new_n11801_ = ~new_n11800_ | ~new_n11799_;
  assign new_n11802_ = ~pi489 | ~new_n11600_;
  assign new_n11803_ = ~pi244 | ~new_n11599_;
  assign new_n11804_ = ~new_n11515_ | ~pi243 | ~new_n11801_;
  assign new_n11805_ = ~pi488 | ~new_n11451_ | ~new_n11514_;
  assign new_n11806_ = ~pi488 | ~new_n11514_;
  assign new_n11807_ = ~pi243 | ~new_n11515_;
  assign new_n11808_ = ~new_n11569_;
  assign new_n11809_ = ~new_n11728_ | ~new_n11808_;
  assign new_n11810_ = ~new_n11569_ | ~new_n11602_;
  assign new_n11811_ = ~pi460 | ~new_n11468_;
  assign new_n11812_ = ~pi215 | ~new_n11466_;
  assign new_n11813_ = ~new_n11570_;
  assign new_n11814_ = ~new_n11629_ | ~new_n11813_;
  assign new_n11815_ = ~new_n11570_ | ~new_n11603_;
  assign new_n11816_ = ~pi487 | ~new_n11513_;
  assign new_n11817_ = ~pi242 | ~new_n11512_;
  assign new_n11818_ = ~new_n11571_;
  assign new_n11819_ = ~new_n11724_ | ~new_n11818_;
  assign new_n11820_ = ~new_n11571_ | ~new_n11604_;
  assign new_n11821_ = ~pi486 | ~new_n11511_;
  assign new_n11822_ = ~pi241 | ~new_n11510_;
  assign new_n11823_ = ~new_n11572_;
  assign new_n11824_ = ~new_n11720_ | ~new_n11823_;
  assign new_n11825_ = ~new_n11572_ | ~new_n11605_;
  assign new_n11826_ = ~pi485 | ~new_n11509_;
  assign new_n11827_ = ~pi240 | ~new_n11508_;
  assign new_n11828_ = ~new_n11573_;
  assign new_n11829_ = ~new_n11716_ | ~new_n11828_;
  assign new_n11830_ = ~new_n11573_ | ~new_n11606_;
  assign new_n11831_ = ~pi484 | ~new_n11507_;
  assign new_n11832_ = ~pi239 | ~new_n11506_;
  assign new_n11833_ = ~new_n11574_;
  assign new_n11834_ = ~new_n11712_ | ~new_n11833_;
  assign new_n11835_ = ~new_n11574_ | ~new_n11607_;
  assign new_n11836_ = ~pi483 | ~new_n11505_;
  assign new_n11837_ = ~pi238 | ~new_n11504_;
  assign new_n11838_ = ~new_n11575_;
  assign new_n11839_ = ~new_n11708_ | ~new_n11838_;
  assign new_n11840_ = ~new_n11575_ | ~new_n11608_;
  assign new_n11841_ = ~pi482 | ~new_n11503_;
  assign new_n11842_ = ~pi237 | ~new_n11502_;
  assign new_n11843_ = ~new_n11576_;
  assign new_n11844_ = ~new_n11704_ | ~new_n11843_;
  assign new_n11845_ = ~new_n11576_ | ~new_n11609_;
  assign new_n11846_ = ~pi481 | ~new_n11501_;
  assign new_n11847_ = ~pi236 | ~new_n11500_;
  assign new_n11848_ = ~new_n11577_;
  assign new_n11849_ = ~new_n11700_ | ~new_n11848_;
  assign new_n11850_ = ~new_n11577_ | ~new_n11610_;
  assign new_n11851_ = ~pi480 | ~new_n11499_;
  assign new_n11852_ = ~pi235 | ~new_n11498_;
  assign new_n11853_ = ~new_n11578_;
  assign new_n11854_ = ~new_n11696_ | ~new_n11853_;
  assign new_n11855_ = ~new_n11578_ | ~new_n11611_;
  assign new_n11856_ = ~pi479 | ~new_n11497_;
  assign new_n11857_ = ~pi234 | ~new_n11496_;
  assign new_n11858_ = ~new_n11579_;
  assign new_n11859_ = ~new_n11692_ | ~new_n11858_;
  assign new_n11860_ = ~new_n11579_ | ~new_n11612_;
  assign new_n11861_ = ~pi478 | ~new_n11495_;
  assign new_n11862_ = ~pi233 | ~new_n11494_;
  assign new_n11863_ = ~new_n11580_;
  assign new_n11864_ = ~new_n11688_ | ~new_n11863_;
  assign new_n11865_ = ~new_n11580_ | ~new_n11613_;
  assign new_n11866_ = ~pi459 | ~new_n11464_;
  assign new_n11867_ = ~pi214 | ~new_n11614_;
  assign new_n11868_ = ~new_n11581_;
  assign new_n11869_ = ~new_n11627_ | ~new_n11868_;
  assign new_n11870_ = ~new_n11581_ | ~new_n11615_;
  assign new_n11871_ = ~pi477 | ~new_n11493_;
  assign new_n11872_ = ~pi232 | ~new_n11492_;
  assign new_n11873_ = ~new_n11582_;
  assign new_n11874_ = ~new_n11684_ | ~new_n11873_;
  assign new_n11875_ = ~new_n11582_ | ~new_n11616_;
  assign new_n11876_ = ~pi476 | ~new_n11491_;
  assign new_n11877_ = ~pi231 | ~new_n11490_;
  assign new_n11878_ = ~new_n11583_;
  assign new_n11879_ = ~new_n11680_ | ~new_n11878_;
  assign new_n11880_ = ~new_n11583_ | ~new_n11617_;
  assign new_n11881_ = ~pi475 | ~new_n11489_;
  assign new_n11882_ = ~pi230 | ~new_n11488_;
  assign new_n11883_ = ~new_n11584_;
  assign new_n11884_ = ~new_n11676_ | ~new_n11883_;
  assign new_n11885_ = ~new_n11584_ | ~new_n11618_;
  assign new_n11886_ = ~pi474 | ~new_n11487_;
  assign new_n11887_ = ~pi229 | ~new_n11486_;
  assign new_n11888_ = ~new_n11585_;
  assign new_n11889_ = ~new_n11672_ | ~new_n11888_;
  assign new_n11890_ = ~new_n11585_ | ~new_n11619_;
  assign new_n11891_ = ~pi473 | ~new_n11485_;
  assign new_n11892_ = ~pi228 | ~new_n11484_;
  assign new_n11893_ = ~new_n11586_;
  assign new_n11894_ = ~new_n11668_ | ~new_n11893_;
  assign new_n11895_ = ~new_n11586_ | ~new_n11620_;
  assign new_n11896_ = ~pi472 | ~new_n11483_;
  assign new_n11897_ = ~pi227 | ~new_n11482_;
  assign new_n11898_ = ~new_n11587_;
  assign new_n11899_ = ~new_n11664_ | ~new_n11898_;
  assign new_n11900_ = ~new_n11587_ | ~new_n11621_;
  assign new_n11901_ = ~pi471 | ~new_n11481_;
  assign new_n11902_ = ~pi226 | ~new_n11480_;
  assign new_n11903_ = ~new_n11588_;
  assign new_n11904_ = ~new_n11660_ | ~new_n11903_;
  assign new_n11905_ = ~new_n11588_ | ~new_n11622_;
  assign new_n11906_ = ~pi470 | ~new_n11473_;
  assign new_n11907_ = ~pi225 | ~new_n11474_;
  assign new_n11908_ = ~new_n11589_;
  assign new_n11909_ = ~new_n11657_ | ~new_n11908_;
  assign new_n11910_ = ~new_n11589_ | ~new_n11623_;
  assign new_n11911_ = ~pi469 | ~new_n11477_;
  assign new_n11912_ = ~pi224 | ~new_n11475_;
  assign new_n11913_ = ~new_n11590_;
  assign new_n11914_ = ~new_n11654_ | ~new_n11913_;
  assign new_n11915_ = ~new_n11590_ | ~new_n11624_;
  assign new_n11916_ = ~pi468 | ~new_n11478_;
  assign new_n11917_ = ~pi223 | ~new_n11476_;
  assign new_n11918_ = ~new_n11591_;
  assign new_n11919_ = ~new_n11651_ | ~new_n11918_;
  assign new_n11920_ = ~new_n11591_ | ~new_n11625_;
  assign new_n11921_ = new_n12123_ & new_n12119_;
  assign new_n11922_ = new_n12131_ & new_n12129_;
  assign new_n11923_ = new_n11922_ & new_n12133_;
  assign new_n11924_ = new_n12139_ & new_n12137_;
  assign new_n11925_ = new_n11924_ & new_n12141_;
  assign new_n11926_ = new_n11925_ & new_n12143_;
  assign new_n11927_ = new_n12116_ & new_n12113_;
  assign new_n11928_ = new_n12308_ & new_n12307_;
  assign new_n11929_ = new_n12045_ & new_n12110_;
  assign new_n11930_ = ~new_n12089_ | ~new_n12254_;
  assign new_n11931_ = ~pi024;
  assign new_n11932_ = ~new_n1628_;
  assign new_n11933_ = ~pi025;
  assign new_n11934_ = ~new_n1629_;
  assign new_n11935_ = ~new_n1629_ | ~pi025;
  assign new_n11936_ = ~pi026;
  assign new_n11937_ = ~new_n1630_;
  assign new_n11938_ = ~pi029;
  assign new_n11939_ = ~new_n1635_;
  assign new_n11940_ = ~pi031;
  assign new_n11941_ = ~pi032;
  assign new_n11942_ = ~new_n1658_;
  assign new_n11943_ = ~new_n1657_;
  assign new_n11944_ = ~pi030;
  assign new_n11945_ = ~new_n1646_;
  assign new_n11946_ = ~new_n1646_ | ~pi030;
  assign new_n11947_ = ~pi027;
  assign new_n11948_ = ~new_n1631_;
  assign new_n11949_ = ~pi028;
  assign new_n11950_ = ~new_n1632_;
  assign new_n11951_ = ~new_n1632_ | ~pi028;
  assign new_n11952_ = ~new_n1627_;
  assign new_n11953_ = ~pi023;
  assign new_n11954_ = ~new_n12211_ | ~new_n12124_;
  assign new_n11955_ = ~pi017;
  assign new_n11956_ = ~new_n1651_;
  assign new_n11957_ = ~pi018;
  assign new_n11958_ = ~new_n1652_;
  assign new_n11959_ = ~pi019;
  assign new_n11960_ = ~new_n1653_;
  assign new_n11961_ = ~pi020;
  assign new_n11962_ = ~new_n1654_;
  assign new_n11963_ = ~pi021;
  assign new_n11964_ = ~new_n1655_;
  assign new_n11965_ = ~new_n1655_ | ~pi021;
  assign new_n11966_ = ~pi022;
  assign new_n11967_ = ~new_n1656_;
  assign new_n11968_ = ~pi016;
  assign new_n11969_ = ~new_n1650_;
  assign new_n11970_ = ~pi015;
  assign new_n11971_ = ~new_n1649_;
  assign new_n11972_ = ~pi014;
  assign new_n11973_ = ~new_n1648_;
  assign new_n11974_ = ~pi013;
  assign new_n11975_ = ~new_n1647_;
  assign new_n11976_ = ~pi012;
  assign new_n11977_ = ~new_n1645_;
  assign new_n11978_ = ~pi011;
  assign new_n11979_ = ~new_n1644_;
  assign new_n11980_ = ~pi010;
  assign new_n11981_ = ~new_n1643_;
  assign new_n11982_ = ~pi009;
  assign new_n11983_ = ~new_n1642_;
  assign new_n11984_ = ~pi008;
  assign new_n11985_ = ~new_n1641_;
  assign new_n11986_ = ~pi007;
  assign new_n11987_ = ~new_n1640_;
  assign new_n11988_ = ~pi006;
  assign new_n11989_ = ~new_n1639_;
  assign new_n11990_ = ~pi005;
  assign new_n11991_ = ~new_n1638_;
  assign new_n11992_ = ~pi004;
  assign new_n11993_ = ~new_n1637_;
  assign new_n11994_ = ~pi003;
  assign new_n11995_ = ~new_n1636_;
  assign new_n11996_ = ~pi002;
  assign new_n11997_ = ~new_n1634_;
  assign new_n11998_ = ~new_n12224_ | ~new_n12144_;
  assign new_n11999_ = ~new_n12222_ | ~new_n12142_;
  assign new_n12000_ = ~new_n12217_ | ~new_n12134_;
  assign new_n12001_ = ~new_n12471_ | ~new_n12470_;
  assign new_n12002_ = ~new_n12261_ | ~new_n12260_;
  assign new_n12003_ = ~new_n12268_ | ~new_n12267_;
  assign new_n12004_ = ~new_n12275_ | ~new_n12274_;
  assign new_n12005_ = ~new_n12282_ | ~new_n12281_;
  assign new_n12006_ = ~new_n12289_ | ~new_n12288_;
  assign new_n12007_ = ~new_n12296_ | ~new_n12295_;
  assign new_n12008_ = ~new_n12303_ | ~new_n12302_;
  assign new_n12009_ = ~new_n12317_ | ~new_n12316_;
  assign new_n12010_ = ~new_n12324_ | ~new_n12323_;
  assign new_n12011_ = ~new_n12331_ | ~new_n12330_;
  assign new_n12012_ = ~new_n12338_ | ~new_n12337_;
  assign new_n12013_ = ~new_n12345_ | ~new_n12344_;
  assign new_n12014_ = ~new_n12352_ | ~new_n12351_;
  assign new_n12015_ = ~new_n12359_ | ~new_n12358_;
  assign new_n12016_ = ~new_n12366_ | ~new_n12365_;
  assign new_n12017_ = ~new_n12373_ | ~new_n12372_;
  assign new_n12018_ = ~new_n12380_ | ~new_n12379_;
  assign new_n12019_ = ~new_n12387_ | ~new_n12386_;
  assign new_n12020_ = ~new_n12394_ | ~new_n12393_;
  assign new_n12021_ = ~new_n12406_ | ~new_n12405_;
  assign new_n12022_ = ~new_n12413_ | ~new_n12412_;
  assign new_n12023_ = ~new_n12420_ | ~new_n12419_;
  assign new_n12024_ = ~new_n12427_ | ~new_n12426_;
  assign new_n12025_ = ~new_n12434_ | ~new_n12433_;
  assign new_n12026_ = ~new_n12441_ | ~new_n12440_;
  assign new_n12027_ = ~new_n12448_ | ~new_n12447_;
  assign new_n12028_ = ~new_n12455_ | ~new_n12454_;
  assign new_n12029_ = ~new_n12462_ | ~new_n12461_;
  assign new_n12030_ = ~new_n12469_ | ~new_n12468_;
  assign new_n12031_ = new_n12209_ & new_n12117_;
  assign new_n12032_ = new_n12126_ & new_n11921_;
  assign new_n12033_ = new_n12214_ & new_n12127_;
  assign new_n12034_ = new_n12215_ & new_n12132_;
  assign new_n12035_ = new_n12209_ & new_n12117_;
  assign new_n12036_ = new_n1657_ & new_n1658_;
  assign new_n12037_ = new_n1658_ & pi032;
  assign new_n12038_ = pi031 & new_n1657_;
  assign new_n12039_ = new_n12135_ & new_n11923_;
  assign new_n12040_ = new_n12219_ & new_n12136_;
  assign new_n12041_ = new_n11926_ & new_n12145_;
  assign new_n12042_ = new_n12226_ & new_n12146_;
  assign new_n12043_ = new_n12204_ & new_n12306_;
  assign new_n12044_ = new_n12201_ & new_n11928_ & new_n12203_;
  assign new_n12045_ = new_n12205_ & new_n12063_;
  assign new_n12046_ = new_n12220_ & new_n12140_;
  assign new_n12047_ = new_n12256_ & new_n12255_;
  assign new_n12048_ = ~new_n12034_ | ~new_n12248_;
  assign new_n12049_ = new_n12263_ & new_n12262_;
  assign new_n12050_ = ~new_n12246_ | ~new_n11935_;
  assign new_n12051_ = new_n12270_ & new_n12269_;
  assign new_n12052_ = ~new_n12033_ | ~new_n12213_;
  assign new_n12053_ = new_n12277_ & new_n12276_;
  assign new_n12054_ = ~new_n12212_ | ~new_n12210_;
  assign new_n12055_ = new_n12284_ & new_n12283_;
  assign new_n12056_ = ~new_n11951_ | ~new_n12120_;
  assign new_n12057_ = new_n12291_ & new_n12290_;
  assign new_n12058_ = ~new_n12035_ | ~new_n12232_;
  assign new_n12059_ = new_n12298_ & new_n12297_;
  assign new_n12060_ = ~new_n12228_ | ~new_n11946_ | ~new_n12227_ | ~new_n12229_;
  assign new_n12061_ = ~new_n1633_;
  assign new_n12062_ = ~pi001;
  assign new_n12063_ = new_n12310_ & new_n12309_;
  assign new_n12064_ = new_n12312_ & new_n12311_;
  assign new_n12065_ = ~new_n12201_ | ~new_n12200_;
  assign new_n12066_ = ~new_n12206_ | ~new_n12207_ | ~new_n12088_;
  assign new_n12067_ = new_n12326_ & new_n12325_;
  assign new_n12068_ = ~new_n12197_ | ~new_n12196_;
  assign new_n12069_ = new_n12333_ & new_n12332_;
  assign new_n12070_ = ~new_n12193_ | ~new_n12192_;
  assign new_n12071_ = new_n12340_ & new_n12339_;
  assign new_n12072_ = ~new_n12189_ | ~new_n12188_;
  assign new_n12073_ = new_n12347_ & new_n12346_;
  assign new_n12074_ = ~new_n12185_ | ~new_n12184_;
  assign new_n12075_ = new_n12354_ & new_n12353_;
  assign new_n12076_ = ~new_n12181_ | ~new_n12180_;
  assign new_n12077_ = new_n12361_ & new_n12360_;
  assign new_n12078_ = ~new_n12177_ | ~new_n12176_;
  assign new_n12079_ = new_n12368_ & new_n12367_;
  assign new_n12080_ = ~new_n12173_ | ~new_n12172_;
  assign new_n12081_ = new_n12375_ & new_n12374_;
  assign new_n12082_ = ~new_n12169_ | ~new_n12168_;
  assign new_n12083_ = new_n12382_ & new_n12381_;
  assign new_n12084_ = ~new_n12165_ | ~new_n12164_;
  assign new_n12085_ = new_n12389_ & new_n12388_;
  assign new_n12086_ = ~new_n12161_ | ~new_n12160_;
  assign new_n12087_ = ~new_n1658_ | ~pi032;
  assign new_n12088_ = ~new_n1658_ | ~pi032 | ~pi031;
  assign new_n12089_ = new_n12399_ & new_n12398_;
  assign new_n12090_ = new_n12401_ & new_n12400_;
  assign new_n12091_ = ~new_n12157_ | ~new_n12156_;
  assign new_n12092_ = new_n12408_ & new_n12407_;
  assign new_n12093_ = ~new_n12153_ | ~new_n12152_;
  assign new_n12094_ = new_n12415_ & new_n12414_;
  assign new_n12095_ = ~new_n12149_ | ~new_n12148_;
  assign new_n12096_ = new_n12422_ & new_n12421_;
  assign new_n12097_ = ~new_n12042_ | ~new_n12244_;
  assign new_n12098_ = new_n12429_ & new_n12428_;
  assign new_n12099_ = ~new_n12225_ | ~new_n12242_;
  assign new_n12100_ = new_n12436_ & new_n12435_;
  assign new_n12101_ = ~new_n12223_ | ~new_n12240_;
  assign new_n12102_ = new_n12443_ & new_n12442_;
  assign new_n12103_ = ~new_n12046_ | ~new_n12238_;
  assign new_n12104_ = new_n12450_ & new_n12449_;
  assign new_n12105_ = ~new_n12236_ | ~new_n11965_;
  assign new_n12106_ = new_n12457_ & new_n12456_;
  assign new_n12107_ = ~new_n12040_ | ~new_n12252_;
  assign new_n12108_ = new_n12464_ & new_n12463_;
  assign new_n12109_ = ~new_n12218_ | ~new_n12250_;
  assign new_n12110_ = ~new_n12043_ | ~new_n12065_;
  assign new_n12111_ = ~new_n12088_;
  assign new_n12112_ = ~new_n12066_;
  assign new_n12113_ = pi030 | new_n1646_;
  assign new_n12114_ = ~new_n11946_;
  assign new_n12115_ = ~new_n12060_;
  assign new_n12116_ = pi029 | new_n1635_;
  assign new_n12117_ = ~new_n1635_ | ~pi029;
  assign new_n12118_ = ~new_n12031_ | ~new_n12208_;
  assign new_n12119_ = pi028 | new_n1632_;
  assign new_n12120_ = ~new_n12119_ | ~new_n12118_;
  assign new_n12121_ = ~new_n11951_;
  assign new_n12122_ = ~new_n12056_;
  assign new_n12123_ = pi027 | new_n1631_;
  assign new_n12124_ = ~new_n1631_ | ~pi027;
  assign new_n12125_ = ~new_n12054_;
  assign new_n12126_ = pi026 | new_n1630_;
  assign new_n12127_ = ~new_n1630_ | ~pi026;
  assign new_n12128_ = ~new_n12052_;
  assign new_n12129_ = pi025 | new_n1629_;
  assign new_n12130_ = ~new_n11935_;
  assign new_n12131_ = pi024 | new_n1628_;
  assign new_n12132_ = ~new_n1628_ | ~pi024;
  assign new_n12133_ = pi023 | new_n1627_;
  assign new_n12134_ = ~pi023 | ~new_n1627_;
  assign new_n12135_ = pi022 | new_n1656_;
  assign new_n12136_ = ~new_n1656_ | ~pi022;
  assign new_n12137_ = pi021 | new_n1655_;
  assign new_n12138_ = ~new_n11965_;
  assign new_n12139_ = pi020 | new_n1654_;
  assign new_n12140_ = ~new_n1654_ | ~pi020;
  assign new_n12141_ = pi019 | new_n1653_;
  assign new_n12142_ = ~new_n1653_ | ~pi019;
  assign new_n12143_ = pi018 | new_n1652_;
  assign new_n12144_ = ~new_n1652_ | ~pi018;
  assign new_n12145_ = pi017 | new_n1651_;
  assign new_n12146_ = ~new_n1651_ | ~pi017;
  assign new_n12147_ = pi016 | new_n1650_;
  assign new_n12148_ = ~new_n12147_ | ~new_n12097_;
  assign new_n12149_ = ~new_n1650_ | ~pi016;
  assign new_n12150_ = ~new_n12095_;
  assign new_n12151_ = pi015 | new_n1649_;
  assign new_n12152_ = ~new_n12151_ | ~new_n12095_;
  assign new_n12153_ = ~new_n1649_ | ~pi015;
  assign new_n12154_ = ~new_n12093_;
  assign new_n12155_ = pi014 | new_n1648_;
  assign new_n12156_ = ~new_n12155_ | ~new_n12093_;
  assign new_n12157_ = ~new_n1648_ | ~pi014;
  assign new_n12158_ = ~new_n12091_;
  assign new_n12159_ = pi013 | new_n1647_;
  assign new_n12160_ = ~new_n12159_ | ~new_n12091_;
  assign new_n12161_ = ~new_n1647_ | ~pi013;
  assign new_n12162_ = ~new_n12086_;
  assign new_n12163_ = pi012 | new_n1645_;
  assign new_n12164_ = ~new_n12163_ | ~new_n12086_;
  assign new_n12165_ = ~new_n1645_ | ~pi012;
  assign new_n12166_ = ~new_n12084_;
  assign new_n12167_ = pi011 | new_n1644_;
  assign new_n12168_ = ~new_n12167_ | ~new_n12084_;
  assign new_n12169_ = ~new_n1644_ | ~pi011;
  assign new_n12170_ = ~new_n12082_;
  assign new_n12171_ = pi010 | new_n1643_;
  assign new_n12172_ = ~new_n12171_ | ~new_n12082_;
  assign new_n12173_ = ~new_n1643_ | ~pi010;
  assign new_n12174_ = ~new_n12080_;
  assign new_n12175_ = pi009 | new_n1642_;
  assign new_n12176_ = ~new_n12175_ | ~new_n12080_;
  assign new_n12177_ = ~new_n1642_ | ~pi009;
  assign new_n12178_ = ~new_n12078_;
  assign new_n12179_ = pi008 | new_n1641_;
  assign new_n12180_ = ~new_n12179_ | ~new_n12078_;
  assign new_n12181_ = ~new_n1641_ | ~pi008;
  assign new_n12182_ = ~new_n12076_;
  assign new_n12183_ = pi007 | new_n1640_;
  assign new_n12184_ = ~new_n12183_ | ~new_n12076_;
  assign new_n12185_ = ~new_n1640_ | ~pi007;
  assign new_n12186_ = ~new_n12074_;
  assign new_n12187_ = pi006 | new_n1639_;
  assign new_n12188_ = ~new_n12187_ | ~new_n12074_;
  assign new_n12189_ = ~new_n1639_ | ~pi006;
  assign new_n12190_ = ~new_n12072_;
  assign new_n12191_ = pi005 | new_n1638_;
  assign new_n12192_ = ~new_n12191_ | ~new_n12072_;
  assign new_n12193_ = ~new_n1638_ | ~pi005;
  assign new_n12194_ = ~new_n12070_;
  assign new_n12195_ = pi004 | new_n1637_;
  assign new_n12196_ = ~new_n12195_ | ~new_n12070_;
  assign new_n12197_ = ~new_n1637_ | ~pi004;
  assign new_n12198_ = ~new_n12068_;
  assign new_n12199_ = pi003 | new_n1636_;
  assign new_n12200_ = ~new_n12199_ | ~new_n12068_;
  assign new_n12201_ = ~new_n1636_ | ~pi003;
  assign new_n12202_ = ~new_n12065_;
  assign new_n12203_ = ~new_n1634_ | ~pi002;
  assign new_n12204_ = new_n1634_ | pi002;
  assign new_n12205_ = ~new_n12200_ | ~new_n12044_;
  assign new_n12206_ = ~new_n1657_ | ~new_n1658_ | ~pi032;
  assign new_n12207_ = ~new_n1657_ | ~pi031;
  assign new_n12208_ = ~new_n11927_ | ~new_n12230_;
  assign new_n12209_ = ~new_n12114_ | ~new_n12116_;
  assign new_n12210_ = ~new_n11921_ | ~new_n12118_;
  assign new_n12211_ = ~new_n12121_ | ~new_n12123_;
  assign new_n12212_ = ~new_n11954_;
  assign new_n12213_ = ~new_n12032_ | ~new_n12118_;
  assign new_n12214_ = ~new_n11954_ | ~new_n12126_;
  assign new_n12215_ = ~new_n12130_ | ~new_n12131_;
  assign new_n12216_ = ~new_n12215_ | ~new_n12132_;
  assign new_n12217_ = ~new_n12216_ | ~new_n12133_;
  assign new_n12218_ = ~new_n12000_;
  assign new_n12219_ = ~new_n12000_ | ~new_n12135_;
  assign new_n12220_ = ~new_n12138_ | ~new_n12139_;
  assign new_n12221_ = ~new_n12220_ | ~new_n12140_;
  assign new_n12222_ = ~new_n12221_ | ~new_n12141_;
  assign new_n12223_ = ~new_n11999_;
  assign new_n12224_ = ~new_n11999_ | ~new_n12143_;
  assign new_n12225_ = ~new_n11998_;
  assign new_n12226_ = ~new_n11998_ | ~new_n12145_;
  assign new_n12227_ = ~new_n12036_ | ~pi032 | ~new_n12113_;
  assign new_n12228_ = ~new_n12037_ | ~pi031 | ~new_n12113_;
  assign new_n12229_ = ~new_n12038_ | ~new_n12113_;
  assign new_n12230_ = ~new_n12206_ | ~new_n12207_ | ~new_n12088_;
  assign new_n12231_ = ~new_n12058_;
  assign new_n12232_ = ~new_n11927_ | ~new_n12233_;
  assign new_n12233_ = ~new_n12234_ | ~new_n12235_ | ~new_n12207_;
  assign new_n12234_ = ~new_n1657_ | ~new_n1658_ | ~pi032;
  assign new_n12235_ = ~new_n1658_ | ~pi032 | ~pi031;
  assign new_n12236_ = ~new_n12137_ | ~new_n12107_;
  assign new_n12237_ = ~new_n12105_;
  assign new_n12238_ = ~new_n11924_ | ~new_n12107_;
  assign new_n12239_ = ~new_n12103_;
  assign new_n12240_ = ~new_n11925_ | ~new_n12107_;
  assign new_n12241_ = ~new_n12101_;
  assign new_n12242_ = ~new_n11926_ | ~new_n12107_;
  assign new_n12243_ = ~new_n12099_;
  assign new_n12244_ = ~new_n12041_ | ~new_n12107_;
  assign new_n12245_ = ~new_n12097_;
  assign new_n12246_ = ~new_n12129_ | ~new_n12052_;
  assign new_n12247_ = ~new_n12050_;
  assign new_n12248_ = ~new_n11922_ | ~new_n12052_;
  assign new_n12249_ = ~new_n12048_;
  assign new_n12250_ = ~new_n11923_ | ~new_n12052_;
  assign new_n12251_ = ~new_n12109_;
  assign new_n12252_ = ~new_n12039_ | ~new_n12052_;
  assign new_n12253_ = ~new_n12107_;
  assign new_n12254_ = ~new_n12397_ | ~new_n11940_;
  assign new_n12255_ = ~new_n1627_ | ~new_n11953_;
  assign new_n12256_ = ~pi023 | ~new_n11952_;
  assign new_n12257_ = ~new_n1627_ | ~new_n11953_;
  assign new_n12258_ = ~pi023 | ~new_n11952_;
  assign new_n12259_ = ~new_n12258_ | ~new_n12257_;
  assign new_n12260_ = ~new_n12047_ | ~new_n12048_;
  assign new_n12261_ = ~new_n12249_ | ~new_n12259_;
  assign new_n12262_ = ~new_n1628_ | ~new_n11931_;
  assign new_n12263_ = ~pi024 | ~new_n11932_;
  assign new_n12264_ = ~new_n1628_ | ~new_n11931_;
  assign new_n12265_ = ~pi024 | ~new_n11932_;
  assign new_n12266_ = ~new_n12265_ | ~new_n12264_;
  assign new_n12267_ = ~new_n12049_ | ~new_n12050_;
  assign new_n12268_ = ~new_n12247_ | ~new_n12266_;
  assign new_n12269_ = ~new_n1629_ | ~new_n11933_;
  assign new_n12270_ = ~pi025 | ~new_n11934_;
  assign new_n12271_ = ~new_n1629_ | ~new_n11933_;
  assign new_n12272_ = ~pi025 | ~new_n11934_;
  assign new_n12273_ = ~new_n12272_ | ~new_n12271_;
  assign new_n12274_ = ~new_n12051_ | ~new_n12052_;
  assign new_n12275_ = ~new_n12128_ | ~new_n12273_;
  assign new_n12276_ = ~new_n1630_ | ~new_n11936_;
  assign new_n12277_ = ~pi026 | ~new_n11937_;
  assign new_n12278_ = ~new_n1630_ | ~new_n11936_;
  assign new_n12279_ = ~pi026 | ~new_n11937_;
  assign new_n12280_ = ~new_n12279_ | ~new_n12278_;
  assign new_n12281_ = ~new_n12053_ | ~new_n12054_;
  assign new_n12282_ = ~new_n12125_ | ~new_n12280_;
  assign new_n12283_ = ~new_n1631_ | ~new_n11947_;
  assign new_n12284_ = ~pi027 | ~new_n11948_;
  assign new_n12285_ = ~new_n1631_ | ~new_n11947_;
  assign new_n12286_ = ~pi027 | ~new_n11948_;
  assign new_n12287_ = ~new_n12286_ | ~new_n12285_;
  assign new_n12288_ = ~new_n12055_ | ~new_n12056_;
  assign new_n12289_ = ~new_n12122_ | ~new_n12287_;
  assign new_n12290_ = ~new_n1632_ | ~new_n11949_;
  assign new_n12291_ = ~pi028 | ~new_n11950_;
  assign new_n12292_ = ~new_n1632_ | ~new_n11949_;
  assign new_n12293_ = ~pi028 | ~new_n11950_;
  assign new_n12294_ = ~new_n12293_ | ~new_n12292_;
  assign new_n12295_ = ~new_n12057_ | ~new_n12058_;
  assign new_n12296_ = ~new_n12231_ | ~new_n12294_;
  assign new_n12297_ = ~new_n1635_ | ~new_n11938_;
  assign new_n12298_ = ~pi029 | ~new_n11939_;
  assign new_n12299_ = ~new_n1635_ | ~new_n11938_;
  assign new_n12300_ = ~pi029 | ~new_n11939_;
  assign new_n12301_ = ~new_n12300_ | ~new_n12299_;
  assign new_n12302_ = ~new_n12059_ | ~new_n12060_;
  assign new_n12303_ = ~new_n12115_ | ~new_n12301_;
  assign new_n12304_ = ~new_n1633_ | ~new_n12062_;
  assign new_n12305_ = ~pi001 | ~new_n12061_;
  assign new_n12306_ = ~new_n12305_ | ~new_n12304_;
  assign new_n12307_ = ~new_n1633_ | ~new_n12062_;
  assign new_n12308_ = ~pi001 | ~new_n12061_;
  assign new_n12309_ = ~new_n11997_ | ~new_n11928_ | ~new_n11996_;
  assign new_n12310_ = ~new_n1634_ | ~pi002 | ~new_n12306_;
  assign new_n12311_ = ~new_n1634_ | ~new_n11996_;
  assign new_n12312_ = ~pi002 | ~new_n11997_;
  assign new_n12313_ = ~new_n1634_ | ~new_n11996_;
  assign new_n12314_ = ~pi002 | ~new_n11997_;
  assign new_n12315_ = ~new_n12314_ | ~new_n12313_;
  assign new_n12316_ = ~new_n12064_ | ~new_n12065_;
  assign new_n12317_ = ~new_n12202_ | ~new_n12315_;
  assign new_n12318_ = ~new_n1646_ | ~new_n11944_;
  assign new_n12319_ = ~pi030 | ~new_n11945_;
  assign new_n12320_ = ~new_n1646_ | ~new_n11944_;
  assign new_n12321_ = ~pi030 | ~new_n11945_;
  assign new_n12322_ = ~new_n12321_ | ~new_n12320_;
  assign new_n12323_ = ~new_n12066_ | ~new_n12319_ | ~new_n12318_;
  assign new_n12324_ = ~new_n12112_ | ~new_n12322_;
  assign new_n12325_ = ~new_n1636_ | ~new_n11994_;
  assign new_n12326_ = ~pi003 | ~new_n11995_;
  assign new_n12327_ = ~new_n1636_ | ~new_n11994_;
  assign new_n12328_ = ~pi003 | ~new_n11995_;
  assign new_n12329_ = ~new_n12328_ | ~new_n12327_;
  assign new_n12330_ = ~new_n12067_ | ~new_n12068_;
  assign new_n12331_ = ~new_n12198_ | ~new_n12329_;
  assign new_n12332_ = ~new_n1637_ | ~new_n11992_;
  assign new_n12333_ = ~pi004 | ~new_n11993_;
  assign new_n12334_ = ~new_n1637_ | ~new_n11992_;
  assign new_n12335_ = ~pi004 | ~new_n11993_;
  assign new_n12336_ = ~new_n12335_ | ~new_n12334_;
  assign new_n12337_ = ~new_n12069_ | ~new_n12070_;
  assign new_n12338_ = ~new_n12194_ | ~new_n12336_;
  assign new_n12339_ = ~new_n1638_ | ~new_n11990_;
  assign new_n12340_ = ~pi005 | ~new_n11991_;
  assign new_n12341_ = ~new_n1638_ | ~new_n11990_;
  assign new_n12342_ = ~pi005 | ~new_n11991_;
  assign new_n12343_ = ~new_n12342_ | ~new_n12341_;
  assign new_n12344_ = ~new_n12071_ | ~new_n12072_;
  assign new_n12345_ = ~new_n12190_ | ~new_n12343_;
  assign new_n12346_ = ~new_n1639_ | ~new_n11988_;
  assign new_n12347_ = ~pi006 | ~new_n11989_;
  assign new_n12348_ = ~new_n1639_ | ~new_n11988_;
  assign new_n12349_ = ~pi006 | ~new_n11989_;
  assign new_n12350_ = ~new_n12349_ | ~new_n12348_;
  assign new_n12351_ = ~new_n12073_ | ~new_n12074_;
  assign new_n12352_ = ~new_n12186_ | ~new_n12350_;
  assign new_n12353_ = ~new_n1640_ | ~new_n11986_;
  assign new_n12354_ = ~pi007 | ~new_n11987_;
  assign new_n12355_ = ~new_n1640_ | ~new_n11986_;
  assign new_n12356_ = ~pi007 | ~new_n11987_;
  assign new_n12357_ = ~new_n12356_ | ~new_n12355_;
  assign new_n12358_ = ~new_n12075_ | ~new_n12076_;
  assign new_n12359_ = ~new_n12182_ | ~new_n12357_;
  assign new_n12360_ = ~new_n1641_ | ~new_n11984_;
  assign new_n12361_ = ~pi008 | ~new_n11985_;
  assign new_n12362_ = ~new_n1641_ | ~new_n11984_;
  assign new_n12363_ = ~pi008 | ~new_n11985_;
  assign new_n12364_ = ~new_n12363_ | ~new_n12362_;
  assign new_n12365_ = ~new_n12077_ | ~new_n12078_;
  assign new_n12366_ = ~new_n12178_ | ~new_n12364_;
  assign new_n12367_ = ~new_n1642_ | ~new_n11982_;
  assign new_n12368_ = ~pi009 | ~new_n11983_;
  assign new_n12369_ = ~new_n1642_ | ~new_n11982_;
  assign new_n12370_ = ~pi009 | ~new_n11983_;
  assign new_n12371_ = ~new_n12370_ | ~new_n12369_;
  assign new_n12372_ = ~new_n12079_ | ~new_n12080_;
  assign new_n12373_ = ~new_n12174_ | ~new_n12371_;
  assign new_n12374_ = ~new_n1643_ | ~new_n11980_;
  assign new_n12375_ = ~pi010 | ~new_n11981_;
  assign new_n12376_ = ~new_n1643_ | ~new_n11980_;
  assign new_n12377_ = ~pi010 | ~new_n11981_;
  assign new_n12378_ = ~new_n12377_ | ~new_n12376_;
  assign new_n12379_ = ~new_n12081_ | ~new_n12082_;
  assign new_n12380_ = ~new_n12170_ | ~new_n12378_;
  assign new_n12381_ = ~new_n1644_ | ~new_n11978_;
  assign new_n12382_ = ~pi011 | ~new_n11979_;
  assign new_n12383_ = ~new_n1644_ | ~new_n11978_;
  assign new_n12384_ = ~pi011 | ~new_n11979_;
  assign new_n12385_ = ~new_n12384_ | ~new_n12383_;
  assign new_n12386_ = ~new_n12083_ | ~new_n12084_;
  assign new_n12387_ = ~new_n12166_ | ~new_n12385_;
  assign new_n12388_ = ~new_n1645_ | ~new_n11976_;
  assign new_n12389_ = ~pi012 | ~new_n11977_;
  assign new_n12390_ = ~new_n1645_ | ~new_n11976_;
  assign new_n12391_ = ~pi012 | ~new_n11977_;
  assign new_n12392_ = ~new_n12391_ | ~new_n12390_;
  assign new_n12393_ = ~new_n12085_ | ~new_n12086_;
  assign new_n12394_ = ~new_n12162_ | ~new_n12392_;
  assign new_n12395_ = ~new_n1657_ | ~new_n12087_;
  assign new_n12396_ = ~new_n12037_ | ~new_n11943_;
  assign new_n12397_ = ~new_n12396_ | ~new_n12395_;
  assign new_n12398_ = ~new_n11943_ | ~pi031 | ~new_n12087_;
  assign new_n12399_ = ~new_n12111_ | ~new_n1657_;
  assign new_n12400_ = ~new_n1647_ | ~new_n11974_;
  assign new_n12401_ = ~pi013 | ~new_n11975_;
  assign new_n12402_ = ~new_n1647_ | ~new_n11974_;
  assign new_n12403_ = ~pi013 | ~new_n11975_;
  assign new_n12404_ = ~new_n12403_ | ~new_n12402_;
  assign new_n12405_ = ~new_n12090_ | ~new_n12091_;
  assign new_n12406_ = ~new_n12158_ | ~new_n12404_;
  assign new_n12407_ = ~new_n1648_ | ~new_n11972_;
  assign new_n12408_ = ~pi014 | ~new_n11973_;
  assign new_n12409_ = ~new_n1648_ | ~new_n11972_;
  assign new_n12410_ = ~pi014 | ~new_n11973_;
  assign new_n12411_ = ~new_n12410_ | ~new_n12409_;
  assign new_n12412_ = ~new_n12092_ | ~new_n12093_;
  assign new_n12413_ = ~new_n12154_ | ~new_n12411_;
  assign new_n12414_ = ~new_n1649_ | ~new_n11970_;
  assign new_n12415_ = ~pi015 | ~new_n11971_;
  assign new_n12416_ = ~new_n1649_ | ~new_n11970_;
  assign new_n12417_ = ~pi015 | ~new_n11971_;
  assign new_n12418_ = ~new_n12417_ | ~new_n12416_;
  assign new_n12419_ = ~new_n12094_ | ~new_n12095_;
  assign new_n12420_ = ~new_n12150_ | ~new_n12418_;
  assign new_n12421_ = ~new_n1650_ | ~new_n11968_;
  assign new_n12422_ = ~pi016 | ~new_n11969_;
  assign new_n12423_ = ~new_n1650_ | ~new_n11968_;
  assign new_n12424_ = ~pi016 | ~new_n11969_;
  assign new_n12425_ = ~new_n12424_ | ~new_n12423_;
  assign new_n12426_ = ~new_n12096_ | ~new_n12097_;
  assign new_n12427_ = ~new_n12245_ | ~new_n12425_;
  assign new_n12428_ = ~new_n1651_ | ~new_n11955_;
  assign new_n12429_ = ~pi017 | ~new_n11956_;
  assign new_n12430_ = ~new_n1651_ | ~new_n11955_;
  assign new_n12431_ = ~pi017 | ~new_n11956_;
  assign new_n12432_ = ~new_n12431_ | ~new_n12430_;
  assign new_n12433_ = ~new_n12098_ | ~new_n12099_;
  assign new_n12434_ = ~new_n12243_ | ~new_n12432_;
  assign new_n12435_ = ~new_n1652_ | ~new_n11957_;
  assign new_n12436_ = ~pi018 | ~new_n11958_;
  assign new_n12437_ = ~new_n1652_ | ~new_n11957_;
  assign new_n12438_ = ~pi018 | ~new_n11958_;
  assign new_n12439_ = ~new_n12438_ | ~new_n12437_;
  assign new_n12440_ = ~new_n12100_ | ~new_n12101_;
  assign new_n12441_ = ~new_n12241_ | ~new_n12439_;
  assign new_n12442_ = ~new_n1653_ | ~new_n11959_;
  assign new_n12443_ = ~pi019 | ~new_n11960_;
  assign new_n12444_ = ~new_n1653_ | ~new_n11959_;
  assign new_n12445_ = ~pi019 | ~new_n11960_;
  assign new_n12446_ = ~new_n12445_ | ~new_n12444_;
  assign new_n12447_ = ~new_n12102_ | ~new_n12103_;
  assign new_n12448_ = ~new_n12239_ | ~new_n12446_;
  assign new_n12449_ = ~new_n1654_ | ~new_n11961_;
  assign new_n12450_ = ~pi020 | ~new_n11962_;
  assign new_n12451_ = ~new_n1654_ | ~new_n11961_;
  assign new_n12452_ = ~pi020 | ~new_n11962_;
  assign new_n12453_ = ~new_n12452_ | ~new_n12451_;
  assign new_n12454_ = ~new_n12104_ | ~new_n12105_;
  assign new_n12455_ = ~new_n12237_ | ~new_n12453_;
  assign new_n12456_ = ~new_n1655_ | ~new_n11963_;
  assign new_n12457_ = ~pi021 | ~new_n11964_;
  assign new_n12458_ = ~new_n1655_ | ~new_n11963_;
  assign new_n12459_ = ~pi021 | ~new_n11964_;
  assign new_n12460_ = ~new_n12459_ | ~new_n12458_;
  assign new_n12461_ = ~new_n12106_ | ~new_n12107_;
  assign new_n12462_ = ~new_n12253_ | ~new_n12460_;
  assign new_n12463_ = ~new_n1656_ | ~new_n11966_;
  assign new_n12464_ = ~pi022 | ~new_n11967_;
  assign new_n12465_ = ~new_n1656_ | ~new_n11966_;
  assign new_n12466_ = ~pi022 | ~new_n11967_;
  assign new_n12467_ = ~new_n12466_ | ~new_n12465_;
  assign new_n12468_ = ~new_n12108_ | ~new_n12109_;
  assign new_n12469_ = ~new_n12251_ | ~new_n12467_;
  assign new_n12470_ = ~new_n1658_ | ~new_n11941_;
  assign new_n12471_ = ~pi032 | ~new_n11942_;
  assign new_n12472_ = ~pi683;
  assign new_n12473_ = ~pi193;
  assign po000 = new_n12629_ & new_n12625_;
  assign po018 = ~new_n12630_ | ~new_n12691_ | ~new_n12690_;
  assign new_n12476_ = ~new_n12763_;
  assign new_n12477_ = ~pi457;
  assign new_n12478_ = ~pi456;
  assign new_n12479_ = ~pi457 | ~new_n12763_;
  assign new_n12480_ = ~new_n12811_;
  assign new_n12481_ = ~new_n12810_;
  assign new_n12482_ = ~pi455;
  assign new_n12483_ = ~new_n12560_ | ~new_n12559_;
  assign new_n12484_ = ~new_n12809_;
  assign new_n12485_ = ~pi454;
  assign new_n12486_ = ~new_n12808_;
  assign new_n12487_ = ~pi453;
  assign new_n12488_ = ~new_n12568_ | ~new_n12567_;
  assign new_n12489_ = ~new_n12807_;
  assign new_n12490_ = ~pi452;
  assign new_n12491_ = ~new_n12806_;
  assign new_n12492_ = ~pi451;
  assign new_n12493_ = ~new_n12805_;
  assign new_n12494_ = ~pi450;
  assign new_n12495_ = ~new_n12580_ | ~new_n12579_;
  assign new_n12496_ = ~new_n12804_;
  assign new_n12497_ = ~pi449;
  assign new_n12498_ = ~pi448;
  assign new_n12499_ = ~new_n12803_;
  assign new_n12500_ = ~new_n12588_ | ~new_n12587_;
  assign new_n12501_ = ~new_n12820_;
  assign new_n12502_ = ~pi447;
  assign new_n12503_ = ~new_n12819_;
  assign new_n12504_ = ~pi446;
  assign new_n12505_ = ~new_n12818_;
  assign new_n12506_ = ~pi445;
  assign new_n12507_ = ~new_n12600_ | ~new_n12599_;
  assign new_n12508_ = ~new_n12817_;
  assign new_n12509_ = ~pi444;
  assign new_n12510_ = ~new_n12604_ | ~new_n12603_;
  assign new_n12511_ = ~new_n12816_;
  assign new_n12512_ = ~pi443;
  assign new_n12513_ = ~new_n12608_ | ~new_n12607_;
  assign new_n12514_ = ~new_n12815_;
  assign new_n12515_ = ~pi442;
  assign new_n12516_ = ~new_n12814_;
  assign new_n12517_ = ~pi441;
  assign new_n12518_ = ~new_n12813_;
  assign new_n12519_ = ~pi440;
  assign new_n12520_ = ~new_n12620_ | ~new_n12619_;
  assign new_n12521_ = ~new_n12812_;
  assign new_n12522_ = ~pi439;
  assign po019 = ~new_n12761_ | ~new_n12760_;
  assign po010 = ~new_n12637_ | ~new_n12636_;
  assign po011 = ~new_n12644_ | ~new_n12643_;
  assign po012 = ~new_n12651_ | ~new_n12650_;
  assign po013 = ~new_n12658_ | ~new_n12657_;
  assign po014 = ~new_n12665_ | ~new_n12664_;
  assign po015 = ~new_n12672_ | ~new_n12671_;
  assign po016 = ~new_n12679_ | ~new_n12678_;
  assign po017 = ~new_n12686_ | ~new_n12685_;
  assign po001 = ~new_n12703_ | ~new_n12702_;
  assign po002 = ~new_n12710_ | ~new_n12709_;
  assign po003 = ~new_n12717_ | ~new_n12716_;
  assign po004 = ~new_n12724_ | ~new_n12723_;
  assign po005 = ~new_n12731_ | ~new_n12730_;
  assign po006 = ~new_n12738_ | ~new_n12737_;
  assign po007 = ~new_n12745_ | ~new_n12744_;
  assign po008 = ~new_n12752_ | ~new_n12751_;
  assign po009 = ~new_n12759_ | ~new_n12758_;
  assign new_n12541_ = ~new_n12584_ | ~new_n12583_;
  assign new_n12542_ = ~new_n12576_ | ~new_n12575_;
  assign new_n12543_ = ~new_n12572_ | ~new_n12571_;
  assign new_n12544_ = ~new_n12564_ | ~new_n12563_;
  assign new_n12545_ = ~new_n12546_ | ~new_n12556_;
  assign new_n12546_ = ~new_n12811_ | ~new_n12554_;
  assign new_n12547_ = ~pi438;
  assign new_n12548_ = ~new_n12762_;
  assign new_n12549_ = ~new_n12616_ | ~new_n12615_;
  assign new_n12550_ = ~new_n12612_ | ~new_n12611_;
  assign new_n12551_ = ~new_n12596_ | ~new_n12595_;
  assign new_n12552_ = ~new_n12592_ | ~new_n12591_;
  assign new_n12553_ = ~new_n12546_;
  assign new_n12554_ = ~new_n12479_;
  assign new_n12555_ = ~new_n12480_ | ~new_n12479_;
  assign new_n12556_ = ~pi456 | ~new_n12555_;
  assign new_n12557_ = ~new_n12545_;
  assign new_n12558_ = new_n12810_ | pi455;
  assign new_n12559_ = ~new_n12558_ | ~new_n12545_;
  assign new_n12560_ = ~pi455 | ~new_n12810_;
  assign new_n12561_ = ~new_n12483_;
  assign new_n12562_ = ~new_n12561_ | ~new_n12485_;
  assign new_n12563_ = ~new_n12809_ | ~new_n12562_;
  assign new_n12564_ = ~pi454 | ~new_n12483_;
  assign new_n12565_ = ~new_n12544_;
  assign new_n12566_ = new_n12808_ | pi453;
  assign new_n12567_ = ~new_n12566_ | ~new_n12544_;
  assign new_n12568_ = ~pi453 | ~new_n12808_;
  assign new_n12569_ = ~new_n12488_;
  assign new_n12570_ = ~new_n12569_ | ~new_n12490_;
  assign new_n12571_ = ~new_n12807_ | ~new_n12570_;
  assign new_n12572_ = ~pi452 | ~new_n12488_;
  assign new_n12573_ = ~new_n12543_;
  assign new_n12574_ = new_n12806_ | pi451;
  assign new_n12575_ = ~new_n12574_ | ~new_n12543_;
  assign new_n12576_ = ~pi451 | ~new_n12806_;
  assign new_n12577_ = ~new_n12542_;
  assign new_n12578_ = new_n12805_ | pi450;
  assign new_n12579_ = ~new_n12578_ | ~new_n12542_;
  assign new_n12580_ = ~pi450 | ~new_n12805_;
  assign new_n12581_ = ~new_n12495_;
  assign new_n12582_ = ~new_n12581_ | ~new_n12497_;
  assign new_n12583_ = ~new_n12804_ | ~new_n12582_;
  assign new_n12584_ = ~pi449 | ~new_n12495_;
  assign new_n12585_ = ~new_n12541_;
  assign new_n12586_ = new_n12803_ | pi448;
  assign new_n12587_ = ~new_n12586_ | ~new_n12541_;
  assign new_n12588_ = ~new_n12803_ | ~pi448;
  assign new_n12589_ = ~new_n12500_;
  assign new_n12590_ = ~new_n12589_ | ~new_n12502_;
  assign new_n12591_ = ~new_n12820_ | ~new_n12590_;
  assign new_n12592_ = ~pi447 | ~new_n12500_;
  assign new_n12593_ = ~new_n12552_;
  assign new_n12594_ = new_n12819_ | pi446;
  assign new_n12595_ = ~new_n12594_ | ~new_n12552_;
  assign new_n12596_ = ~pi446 | ~new_n12819_;
  assign new_n12597_ = ~new_n12551_;
  assign new_n12598_ = new_n12818_ | pi445;
  assign new_n12599_ = ~new_n12598_ | ~new_n12551_;
  assign new_n12600_ = ~pi445 | ~new_n12818_;
  assign new_n12601_ = ~new_n12507_;
  assign new_n12602_ = ~new_n12601_ | ~new_n12509_;
  assign new_n12603_ = ~new_n12817_ | ~new_n12602_;
  assign new_n12604_ = ~pi444 | ~new_n12507_;
  assign new_n12605_ = ~new_n12510_;
  assign new_n12606_ = ~new_n12605_ | ~new_n12512_;
  assign new_n12607_ = ~new_n12816_ | ~new_n12606_;
  assign new_n12608_ = ~pi443 | ~new_n12510_;
  assign new_n12609_ = ~new_n12513_;
  assign new_n12610_ = ~new_n12609_ | ~new_n12515_;
  assign new_n12611_ = ~new_n12815_ | ~new_n12610_;
  assign new_n12612_ = ~pi442 | ~new_n12513_;
  assign new_n12613_ = ~new_n12550_;
  assign new_n12614_ = new_n12814_ | pi441;
  assign new_n12615_ = ~new_n12614_ | ~new_n12550_;
  assign new_n12616_ = ~pi441 | ~new_n12814_;
  assign new_n12617_ = ~new_n12549_;
  assign new_n12618_ = new_n12813_ | pi440;
  assign new_n12619_ = ~new_n12618_ | ~new_n12549_;
  assign new_n12620_ = ~pi440 | ~new_n12813_;
  assign new_n12621_ = ~new_n12520_;
  assign new_n12622_ = ~new_n12621_ | ~new_n12522_;
  assign new_n12623_ = ~new_n12812_ | ~new_n12622_;
  assign new_n12624_ = ~pi439 | ~new_n12520_;
  assign new_n12625_ = ~new_n12623_ | ~new_n12692_ | ~new_n12693_ | ~new_n12624_;
  assign new_n12626_ = ~pi439 | ~new_n12520_;
  assign new_n12627_ = ~new_n12626_ | ~new_n12521_;
  assign new_n12628_ = ~new_n12621_ | ~new_n12522_;
  assign new_n12629_ = ~new_n12696_ | ~new_n12628_ | ~new_n12627_;
  assign new_n12630_ = ~new_n12689_ | ~new_n12480_;
  assign new_n12631_ = ~pi448 | ~new_n12499_;
  assign new_n12632_ = ~new_n12803_ | ~new_n12498_;
  assign new_n12633_ = ~pi448 | ~new_n12499_;
  assign new_n12634_ = ~new_n12803_ | ~new_n12498_;
  assign new_n12635_ = ~new_n12634_ | ~new_n12633_;
  assign new_n12636_ = ~new_n12541_ | ~new_n12632_ | ~new_n12631_;
  assign new_n12637_ = ~new_n12585_ | ~new_n12635_;
  assign new_n12638_ = ~pi449 | ~new_n12495_;
  assign new_n12639_ = ~new_n12581_ | ~new_n12497_;
  assign new_n12640_ = ~pi449 | ~new_n12495_;
  assign new_n12641_ = ~new_n12581_ | ~new_n12497_;
  assign new_n12642_ = ~new_n12641_ | ~new_n12640_;
  assign new_n12643_ = ~new_n12496_ | ~new_n12639_ | ~new_n12638_;
  assign new_n12644_ = ~new_n12642_ | ~new_n12804_;
  assign new_n12645_ = ~pi450 | ~new_n12493_;
  assign new_n12646_ = ~new_n12805_ | ~new_n12494_;
  assign new_n12647_ = ~pi450 | ~new_n12493_;
  assign new_n12648_ = ~new_n12805_ | ~new_n12494_;
  assign new_n12649_ = ~new_n12648_ | ~new_n12647_;
  assign new_n12650_ = ~new_n12542_ | ~new_n12646_ | ~new_n12645_;
  assign new_n12651_ = ~new_n12577_ | ~new_n12649_;
  assign new_n12652_ = ~pi451 | ~new_n12491_;
  assign new_n12653_ = ~new_n12806_ | ~new_n12492_;
  assign new_n12654_ = ~pi451 | ~new_n12491_;
  assign new_n12655_ = ~new_n12806_ | ~new_n12492_;
  assign new_n12656_ = ~new_n12655_ | ~new_n12654_;
  assign new_n12657_ = ~new_n12543_ | ~new_n12653_ | ~new_n12652_;
  assign new_n12658_ = ~new_n12573_ | ~new_n12656_;
  assign new_n12659_ = ~pi452 | ~new_n12488_;
  assign new_n12660_ = ~new_n12569_ | ~new_n12490_;
  assign new_n12661_ = ~pi452 | ~new_n12488_;
  assign new_n12662_ = ~new_n12569_ | ~new_n12490_;
  assign new_n12663_ = ~new_n12662_ | ~new_n12661_;
  assign new_n12664_ = ~new_n12489_ | ~new_n12660_ | ~new_n12659_;
  assign new_n12665_ = ~new_n12663_ | ~new_n12807_;
  assign new_n12666_ = ~pi453 | ~new_n12486_;
  assign new_n12667_ = ~new_n12808_ | ~new_n12487_;
  assign new_n12668_ = ~pi453 | ~new_n12486_;
  assign new_n12669_ = ~new_n12808_ | ~new_n12487_;
  assign new_n12670_ = ~new_n12669_ | ~new_n12668_;
  assign new_n12671_ = ~new_n12544_ | ~new_n12667_ | ~new_n12666_;
  assign new_n12672_ = ~new_n12565_ | ~new_n12670_;
  assign new_n12673_ = ~pi454 | ~new_n12483_;
  assign new_n12674_ = ~new_n12561_ | ~new_n12485_;
  assign new_n12675_ = ~pi454 | ~new_n12483_;
  assign new_n12676_ = ~new_n12561_ | ~new_n12485_;
  assign new_n12677_ = ~new_n12676_ | ~new_n12675_;
  assign new_n12678_ = ~new_n12484_ | ~new_n12674_ | ~new_n12673_;
  assign new_n12679_ = ~new_n12677_ | ~new_n12809_;
  assign new_n12680_ = ~pi455 | ~new_n12481_;
  assign new_n12681_ = ~new_n12810_ | ~new_n12482_;
  assign new_n12682_ = ~pi455 | ~new_n12481_;
  assign new_n12683_ = ~new_n12810_ | ~new_n12482_;
  assign new_n12684_ = ~new_n12683_ | ~new_n12682_;
  assign new_n12685_ = ~new_n12545_ | ~new_n12681_ | ~new_n12680_;
  assign new_n12686_ = ~new_n12557_ | ~new_n12684_;
  assign new_n12687_ = ~pi456 | ~new_n12479_;
  assign new_n12688_ = ~new_n12554_ | ~new_n12478_;
  assign new_n12689_ = ~new_n12688_ | ~new_n12687_;
  assign new_n12690_ = ~new_n12478_ | ~new_n12811_ | ~new_n12479_;
  assign new_n12691_ = ~new_n12553_ | ~pi456;
  assign new_n12692_ = ~pi438 | ~new_n12548_;
  assign new_n12693_ = ~new_n12762_ | ~new_n12547_;
  assign new_n12694_ = ~pi438 | ~new_n12548_;
  assign new_n12695_ = ~new_n12762_ | ~new_n12547_;
  assign new_n12696_ = ~new_n12695_ | ~new_n12694_;
  assign new_n12697_ = ~pi439 | ~new_n12520_;
  assign new_n12698_ = ~new_n12621_ | ~new_n12522_;
  assign new_n12699_ = ~pi439 | ~new_n12520_;
  assign new_n12700_ = ~new_n12621_ | ~new_n12522_;
  assign new_n12701_ = ~new_n12700_ | ~new_n12699_;
  assign new_n12702_ = ~new_n12521_ | ~new_n12698_ | ~new_n12697_;
  assign new_n12703_ = ~new_n12701_ | ~new_n12812_;
  assign new_n12704_ = ~pi440 | ~new_n12518_;
  assign new_n12705_ = ~new_n12813_ | ~new_n12519_;
  assign new_n12706_ = ~pi440 | ~new_n12518_;
  assign new_n12707_ = ~new_n12813_ | ~new_n12519_;
  assign new_n12708_ = ~new_n12707_ | ~new_n12706_;
  assign new_n12709_ = ~new_n12549_ | ~new_n12705_ | ~new_n12704_;
  assign new_n12710_ = ~new_n12617_ | ~new_n12708_;
  assign new_n12711_ = ~pi441 | ~new_n12516_;
  assign new_n12712_ = ~new_n12814_ | ~new_n12517_;
  assign new_n12713_ = ~pi441 | ~new_n12516_;
  assign new_n12714_ = ~new_n12814_ | ~new_n12517_;
  assign new_n12715_ = ~new_n12714_ | ~new_n12713_;
  assign new_n12716_ = ~new_n12550_ | ~new_n12712_ | ~new_n12711_;
  assign new_n12717_ = ~new_n12613_ | ~new_n12715_;
  assign new_n12718_ = ~pi442 | ~new_n12513_;
  assign new_n12719_ = ~new_n12609_ | ~new_n12515_;
  assign new_n12720_ = ~pi442 | ~new_n12513_;
  assign new_n12721_ = ~new_n12609_ | ~new_n12515_;
  assign new_n12722_ = ~new_n12721_ | ~new_n12720_;
  assign new_n12723_ = ~new_n12514_ | ~new_n12719_ | ~new_n12718_;
  assign new_n12724_ = ~new_n12722_ | ~new_n12815_;
  assign new_n12725_ = ~pi443 | ~new_n12510_;
  assign new_n12726_ = ~new_n12605_ | ~new_n12512_;
  assign new_n12727_ = ~pi443 | ~new_n12510_;
  assign new_n12728_ = ~new_n12605_ | ~new_n12512_;
  assign new_n12729_ = ~new_n12728_ | ~new_n12727_;
  assign new_n12730_ = ~new_n12511_ | ~new_n12726_ | ~new_n12725_;
  assign new_n12731_ = ~new_n12729_ | ~new_n12816_;
  assign new_n12732_ = ~pi444 | ~new_n12507_;
  assign new_n12733_ = ~new_n12601_ | ~new_n12509_;
  assign new_n12734_ = ~pi444 | ~new_n12507_;
  assign new_n12735_ = ~new_n12601_ | ~new_n12509_;
  assign new_n12736_ = ~new_n12735_ | ~new_n12734_;
  assign new_n12737_ = ~new_n12508_ | ~new_n12733_ | ~new_n12732_;
  assign new_n12738_ = ~new_n12736_ | ~new_n12817_;
  assign new_n12739_ = ~pi445 | ~new_n12505_;
  assign new_n12740_ = ~new_n12818_ | ~new_n12506_;
  assign new_n12741_ = ~pi445 | ~new_n12505_;
  assign new_n12742_ = ~new_n12818_ | ~new_n12506_;
  assign new_n12743_ = ~new_n12742_ | ~new_n12741_;
  assign new_n12744_ = ~new_n12551_ | ~new_n12740_ | ~new_n12739_;
  assign new_n12745_ = ~new_n12597_ | ~new_n12743_;
  assign new_n12746_ = ~pi446 | ~new_n12503_;
  assign new_n12747_ = ~new_n12819_ | ~new_n12504_;
  assign new_n12748_ = ~pi446 | ~new_n12503_;
  assign new_n12749_ = ~new_n12819_ | ~new_n12504_;
  assign new_n12750_ = ~new_n12749_ | ~new_n12748_;
  assign new_n12751_ = ~new_n12552_ | ~new_n12747_ | ~new_n12746_;
  assign new_n12752_ = ~new_n12593_ | ~new_n12750_;
  assign new_n12753_ = ~pi447 | ~new_n12500_;
  assign new_n12754_ = ~new_n12589_ | ~new_n12502_;
  assign new_n12755_ = ~pi447 | ~new_n12500_;
  assign new_n12756_ = ~new_n12589_ | ~new_n12502_;
  assign new_n12757_ = ~new_n12756_ | ~new_n12755_;
  assign new_n12758_ = ~new_n12501_ | ~new_n12754_ | ~new_n12753_;
  assign new_n12759_ = ~new_n12757_ | ~new_n12820_;
  assign new_n12760_ = ~pi457 | ~new_n12476_;
  assign new_n12761_ = ~new_n12763_ | ~new_n12477_;
  assign new_n12762_ = ~new_n12930_ | ~new_n12934_;
  assign new_n12763_ = ~new_n12765_ | ~new_n12935_;
  assign new_n12764_ = ~pi702;
  assign new_n12765_ = ~pi702 | ~new_n12802_;
  assign new_n12766_ = ~pi211;
  assign new_n12767_ = ~pi700;
  assign new_n12768_ = ~pi210;
  assign new_n12769_ = ~pi699;
  assign new_n12770_ = ~pi209;
  assign new_n12771_ = ~pi698;
  assign new_n12772_ = ~pi208;
  assign new_n12773_ = ~pi697;
  assign new_n12774_ = ~pi207;
  assign new_n12775_ = ~pi696;
  assign new_n12776_ = ~pi206;
  assign new_n12777_ = ~pi695;
  assign new_n12778_ = ~pi205;
  assign new_n12779_ = ~pi694;
  assign new_n12780_ = ~pi204;
  assign new_n12781_ = ~pi693;
  assign new_n12782_ = ~pi203;
  assign new_n12783_ = ~pi692;
  assign new_n12784_ = ~pi202;
  assign new_n12785_ = ~pi691;
  assign new_n12786_ = ~pi201;
  assign new_n12787_ = ~pi690;
  assign new_n12788_ = ~pi200;
  assign new_n12789_ = ~pi689;
  assign new_n12790_ = ~pi199;
  assign new_n12791_ = ~pi688;
  assign new_n12792_ = ~pi198;
  assign new_n12793_ = ~pi687;
  assign new_n12794_ = ~pi197;
  assign new_n12795_ = ~pi686;
  assign new_n12796_ = ~pi196;
  assign new_n12797_ = ~pi685;
  assign new_n12798_ = ~pi195;
  assign new_n12799_ = ~pi684;
  assign new_n12800_ = ~pi194;
  assign new_n12801_ = ~new_n12925_ | ~new_n12924_;
  assign new_n12802_ = ~pi212;
  assign new_n12803_ = ~new_n12940_ | ~new_n12939_;
  assign new_n12804_ = ~new_n12945_ | ~new_n12944_;
  assign new_n12805_ = ~new_n12950_ | ~new_n12949_;
  assign new_n12806_ = ~new_n12955_ | ~new_n12954_;
  assign new_n12807_ = ~new_n12960_ | ~new_n12959_;
  assign new_n12808_ = ~new_n12965_ | ~new_n12964_;
  assign new_n12809_ = ~new_n12970_ | ~new_n12969_;
  assign new_n12810_ = ~new_n12975_ | ~new_n12974_;
  assign new_n12811_ = ~new_n12980_ | ~new_n12979_;
  assign new_n12812_ = ~new_n12990_ | ~new_n12989_;
  assign new_n12813_ = ~new_n12995_ | ~new_n12994_;
  assign new_n12814_ = ~new_n13000_ | ~new_n12999_;
  assign new_n12815_ = ~new_n13005_ | ~new_n13004_;
  assign new_n12816_ = ~new_n13010_ | ~new_n13009_;
  assign new_n12817_ = ~new_n13015_ | ~new_n13014_;
  assign new_n12818_ = ~new_n13020_ | ~new_n13019_;
  assign new_n12819_ = ~new_n13025_ | ~new_n13024_;
  assign new_n12820_ = ~new_n13030_ | ~new_n13029_;
  assign new_n12821_ = ~new_n12937_ | ~new_n12936_;
  assign new_n12822_ = ~new_n12942_ | ~new_n12941_;
  assign new_n12823_ = ~new_n12947_ | ~new_n12946_;
  assign new_n12824_ = ~new_n12952_ | ~new_n12951_;
  assign new_n12825_ = ~new_n12957_ | ~new_n12956_;
  assign new_n12826_ = ~new_n12962_ | ~new_n12961_;
  assign new_n12827_ = ~new_n12967_ | ~new_n12966_;
  assign new_n12828_ = ~new_n12972_ | ~new_n12971_;
  assign new_n12829_ = ~new_n12977_ | ~new_n12976_;
  assign new_n12830_ = ~new_n12987_ | ~new_n12986_;
  assign new_n12831_ = ~new_n12992_ | ~new_n12991_;
  assign new_n12832_ = ~new_n12997_ | ~new_n12996_;
  assign new_n12833_ = ~new_n13002_ | ~new_n13001_;
  assign new_n12834_ = ~new_n13007_ | ~new_n13006_;
  assign new_n12835_ = ~new_n13012_ | ~new_n13011_;
  assign new_n12836_ = ~new_n13017_ | ~new_n13016_;
  assign new_n12837_ = ~new_n13022_ | ~new_n13021_;
  assign new_n12838_ = ~new_n13027_ | ~new_n13026_;
  assign new_n12839_ = ~new_n12889_ | ~new_n12888_;
  assign new_n12840_ = ~new_n12885_ | ~new_n12884_;
  assign new_n12841_ = ~new_n12881_ | ~new_n12880_;
  assign new_n12842_ = ~new_n12877_ | ~new_n12876_;
  assign new_n12843_ = ~new_n12873_ | ~new_n12872_;
  assign new_n12844_ = ~new_n12869_ | ~new_n12868_;
  assign new_n12845_ = ~new_n12865_ | ~new_n12864_;
  assign new_n12846_ = ~new_n12861_ | ~new_n12860_;
  assign new_n12847_ = ~pi701;
  assign new_n12848_ = ~pi683;
  assign new_n12849_ = ~pi193;
  assign new_n12850_ = ~new_n12921_ | ~new_n12920_;
  assign new_n12851_ = ~new_n12917_ | ~new_n12916_;
  assign new_n12852_ = ~new_n12913_ | ~new_n12912_;
  assign new_n12853_ = ~new_n12909_ | ~new_n12908_;
  assign new_n12854_ = ~new_n12905_ | ~new_n12904_;
  assign new_n12855_ = ~new_n12901_ | ~new_n12900_;
  assign new_n12856_ = ~new_n12897_ | ~new_n12896_;
  assign new_n12857_ = ~new_n12893_ | ~new_n12892_;
  assign new_n12858_ = ~new_n12765_;
  assign new_n12859_ = ~new_n12858_ | ~new_n12766_;
  assign new_n12860_ = ~new_n12859_ | ~new_n12847_;
  assign new_n12861_ = ~pi211 | ~new_n12765_;
  assign new_n12862_ = ~new_n12846_;
  assign new_n12863_ = ~pi700 | ~new_n12768_;
  assign new_n12864_ = ~new_n12863_ | ~new_n12846_;
  assign new_n12865_ = ~pi210 | ~new_n12767_;
  assign new_n12866_ = ~new_n12845_;
  assign new_n12867_ = ~pi699 | ~new_n12770_;
  assign new_n12868_ = ~new_n12867_ | ~new_n12845_;
  assign new_n12869_ = ~pi209 | ~new_n12769_;
  assign new_n12870_ = ~new_n12844_;
  assign new_n12871_ = ~pi698 | ~new_n12772_;
  assign new_n12872_ = ~new_n12871_ | ~new_n12844_;
  assign new_n12873_ = ~pi208 | ~new_n12771_;
  assign new_n12874_ = ~new_n12843_;
  assign new_n12875_ = ~pi697 | ~new_n12774_;
  assign new_n12876_ = ~new_n12875_ | ~new_n12843_;
  assign new_n12877_ = ~pi207 | ~new_n12773_;
  assign new_n12878_ = ~new_n12842_;
  assign new_n12879_ = ~pi696 | ~new_n12776_;
  assign new_n12880_ = ~new_n12879_ | ~new_n12842_;
  assign new_n12881_ = ~pi206 | ~new_n12775_;
  assign new_n12882_ = ~new_n12841_;
  assign new_n12883_ = ~pi695 | ~new_n12778_;
  assign new_n12884_ = ~new_n12883_ | ~new_n12841_;
  assign new_n12885_ = ~pi205 | ~new_n12777_;
  assign new_n12886_ = ~new_n12840_;
  assign new_n12887_ = ~pi694 | ~new_n12780_;
  assign new_n12888_ = ~new_n12887_ | ~new_n12840_;
  assign new_n12889_ = ~pi204 | ~new_n12779_;
  assign new_n12890_ = ~new_n12839_;
  assign new_n12891_ = ~pi693 | ~new_n12782_;
  assign new_n12892_ = ~new_n12891_ | ~new_n12839_;
  assign new_n12893_ = ~pi203 | ~new_n12781_;
  assign new_n12894_ = ~new_n12857_;
  assign new_n12895_ = ~pi692 | ~new_n12784_;
  assign new_n12896_ = ~new_n12895_ | ~new_n12857_;
  assign new_n12897_ = ~pi202 | ~new_n12783_;
  assign new_n12898_ = ~new_n12856_;
  assign new_n12899_ = ~pi691 | ~new_n12786_;
  assign new_n12900_ = ~new_n12899_ | ~new_n12856_;
  assign new_n12901_ = ~pi201 | ~new_n12785_;
  assign new_n12902_ = ~new_n12855_;
  assign new_n12903_ = ~pi690 | ~new_n12788_;
  assign new_n12904_ = ~new_n12903_ | ~new_n12855_;
  assign new_n12905_ = ~pi200 | ~new_n12787_;
  assign new_n12906_ = ~new_n12854_;
  assign new_n12907_ = ~pi689 | ~new_n12790_;
  assign new_n12908_ = ~new_n12907_ | ~new_n12854_;
  assign new_n12909_ = ~pi199 | ~new_n12789_;
  assign new_n12910_ = ~new_n12853_;
  assign new_n12911_ = ~pi688 | ~new_n12792_;
  assign new_n12912_ = ~new_n12911_ | ~new_n12853_;
  assign new_n12913_ = ~pi198 | ~new_n12791_;
  assign new_n12914_ = ~new_n12852_;
  assign new_n12915_ = ~pi687 | ~new_n12794_;
  assign new_n12916_ = ~new_n12915_ | ~new_n12852_;
  assign new_n12917_ = ~pi197 | ~new_n12793_;
  assign new_n12918_ = ~new_n12851_;
  assign new_n12919_ = ~pi686 | ~new_n12796_;
  assign new_n12920_ = ~new_n12919_ | ~new_n12851_;
  assign new_n12921_ = ~pi196 | ~new_n12795_;
  assign new_n12922_ = ~new_n12850_;
  assign new_n12923_ = ~pi685 | ~new_n12798_;
  assign new_n12924_ = ~new_n12923_ | ~new_n12850_;
  assign new_n12925_ = ~pi195 | ~new_n12797_;
  assign new_n12926_ = ~new_n12801_;
  assign new_n12927_ = ~pi194 | ~new_n12799_;
  assign new_n12928_ = ~new_n12926_ | ~new_n12927_;
  assign new_n12929_ = ~pi684 | ~new_n12800_;
  assign new_n12930_ = ~new_n12928_ | ~new_n12929_ | ~new_n12985_;
  assign new_n12931_ = ~pi684 | ~new_n12800_;
  assign new_n12932_ = ~new_n12931_ | ~new_n12801_;
  assign new_n12933_ = ~pi194 | ~new_n12799_;
  assign new_n12934_ = ~new_n12981_ | ~new_n12932_ | ~new_n12933_ | ~new_n12982_;
  assign new_n12935_ = ~pi212 | ~new_n12764_;
  assign new_n12936_ = ~pi693 | ~new_n12782_;
  assign new_n12937_ = ~pi203 | ~new_n12781_;
  assign new_n12938_ = ~new_n12821_;
  assign new_n12939_ = ~new_n12890_ | ~new_n12938_;
  assign new_n12940_ = ~new_n12821_ | ~new_n12839_;
  assign new_n12941_ = ~pi694 | ~new_n12780_;
  assign new_n12942_ = ~pi204 | ~new_n12779_;
  assign new_n12943_ = ~new_n12822_;
  assign new_n12944_ = ~new_n12886_ | ~new_n12943_;
  assign new_n12945_ = ~new_n12822_ | ~new_n12840_;
  assign new_n12946_ = ~pi695 | ~new_n12778_;
  assign new_n12947_ = ~pi205 | ~new_n12777_;
  assign new_n12948_ = ~new_n12823_;
  assign new_n12949_ = ~new_n12882_ | ~new_n12948_;
  assign new_n12950_ = ~new_n12823_ | ~new_n12841_;
  assign new_n12951_ = ~pi696 | ~new_n12776_;
  assign new_n12952_ = ~pi206 | ~new_n12775_;
  assign new_n12953_ = ~new_n12824_;
  assign new_n12954_ = ~new_n12878_ | ~new_n12953_;
  assign new_n12955_ = ~new_n12824_ | ~new_n12842_;
  assign new_n12956_ = ~pi697 | ~new_n12774_;
  assign new_n12957_ = ~pi207 | ~new_n12773_;
  assign new_n12958_ = ~new_n12825_;
  assign new_n12959_ = ~new_n12874_ | ~new_n12958_;
  assign new_n12960_ = ~new_n12825_ | ~new_n12843_;
  assign new_n12961_ = ~pi698 | ~new_n12772_;
  assign new_n12962_ = ~pi208 | ~new_n12771_;
  assign new_n12963_ = ~new_n12826_;
  assign new_n12964_ = ~new_n12870_ | ~new_n12963_;
  assign new_n12965_ = ~new_n12826_ | ~new_n12844_;
  assign new_n12966_ = ~pi699 | ~new_n12770_;
  assign new_n12967_ = ~pi209 | ~new_n12769_;
  assign new_n12968_ = ~new_n12827_;
  assign new_n12969_ = ~new_n12866_ | ~new_n12968_;
  assign new_n12970_ = ~new_n12827_ | ~new_n12845_;
  assign new_n12971_ = ~pi700 | ~new_n12768_;
  assign new_n12972_ = ~pi210 | ~new_n12767_;
  assign new_n12973_ = ~new_n12828_;
  assign new_n12974_ = ~new_n12862_ | ~new_n12973_;
  assign new_n12975_ = ~new_n12828_ | ~new_n12846_;
  assign new_n12976_ = ~pi701 | ~new_n12766_;
  assign new_n12977_ = ~pi211 | ~new_n12847_;
  assign new_n12978_ = ~new_n12829_;
  assign new_n12979_ = ~new_n12978_ | ~new_n12858_;
  assign new_n12980_ = ~new_n12829_ | ~new_n12765_;
  assign new_n12981_ = ~pi683 | ~new_n12849_;
  assign new_n12982_ = ~pi193 | ~new_n12848_;
  assign new_n12983_ = ~pi683 | ~new_n12849_;
  assign new_n12984_ = ~pi193 | ~new_n12848_;
  assign new_n12985_ = ~new_n12984_ | ~new_n12983_;
  assign new_n12986_ = ~pi684 | ~new_n12800_;
  assign new_n12987_ = ~pi194 | ~new_n12799_;
  assign new_n12988_ = ~new_n12830_;
  assign new_n12989_ = ~new_n12988_ | ~new_n12926_;
  assign new_n12990_ = ~new_n12830_ | ~new_n12801_;
  assign new_n12991_ = ~pi685 | ~new_n12798_;
  assign new_n12992_ = ~pi195 | ~new_n12797_;
  assign new_n12993_ = ~new_n12831_;
  assign new_n12994_ = ~new_n12922_ | ~new_n12993_;
  assign new_n12995_ = ~new_n12831_ | ~new_n12850_;
  assign new_n12996_ = ~pi686 | ~new_n12796_;
  assign new_n12997_ = ~pi196 | ~new_n12795_;
  assign new_n12998_ = ~new_n12832_;
  assign new_n12999_ = ~new_n12918_ | ~new_n12998_;
  assign new_n13000_ = ~new_n12832_ | ~new_n12851_;
  assign new_n13001_ = ~pi687 | ~new_n12794_;
  assign new_n13002_ = ~pi197 | ~new_n12793_;
  assign new_n13003_ = ~new_n12833_;
  assign new_n13004_ = ~new_n12914_ | ~new_n13003_;
  assign new_n13005_ = ~new_n12833_ | ~new_n12852_;
  assign new_n13006_ = ~pi688 | ~new_n12792_;
  assign new_n13007_ = ~pi198 | ~new_n12791_;
  assign new_n13008_ = ~new_n12834_;
  assign new_n13009_ = ~new_n12910_ | ~new_n13008_;
  assign new_n13010_ = ~new_n12834_ | ~new_n12853_;
  assign new_n13011_ = ~pi689 | ~new_n12790_;
  assign new_n13012_ = ~pi199 | ~new_n12789_;
  assign new_n13013_ = ~new_n12835_;
  assign new_n13014_ = ~new_n12906_ | ~new_n13013_;
  assign new_n13015_ = ~new_n12835_ | ~new_n12854_;
  assign new_n13016_ = ~pi690 | ~new_n12788_;
  assign new_n13017_ = ~pi200 | ~new_n12787_;
  assign new_n13018_ = ~new_n12836_;
  assign new_n13019_ = ~new_n12902_ | ~new_n13018_;
  assign new_n13020_ = ~new_n12836_ | ~new_n12855_;
  assign new_n13021_ = ~pi691 | ~new_n12786_;
  assign new_n13022_ = ~pi201 | ~new_n12785_;
  assign new_n13023_ = ~new_n12837_;
  assign new_n13024_ = ~new_n12898_ | ~new_n13023_;
  assign new_n13025_ = ~new_n12837_ | ~new_n12856_;
  assign new_n13026_ = ~pi692 | ~new_n12784_;
  assign new_n13027_ = ~pi202 | ~new_n12783_;
  assign new_n13028_ = ~new_n12838_;
  assign new_n13029_ = ~new_n12894_ | ~new_n13028_;
  assign new_n13030_ = ~new_n12838_ | ~new_n12857_;
  assign new_n13031_ = ~pi438;
  assign new_n13032_ = ~pi269;
  assign new_n13033_ = new_n13130_ & pi267 & pi273;
  assign new_n13034_ = ~pi257;
  assign new_n13035_ = ~pi257 | ~pi269;
  assign new_n13036_ = ~pi260;
  assign new_n13037_ = ~pi260 | ~new_n13108_;
  assign new_n13038_ = ~pi248;
  assign new_n13039_ = ~pi248 | ~new_n13109_;
  assign new_n13040_ = ~pi274;
  assign new_n13041_ = ~pi274 | ~new_n13110_;
  assign new_n13042_ = ~pi266;
  assign new_n13043_ = ~pi256;
  assign new_n13044_ = ~pi266 | ~new_n13111_;
  assign new_n13045_ = ~new_n13112_ | ~pi256;
  assign new_n13046_ = ~pi270;
  assign new_n13047_ = ~pi270 | ~new_n13113_;
  assign new_n13048_ = ~pi251;
  assign new_n13049_ = ~pi251 | ~new_n13114_;
  assign new_n13050_ = ~pi263;
  assign new_n13051_ = ~pi263 | ~new_n13115_;
  assign new_n13052_ = ~pi253;
  assign new_n13053_ = ~pi253 | ~new_n13116_;
  assign new_n13054_ = ~pi272;
  assign new_n13055_ = ~pi272 | ~new_n13117_;
  assign new_n13056_ = ~pi246;
  assign new_n13057_ = ~pi246 | ~new_n13118_;
  assign new_n13058_ = ~pi261;
  assign new_n13059_ = ~pi261 | ~new_n13119_;
  assign new_n13060_ = ~pi259;
  assign new_n13061_ = ~pi259 | ~new_n13120_;
  assign new_n13062_ = ~pi249;
  assign new_n13063_ = ~pi249 | ~new_n13121_;
  assign new_n13064_ = ~pi268;
  assign new_n13065_ = ~pi268 | ~new_n13122_;
  assign new_n13066_ = ~pi254;
  assign new_n13067_ = ~pi254 | ~new_n13123_;
  assign new_n13068_ = ~pi264;
  assign new_n13069_ = ~pi264 | ~new_n13124_;
  assign new_n13070_ = ~pi252;
  assign new_n13071_ = ~pi252 | ~new_n13125_;
  assign new_n13072_ = ~pi271;
  assign new_n13073_ = ~pi271 | ~new_n13126_;
  assign new_n13074_ = ~pi258;
  assign new_n13075_ = ~pi258 | ~new_n13127_;
  assign new_n13076_ = ~pi262;
  assign new_n13077_ = ~pi262 | ~new_n13128_;
  assign new_n13078_ = ~pi247;
  assign new_n13079_ = ~pi247 | ~new_n13129_;
  assign new_n13080_ = ~pi267;
  assign new_n13081_ = ~pi273;
  assign new_n13082_ = ~new_n13133_ | ~new_n13132_;
  assign new_n13083_ = ~new_n13135_ | ~new_n13134_;
  assign new_n13084_ = ~new_n13137_ | ~new_n13136_;
  assign new_n13085_ = ~new_n13139_ | ~new_n13138_;
  assign new_n13086_ = ~new_n13141_ | ~new_n13140_;
  assign new_n13087_ = ~new_n13143_ | ~new_n13142_;
  assign new_n13088_ = ~new_n13145_ | ~new_n13144_;
  assign new_n13089_ = ~new_n13147_ | ~new_n13146_;
  assign new_n13090_ = ~new_n13149_ | ~new_n13148_;
  assign new_n13091_ = ~new_n13151_ | ~new_n13150_;
  assign new_n13092_ = ~new_n13153_ | ~new_n13152_;
  assign new_n13093_ = ~new_n13155_ | ~new_n13154_;
  assign new_n13094_ = ~new_n13157_ | ~new_n13156_;
  assign new_n13095_ = ~new_n13159_ | ~new_n13158_;
  assign new_n13096_ = ~new_n13161_ | ~new_n13160_;
  assign new_n13097_ = ~new_n13163_ | ~new_n13162_;
  assign new_n13098_ = ~new_n13165_ | ~new_n13164_;
  assign new_n13099_ = ~new_n13167_ | ~new_n13166_;
  assign new_n13100_ = ~new_n13169_ | ~new_n13168_;
  assign new_n13101_ = ~new_n13171_ | ~new_n13170_;
  assign new_n13102_ = ~new_n13173_ | ~new_n13172_;
  assign new_n13103_ = ~new_n13175_ | ~new_n13174_;
  assign new_n13104_ = ~new_n13177_ | ~new_n13176_;
  assign new_n13105_ = ~new_n13179_ | ~new_n13178_;
  assign new_n13106_ = ~new_n13181_ | ~new_n13180_;
  assign new_n13107_ = ~pi273 | ~new_n13130_;
  assign new_n13108_ = ~new_n13035_;
  assign new_n13109_ = ~new_n13037_;
  assign new_n13110_ = ~new_n13039_;
  assign new_n13111_ = ~new_n13041_;
  assign new_n13112_ = ~new_n13044_;
  assign new_n13113_ = ~new_n13045_;
  assign new_n13114_ = ~new_n13047_;
  assign new_n13115_ = ~new_n13049_;
  assign new_n13116_ = ~new_n13051_;
  assign new_n13117_ = ~new_n13053_;
  assign new_n13118_ = ~new_n13055_;
  assign new_n13119_ = ~new_n13057_;
  assign new_n13120_ = ~new_n13059_;
  assign new_n13121_ = ~new_n13061_;
  assign new_n13122_ = ~new_n13063_;
  assign new_n13123_ = ~new_n13065_;
  assign new_n13124_ = ~new_n13067_;
  assign new_n13125_ = ~new_n13069_;
  assign new_n13126_ = ~new_n13071_;
  assign new_n13127_ = ~new_n13073_;
  assign new_n13128_ = ~new_n13075_;
  assign new_n13129_ = ~new_n13077_;
  assign new_n13130_ = ~new_n13079_;
  assign new_n13131_ = ~new_n13107_;
  assign new_n13132_ = ~pi256 | ~new_n13044_;
  assign new_n13133_ = ~new_n13112_ | ~new_n13043_;
  assign new_n13134_ = ~pi266 | ~new_n13041_;
  assign new_n13135_ = ~new_n13111_ | ~new_n13042_;
  assign new_n13136_ = ~pi274 | ~new_n13039_;
  assign new_n13137_ = ~new_n13110_ | ~new_n13040_;
  assign new_n13138_ = ~pi248 | ~new_n13037_;
  assign new_n13139_ = ~new_n13109_ | ~new_n13038_;
  assign new_n13140_ = ~pi260 | ~new_n13035_;
  assign new_n13141_ = ~new_n13108_ | ~new_n13036_;
  assign new_n13142_ = ~pi257 | ~new_n13032_;
  assign new_n13143_ = ~pi269 | ~new_n13034_;
  assign new_n13144_ = ~pi267 | ~new_n13107_;
  assign new_n13145_ = ~new_n13131_ | ~new_n13080_;
  assign new_n13146_ = ~pi273 | ~new_n13079_;
  assign new_n13147_ = ~new_n13130_ | ~new_n13081_;
  assign new_n13148_ = ~pi247 | ~new_n13077_;
  assign new_n13149_ = ~new_n13129_ | ~new_n13078_;
  assign new_n13150_ = ~pi262 | ~new_n13075_;
  assign new_n13151_ = ~new_n13128_ | ~new_n13076_;
  assign new_n13152_ = ~pi258 | ~new_n13073_;
  assign new_n13153_ = ~new_n13127_ | ~new_n13074_;
  assign new_n13154_ = ~pi271 | ~new_n13071_;
  assign new_n13155_ = ~new_n13126_ | ~new_n13072_;
  assign new_n13156_ = ~pi252 | ~new_n13069_;
  assign new_n13157_ = ~new_n13125_ | ~new_n13070_;
  assign new_n13158_ = ~pi264 | ~new_n13067_;
  assign new_n13159_ = ~new_n13124_ | ~new_n13068_;
  assign new_n13160_ = ~pi254 | ~new_n13065_;
  assign new_n13161_ = ~new_n13123_ | ~new_n13066_;
  assign new_n13162_ = ~pi268 | ~new_n13063_;
  assign new_n13163_ = ~new_n13122_ | ~new_n13064_;
  assign new_n13164_ = ~pi249 | ~new_n13061_;
  assign new_n13165_ = ~new_n13121_ | ~new_n13062_;
  assign new_n13166_ = ~pi259 | ~new_n13059_;
  assign new_n13167_ = ~new_n13120_ | ~new_n13060_;
  assign new_n13168_ = ~pi261 | ~new_n13057_;
  assign new_n13169_ = ~new_n13119_ | ~new_n13058_;
  assign new_n13170_ = ~pi246 | ~new_n13055_;
  assign new_n13171_ = ~new_n13118_ | ~new_n13056_;
  assign new_n13172_ = ~pi272 | ~new_n13053_;
  assign new_n13173_ = ~new_n13117_ | ~new_n13054_;
  assign new_n13174_ = ~pi253 | ~new_n13051_;
  assign new_n13175_ = ~new_n13116_ | ~new_n13052_;
  assign new_n13176_ = ~pi263 | ~new_n13049_;
  assign new_n13177_ = ~new_n13115_ | ~new_n13050_;
  assign new_n13178_ = ~pi251 | ~new_n13047_;
  assign new_n13179_ = ~new_n13114_ | ~new_n13048_;
  assign new_n13180_ = ~pi270 | ~new_n13045_;
  assign new_n13181_ = ~new_n13113_ | ~new_n13046_;
  assign new_n13182_ = new_n13273_ & new_n13272_;
  assign new_n13183_ = new_n13274_ & new_n13275_;
  assign new_n13184_ = new_n13291_ & new_n13290_;
  assign new_n13185_ = new_n13333_ & new_n13332_;
  assign new_n13186_ = new_n13342_ & new_n13341_;
  assign new_n13187_ = new_n13360_ & new_n13359_;
  assign new_n13188_ = new_n13396_ & new_n13393_;
  assign new_n13189_ = new_n13389_ & new_n13386_;
  assign new_n13190_ = new_n13380_ & new_n13377_;
  assign new_n13191_ = new_n13374_ & new_n13370_;
  assign new_n13192_ = new_n13329_ & new_n13326_;
  assign new_n13193_ = new_n13321_ & new_n13318_;
  assign new_n13194_ = new_n13307_ & new_n13304_;
  assign new_n13195_ = ~pi167;
  assign new_n13196_ = ~new_n2402_;
  assign new_n13197_ = ~new_n2405_;
  assign new_n13198_ = ~new_n2402_ | ~pi167;
  assign new_n13199_ = ~pi168;
  assign new_n13200_ = ~pi165;
  assign new_n13201_ = ~new_n2396_;
  assign new_n13202_ = ~new_n2399_;
  assign new_n13203_ = ~pi163;
  assign new_n13204_ = ~new_n2390_;
  assign new_n13205_ = ~pi161;
  assign new_n13206_ = ~new_n2381_;
  assign new_n13207_ = ~new_n2381_ | ~pi161;
  assign new_n13208_ = ~pi164;
  assign new_n13209_ = ~new_n2393_;
  assign new_n13210_ = ~new_n2396_ | ~pi165;
  assign new_n13211_ = ~pi166;
  assign new_n13212_ = ~pi169;
  assign new_n13213_ = ~new_n2408_;
  assign new_n13214_ = ~new_n2411_;
  assign new_n13215_ = ~pi170;
  assign new_n13216_ = ~new_n13227_ | ~new_n13299_;
  assign new_n13217_ = ~new_n13287_ | ~new_n13288_ | ~new_n13286_;
  assign new_n13218_ = ~new_n13276_ | ~new_n13277_;
  assign new_n13219_ = ~pi162 | ~new_n2387_;
  assign new_n13220_ = ~new_n13313_ | ~new_n13314_ | ~new_n13312_;
  assign new_n13221_ = ~new_n13310_ | ~new_n13309_;
  assign new_n13222_ = ~pi177;
  assign new_n13223_ = ~new_n2432_;
  assign new_n13224_ = ~new_n2435_;
  assign new_n13225_ = ~new_n2432_ | ~pi177;
  assign new_n13226_ = ~pi178;
  assign new_n13227_ = ~new_n2408_ | ~pi169;
  assign new_n13228_ = ~pi171;
  assign new_n13229_ = ~new_n2414_;
  assign new_n13230_ = ~pi173;
  assign new_n13231_ = ~new_n2420_;
  assign new_n13232_ = ~pi172;
  assign new_n13233_ = ~new_n2417_;
  assign new_n13234_ = ~new_n2417_ | ~pi172;
  assign new_n13235_ = ~pi174;
  assign new_n13236_ = ~new_n2423_;
  assign new_n13237_ = ~pi175;
  assign new_n13238_ = ~new_n2426_;
  assign new_n13239_ = ~pi176;
  assign new_n13240_ = ~new_n2429_;
  assign new_n13241_ = ~pi179;
  assign new_n13242_ = ~new_n2438_;
  assign new_n13243_ = ~new_n13365_ | ~new_n13364_ | ~new_n13363_;
  assign new_n13244_ = ~new_n13357_ | ~new_n13356_;
  assign new_n13245_ = ~new_n13234_ | ~new_n13382_;
  assign new_n13246_ = ~new_n13437_ | ~new_n13436_;
  assign new_n13247_ = ~new_n13486_ | ~new_n13485_;
  assign new_n13248_ = ~new_n13409_ | ~new_n13408_;
  assign new_n13249_ = ~new_n13414_ | ~new_n13413_;
  assign new_n13250_ = ~new_n13421_ | ~new_n13420_;
  assign new_n13251_ = ~new_n13428_ | ~new_n13427_;
  assign new_n13252_ = ~new_n13433_ | ~new_n13432_;
  assign new_n13253_ = ~new_n13449_ | ~new_n13448_;
  assign new_n13254_ = ~new_n13456_ | ~new_n13455_;
  assign new_n13255_ = ~new_n13463_ | ~new_n13462_;
  assign new_n13256_ = ~new_n13470_ | ~new_n13469_;
  assign new_n13257_ = ~new_n13477_ | ~new_n13476_;
  assign new_n13258_ = ~new_n13482_ | ~new_n13481_;
  assign new_n13259_ = ~new_n13296_ | ~new_n13295_ | ~new_n13294_;
  assign new_n13260_ = ~new_n13311_ | ~new_n13323_;
  assign new_n13261_ = ~new_n13219_ | ~new_n13330_;
  assign new_n13262_ = ~new_n2379_;
  assign new_n13263_ = ~pi180;
  assign new_n13264_ = ~new_n13353_ | ~new_n13352_;
  assign new_n13265_ = ~new_n13349_ | ~new_n13348_;
  assign new_n13266_ = ~new_n13339_ | ~new_n13338_;
  assign new_n13267_ = ~new_n13210_;
  assign new_n13268_ = ~pi170 | ~new_n2411_;
  assign new_n13269_ = ~new_n2420_ | ~pi173;
  assign new_n13270_ = ~new_n13234_;
  assign new_n13271_ = ~new_n13227_;
  assign new_n13272_ = new_n2399_ | pi166;
  assign new_n13273_ = new_n2396_ | pi165;
  assign new_n13274_ = pi164 | new_n2393_;
  assign new_n13275_ = pi163 | new_n2390_;
  assign new_n13276_ = ~new_n13207_;
  assign new_n13277_ = pi162 | new_n2387_;
  assign new_n13278_ = ~new_n13218_;
  assign new_n13279_ = ~new_n13219_;
  assign new_n13280_ = ~new_n13218_ | ~new_n13219_;
  assign new_n13281_ = ~new_n13274_ | ~pi163 | ~new_n2390_;
  assign new_n13282_ = ~new_n13183_ | ~new_n13280_;
  assign new_n13283_ = ~new_n2393_ | ~pi164;
  assign new_n13284_ = ~new_n13282_ | ~new_n13283_ | ~new_n13281_;
  assign new_n13285_ = ~new_n13211_ | ~new_n13210_;
  assign new_n13286_ = ~new_n2399_ | ~new_n13285_;
  assign new_n13287_ = ~new_n13182_ | ~new_n13284_;
  assign new_n13288_ = ~pi166 | ~new_n13267_;
  assign new_n13289_ = ~new_n13217_;
  assign new_n13290_ = new_n2405_ | pi168;
  assign new_n13291_ = new_n2402_ | pi167;
  assign new_n13292_ = ~new_n13198_;
  assign new_n13293_ = ~new_n13199_ | ~new_n13198_;
  assign new_n13294_ = ~new_n2405_ | ~new_n13293_;
  assign new_n13295_ = ~pi168 | ~new_n13292_;
  assign new_n13296_ = ~new_n13184_ | ~new_n13217_;
  assign new_n13297_ = ~new_n13259_;
  assign new_n13298_ = pi169 | new_n2408_;
  assign new_n13299_ = ~new_n13298_ | ~new_n13259_;
  assign new_n13300_ = ~new_n13216_;
  assign new_n13301_ = new_n2411_ | pi170;
  assign new_n13302_ = pi167 | new_n2402_;
  assign new_n13303_ = ~new_n13302_ | ~new_n13217_;
  assign new_n13304_ = ~new_n13415_ | ~new_n13303_ | ~new_n13198_ | ~new_n13416_;
  assign new_n13305_ = ~new_n13289_ | ~new_n13198_;
  assign new_n13306_ = ~pi168 | ~new_n2405_;
  assign new_n13307_ = ~new_n13305_ | ~new_n13306_ | ~new_n13184_;
  assign new_n13308_ = new_n2402_ | pi167;
  assign new_n13309_ = ~new_n13279_ | ~new_n13275_;
  assign new_n13310_ = ~new_n2390_ | ~pi163;
  assign new_n13311_ = ~new_n13221_;
  assign new_n13312_ = ~new_n13278_ | ~new_n13183_;
  assign new_n13313_ = ~new_n13221_ | ~new_n13274_;
  assign new_n13314_ = ~new_n2393_ | ~pi164;
  assign new_n13315_ = ~new_n13220_;
  assign new_n13316_ = pi165 | new_n2396_;
  assign new_n13317_ = ~new_n13316_ | ~new_n13220_;
  assign new_n13318_ = ~new_n13422_ | ~new_n13317_ | ~new_n13210_ | ~new_n13423_;
  assign new_n13319_ = ~new_n13315_ | ~new_n13210_;
  assign new_n13320_ = ~pi166 | ~new_n2399_;
  assign new_n13321_ = ~new_n13319_ | ~new_n13320_ | ~new_n13182_;
  assign new_n13322_ = new_n2396_ | pi165;
  assign new_n13323_ = ~new_n13278_ | ~new_n13275_;
  assign new_n13324_ = ~new_n13260_;
  assign new_n13325_ = ~new_n2393_ | ~pi164;
  assign new_n13326_ = ~new_n13218_ | ~new_n13434_ | ~new_n13435_ | ~new_n13219_;
  assign new_n13327_ = ~new_n13219_ | ~new_n13218_;
  assign new_n13328_ = ~new_n2390_ | ~pi163;
  assign new_n13329_ = ~new_n13327_ | ~new_n13328_ | ~new_n13275_;
  assign new_n13330_ = pi162 | new_n2387_;
  assign new_n13331_ = ~new_n13261_;
  assign new_n13332_ = new_n2411_ | pi170;
  assign new_n13333_ = new_n2414_ | pi171;
  assign new_n13334_ = ~new_n13271_ | ~new_n13185_;
  assign new_n13335_ = ~new_n2414_ | ~pi171;
  assign new_n13336_ = ~new_n13334_ | ~new_n13335_ | ~new_n13268_;
  assign new_n13337_ = pi171 | new_n2414_;
  assign new_n13338_ = ~new_n13259_ | ~new_n13298_ | ~new_n13185_;
  assign new_n13339_ = ~new_n13337_ | ~new_n13336_;
  assign new_n13340_ = ~new_n13266_;
  assign new_n13341_ = new_n2423_ | pi174;
  assign new_n13342_ = new_n2420_ | pi173;
  assign new_n13343_ = ~new_n13270_ | ~new_n13186_;
  assign new_n13344_ = ~new_n2423_ | ~pi174;
  assign new_n13345_ = ~new_n13343_ | ~new_n13344_ | ~new_n13269_;
  assign new_n13346_ = pi172 | new_n2417_;
  assign new_n13347_ = pi174 | new_n2423_;
  assign new_n13348_ = ~new_n13266_ | ~new_n13346_ | ~new_n13186_;
  assign new_n13349_ = ~new_n13347_ | ~new_n13345_;
  assign new_n13350_ = ~new_n13265_;
  assign new_n13351_ = pi175 | new_n2426_;
  assign new_n13352_ = ~new_n13351_ | ~new_n13265_;
  assign new_n13353_ = ~new_n2426_ | ~pi175;
  assign new_n13354_ = ~new_n13264_;
  assign new_n13355_ = pi176 | new_n2429_;
  assign new_n13356_ = ~new_n13355_ | ~new_n13264_;
  assign new_n13357_ = ~new_n2429_ | ~pi176;
  assign new_n13358_ = ~new_n13244_;
  assign new_n13359_ = new_n2435_ | pi178;
  assign new_n13360_ = new_n2432_ | pi177;
  assign new_n13361_ = ~new_n13225_;
  assign new_n13362_ = ~new_n13226_ | ~new_n13225_;
  assign new_n13363_ = ~new_n2435_ | ~new_n13362_;
  assign new_n13364_ = ~pi178 | ~new_n13361_;
  assign new_n13365_ = ~new_n13187_ | ~new_n13244_;
  assign new_n13366_ = ~new_n13243_;
  assign new_n13367_ = pi179 | new_n2438_;
  assign new_n13368_ = ~new_n13367_ | ~new_n13243_;
  assign new_n13369_ = ~new_n2438_ | ~pi179;
  assign new_n13370_ = ~new_n13438_ | ~new_n13368_ | ~new_n13369_ | ~new_n13439_;
  assign new_n13371_ = ~new_n2438_ | ~pi179;
  assign new_n13372_ = ~new_n13366_ | ~new_n13371_;
  assign new_n13373_ = new_n2438_ | pi179;
  assign new_n13374_ = ~new_n13372_ | ~new_n13373_ | ~new_n13442_;
  assign new_n13375_ = pi177 | new_n2432_;
  assign new_n13376_ = ~new_n13375_ | ~new_n13244_;
  assign new_n13377_ = ~new_n13450_ | ~new_n13376_ | ~new_n13225_ | ~new_n13451_;
  assign new_n13378_ = ~new_n13358_ | ~new_n13225_;
  assign new_n13379_ = ~pi178 | ~new_n2435_;
  assign new_n13380_ = ~new_n13378_ | ~new_n13379_ | ~new_n13187_;
  assign new_n13381_ = new_n2432_ | pi177;
  assign new_n13382_ = ~new_n13346_ | ~new_n13266_;
  assign new_n13383_ = ~new_n13245_;
  assign new_n13384_ = pi173 | new_n2420_;
  assign new_n13385_ = ~new_n13384_ | ~new_n13245_;
  assign new_n13386_ = ~new_n13471_ | ~new_n13385_ | ~new_n13269_ | ~new_n13472_;
  assign new_n13387_ = ~new_n13383_ | ~new_n13269_;
  assign new_n13388_ = ~new_n2423_ | ~pi174;
  assign new_n13389_ = ~new_n13387_ | ~new_n13388_ | ~new_n13186_;
  assign new_n13390_ = new_n2420_ | pi173;
  assign new_n13391_ = pi170 | new_n2411_;
  assign new_n13392_ = ~new_n13391_ | ~new_n13216_;
  assign new_n13393_ = ~new_n13483_ | ~new_n13392_ | ~new_n13268_ | ~new_n13484_;
  assign new_n13394_ = ~new_n13300_ | ~new_n13268_;
  assign new_n13395_ = ~new_n2414_ | ~pi171;
  assign new_n13396_ = ~new_n13394_ | ~new_n13395_ | ~new_n13185_;
  assign new_n13397_ = ~new_n13301_ | ~new_n13268_;
  assign new_n13398_ = ~new_n13298_ | ~new_n13227_;
  assign new_n13399_ = ~new_n13308_ | ~new_n13198_;
  assign new_n13400_ = ~new_n13322_ | ~new_n13210_;
  assign new_n13401_ = ~new_n13325_ | ~new_n13274_;
  assign new_n13402_ = ~new_n13381_ | ~new_n13225_;
  assign new_n13403_ = ~new_n13390_ | ~new_n13269_;
  assign new_n13404_ = ~new_n13346_ | ~new_n13234_;
  assign new_n13405_ = ~new_n2411_ | ~new_n13215_;
  assign new_n13406_ = ~pi170 | ~new_n13214_;
  assign new_n13407_ = ~new_n13406_ | ~new_n13405_;
  assign new_n13408_ = ~new_n13397_ | ~new_n13216_;
  assign new_n13409_ = ~new_n13407_ | ~new_n13300_;
  assign new_n13410_ = ~new_n2408_ | ~new_n13212_;
  assign new_n13411_ = ~pi169 | ~new_n13213_;
  assign new_n13412_ = ~new_n13411_ | ~new_n13410_;
  assign new_n13413_ = ~new_n13398_ | ~new_n13259_;
  assign new_n13414_ = ~new_n13297_ | ~new_n13412_;
  assign new_n13415_ = ~new_n2405_ | ~new_n13199_;
  assign new_n13416_ = ~pi168 | ~new_n13197_;
  assign new_n13417_ = ~new_n2402_ | ~new_n13195_;
  assign new_n13418_ = ~pi167 | ~new_n13196_;
  assign new_n13419_ = ~new_n13418_ | ~new_n13417_;
  assign new_n13420_ = ~new_n13399_ | ~new_n13217_;
  assign new_n13421_ = ~new_n13419_ | ~new_n13289_;
  assign new_n13422_ = ~new_n2399_ | ~new_n13211_;
  assign new_n13423_ = ~pi166 | ~new_n13202_;
  assign new_n13424_ = ~new_n2396_ | ~new_n13200_;
  assign new_n13425_ = ~pi165 | ~new_n13201_;
  assign new_n13426_ = ~new_n13425_ | ~new_n13424_;
  assign new_n13427_ = ~new_n13400_ | ~new_n13220_;
  assign new_n13428_ = ~new_n13426_ | ~new_n13315_;
  assign new_n13429_ = ~new_n2393_ | ~new_n13208_;
  assign new_n13430_ = ~pi164 | ~new_n13209_;
  assign new_n13431_ = ~new_n13430_ | ~new_n13429_;
  assign new_n13432_ = ~new_n13401_ | ~new_n13260_;
  assign new_n13433_ = ~new_n13324_ | ~new_n13431_;
  assign new_n13434_ = ~new_n2390_ | ~new_n13203_;
  assign new_n13435_ = ~pi163 | ~new_n13204_;
  assign new_n13436_ = ~new_n13276_ | ~new_n13261_;
  assign new_n13437_ = ~new_n13331_ | ~new_n13207_;
  assign new_n13438_ = ~new_n2379_ | ~new_n13263_;
  assign new_n13439_ = ~pi180 | ~new_n13262_;
  assign new_n13440_ = ~new_n2379_ | ~new_n13263_;
  assign new_n13441_ = ~pi180 | ~new_n13262_;
  assign new_n13442_ = ~new_n13441_ | ~new_n13440_;
  assign new_n13443_ = ~new_n2438_ | ~new_n13241_;
  assign new_n13444_ = ~pi179 | ~new_n13242_;
  assign new_n13445_ = ~new_n2438_ | ~new_n13241_;
  assign new_n13446_ = ~pi179 | ~new_n13242_;
  assign new_n13447_ = ~new_n13446_ | ~new_n13445_;
  assign new_n13448_ = ~new_n13243_ | ~new_n13444_ | ~new_n13443_;
  assign new_n13449_ = ~new_n13447_ | ~new_n13366_;
  assign new_n13450_ = ~new_n2435_ | ~new_n13226_;
  assign new_n13451_ = ~pi178 | ~new_n13224_;
  assign new_n13452_ = ~new_n2432_ | ~new_n13222_;
  assign new_n13453_ = ~pi177 | ~new_n13223_;
  assign new_n13454_ = ~new_n13453_ | ~new_n13452_;
  assign new_n13455_ = ~new_n13402_ | ~new_n13244_;
  assign new_n13456_ = ~new_n13454_ | ~new_n13358_;
  assign new_n13457_ = ~new_n2429_ | ~new_n13239_;
  assign new_n13458_ = ~pi176 | ~new_n13240_;
  assign new_n13459_ = ~new_n2429_ | ~new_n13239_;
  assign new_n13460_ = ~pi176 | ~new_n13240_;
  assign new_n13461_ = ~new_n13460_ | ~new_n13459_;
  assign new_n13462_ = ~new_n13264_ | ~new_n13458_ | ~new_n13457_;
  assign new_n13463_ = ~new_n13354_ | ~new_n13461_;
  assign new_n13464_ = ~new_n2426_ | ~new_n13237_;
  assign new_n13465_ = ~pi175 | ~new_n13238_;
  assign new_n13466_ = ~new_n2426_ | ~new_n13237_;
  assign new_n13467_ = ~pi175 | ~new_n13238_;
  assign new_n13468_ = ~new_n13467_ | ~new_n13466_;
  assign new_n13469_ = ~new_n13265_ | ~new_n13465_ | ~new_n13464_;
  assign new_n13470_ = ~new_n13350_ | ~new_n13468_;
  assign new_n13471_ = ~new_n2423_ | ~new_n13235_;
  assign new_n13472_ = ~pi174 | ~new_n13236_;
  assign new_n13473_ = ~new_n2420_ | ~new_n13230_;
  assign new_n13474_ = ~pi173 | ~new_n13231_;
  assign new_n13475_ = ~new_n13474_ | ~new_n13473_;
  assign new_n13476_ = ~new_n13403_ | ~new_n13245_;
  assign new_n13477_ = ~new_n13475_ | ~new_n13383_;
  assign new_n13478_ = ~new_n2417_ | ~new_n13232_;
  assign new_n13479_ = ~pi172 | ~new_n13233_;
  assign new_n13480_ = ~new_n13479_ | ~new_n13478_;
  assign new_n13481_ = ~new_n13404_ | ~new_n13266_;
  assign new_n13482_ = ~new_n13340_ | ~new_n13480_;
  assign new_n13483_ = ~new_n2414_ | ~new_n13228_;
  assign new_n13484_ = ~pi171 | ~new_n13229_;
  assign new_n13485_ = ~new_n2381_ | ~new_n13205_;
  assign new_n13486_ = ~pi161 | ~new_n13206_;
  assign new_n13487_ = new_n13708_ & new_n13519_;
  assign new_n13488_ = new_n13706_ & new_n13673_;
  assign new_n13489_ = new_n13705_ & new_n13516_;
  assign new_n13490_ = new_n13704_ & new_n13517_;
  assign new_n13491_ = new_n13702_ & new_n13676_;
  assign new_n13492_ = new_n13701_ & new_n13515_;
  assign new_n13493_ = new_n13700_ & new_n13678_;
  assign new_n13494_ = new_n13698_ & new_n13679_;
  assign new_n13495_ = new_n13697_ & new_n13653_;
  assign new_n13496_ = new_n13696_ & new_n13681_;
  assign new_n13497_ = new_n13694_ & new_n13682_;
  assign new_n13498_ = new_n13693_ & new_n13650_;
  assign new_n13499_ = new_n13692_ & new_n13648_;
  assign new_n13500_ = new_n13690_ & new_n13685_;
  assign new_n13501_ = new_n13689_ & new_n13514_;
  assign new_n13502_ = new_n13688_ & new_n13508_;
  assign new_n13503_ = new_n13671_ & new_n13661_;
  assign new_n13504_ = new_n13670_ & new_n13510_;
  assign new_n13505_ = new_n13669_ & new_n13511_;
  assign new_n13506_ = new_n13667_ & new_n13664_;
  assign new_n13507_ = new_n13666_ & new_n13509_;
  assign new_n13508_ = pi035 | pi034 | pi033;
  assign new_n13509_ = ~new_n13524_ | ~new_n13525_ | ~new_n13711_;
  assign new_n13510_ = ~new_n13526_ | ~new_n13711_;
  assign new_n13511_ = ~new_n13527_ | ~new_n13662_;
  assign new_n13512_ = ~pi040;
  assign new_n13513_ = ~pi036;
  assign new_n13514_ = ~new_n13537_ | ~new_n13532_;
  assign new_n13515_ = ~new_n13610_ | ~new_n13608_ | ~new_n13609_ | ~new_n13611_;
  assign new_n13516_ = ~new_n13637_ | ~new_n13665_;
  assign new_n13517_ = ~new_n13638_ | ~new_n13674_;
  assign new_n13518_ = ~pi048;
  assign new_n13519_ = ~new_n13639_ | ~new_n13665_;
  assign new_n13520_ = ~pi044;
  assign new_n13521_ = ~new_n13728_ | ~new_n13727_;
  assign new_n13522_ = ~new_n13718_ | ~new_n13717_;
  assign new_n13523_ = ~new_n13722_ | ~new_n13721_;
  assign new_n13524_ = ~pi037 & ~pi039 & ~pi038 & ~pi036;
  assign new_n13525_ = ~pi040 & ~pi041;
  assign new_n13526_ = ~pi036 & ~pi037;
  assign new_n13527_ = ~pi038 & ~pi039;
  assign new_n13528_ = ~pi044 & ~pi046 & ~pi045 & ~pi043;
  assign new_n13529_ = ~pi048 & ~pi050 & ~pi049 & ~pi047;
  assign new_n13530_ = ~pi052 & ~pi033 & ~pi034 & ~pi051;
  assign new_n13531_ = ~pi054 & ~pi055 & ~pi053;
  assign new_n13532_ = new_n13530_ & new_n13528_ & new_n13529_ & new_n13531_;
  assign new_n13533_ = ~pi057 & ~pi059 & ~pi058 & ~pi056;
  assign new_n13534_ = ~pi061 & ~pi035 & ~pi062 & ~pi060;
  assign new_n13535_ = ~pi037 & ~pi039 & ~pi038 & ~pi036;
  assign new_n13536_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13537_ = new_n13535_ & new_n13533_ & new_n13534_ & new_n13536_;
  assign new_n13538_ = ~pi044 & ~pi046 & ~pi045 & ~pi043;
  assign new_n13539_ = ~pi048 & ~pi050 & ~pi049 & ~pi047;
  assign new_n13540_ = ~pi052 & ~pi033 & ~pi034 & ~pi051;
  assign new_n13541_ = ~pi054 & ~pi055 & ~pi053;
  assign new_n13542_ = new_n13540_ & new_n13538_ & new_n13539_ & new_n13541_;
  assign new_n13543_ = ~pi057 & ~pi059 & ~pi058 & ~pi056;
  assign new_n13544_ = ~pi061 & ~pi035 & ~pi060;
  assign new_n13545_ = ~pi037 & ~pi039 & ~pi038 & ~pi036;
  assign new_n13546_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13547_ = new_n13545_ & new_n13543_ & new_n13544_ & new_n13546_;
  assign new_n13548_ = ~pi044 & ~pi046 & ~pi045 & ~pi043;
  assign new_n13549_ = ~pi048 & ~pi049 & ~pi047;
  assign new_n13550_ = ~pi051 & ~pi034 & ~pi052 & ~pi050;
  assign new_n13551_ = ~pi053 & ~pi054 & ~pi033;
  assign new_n13552_ = new_n13550_ & new_n13548_ & new_n13549_ & new_n13551_;
  assign new_n13553_ = ~pi056 & ~pi058 & ~pi057 & ~pi055;
  assign new_n13554_ = ~pi060 & ~pi035 & ~pi059;
  assign new_n13555_ = ~pi037 & ~pi039 & ~pi038 & ~pi036;
  assign new_n13556_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13557_ = new_n13555_ & new_n13553_ & new_n13554_ & new_n13556_;
  assign new_n13558_ = ~pi044 & ~pi046 & ~pi045 & ~pi043;
  assign new_n13559_ = ~pi048 & ~pi049 & ~pi047;
  assign new_n13560_ = ~pi051 & ~pi034 & ~pi052 & ~pi050;
  assign new_n13561_ = ~pi053 & ~pi054 & ~pi033;
  assign new_n13562_ = new_n13560_ & new_n13558_ & new_n13559_ & new_n13561_;
  assign new_n13563_ = ~pi056 & ~pi058 & ~pi057 & ~pi055;
  assign new_n13564_ = ~pi035 & ~pi036 & ~pi059;
  assign new_n13565_ = ~pi038 & ~pi039 & ~pi037;
  assign new_n13566_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13567_ = new_n13565_ & new_n13563_ & new_n13564_ & new_n13566_;
  assign new_n13568_ = ~pi044 & ~pi046 & ~pi045 & ~pi043;
  assign new_n13569_ = ~pi048 & ~pi049 & ~pi047;
  assign new_n13570_ = ~pi051 & ~pi034 & ~pi052 & ~pi050;
  assign new_n13571_ = ~pi053 & ~pi054 & ~pi033;
  assign new_n13572_ = new_n13570_ & new_n13568_ & new_n13569_ & new_n13571_;
  assign new_n13573_ = ~pi056 & ~pi058 & ~pi057 & ~pi055;
  assign new_n13574_ = ~pi035 & ~pi036 & ~pi059;
  assign new_n13575_ = ~pi038 & ~pi039 & ~pi037;
  assign new_n13576_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13577_ = new_n13575_ & new_n13573_ & new_n13574_ & new_n13576_;
  assign new_n13578_ = ~pi044 & ~pi046 & ~pi045 & ~pi043;
  assign new_n13579_ = ~pi048 & ~pi049 & ~pi047;
  assign new_n13580_ = ~pi051 & ~pi052 & ~pi050;
  assign new_n13581_ = ~pi033 & ~pi053 & ~pi034;
  assign new_n13582_ = new_n13580_ & new_n13578_ & new_n13579_ & new_n13581_;
  assign new_n13583_ = ~pi055 & ~pi057 & ~pi056 & ~pi054;
  assign new_n13584_ = ~pi035 & ~pi036 & ~pi058;
  assign new_n13585_ = ~pi038 & ~pi039 & ~pi037;
  assign new_n13586_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13587_ = new_n13585_ & new_n13583_ & new_n13584_ & new_n13586_;
  assign new_n13588_ = ~pi044 & ~pi046 & ~pi045 & ~pi043;
  assign new_n13589_ = ~pi048 & ~pi049 & ~pi047;
  assign new_n13590_ = ~pi051 & ~pi052 & ~pi050;
  assign new_n13591_ = ~pi033 & ~pi053 & ~pi034;
  assign new_n13592_ = new_n13590_ & new_n13588_ & new_n13589_ & new_n13591_;
  assign new_n13593_ = ~pi055 & ~pi056 & ~pi054;
  assign new_n13594_ = ~pi035 & ~pi036 & ~pi057;
  assign new_n13595_ = ~pi038 & ~pi039 & ~pi037;
  assign new_n13596_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13597_ = new_n13595_ & new_n13593_ & new_n13594_ & new_n13596_;
  assign new_n13598_ = ~pi044 & ~pi045 & ~pi043;
  assign new_n13599_ = ~pi047 & ~pi048 & ~pi046;
  assign new_n13600_ = ~pi050 & ~pi051 & ~pi049;
  assign new_n13601_ = ~pi034 & ~pi033 & ~pi052;
  assign new_n13602_ = new_n13600_ & new_n13598_ & new_n13599_ & new_n13601_;
  assign new_n13603_ = ~pi054 & ~pi055 & ~pi053;
  assign new_n13604_ = ~pi035 & ~pi036 & ~pi056;
  assign new_n13605_ = ~pi038 & ~pi039 & ~pi037;
  assign new_n13606_ = ~pi041 & ~pi042 & ~pi040;
  assign new_n13607_ = new_n13605_ & new_n13603_ & new_n13604_ & new_n13606_;
  assign new_n13608_ = ~pi047 & ~pi046 & ~pi044 & ~pi043 & ~pi045;
  assign new_n13609_ = ~pi049 & ~pi033 & ~pi034 & ~pi048;
  assign new_n13610_ = ~pi036 & ~pi038 & ~pi037 & ~pi035;
  assign new_n13611_ = ~pi040 & ~pi042 & ~pi041 & ~pi039;
  assign new_n13612_ = ~pi050 & ~pi051;
  assign new_n13613_ = ~pi052 & ~pi053;
  assign new_n13614_ = ~pi054 & ~pi055;
  assign new_n13615_ = new_n13614_ & new_n13613_ & new_n13612_;
  assign new_n13616_ = ~pi044 & ~pi045 & ~pi043;
  assign new_n13617_ = ~pi047 & ~pi048 & ~pi046;
  assign new_n13618_ = new_n13617_ & new_n13616_;
  assign new_n13619_ = ~pi034 & ~pi052 & ~pi050 & ~pi049 & ~pi051;
  assign new_n13620_ = ~pi053 & ~pi054 & ~pi033;
  assign new_n13621_ = ~pi036 & ~pi037 & ~pi035;
  assign new_n13622_ = new_n13621_ & new_n13620_;
  assign new_n13623_ = ~pi042 & ~pi041 & ~pi039 & ~pi038 & ~pi040;
  assign new_n13624_ = ~pi044 & ~pi045 & ~pi043;
  assign new_n13625_ = ~pi047 & ~pi048 & ~pi046;
  assign new_n13626_ = ~pi034 & ~pi052 & ~pi050 & ~pi049 & ~pi051;
  assign new_n13627_ = ~pi037 & ~pi036 & ~pi053 & ~pi033 & ~pi035;
  assign new_n13628_ = ~pi042 & ~pi041 & ~pi039 & ~pi038 & ~pi040;
  assign new_n13629_ = ~pi047 & ~pi046 & ~pi044 & ~pi043 & ~pi045;
  assign new_n13630_ = ~pi052 & ~pi051 & ~pi049 & ~pi048 & ~pi050;
  assign new_n13631_ = ~pi037 & ~pi036 & ~pi033 & ~pi034 & ~pi035;
  assign new_n13632_ = ~pi042 & ~pi041 & ~pi039 & ~pi038 & ~pi040;
  assign new_n13633_ = ~pi047 & ~pi046 & ~pi044 & ~pi043 & ~pi045;
  assign new_n13634_ = ~pi034 & ~pi051 & ~pi049 & ~pi048 & ~pi050;
  assign new_n13635_ = ~pi038 & ~pi037 & ~pi035 & ~pi033 & ~pi036;
  assign new_n13636_ = ~pi040 & ~pi042 & ~pi041 & ~pi039;
  assign new_n13637_ = ~pi044 & ~pi042 & ~pi045 & ~pi043;
  assign new_n13638_ = ~pi046 & ~pi047;
  assign new_n13639_ = ~pi043 & ~pi042;
  assign new_n13640_ = ~pi042;
  assign new_n13641_ = new_n13714_ & new_n13713_;
  assign new_n13642_ = ~pi038;
  assign new_n13643_ = new_n13716_ & new_n13715_;
  assign new_n13644_ = ~pi064;
  assign new_n13645_ = ~pi063;
  assign new_n13646_ = new_n13720_ & new_n13719_;
  assign new_n13647_ = ~pi060;
  assign new_n13648_ = ~new_n13577_ | ~new_n13572_;
  assign new_n13649_ = ~pi058;
  assign new_n13650_ = ~new_n13597_ | ~new_n13592_;
  assign new_n13651_ = new_n13724_ & new_n13723_;
  assign new_n13652_ = ~pi054;
  assign new_n13653_ = ~new_n13625_ | ~new_n13627_ | ~new_n13628_ | ~new_n13626_ | ~new_n13624_;
  assign new_n13654_ = new_n13726_ & new_n13725_;
  assign new_n13655_ = ~pi034;
  assign new_n13656_ = ~pi033;
  assign new_n13657_ = ~pi050;
  assign new_n13658_ = new_n13730_ & new_n13729_;
  assign new_n13659_ = ~pi046;
  assign new_n13660_ = new_n13732_ & new_n13731_;
  assign new_n13661_ = ~new_n13711_ | ~new_n13513_;
  assign new_n13662_ = ~new_n13510_;
  assign new_n13663_ = ~new_n13511_;
  assign new_n13664_ = ~new_n13663_ | ~new_n13512_;
  assign new_n13665_ = ~new_n13509_;
  assign new_n13666_ = ~pi041 | ~new_n13664_;
  assign new_n13667_ = ~pi040 | ~new_n13511_;
  assign new_n13668_ = ~new_n13662_ | ~new_n13642_;
  assign new_n13669_ = ~pi039 | ~new_n13668_;
  assign new_n13670_ = ~pi037 | ~new_n13661_;
  assign new_n13671_ = ~pi036 | ~new_n13508_;
  assign new_n13672_ = ~new_n13519_;
  assign new_n13673_ = ~new_n13672_ | ~new_n13520_;
  assign new_n13674_ = ~new_n13516_;
  assign new_n13675_ = ~new_n13517_;
  assign new_n13676_ = ~new_n13675_ | ~new_n13518_;
  assign new_n13677_ = ~new_n13515_;
  assign new_n13678_ = ~new_n13635_ | ~new_n13633_ | ~new_n13634_ | ~new_n13636_;
  assign new_n13679_ = ~new_n13631_ | ~new_n13629_ | ~new_n13630_ | ~new_n13632_;
  assign new_n13680_ = ~new_n13653_;
  assign new_n13681_ = ~new_n13615_ | ~new_n13677_;
  assign new_n13682_ = ~new_n13607_ | ~new_n13602_;
  assign new_n13683_ = ~new_n13650_;
  assign new_n13684_ = ~new_n13648_;
  assign new_n13685_ = ~new_n13547_ | ~new_n13542_;
  assign new_n13686_ = ~new_n13514_;
  assign new_n13687_ = pi034 | pi033;
  assign new_n13688_ = ~pi035 | ~new_n13687_;
  assign new_n13689_ = ~pi062 | ~new_n13685_;
  assign new_n13690_ = ~pi061 | ~new_n13710_;
  assign new_n13691_ = ~new_n13587_ | ~new_n13582_;
  assign new_n13692_ = ~pi059 | ~new_n13691_;
  assign new_n13693_ = ~pi057 | ~new_n13682_;
  assign new_n13694_ = ~pi056 | ~new_n13681_;
  assign new_n13695_ = ~new_n13622_ | ~new_n13618_ | ~new_n13619_ | ~new_n13623_;
  assign new_n13696_ = ~pi055 | ~new_n13695_;
  assign new_n13697_ = ~pi053 | ~new_n13679_;
  assign new_n13698_ = ~pi052 | ~new_n13678_;
  assign new_n13699_ = ~new_n13677_ | ~new_n13657_;
  assign new_n13700_ = ~pi051 | ~new_n13699_;
  assign new_n13701_ = ~pi049 | ~new_n13676_;
  assign new_n13702_ = ~pi048 | ~new_n13517_;
  assign new_n13703_ = ~new_n13674_ | ~new_n13659_;
  assign new_n13704_ = ~pi047 | ~new_n13703_;
  assign new_n13705_ = ~pi045 | ~new_n13673_;
  assign new_n13706_ = ~pi044 | ~new_n13519_;
  assign new_n13707_ = ~new_n13665_ | ~new_n13640_;
  assign new_n13708_ = ~pi043 | ~new_n13707_;
  assign new_n13709_ = ~new_n13686_ | ~new_n13645_;
  assign new_n13710_ = ~new_n13557_ | ~new_n13552_;
  assign new_n13711_ = ~new_n13508_;
  assign new_n13712_ = ~new_n13567_ | ~new_n13562_;
  assign new_n13713_ = ~pi042 | ~new_n13509_;
  assign new_n13714_ = ~new_n13665_ | ~new_n13640_;
  assign new_n13715_ = ~pi038 | ~new_n13510_;
  assign new_n13716_ = ~new_n13662_ | ~new_n13642_;
  assign new_n13717_ = ~new_n13709_ | ~new_n13644_;
  assign new_n13718_ = ~pi064 | ~new_n13686_ | ~new_n13645_;
  assign new_n13719_ = ~pi063 | ~new_n13514_;
  assign new_n13720_ = ~new_n13686_ | ~new_n13645_;
  assign new_n13721_ = ~new_n13684_ | ~pi060;
  assign new_n13722_ = ~new_n13712_ | ~new_n13647_;
  assign new_n13723_ = ~pi058 | ~new_n13650_;
  assign new_n13724_ = ~new_n13683_ | ~new_n13649_;
  assign new_n13725_ = ~pi054 | ~new_n13653_;
  assign new_n13726_ = ~new_n13680_ | ~new_n13652_;
  assign new_n13727_ = ~pi034 | ~new_n13656_;
  assign new_n13728_ = ~pi033 | ~new_n13655_;
  assign new_n13729_ = ~pi050 | ~new_n13515_;
  assign new_n13730_ = ~new_n13677_ | ~new_n13657_;
  assign new_n13731_ = ~pi046 | ~new_n13516_;
  assign new_n13732_ = ~new_n13674_ | ~new_n13659_;
  assign new_n13733_ = ~new_n1986_;
  assign new_n13734_ = ~new_n1983_;
  assign new_n13735_ = new_n13737_ & new_n13736_;
  assign new_n13736_ = ~new_n1983_ | ~new_n13733_;
  assign new_n13737_ = ~new_n1986_ | ~new_n13734_;
  assign new_n13738_ = new_n13867_ & new_n13767_;
  assign new_n13739_ = new_n13865_ & new_n13768_;
  assign new_n13740_ = new_n13864_ & new_n13769_;
  assign new_n13741_ = new_n13863_ & new_n13770_;
  assign new_n13742_ = new_n13861_ & new_n13771_;
  assign new_n13743_ = new_n13860_ & new_n13772_;
  assign new_n13744_ = new_n13859_ & new_n13773_;
  assign new_n13745_ = new_n13857_ & new_n13774_;
  assign new_n13746_ = new_n13855_ & new_n13775_;
  assign new_n13747_ = new_n13853_ & new_n13776_;
  assign new_n13748_ = new_n13851_ & new_n13777_;
  assign new_n13749_ = new_n13849_ & new_n13778_;
  assign new_n13750_ = new_n13847_ & new_n13757_;
  assign new_n13751_ = new_n13845_ & new_n13799_;
  assign new_n13752_ = new_n13830_ & new_n13758_;
  assign new_n13753_ = new_n13829_ & new_n13759_;
  assign new_n13754_ = new_n13828_ & new_n13760_;
  assign new_n13755_ = new_n13826_ & new_n13761_;
  assign new_n13756_ = new_n13825_ & new_n13762_;
  assign new_n13757_ = new_n2391_ | new_n2388_ | new_n2383_;
  assign new_n13758_ = ~new_n13819_ | ~new_n13766_;
  assign new_n13759_ = ~new_n13820_ | ~new_n13765_;
  assign new_n13760_ = ~new_n13789_ | ~new_n13821_;
  assign new_n13761_ = ~new_n13822_ | ~new_n13764_;
  assign new_n13762_ = ~new_n13823_ | ~new_n13763_;
  assign new_n13763_ = ~new_n2409_;
  assign new_n13764_ = ~new_n2406_;
  assign new_n13765_ = ~new_n2397_;
  assign new_n13766_ = ~new_n2394_;
  assign new_n13767_ = ~new_n13790_ | ~new_n13824_;
  assign new_n13768_ = ~new_n13831_ | ~new_n13787_;
  assign new_n13769_ = ~new_n13832_ | ~new_n13786_;
  assign new_n13770_ = ~new_n13791_ | ~new_n13833_;
  assign new_n13771_ = ~new_n13834_ | ~new_n13785_;
  assign new_n13772_ = ~new_n13835_ | ~new_n13784_;
  assign new_n13773_ = ~new_n13792_ | ~new_n13836_;
  assign new_n13774_ = ~new_n13793_ | ~new_n13837_;
  assign new_n13775_ = ~new_n13783_ | ~new_n13838_ | ~new_n13809_;
  assign new_n13776_ = ~new_n13782_ | ~new_n13839_ | ~new_n13807_;
  assign new_n13777_ = ~new_n13781_ | ~new_n13840_ | ~new_n13805_;
  assign new_n13778_ = ~new_n13780_ | ~new_n13841_ | ~new_n13803_;
  assign new_n13779_ = ~new_n2954_;
  assign new_n13780_ = ~new_n2944_;
  assign new_n13781_ = ~new_n2946_;
  assign new_n13782_ = ~new_n2948_;
  assign new_n13783_ = ~new_n2950_;
  assign new_n13784_ = ~new_n2433_;
  assign new_n13785_ = ~new_n2430_;
  assign new_n13786_ = ~new_n2421_;
  assign new_n13787_ = ~new_n2418_;
  assign new_n13788_ = ~new_n13885_ | ~new_n13884_;
  assign new_n13789_ = ~new_n2400_ & ~new_n2403_;
  assign new_n13790_ = ~new_n2415_ & ~new_n2412_;
  assign new_n13791_ = ~new_n2424_ & ~new_n2427_;
  assign new_n13792_ = ~new_n2436_ & ~new_n2439_;
  assign new_n13793_ = ~new_n2441_ & ~new_n2952_;
  assign new_n13794_ = ~new_n2412_;
  assign new_n13795_ = new_n13869_ & new_n13868_;
  assign new_n13796_ = ~new_n2400_;
  assign new_n13797_ = new_n13871_ & new_n13870_;
  assign new_n13798_ = ~new_n2953_;
  assign new_n13799_ = ~new_n13779_ | ~new_n13842_ | ~new_n13801_;
  assign new_n13800_ = new_n13873_ & new_n13872_;
  assign new_n13801_ = ~new_n2955_;
  assign new_n13802_ = new_n13875_ & new_n13874_;
  assign new_n13803_ = ~new_n2945_;
  assign new_n13804_ = new_n13877_ & new_n13876_;
  assign new_n13805_ = ~new_n2947_;
  assign new_n13806_ = new_n13879_ & new_n13878_;
  assign new_n13807_ = ~new_n2949_;
  assign new_n13808_ = new_n13881_ & new_n13880_;
  assign new_n13809_ = ~new_n2951_;
  assign new_n13810_ = new_n13883_ & new_n13882_;
  assign new_n13811_ = ~new_n2388_;
  assign new_n13812_ = ~new_n2383_;
  assign new_n13813_ = ~new_n2441_;
  assign new_n13814_ = new_n13887_ & new_n13886_;
  assign new_n13815_ = ~new_n2436_;
  assign new_n13816_ = new_n13889_ & new_n13888_;
  assign new_n13817_ = ~new_n2424_;
  assign new_n13818_ = new_n13891_ & new_n13890_;
  assign new_n13819_ = ~new_n13757_;
  assign new_n13820_ = ~new_n13758_;
  assign new_n13821_ = ~new_n13759_;
  assign new_n13822_ = ~new_n13760_;
  assign new_n13823_ = ~new_n13761_;
  assign new_n13824_ = ~new_n13762_;
  assign new_n13825_ = ~new_n2409_ | ~new_n13761_;
  assign new_n13826_ = ~new_n2406_ | ~new_n13760_;
  assign new_n13827_ = ~new_n13821_ | ~new_n13796_;
  assign new_n13828_ = ~new_n2403_ | ~new_n13827_;
  assign new_n13829_ = ~new_n2397_ | ~new_n13758_;
  assign new_n13830_ = ~new_n2394_ | ~new_n13757_;
  assign new_n13831_ = ~new_n13767_;
  assign new_n13832_ = ~new_n13768_;
  assign new_n13833_ = ~new_n13769_;
  assign new_n13834_ = ~new_n13770_;
  assign new_n13835_ = ~new_n13771_;
  assign new_n13836_ = ~new_n13772_;
  assign new_n13837_ = ~new_n13773_;
  assign new_n13838_ = ~new_n13774_;
  assign new_n13839_ = ~new_n13775_;
  assign new_n13840_ = ~new_n13776_;
  assign new_n13841_ = ~new_n13777_;
  assign new_n13842_ = ~new_n13778_;
  assign new_n13843_ = ~new_n13799_;
  assign new_n13844_ = ~new_n13842_ | ~new_n13801_;
  assign new_n13845_ = ~new_n2954_ | ~new_n13844_;
  assign new_n13846_ = new_n2388_ | new_n2383_;
  assign new_n13847_ = ~new_n2391_ | ~new_n13846_;
  assign new_n13848_ = ~new_n13841_ | ~new_n13803_;
  assign new_n13849_ = ~new_n2944_ | ~new_n13848_;
  assign new_n13850_ = ~new_n13840_ | ~new_n13805_;
  assign new_n13851_ = ~new_n2946_ | ~new_n13850_;
  assign new_n13852_ = ~new_n13839_ | ~new_n13807_;
  assign new_n13853_ = ~new_n2948_ | ~new_n13852_;
  assign new_n13854_ = ~new_n13838_ | ~new_n13809_;
  assign new_n13855_ = ~new_n2950_ | ~new_n13854_;
  assign new_n13856_ = ~new_n13837_ | ~new_n13813_;
  assign new_n13857_ = ~new_n2952_ | ~new_n13856_;
  assign new_n13858_ = ~new_n13836_ | ~new_n13815_;
  assign new_n13859_ = ~new_n2439_ | ~new_n13858_;
  assign new_n13860_ = ~new_n2433_ | ~new_n13771_;
  assign new_n13861_ = ~new_n2430_ | ~new_n13770_;
  assign new_n13862_ = ~new_n13833_ | ~new_n13817_;
  assign new_n13863_ = ~new_n2427_ | ~new_n13862_;
  assign new_n13864_ = ~new_n2421_ | ~new_n13768_;
  assign new_n13865_ = ~new_n2418_ | ~new_n13767_;
  assign new_n13866_ = ~new_n13824_ | ~new_n13794_;
  assign new_n13867_ = ~new_n2415_ | ~new_n13866_;
  assign new_n13868_ = ~new_n2412_ | ~new_n13762_;
  assign new_n13869_ = ~new_n13824_ | ~new_n13794_;
  assign new_n13870_ = ~new_n2400_ | ~new_n13759_;
  assign new_n13871_ = ~new_n13821_ | ~new_n13796_;
  assign new_n13872_ = ~new_n2953_ | ~new_n13799_;
  assign new_n13873_ = ~new_n13843_ | ~new_n13798_;
  assign new_n13874_ = ~new_n2955_ | ~new_n13778_;
  assign new_n13875_ = ~new_n13842_ | ~new_n13801_;
  assign new_n13876_ = ~new_n2945_ | ~new_n13777_;
  assign new_n13877_ = ~new_n13841_ | ~new_n13803_;
  assign new_n13878_ = ~new_n2947_ | ~new_n13776_;
  assign new_n13879_ = ~new_n13840_ | ~new_n13805_;
  assign new_n13880_ = ~new_n2949_ | ~new_n13775_;
  assign new_n13881_ = ~new_n13839_ | ~new_n13807_;
  assign new_n13882_ = ~new_n2951_ | ~new_n13774_;
  assign new_n13883_ = ~new_n13838_ | ~new_n13809_;
  assign new_n13884_ = ~new_n2388_ | ~new_n13812_;
  assign new_n13885_ = ~new_n2383_ | ~new_n13811_;
  assign new_n13886_ = ~new_n2441_ | ~new_n13773_;
  assign new_n13887_ = ~new_n13837_ | ~new_n13813_;
  assign new_n13888_ = ~new_n2436_ | ~new_n13772_;
  assign new_n13889_ = ~new_n13836_ | ~new_n13815_;
  assign new_n13890_ = ~new_n2424_ | ~new_n13769_;
  assign new_n13891_ = ~new_n13833_ | ~new_n13817_;
  assign new_n13892_ = new_n14064_ & new_n14063_;
  assign new_n13893_ = new_n14065_ & new_n14066_;
  assign new_n13894_ = new_n14082_ & new_n14081_;
  assign new_n13895_ = new_n14122_ & new_n14121_;
  assign new_n13896_ = new_n14131_ & new_n14130_;
  assign new_n13897_ = new_n14149_ & new_n14148_;
  assign new_n13898_ = new_n14157_ & new_n14156_;
  assign new_n13899_ = new_n14236_ & new_n14233_;
  assign new_n13900_ = new_n14229_ & new_n14226_;
  assign new_n13901_ = new_n14220_ & new_n14217_;
  assign new_n13902_ = new_n14211_ & new_n14208_;
  assign new_n13903_ = new_n14205_ & new_n14203_;
  assign new_n13904_ = new_n14198_ & new_n14195_;
  assign new_n13905_ = new_n14120_ & new_n14117_;
  assign new_n13906_ = new_n14112_ & new_n14109_;
  assign new_n13907_ = new_n14098_ & new_n14095_;
  assign new_n13908_ = ~new_n2403_;
  assign new_n13909_ = ~new_n1998_;
  assign new_n13910_ = ~new_n1997_;
  assign new_n13911_ = ~new_n1998_ | ~new_n2403_;
  assign new_n13912_ = ~new_n2406_;
  assign new_n13913_ = ~new_n2397_;
  assign new_n13914_ = ~new_n1987_;
  assign new_n13915_ = ~new_n1994_;
  assign new_n13916_ = ~new_n2391_;
  assign new_n13917_ = ~new_n1995_;
  assign new_n13918_ = ~new_n2383_;
  assign new_n13919_ = ~new_n2004_;
  assign new_n13920_ = ~new_n2004_ | ~new_n2383_;
  assign new_n13921_ = ~new_n2394_;
  assign new_n13922_ = ~new_n1991_;
  assign new_n13923_ = ~new_n1987_ | ~new_n2397_;
  assign new_n13924_ = ~new_n2400_;
  assign new_n13925_ = ~new_n2409_;
  assign new_n13926_ = ~new_n2011_;
  assign new_n13927_ = ~new_n2010_;
  assign new_n13928_ = ~new_n2412_;
  assign new_n13929_ = ~new_n13950_ | ~new_n14090_;
  assign new_n13930_ = ~new_n14006_ | ~new_n14078_;
  assign new_n13931_ = ~new_n14067_ | ~new_n14068_;
  assign new_n13932_ = ~new_n2388_ | ~new_n2005_;
  assign new_n13933_ = ~new_n14010_ | ~new_n14104_;
  assign new_n13934_ = ~new_n14101_ | ~new_n14100_;
  assign new_n13935_ = ~new_n2945_;
  assign new_n13936_ = ~new_n1980_;
  assign new_n13937_ = ~new_n1984_;
  assign new_n13938_ = ~new_n2946_;
  assign new_n13939_ = ~new_n2947_;
  assign new_n13940_ = ~new_n1985_;
  assign new_n13941_ = ~new_n2948_;
  assign new_n13942_ = ~new_n1992_;
  assign new_n13943_ = ~new_n2951_;
  assign new_n13944_ = ~new_n2002_;
  assign new_n13945_ = ~new_n2433_;
  assign new_n13946_ = ~new_n2000_;
  assign new_n13947_ = ~new_n1996_;
  assign new_n13948_ = ~new_n2000_ | ~new_n2433_;
  assign new_n13949_ = ~new_n2436_;
  assign new_n13950_ = ~new_n2011_ | ~new_n2409_;
  assign new_n13951_ = ~new_n2415_;
  assign new_n13952_ = ~new_n1989_;
  assign new_n13953_ = ~new_n2421_;
  assign new_n13954_ = ~new_n1999_;
  assign new_n13955_ = ~new_n2418_;
  assign new_n13956_ = ~new_n1990_;
  assign new_n13957_ = ~new_n1990_ | ~new_n2418_;
  assign new_n13958_ = ~new_n2424_;
  assign new_n13959_ = ~new_n2007_;
  assign new_n13960_ = ~new_n2427_;
  assign new_n13961_ = ~new_n2006_;
  assign new_n13962_ = ~new_n2430_;
  assign new_n13963_ = ~new_n2001_;
  assign new_n13964_ = ~new_n2439_;
  assign new_n13965_ = ~new_n2009_;
  assign new_n13966_ = ~new_n2009_ | ~new_n2439_;
  assign new_n13967_ = ~new_n2441_;
  assign new_n13968_ = ~new_n2008_;
  assign new_n13969_ = ~new_n2008_ | ~new_n2441_;
  assign new_n13970_ = ~new_n2952_;
  assign new_n13971_ = ~new_n2950_;
  assign new_n13972_ = ~new_n1988_;
  assign new_n13973_ = ~new_n2949_;
  assign new_n13974_ = ~new_n1993_;
  assign new_n13975_ = ~new_n2946_ | ~new_n1984_;
  assign new_n13976_ = ~new_n1981_;
  assign new_n13977_ = ~new_n2944_;
  assign new_n13978_ = ~new_n14191_ | ~new_n14061_;
  assign new_n13979_ = ~new_n2003_;
  assign new_n13980_ = ~new_n13966_ | ~new_n14200_;
  assign new_n13981_ = ~new_n14146_ | ~new_n14145_;
  assign new_n13982_ = ~new_n13957_ | ~new_n14222_;
  assign new_n13983_ = ~new_n14342_ | ~new_n14341_;
  assign new_n13984_ = ~new_n14389_ | ~new_n14388_;
  assign new_n13985_ = ~new_n14260_ | ~new_n14259_;
  assign new_n13986_ = ~new_n14265_ | ~new_n14264_;
  assign new_n13987_ = ~new_n14272_ | ~new_n14271_;
  assign new_n13988_ = ~new_n14279_ | ~new_n14278_;
  assign new_n13989_ = ~new_n14284_ | ~new_n14283_;
  assign new_n13990_ = ~new_n14293_ | ~new_n14292_;
  assign new_n13991_ = ~new_n14300_ | ~new_n14299_;
  assign new_n13992_ = ~new_n14307_ | ~new_n14306_;
  assign new_n13993_ = ~new_n14314_ | ~new_n14313_;
  assign new_n13994_ = ~new_n14319_ | ~new_n14318_;
  assign new_n13995_ = ~new_n14326_ | ~new_n14325_;
  assign new_n13996_ = ~new_n14333_ | ~new_n14332_;
  assign new_n13997_ = ~new_n14347_ | ~new_n14346_;
  assign new_n13998_ = ~new_n14352_ | ~new_n14351_;
  assign new_n13999_ = ~new_n14359_ | ~new_n14358_;
  assign new_n14000_ = ~new_n14366_ | ~new_n14365_;
  assign new_n14001_ = ~new_n14373_ | ~new_n14372_;
  assign new_n14002_ = ~new_n14380_ | ~new_n14379_;
  assign new_n14003_ = ~new_n14385_ | ~new_n14384_;
  assign new_n14004_ = new_n2391_ & new_n1995_;
  assign new_n14005_ = new_n14074_ & new_n14072_;
  assign new_n14006_ = new_n14079_ & new_n14077_;
  assign new_n14007_ = new_n14086_ & new_n14085_;
  assign new_n14008_ = new_n13911_ & new_n14267_ & new_n14266_;
  assign new_n14009_ = new_n14097_ & new_n13894_;
  assign new_n14010_ = new_n14105_ & new_n14103_;
  assign new_n14011_ = new_n13923_ & new_n14274_ & new_n14273_;
  assign new_n14012_ = new_n14111_ & new_n13892_;
  assign new_n14013_ = new_n14119_ & new_n14066_;
  assign new_n14014_ = new_n14089_ & new_n13895_;
  assign new_n14015_ = new_n14124_ & new_n14056_;
  assign new_n14016_ = new_n14133_ & new_n14057_;
  assign new_n14017_ = new_n14153_ & new_n14152_;
  assign new_n14018_ = new_n13898_ & new_n14167_;
  assign new_n14019_ = new_n14170_ & new_n14165_;
  assign new_n14020_ = new_n14186_ & new_n14183_;
  assign new_n14021_ = new_n14253_ & new_n14187_;
  assign new_n14022_ = new_n14044_ & new_n14163_;
  assign new_n14023_ = new_n13948_ & new_n14354_ & new_n14353_;
  assign new_n14024_ = new_n14057_ & new_n14375_ & new_n14374_;
  assign new_n14025_ = new_n14228_ & new_n13896_;
  assign new_n14026_ = new_n14056_ & new_n14387_ & new_n14386_;
  assign new_n14027_ = new_n14235_ & new_n13895_;
  assign new_n14028_ = ~new_n14007_ | ~new_n14087_;
  assign new_n14029_ = ~new_n14102_ | ~new_n14114_;
  assign new_n14030_ = ~new_n1982_;
  assign new_n14031_ = ~new_n2955_;
  assign new_n14032_ = new_n14288_ & new_n14287_;
  assign new_n14033_ = ~new_n14249_ | ~new_n14189_ | ~new_n14054_;
  assign new_n14034_ = new_n14295_ & new_n14294_;
  assign new_n14035_ = ~new_n14021_ | ~new_n14255_ | ~new_n14254_;
  assign new_n14036_ = new_n14302_ & new_n14301_;
  assign new_n14037_ = ~new_n13975_ | ~new_n14250_ | ~new_n14184_;
  assign new_n14038_ = new_n14309_ & new_n14308_;
  assign new_n14039_ = ~new_n14178_ | ~new_n14177_;
  assign new_n14040_ = new_n14321_ & new_n14320_;
  assign new_n14041_ = ~new_n14174_ | ~new_n14173_;
  assign new_n14042_ = new_n14328_ & new_n14327_;
  assign new_n14043_ = ~new_n14019_ | ~new_n14169_;
  assign new_n14044_ = new_n14335_ & new_n14334_;
  assign new_n14045_ = new_n14340_ & new_n14339_;
  assign new_n14046_ = ~new_n13932_ | ~new_n14212_;
  assign new_n14047_ = ~new_n14017_ | ~new_n14154_;
  assign new_n14048_ = new_n14361_ & new_n14360_;
  assign new_n14049_ = ~new_n14142_ | ~new_n14141_;
  assign new_n14050_ = new_n14368_ & new_n14367_;
  assign new_n14051_ = ~new_n14138_ | ~new_n14137_;
  assign new_n14052_ = ~new_n14128_ | ~new_n14127_;
  assign new_n14053_ = ~new_n14252_ | ~new_n14251_;
  assign new_n14054_ = ~new_n1981_ | ~new_n14035_;
  assign new_n14055_ = ~new_n13923_;
  assign new_n14056_ = ~new_n2412_ | ~new_n2010_;
  assign new_n14057_ = ~new_n1999_ | ~new_n2421_;
  assign new_n14058_ = ~new_n1985_ | ~new_n2947_;
  assign new_n14059_ = ~new_n13957_;
  assign new_n14060_ = ~new_n13966_;
  assign new_n14061_ = ~new_n1992_ | ~new_n2948_;
  assign new_n14062_ = ~new_n13950_;
  assign new_n14063_ = new_n1994_ | new_n2400_;
  assign new_n14064_ = new_n1987_ | new_n2397_;
  assign new_n14065_ = new_n2394_ | new_n1991_;
  assign new_n14066_ = new_n2391_ | new_n1995_;
  assign new_n14067_ = ~new_n13920_;
  assign new_n14068_ = new_n2388_ | new_n2005_;
  assign new_n14069_ = ~new_n13931_;
  assign new_n14070_ = ~new_n13932_;
  assign new_n14071_ = ~new_n13931_ | ~new_n13932_;
  assign new_n14072_ = ~new_n14004_ | ~new_n14065_;
  assign new_n14073_ = ~new_n13893_ | ~new_n14071_;
  assign new_n14074_ = ~new_n1991_ | ~new_n2394_;
  assign new_n14075_ = ~new_n14005_ | ~new_n14073_;
  assign new_n14076_ = ~new_n13924_ | ~new_n13923_;
  assign new_n14077_ = ~new_n1994_ | ~new_n14076_;
  assign new_n14078_ = ~new_n13892_ | ~new_n14075_;
  assign new_n14079_ = ~new_n2400_ | ~new_n14055_;
  assign new_n14080_ = ~new_n13930_;
  assign new_n14081_ = new_n1997_ | new_n2406_;
  assign new_n14082_ = new_n1998_ | new_n2403_;
  assign new_n14083_ = ~new_n13911_;
  assign new_n14084_ = ~new_n13912_ | ~new_n13911_;
  assign new_n14085_ = ~new_n1997_ | ~new_n14084_;
  assign new_n14086_ = ~new_n2406_ | ~new_n14083_;
  assign new_n14087_ = ~new_n13894_ | ~new_n13930_;
  assign new_n14088_ = ~new_n14028_;
  assign new_n14089_ = new_n2409_ | new_n2011_;
  assign new_n14090_ = ~new_n14089_ | ~new_n14028_;
  assign new_n14091_ = ~new_n13929_;
  assign new_n14092_ = new_n2010_ | new_n2412_;
  assign new_n14093_ = new_n2403_ | new_n1998_;
  assign new_n14094_ = ~new_n14093_ | ~new_n13930_;
  assign new_n14095_ = ~new_n14008_ | ~new_n14094_;
  assign new_n14096_ = ~new_n14080_ | ~new_n13911_;
  assign new_n14097_ = ~new_n2406_ | ~new_n1997_;
  assign new_n14098_ = ~new_n14009_ | ~new_n14096_;
  assign new_n14099_ = new_n1998_ | new_n2403_;
  assign new_n14100_ = ~new_n14070_ | ~new_n14066_;
  assign new_n14101_ = ~new_n1995_ | ~new_n2391_;
  assign new_n14102_ = ~new_n13934_;
  assign new_n14103_ = ~new_n14069_ | ~new_n13893_;
  assign new_n14104_ = ~new_n13934_ | ~new_n14065_;
  assign new_n14105_ = ~new_n1991_ | ~new_n2394_;
  assign new_n14106_ = ~new_n13933_;
  assign new_n14107_ = new_n2397_ | new_n1987_;
  assign new_n14108_ = ~new_n14107_ | ~new_n13933_;
  assign new_n14109_ = ~new_n14011_ | ~new_n14108_;
  assign new_n14110_ = ~new_n14106_ | ~new_n13923_;
  assign new_n14111_ = ~new_n2400_ | ~new_n1994_;
  assign new_n14112_ = ~new_n14012_ | ~new_n14110_;
  assign new_n14113_ = new_n1987_ | new_n2397_;
  assign new_n14114_ = ~new_n14069_ | ~new_n14066_;
  assign new_n14115_ = ~new_n14029_;
  assign new_n14116_ = ~new_n1991_ | ~new_n2394_;
  assign new_n14117_ = ~new_n14285_ | ~new_n13931_ | ~new_n13932_ | ~new_n14286_;
  assign new_n14118_ = ~new_n13932_ | ~new_n13931_;
  assign new_n14119_ = ~new_n1995_ | ~new_n2391_;
  assign new_n14120_ = ~new_n14013_ | ~new_n14118_;
  assign new_n14121_ = new_n2010_ | new_n2412_;
  assign new_n14122_ = new_n1989_ | new_n2415_;
  assign new_n14123_ = ~new_n14062_ | ~new_n13895_;
  assign new_n14124_ = ~new_n1989_ | ~new_n2415_;
  assign new_n14125_ = ~new_n14015_ | ~new_n14123_;
  assign new_n14126_ = new_n2415_ | new_n1989_;
  assign new_n14127_ = ~new_n14014_ | ~new_n14028_;
  assign new_n14128_ = ~new_n14126_ | ~new_n14125_;
  assign new_n14129_ = ~new_n14052_;
  assign new_n14130_ = new_n2007_ | new_n2424_;
  assign new_n14131_ = new_n1999_ | new_n2421_;
  assign new_n14132_ = ~new_n14059_ | ~new_n13896_;
  assign new_n14133_ = ~new_n2007_ | ~new_n2424_;
  assign new_n14134_ = ~new_n14016_ | ~new_n14132_;
  assign new_n14135_ = new_n2418_ | new_n1990_;
  assign new_n14136_ = new_n2424_ | new_n2007_;
  assign new_n14137_ = ~new_n13896_ | ~new_n14135_ | ~new_n14052_;
  assign new_n14138_ = ~new_n14136_ | ~new_n14134_;
  assign new_n14139_ = ~new_n14051_;
  assign new_n14140_ = new_n2427_ | new_n2006_;
  assign new_n14141_ = ~new_n14140_ | ~new_n14051_;
  assign new_n14142_ = ~new_n2006_ | ~new_n2427_;
  assign new_n14143_ = ~new_n14049_;
  assign new_n14144_ = new_n2430_ | new_n2001_;
  assign new_n14145_ = ~new_n14144_ | ~new_n14049_;
  assign new_n14146_ = ~new_n2001_ | ~new_n2430_;
  assign new_n14147_ = ~new_n13981_;
  assign new_n14148_ = new_n1996_ | new_n2436_;
  assign new_n14149_ = new_n2000_ | new_n2433_;
  assign new_n14150_ = ~new_n13948_;
  assign new_n14151_ = ~new_n13949_ | ~new_n13948_;
  assign new_n14152_ = ~new_n1996_ | ~new_n14151_;
  assign new_n14153_ = ~new_n2436_ | ~new_n14150_;
  assign new_n14154_ = ~new_n13897_ | ~new_n13981_;
  assign new_n14155_ = ~new_n14047_;
  assign new_n14156_ = new_n2003_ | new_n2952_;
  assign new_n14157_ = new_n2008_ | new_n2441_;
  assign new_n14158_ = new_n2002_ | new_n2951_;
  assign new_n14159_ = ~new_n13969_;
  assign new_n14160_ = ~new_n2952_ | ~new_n14159_;
  assign new_n14161_ = ~new_n14160_ | ~new_n13979_;
  assign new_n14162_ = ~new_n13969_ | ~new_n13970_;
  assign new_n14163_ = ~new_n14162_ | ~new_n14161_;
  assign new_n14164_ = ~new_n14060_ | ~new_n13898_;
  assign new_n14165_ = ~new_n2002_ | ~new_n2951_;
  assign new_n14166_ = ~new_n14163_ | ~new_n14164_;
  assign new_n14167_ = new_n2439_ | new_n2009_;
  assign new_n14168_ = new_n2951_ | new_n2002_;
  assign new_n14169_ = ~new_n14018_ | ~new_n14158_ | ~new_n14047_;
  assign new_n14170_ = ~new_n14168_ | ~new_n14166_;
  assign new_n14171_ = ~new_n14043_;
  assign new_n14172_ = new_n2950_ | new_n1988_;
  assign new_n14173_ = ~new_n14172_ | ~new_n14043_;
  assign new_n14174_ = ~new_n1988_ | ~new_n2950_;
  assign new_n14175_ = ~new_n14041_;
  assign new_n14176_ = new_n2949_ | new_n1993_;
  assign new_n14177_ = ~new_n14176_ | ~new_n14041_;
  assign new_n14178_ = ~new_n1993_ | ~new_n2949_;
  assign new_n14179_ = ~new_n14039_;
  assign new_n14180_ = new_n1985_ | new_n2947_;
  assign new_n14181_ = ~new_n14061_ | ~new_n14058_;
  assign new_n14182_ = ~new_n13975_;
  assign new_n14183_ = new_n2948_ | new_n1992_;
  assign new_n14184_ = ~new_n14053_ | ~new_n14039_ | ~new_n14183_;
  assign new_n14185_ = ~new_n14037_;
  assign new_n14186_ = new_n2945_ | new_n1980_;
  assign new_n14187_ = ~new_n1980_ | ~new_n2945_;
  assign new_n14188_ = ~new_n14035_;
  assign new_n14189_ = ~new_n2944_ | ~new_n14035_;
  assign new_n14190_ = ~new_n14033_;
  assign new_n14191_ = ~new_n14183_ | ~new_n14039_;
  assign new_n14192_ = ~new_n13978_;
  assign new_n14193_ = new_n2947_ | new_n1985_;
  assign new_n14194_ = ~new_n14193_ | ~new_n13978_;
  assign new_n14195_ = ~new_n14038_ | ~new_n14194_ | ~new_n14058_;
  assign new_n14196_ = ~new_n14192_ | ~new_n14058_;
  assign new_n14197_ = ~new_n2946_ | ~new_n1984_;
  assign new_n14198_ = ~new_n14053_ | ~new_n14196_ | ~new_n14197_;
  assign new_n14199_ = new_n1985_ | new_n2947_;
  assign new_n14200_ = ~new_n14167_ | ~new_n14047_;
  assign new_n14201_ = ~new_n13980_;
  assign new_n14202_ = ~new_n13898_ | ~new_n13980_;
  assign new_n14203_ = ~new_n14022_ | ~new_n14202_;
  assign new_n14204_ = ~new_n14202_ | ~new_n14163_;
  assign new_n14205_ = ~new_n14338_ | ~new_n14204_;
  assign new_n14206_ = new_n2441_ | new_n2008_;
  assign new_n14207_ = ~new_n14206_ | ~new_n13980_;
  assign new_n14208_ = ~new_n14045_ | ~new_n14207_ | ~new_n13969_;
  assign new_n14209_ = ~new_n14201_ | ~new_n13969_;
  assign new_n14210_ = ~new_n2003_ | ~new_n2952_;
  assign new_n14211_ = ~new_n13898_ | ~new_n14210_ | ~new_n14209_;
  assign new_n14212_ = new_n2388_ | new_n2005_;
  assign new_n14213_ = ~new_n14046_;
  assign new_n14214_ = new_n2008_ | new_n2441_;
  assign new_n14215_ = new_n2433_ | new_n2000_;
  assign new_n14216_ = ~new_n14215_ | ~new_n13981_;
  assign new_n14217_ = ~new_n14023_ | ~new_n14216_;
  assign new_n14218_ = ~new_n14147_ | ~new_n13948_;
  assign new_n14219_ = ~new_n2436_ | ~new_n1996_;
  assign new_n14220_ = ~new_n13897_ | ~new_n14219_ | ~new_n14218_;
  assign new_n14221_ = new_n2000_ | new_n2433_;
  assign new_n14222_ = ~new_n14135_ | ~new_n14052_;
  assign new_n14223_ = ~new_n13982_;
  assign new_n14224_ = new_n2421_ | new_n1999_;
  assign new_n14225_ = ~new_n14224_ | ~new_n13982_;
  assign new_n14226_ = ~new_n14024_ | ~new_n14225_;
  assign new_n14227_ = ~new_n14223_ | ~new_n14057_;
  assign new_n14228_ = ~new_n2007_ | ~new_n2424_;
  assign new_n14229_ = ~new_n14025_ | ~new_n14227_;
  assign new_n14230_ = new_n1999_ | new_n2421_;
  assign new_n14231_ = new_n2412_ | new_n2010_;
  assign new_n14232_ = ~new_n14231_ | ~new_n13929_;
  assign new_n14233_ = ~new_n14026_ | ~new_n14232_;
  assign new_n14234_ = ~new_n14091_ | ~new_n14056_;
  assign new_n14235_ = ~new_n1989_ | ~new_n2415_;
  assign new_n14236_ = ~new_n14027_ | ~new_n14234_;
  assign new_n14237_ = ~new_n14092_ | ~new_n14056_;
  assign new_n14238_ = ~new_n14089_ | ~new_n13950_;
  assign new_n14239_ = ~new_n14099_ | ~new_n13911_;
  assign new_n14240_ = ~new_n14113_ | ~new_n13923_;
  assign new_n14241_ = ~new_n14116_ | ~new_n14065_;
  assign new_n14242_ = ~new_n14199_ | ~new_n14058_;
  assign new_n14243_ = ~new_n14183_ | ~new_n14061_;
  assign new_n14244_ = ~new_n14214_ | ~new_n13969_;
  assign new_n14245_ = ~new_n14167_ | ~new_n13966_;
  assign new_n14246_ = ~new_n14221_ | ~new_n13948_;
  assign new_n14247_ = ~new_n14230_ | ~new_n14057_;
  assign new_n14248_ = ~new_n14135_ | ~new_n13957_;
  assign new_n14249_ = ~new_n2944_ | ~new_n1981_;
  assign new_n14250_ = ~new_n14181_ | ~new_n14053_;
  assign new_n14251_ = ~new_n1984_ | ~new_n14180_;
  assign new_n14252_ = ~new_n2946_ | ~new_n14180_;
  assign new_n14253_ = ~new_n14186_ | ~new_n14181_ | ~new_n14053_;
  assign new_n14254_ = ~new_n14020_ | ~new_n14039_ | ~new_n14053_;
  assign new_n14255_ = ~new_n14182_ | ~new_n14186_;
  assign new_n14256_ = ~new_n2010_ | ~new_n13928_;
  assign new_n14257_ = ~new_n2412_ | ~new_n13927_;
  assign new_n14258_ = ~new_n14257_ | ~new_n14256_;
  assign new_n14259_ = ~new_n14237_ | ~new_n13929_;
  assign new_n14260_ = ~new_n14258_ | ~new_n14091_;
  assign new_n14261_ = ~new_n2011_ | ~new_n13925_;
  assign new_n14262_ = ~new_n2409_ | ~new_n13926_;
  assign new_n14263_ = ~new_n14262_ | ~new_n14261_;
  assign new_n14264_ = ~new_n14238_ | ~new_n14028_;
  assign new_n14265_ = ~new_n14088_ | ~new_n14263_;
  assign new_n14266_ = ~new_n1997_ | ~new_n13912_;
  assign new_n14267_ = ~new_n2406_ | ~new_n13910_;
  assign new_n14268_ = ~new_n1998_ | ~new_n13908_;
  assign new_n14269_ = ~new_n2403_ | ~new_n13909_;
  assign new_n14270_ = ~new_n14269_ | ~new_n14268_;
  assign new_n14271_ = ~new_n14239_ | ~new_n13930_;
  assign new_n14272_ = ~new_n14270_ | ~new_n14080_;
  assign new_n14273_ = ~new_n1994_ | ~new_n13924_;
  assign new_n14274_ = ~new_n2400_ | ~new_n13915_;
  assign new_n14275_ = ~new_n1987_ | ~new_n13913_;
  assign new_n14276_ = ~new_n2397_ | ~new_n13914_;
  assign new_n14277_ = ~new_n14276_ | ~new_n14275_;
  assign new_n14278_ = ~new_n14240_ | ~new_n13933_;
  assign new_n14279_ = ~new_n14277_ | ~new_n14106_;
  assign new_n14280_ = ~new_n1991_ | ~new_n13921_;
  assign new_n14281_ = ~new_n2394_ | ~new_n13922_;
  assign new_n14282_ = ~new_n14281_ | ~new_n14280_;
  assign new_n14283_ = ~new_n14241_ | ~new_n14029_;
  assign new_n14284_ = ~new_n14115_ | ~new_n14282_;
  assign new_n14285_ = ~new_n1995_ | ~new_n13916_;
  assign new_n14286_ = ~new_n2391_ | ~new_n13917_;
  assign new_n14287_ = ~new_n1982_ | ~new_n14031_;
  assign new_n14288_ = ~new_n2955_ | ~new_n14030_;
  assign new_n14289_ = ~new_n1982_ | ~new_n14031_;
  assign new_n14290_ = ~new_n2955_ | ~new_n14030_;
  assign new_n14291_ = ~new_n14290_ | ~new_n14289_;
  assign new_n14292_ = ~new_n14032_ | ~new_n14033_;
  assign new_n14293_ = ~new_n14190_ | ~new_n14291_;
  assign new_n14294_ = ~new_n1981_ | ~new_n13977_;
  assign new_n14295_ = ~new_n2944_ | ~new_n13976_;
  assign new_n14296_ = ~new_n1981_ | ~new_n13977_;
  assign new_n14297_ = ~new_n2944_ | ~new_n13976_;
  assign new_n14298_ = ~new_n14297_ | ~new_n14296_;
  assign new_n14299_ = ~new_n14034_ | ~new_n14035_;
  assign new_n14300_ = ~new_n14188_ | ~new_n14298_;
  assign new_n14301_ = ~new_n1980_ | ~new_n13935_;
  assign new_n14302_ = ~new_n2945_ | ~new_n13936_;
  assign new_n14303_ = ~new_n1980_ | ~new_n13935_;
  assign new_n14304_ = ~new_n2945_ | ~new_n13936_;
  assign new_n14305_ = ~new_n14304_ | ~new_n14303_;
  assign new_n14306_ = ~new_n14036_ | ~new_n14037_;
  assign new_n14307_ = ~new_n14185_ | ~new_n14305_;
  assign new_n14308_ = ~new_n1984_ | ~new_n13938_;
  assign new_n14309_ = ~new_n2946_ | ~new_n13937_;
  assign new_n14310_ = ~new_n1985_ | ~new_n13939_;
  assign new_n14311_ = ~new_n2947_ | ~new_n13940_;
  assign new_n14312_ = ~new_n14311_ | ~new_n14310_;
  assign new_n14313_ = ~new_n14242_ | ~new_n13978_;
  assign new_n14314_ = ~new_n14312_ | ~new_n14192_;
  assign new_n14315_ = ~new_n1992_ | ~new_n13941_;
  assign new_n14316_ = ~new_n2948_ | ~new_n13942_;
  assign new_n14317_ = ~new_n14316_ | ~new_n14315_;
  assign new_n14318_ = ~new_n14243_ | ~new_n14039_;
  assign new_n14319_ = ~new_n14179_ | ~new_n14317_;
  assign new_n14320_ = ~new_n1993_ | ~new_n13973_;
  assign new_n14321_ = ~new_n2949_ | ~new_n13974_;
  assign new_n14322_ = ~new_n1993_ | ~new_n13973_;
  assign new_n14323_ = ~new_n2949_ | ~new_n13974_;
  assign new_n14324_ = ~new_n14323_ | ~new_n14322_;
  assign new_n14325_ = ~new_n14040_ | ~new_n14041_;
  assign new_n14326_ = ~new_n14175_ | ~new_n14324_;
  assign new_n14327_ = ~new_n1988_ | ~new_n13971_;
  assign new_n14328_ = ~new_n2950_ | ~new_n13972_;
  assign new_n14329_ = ~new_n1988_ | ~new_n13971_;
  assign new_n14330_ = ~new_n2950_ | ~new_n13972_;
  assign new_n14331_ = ~new_n14330_ | ~new_n14329_;
  assign new_n14332_ = ~new_n14042_ | ~new_n14043_;
  assign new_n14333_ = ~new_n14171_ | ~new_n14331_;
  assign new_n14334_ = ~new_n2002_ | ~new_n13943_;
  assign new_n14335_ = ~new_n2951_ | ~new_n13944_;
  assign new_n14336_ = ~new_n2002_ | ~new_n13943_;
  assign new_n14337_ = ~new_n2951_ | ~new_n13944_;
  assign new_n14338_ = ~new_n14337_ | ~new_n14336_;
  assign new_n14339_ = ~new_n2003_ | ~new_n13970_;
  assign new_n14340_ = ~new_n2952_ | ~new_n13979_;
  assign new_n14341_ = ~new_n14067_ | ~new_n14046_;
  assign new_n14342_ = ~new_n14213_ | ~new_n13920_;
  assign new_n14343_ = ~new_n2008_ | ~new_n13967_;
  assign new_n14344_ = ~new_n2441_ | ~new_n13968_;
  assign new_n14345_ = ~new_n14344_ | ~new_n14343_;
  assign new_n14346_ = ~new_n14244_ | ~new_n13980_;
  assign new_n14347_ = ~new_n14345_ | ~new_n14201_;
  assign new_n14348_ = ~new_n2009_ | ~new_n13964_;
  assign new_n14349_ = ~new_n2439_ | ~new_n13965_;
  assign new_n14350_ = ~new_n14349_ | ~new_n14348_;
  assign new_n14351_ = ~new_n14245_ | ~new_n14047_;
  assign new_n14352_ = ~new_n14155_ | ~new_n14350_;
  assign new_n14353_ = ~new_n1996_ | ~new_n13949_;
  assign new_n14354_ = ~new_n2436_ | ~new_n13947_;
  assign new_n14355_ = ~new_n2000_ | ~new_n13945_;
  assign new_n14356_ = ~new_n2433_ | ~new_n13946_;
  assign new_n14357_ = ~new_n14356_ | ~new_n14355_;
  assign new_n14358_ = ~new_n14246_ | ~new_n13981_;
  assign new_n14359_ = ~new_n14357_ | ~new_n14147_;
  assign new_n14360_ = ~new_n2001_ | ~new_n13962_;
  assign new_n14361_ = ~new_n2430_ | ~new_n13963_;
  assign new_n14362_ = ~new_n2001_ | ~new_n13962_;
  assign new_n14363_ = ~new_n2430_ | ~new_n13963_;
  assign new_n14364_ = ~new_n14363_ | ~new_n14362_;
  assign new_n14365_ = ~new_n14048_ | ~new_n14049_;
  assign new_n14366_ = ~new_n14143_ | ~new_n14364_;
  assign new_n14367_ = ~new_n2006_ | ~new_n13960_;
  assign new_n14368_ = ~new_n2427_ | ~new_n13961_;
  assign new_n14369_ = ~new_n2006_ | ~new_n13960_;
  assign new_n14370_ = ~new_n2427_ | ~new_n13961_;
  assign new_n14371_ = ~new_n14370_ | ~new_n14369_;
  assign new_n14372_ = ~new_n14050_ | ~new_n14051_;
  assign new_n14373_ = ~new_n14139_ | ~new_n14371_;
  assign new_n14374_ = ~new_n2007_ | ~new_n13958_;
  assign new_n14375_ = ~new_n2424_ | ~new_n13959_;
  assign new_n14376_ = ~new_n1999_ | ~new_n13953_;
  assign new_n14377_ = ~new_n2421_ | ~new_n13954_;
  assign new_n14378_ = ~new_n14377_ | ~new_n14376_;
  assign new_n14379_ = ~new_n14247_ | ~new_n13982_;
  assign new_n14380_ = ~new_n14378_ | ~new_n14223_;
  assign new_n14381_ = ~new_n1990_ | ~new_n13955_;
  assign new_n14382_ = ~new_n2418_ | ~new_n13956_;
  assign new_n14383_ = ~new_n14382_ | ~new_n14381_;
  assign new_n14384_ = ~new_n14248_ | ~new_n14052_;
  assign new_n14385_ = ~new_n14129_ | ~new_n14383_;
  assign new_n14386_ = ~new_n1989_ | ~new_n13951_;
  assign new_n14387_ = ~new_n2415_ | ~new_n13952_;
  assign new_n14388_ = ~new_n2004_ | ~new_n13918_;
  assign new_n14389_ = ~new_n2383_ | ~new_n13919_;
  assign new_n14390_ = new_n14481_ & new_n14480_;
  assign new_n14391_ = new_n14482_ & new_n14483_;
  assign new_n14392_ = new_n14499_ & new_n14498_;
  assign new_n14393_ = new_n14541_ & new_n14540_;
  assign new_n14394_ = new_n14550_ & new_n14549_;
  assign new_n14395_ = new_n14568_ & new_n14567_;
  assign new_n14396_ = new_n14604_ & new_n14601_;
  assign new_n14397_ = new_n14597_ & new_n14594_;
  assign new_n14398_ = new_n14588_ & new_n14585_;
  assign new_n14399_ = new_n14582_ & new_n14578_;
  assign new_n14400_ = new_n14537_ & new_n14534_;
  assign new_n14401_ = new_n14529_ & new_n14526_;
  assign new_n14402_ = new_n14515_ & new_n14512_;
  assign new_n14403_ = ~pi135;
  assign new_n14404_ = ~new_n2402_;
  assign new_n14405_ = ~new_n2405_;
  assign new_n14406_ = ~new_n2402_ | ~pi135;
  assign new_n14407_ = ~pi136;
  assign new_n14408_ = ~pi133;
  assign new_n14409_ = ~new_n2396_;
  assign new_n14410_ = ~new_n2399_;
  assign new_n14411_ = ~pi131;
  assign new_n14412_ = ~new_n2390_;
  assign new_n14413_ = ~pi129;
  assign new_n14414_ = ~new_n2381_;
  assign new_n14415_ = ~new_n2381_ | ~pi129;
  assign new_n14416_ = ~pi132;
  assign new_n14417_ = ~new_n2393_;
  assign new_n14418_ = ~new_n2396_ | ~pi133;
  assign new_n14419_ = ~pi134;
  assign new_n14420_ = ~pi137;
  assign new_n14421_ = ~new_n2408_;
  assign new_n14422_ = ~new_n2411_;
  assign new_n14423_ = ~pi138;
  assign new_n14424_ = ~new_n14435_ | ~new_n14507_;
  assign new_n14425_ = ~new_n14495_ | ~new_n14496_ | ~new_n14494_;
  assign new_n14426_ = ~new_n14484_ | ~new_n14485_;
  assign new_n14427_ = ~pi130 | ~new_n2387_;
  assign new_n14428_ = ~new_n14521_ | ~new_n14522_ | ~new_n14520_;
  assign new_n14429_ = ~new_n14518_ | ~new_n14517_;
  assign new_n14430_ = ~pi145;
  assign new_n14431_ = ~new_n2432_;
  assign new_n14432_ = ~new_n2435_;
  assign new_n14433_ = ~new_n2432_ | ~pi145;
  assign new_n14434_ = ~pi146;
  assign new_n14435_ = ~new_n2408_ | ~pi137;
  assign new_n14436_ = ~pi139;
  assign new_n14437_ = ~new_n2414_;
  assign new_n14438_ = ~pi141;
  assign new_n14439_ = ~new_n2420_;
  assign new_n14440_ = ~pi140;
  assign new_n14441_ = ~new_n2417_;
  assign new_n14442_ = ~new_n2417_ | ~pi140;
  assign new_n14443_ = ~pi142;
  assign new_n14444_ = ~new_n2423_;
  assign new_n14445_ = ~pi143;
  assign new_n14446_ = ~new_n2426_;
  assign new_n14447_ = ~pi144;
  assign new_n14448_ = ~new_n2429_;
  assign new_n14449_ = ~pi147;
  assign new_n14450_ = ~new_n2438_;
  assign new_n14451_ = ~new_n14573_ | ~new_n14572_ | ~new_n14571_;
  assign new_n14452_ = ~new_n14565_ | ~new_n14564_;
  assign new_n14453_ = ~new_n14442_ | ~new_n14590_;
  assign new_n14454_ = ~new_n14645_ | ~new_n14644_;
  assign new_n14455_ = ~new_n14694_ | ~new_n14693_;
  assign new_n14456_ = ~new_n14617_ | ~new_n14616_;
  assign new_n14457_ = ~new_n14622_ | ~new_n14621_;
  assign new_n14458_ = ~new_n14629_ | ~new_n14628_;
  assign new_n14459_ = ~new_n14636_ | ~new_n14635_;
  assign new_n14460_ = ~new_n14641_ | ~new_n14640_;
  assign new_n14461_ = ~new_n14657_ | ~new_n14656_;
  assign new_n14462_ = ~new_n14664_ | ~new_n14663_;
  assign new_n14463_ = ~new_n14671_ | ~new_n14670_;
  assign new_n14464_ = ~new_n14678_ | ~new_n14677_;
  assign new_n14465_ = ~new_n14685_ | ~new_n14684_;
  assign new_n14466_ = ~new_n14690_ | ~new_n14689_;
  assign new_n14467_ = ~new_n14504_ | ~new_n14503_ | ~new_n14502_;
  assign new_n14468_ = ~new_n14519_ | ~new_n14531_;
  assign new_n14469_ = ~new_n14427_ | ~new_n14538_;
  assign new_n14470_ = ~new_n2379_;
  assign new_n14471_ = ~pi148;
  assign new_n14472_ = ~new_n14561_ | ~new_n14560_;
  assign new_n14473_ = ~new_n14557_ | ~new_n14556_;
  assign new_n14474_ = ~new_n14547_ | ~new_n14546_;
  assign new_n14475_ = ~new_n14418_;
  assign new_n14476_ = ~pi138 | ~new_n2411_;
  assign new_n14477_ = ~new_n2420_ | ~pi141;
  assign new_n14478_ = ~new_n14442_;
  assign new_n14479_ = ~new_n14435_;
  assign new_n14480_ = new_n2399_ | pi134;
  assign new_n14481_ = new_n2396_ | pi133;
  assign new_n14482_ = pi132 | new_n2393_;
  assign new_n14483_ = pi131 | new_n2390_;
  assign new_n14484_ = ~new_n14415_;
  assign new_n14485_ = pi130 | new_n2387_;
  assign new_n14486_ = ~new_n14426_;
  assign new_n14487_ = ~new_n14427_;
  assign new_n14488_ = ~new_n14426_ | ~new_n14427_;
  assign new_n14489_ = ~new_n14482_ | ~pi131 | ~new_n2390_;
  assign new_n14490_ = ~new_n14391_ | ~new_n14488_;
  assign new_n14491_ = ~new_n2393_ | ~pi132;
  assign new_n14492_ = ~new_n14490_ | ~new_n14491_ | ~new_n14489_;
  assign new_n14493_ = ~new_n14419_ | ~new_n14418_;
  assign new_n14494_ = ~new_n2399_ | ~new_n14493_;
  assign new_n14495_ = ~new_n14390_ | ~new_n14492_;
  assign new_n14496_ = ~pi134 | ~new_n14475_;
  assign new_n14497_ = ~new_n14425_;
  assign new_n14498_ = new_n2405_ | pi136;
  assign new_n14499_ = new_n2402_ | pi135;
  assign new_n14500_ = ~new_n14406_;
  assign new_n14501_ = ~new_n14407_ | ~new_n14406_;
  assign new_n14502_ = ~new_n2405_ | ~new_n14501_;
  assign new_n14503_ = ~pi136 | ~new_n14500_;
  assign new_n14504_ = ~new_n14392_ | ~new_n14425_;
  assign new_n14505_ = ~new_n14467_;
  assign new_n14506_ = pi137 | new_n2408_;
  assign new_n14507_ = ~new_n14506_ | ~new_n14467_;
  assign new_n14508_ = ~new_n14424_;
  assign new_n14509_ = new_n2411_ | pi138;
  assign new_n14510_ = pi135 | new_n2402_;
  assign new_n14511_ = ~new_n14510_ | ~new_n14425_;
  assign new_n14512_ = ~new_n14623_ | ~new_n14511_ | ~new_n14406_ | ~new_n14624_;
  assign new_n14513_ = ~new_n14497_ | ~new_n14406_;
  assign new_n14514_ = ~pi136 | ~new_n2405_;
  assign new_n14515_ = ~new_n14513_ | ~new_n14514_ | ~new_n14392_;
  assign new_n14516_ = new_n2402_ | pi135;
  assign new_n14517_ = ~new_n14487_ | ~new_n14483_;
  assign new_n14518_ = ~new_n2390_ | ~pi131;
  assign new_n14519_ = ~new_n14429_;
  assign new_n14520_ = ~new_n14486_ | ~new_n14391_;
  assign new_n14521_ = ~new_n14429_ | ~new_n14482_;
  assign new_n14522_ = ~new_n2393_ | ~pi132;
  assign new_n14523_ = ~new_n14428_;
  assign new_n14524_ = pi133 | new_n2396_;
  assign new_n14525_ = ~new_n14524_ | ~new_n14428_;
  assign new_n14526_ = ~new_n14630_ | ~new_n14525_ | ~new_n14418_ | ~new_n14631_;
  assign new_n14527_ = ~new_n14523_ | ~new_n14418_;
  assign new_n14528_ = ~pi134 | ~new_n2399_;
  assign new_n14529_ = ~new_n14527_ | ~new_n14528_ | ~new_n14390_;
  assign new_n14530_ = new_n2396_ | pi133;
  assign new_n14531_ = ~new_n14486_ | ~new_n14483_;
  assign new_n14532_ = ~new_n14468_;
  assign new_n14533_ = ~new_n2393_ | ~pi132;
  assign new_n14534_ = ~new_n14642_ | ~new_n14426_ | ~new_n14427_ | ~new_n14643_;
  assign new_n14535_ = ~new_n14427_ | ~new_n14426_;
  assign new_n14536_ = ~new_n2390_ | ~pi131;
  assign new_n14537_ = ~new_n14535_ | ~new_n14536_ | ~new_n14483_;
  assign new_n14538_ = pi130 | new_n2387_;
  assign new_n14539_ = ~new_n14469_;
  assign new_n14540_ = new_n2411_ | pi138;
  assign new_n14541_ = new_n2414_ | pi139;
  assign new_n14542_ = ~new_n14479_ | ~new_n14393_;
  assign new_n14543_ = ~new_n2414_ | ~pi139;
  assign new_n14544_ = ~new_n14542_ | ~new_n14543_ | ~new_n14476_;
  assign new_n14545_ = pi139 | new_n2414_;
  assign new_n14546_ = ~new_n14467_ | ~new_n14506_ | ~new_n14393_;
  assign new_n14547_ = ~new_n14545_ | ~new_n14544_;
  assign new_n14548_ = ~new_n14474_;
  assign new_n14549_ = new_n2423_ | pi142;
  assign new_n14550_ = new_n2420_ | pi141;
  assign new_n14551_ = ~new_n14478_ | ~new_n14394_;
  assign new_n14552_ = ~new_n2423_ | ~pi142;
  assign new_n14553_ = ~new_n14551_ | ~new_n14552_ | ~new_n14477_;
  assign new_n14554_ = pi140 | new_n2417_;
  assign new_n14555_ = pi142 | new_n2423_;
  assign new_n14556_ = ~new_n14474_ | ~new_n14554_ | ~new_n14394_;
  assign new_n14557_ = ~new_n14555_ | ~new_n14553_;
  assign new_n14558_ = ~new_n14473_;
  assign new_n14559_ = pi143 | new_n2426_;
  assign new_n14560_ = ~new_n14559_ | ~new_n14473_;
  assign new_n14561_ = ~new_n2426_ | ~pi143;
  assign new_n14562_ = ~new_n14472_;
  assign new_n14563_ = pi144 | new_n2429_;
  assign new_n14564_ = ~new_n14563_ | ~new_n14472_;
  assign new_n14565_ = ~new_n2429_ | ~pi144;
  assign new_n14566_ = ~new_n14452_;
  assign new_n14567_ = new_n2435_ | pi146;
  assign new_n14568_ = new_n2432_ | pi145;
  assign new_n14569_ = ~new_n14433_;
  assign new_n14570_ = ~new_n14434_ | ~new_n14433_;
  assign new_n14571_ = ~new_n2435_ | ~new_n14570_;
  assign new_n14572_ = ~pi146 | ~new_n14569_;
  assign new_n14573_ = ~new_n14395_ | ~new_n14452_;
  assign new_n14574_ = ~new_n14451_;
  assign new_n14575_ = pi147 | new_n2438_;
  assign new_n14576_ = ~new_n14575_ | ~new_n14451_;
  assign new_n14577_ = ~new_n2438_ | ~pi147;
  assign new_n14578_ = ~new_n14646_ | ~new_n14576_ | ~new_n14577_ | ~new_n14647_;
  assign new_n14579_ = ~new_n2438_ | ~pi147;
  assign new_n14580_ = ~new_n14574_ | ~new_n14579_;
  assign new_n14581_ = new_n2438_ | pi147;
  assign new_n14582_ = ~new_n14580_ | ~new_n14581_ | ~new_n14650_;
  assign new_n14583_ = pi145 | new_n2432_;
  assign new_n14584_ = ~new_n14583_ | ~new_n14452_;
  assign new_n14585_ = ~new_n14658_ | ~new_n14584_ | ~new_n14433_ | ~new_n14659_;
  assign new_n14586_ = ~new_n14566_ | ~new_n14433_;
  assign new_n14587_ = ~pi146 | ~new_n2435_;
  assign new_n14588_ = ~new_n14586_ | ~new_n14587_ | ~new_n14395_;
  assign new_n14589_ = new_n2432_ | pi145;
  assign new_n14590_ = ~new_n14554_ | ~new_n14474_;
  assign new_n14591_ = ~new_n14453_;
  assign new_n14592_ = pi141 | new_n2420_;
  assign new_n14593_ = ~new_n14592_ | ~new_n14453_;
  assign new_n14594_ = ~new_n14679_ | ~new_n14593_ | ~new_n14477_ | ~new_n14680_;
  assign new_n14595_ = ~new_n14591_ | ~new_n14477_;
  assign new_n14596_ = ~new_n2423_ | ~pi142;
  assign new_n14597_ = ~new_n14595_ | ~new_n14596_ | ~new_n14394_;
  assign new_n14598_ = new_n2420_ | pi141;
  assign new_n14599_ = pi138 | new_n2411_;
  assign new_n14600_ = ~new_n14599_ | ~new_n14424_;
  assign new_n14601_ = ~new_n14691_ | ~new_n14600_ | ~new_n14476_ | ~new_n14692_;
  assign new_n14602_ = ~new_n14508_ | ~new_n14476_;
  assign new_n14603_ = ~new_n2414_ | ~pi139;
  assign new_n14604_ = ~new_n14602_ | ~new_n14603_ | ~new_n14393_;
  assign new_n14605_ = ~new_n14509_ | ~new_n14476_;
  assign new_n14606_ = ~new_n14506_ | ~new_n14435_;
  assign new_n14607_ = ~new_n14516_ | ~new_n14406_;
  assign new_n14608_ = ~new_n14530_ | ~new_n14418_;
  assign new_n14609_ = ~new_n14533_ | ~new_n14482_;
  assign new_n14610_ = ~new_n14589_ | ~new_n14433_;
  assign new_n14611_ = ~new_n14598_ | ~new_n14477_;
  assign new_n14612_ = ~new_n14554_ | ~new_n14442_;
  assign new_n14613_ = ~new_n2411_ | ~new_n14423_;
  assign new_n14614_ = ~pi138 | ~new_n14422_;
  assign new_n14615_ = ~new_n14614_ | ~new_n14613_;
  assign new_n14616_ = ~new_n14605_ | ~new_n14424_;
  assign new_n14617_ = ~new_n14615_ | ~new_n14508_;
  assign new_n14618_ = ~new_n2408_ | ~new_n14420_;
  assign new_n14619_ = ~pi137 | ~new_n14421_;
  assign new_n14620_ = ~new_n14619_ | ~new_n14618_;
  assign new_n14621_ = ~new_n14606_ | ~new_n14467_;
  assign new_n14622_ = ~new_n14505_ | ~new_n14620_;
  assign new_n14623_ = ~new_n2405_ | ~new_n14407_;
  assign new_n14624_ = ~pi136 | ~new_n14405_;
  assign new_n14625_ = ~new_n2402_ | ~new_n14403_;
  assign new_n14626_ = ~pi135 | ~new_n14404_;
  assign new_n14627_ = ~new_n14626_ | ~new_n14625_;
  assign new_n14628_ = ~new_n14607_ | ~new_n14425_;
  assign new_n14629_ = ~new_n14627_ | ~new_n14497_;
  assign new_n14630_ = ~new_n2399_ | ~new_n14419_;
  assign new_n14631_ = ~pi134 | ~new_n14410_;
  assign new_n14632_ = ~new_n2396_ | ~new_n14408_;
  assign new_n14633_ = ~pi133 | ~new_n14409_;
  assign new_n14634_ = ~new_n14633_ | ~new_n14632_;
  assign new_n14635_ = ~new_n14608_ | ~new_n14428_;
  assign new_n14636_ = ~new_n14634_ | ~new_n14523_;
  assign new_n14637_ = ~new_n2393_ | ~new_n14416_;
  assign new_n14638_ = ~pi132 | ~new_n14417_;
  assign new_n14639_ = ~new_n14638_ | ~new_n14637_;
  assign new_n14640_ = ~new_n14609_ | ~new_n14468_;
  assign new_n14641_ = ~new_n14532_ | ~new_n14639_;
  assign new_n14642_ = ~new_n2390_ | ~new_n14411_;
  assign new_n14643_ = ~pi131 | ~new_n14412_;
  assign new_n14644_ = ~new_n14484_ | ~new_n14469_;
  assign new_n14645_ = ~new_n14539_ | ~new_n14415_;
  assign new_n14646_ = ~new_n2379_ | ~new_n14471_;
  assign new_n14647_ = ~pi148 | ~new_n14470_;
  assign new_n14648_ = ~new_n2379_ | ~new_n14471_;
  assign new_n14649_ = ~pi148 | ~new_n14470_;
  assign new_n14650_ = ~new_n14649_ | ~new_n14648_;
  assign new_n14651_ = ~new_n2438_ | ~new_n14449_;
  assign new_n14652_ = ~pi147 | ~new_n14450_;
  assign new_n14653_ = ~new_n2438_ | ~new_n14449_;
  assign new_n14654_ = ~pi147 | ~new_n14450_;
  assign new_n14655_ = ~new_n14654_ | ~new_n14653_;
  assign new_n14656_ = ~new_n14451_ | ~new_n14652_ | ~new_n14651_;
  assign new_n14657_ = ~new_n14655_ | ~new_n14574_;
  assign new_n14658_ = ~new_n2435_ | ~new_n14434_;
  assign new_n14659_ = ~pi146 | ~new_n14432_;
  assign new_n14660_ = ~new_n2432_ | ~new_n14430_;
  assign new_n14661_ = ~pi145 | ~new_n14431_;
  assign new_n14662_ = ~new_n14661_ | ~new_n14660_;
  assign new_n14663_ = ~new_n14610_ | ~new_n14452_;
  assign new_n14664_ = ~new_n14662_ | ~new_n14566_;
  assign new_n14665_ = ~new_n2429_ | ~new_n14447_;
  assign new_n14666_ = ~pi144 | ~new_n14448_;
  assign new_n14667_ = ~new_n2429_ | ~new_n14447_;
  assign new_n14668_ = ~pi144 | ~new_n14448_;
  assign new_n14669_ = ~new_n14668_ | ~new_n14667_;
  assign new_n14670_ = ~new_n14472_ | ~new_n14666_ | ~new_n14665_;
  assign new_n14671_ = ~new_n14562_ | ~new_n14669_;
  assign new_n14672_ = ~new_n2426_ | ~new_n14445_;
  assign new_n14673_ = ~pi143 | ~new_n14446_;
  assign new_n14674_ = ~new_n2426_ | ~new_n14445_;
  assign new_n14675_ = ~pi143 | ~new_n14446_;
  assign new_n14676_ = ~new_n14675_ | ~new_n14674_;
  assign new_n14677_ = ~new_n14473_ | ~new_n14673_ | ~new_n14672_;
  assign new_n14678_ = ~new_n14558_ | ~new_n14676_;
  assign new_n14679_ = ~new_n2423_ | ~new_n14443_;
  assign new_n14680_ = ~pi142 | ~new_n14444_;
  assign new_n14681_ = ~new_n2420_ | ~new_n14438_;
  assign new_n14682_ = ~pi141 | ~new_n14439_;
  assign new_n14683_ = ~new_n14682_ | ~new_n14681_;
  assign new_n14684_ = ~new_n14611_ | ~new_n14453_;
  assign new_n14685_ = ~new_n14683_ | ~new_n14591_;
  assign new_n14686_ = ~new_n2417_ | ~new_n14440_;
  assign new_n14687_ = ~pi140 | ~new_n14441_;
  assign new_n14688_ = ~new_n14687_ | ~new_n14686_;
  assign new_n14689_ = ~new_n14612_ | ~new_n14474_;
  assign new_n14690_ = ~new_n14548_ | ~new_n14688_;
  assign new_n14691_ = ~new_n2414_ | ~new_n14436_;
  assign new_n14692_ = ~pi139 | ~new_n14437_;
  assign new_n14693_ = ~new_n2381_ | ~new_n14413_;
  assign new_n14694_ = ~pi129 | ~new_n14414_;
  assign new_n14695_ = new_n14873_ & new_n14890_;
  assign new_n14696_ = new_n14892_ & new_n14891_;
  assign new_n14697_ = new_n14868_ & new_n14929_;
  assign new_n14698_ = new_n14931_ & new_n14930_;
  assign new_n14699_ = new_n14948_ & new_n14947_;
  assign new_n14700_ = new_n14974_ & new_n14973_;
  assign new_n14701_ = new_n15072_ & new_n15071_;
  assign new_n14702_ = ~new_n15029_ | ~new_n15032_;
  assign new_n14703_ = ~new_n15018_ | ~new_n15021_;
  assign new_n14704_ = ~new_n15007_ | ~new_n15010_;
  assign new_n14705_ = ~new_n14999_ | ~new_n15001_;
  assign new_n14706_ = ~new_n15037_ | ~new_n14845_ | ~new_n14864_;
  assign new_n14707_ = ~new_n14925_ | ~new_n14927_;
  assign new_n14708_ = ~new_n14917_ | ~new_n14920_;
  assign new_n14709_ = ~new_n14909_ | ~new_n14911_;
  assign new_n14710_ = ~new_n14714_ | ~new_n15035_;
  assign new_n14711_ = ~new_n2406_;
  assign new_n14712_ = ~new_n2391_;
  assign new_n14713_ = ~new_n2383_;
  assign new_n14714_ = ~new_n2383_ | ~new_n14782_;
  assign new_n14715_ = ~new_n2005_;
  assign new_n14716_ = ~new_n2394_;
  assign new_n14717_ = ~new_n1995_;
  assign new_n14718_ = ~new_n1995_ | ~new_n14712_;
  assign new_n14719_ = ~new_n1991_;
  assign new_n14720_ = ~new_n2403_;
  assign new_n14721_ = ~new_n2400_;
  assign new_n14722_ = ~new_n2397_;
  assign new_n14723_ = ~new_n1998_;
  assign new_n14724_ = ~new_n1994_;
  assign new_n14725_ = ~new_n1987_;
  assign new_n14726_ = ~new_n1987_ | ~new_n14722_;
  assign new_n14727_ = ~new_n2409_;
  assign new_n14728_ = ~new_n1997_;
  assign new_n14729_ = ~new_n1997_ | ~new_n14711_;
  assign new_n14730_ = ~new_n2011_;
  assign new_n14731_ = ~new_n2412_;
  assign new_n14732_ = ~new_n2010_;
  assign new_n14733_ = ~new_n14898_ | ~new_n14897_;
  assign new_n14734_ = ~new_n14726_ | ~new_n14913_;
  assign new_n14735_ = ~new_n14882_ | ~new_n14881_;
  assign new_n14736_ = ~new_n2946_;
  assign new_n14737_ = ~new_n2950_;
  assign new_n14738_ = ~new_n2430_;
  assign new_n14739_ = ~new_n2418_;
  assign new_n14740_ = ~new_n2415_;
  assign new_n14741_ = ~new_n1990_;
  assign new_n14742_ = ~new_n1989_;
  assign new_n14743_ = ~new_n2010_ | ~new_n14731_;
  assign new_n14744_ = ~new_n2421_;
  assign new_n14745_ = ~new_n1999_;
  assign new_n14746_ = ~new_n2424_;
  assign new_n14747_ = ~new_n2007_;
  assign new_n14748_ = ~new_n2433_;
  assign new_n14749_ = ~new_n2427_;
  assign new_n14750_ = ~new_n2000_;
  assign new_n14751_ = ~new_n2001_;
  assign new_n14752_ = ~new_n2006_;
  assign new_n14753_ = ~new_n2006_ | ~new_n14749_;
  assign new_n14754_ = ~new_n2436_;
  assign new_n14755_ = ~new_n1996_;
  assign new_n14756_ = ~new_n14958_ | ~new_n14957_;
  assign new_n14757_ = ~new_n2009_;
  assign new_n14758_ = ~new_n2441_;
  assign new_n14759_ = ~new_n2008_;
  assign new_n14760_ = ~new_n2952_;
  assign new_n14761_ = ~new_n2003_;
  assign new_n14762_ = ~new_n2949_;
  assign new_n14763_ = ~new_n2951_;
  assign new_n14764_ = ~new_n1993_;
  assign new_n14765_ = ~new_n1988_;
  assign new_n14766_ = ~new_n2002_;
  assign new_n14767_ = ~new_n2002_ | ~new_n14763_;
  assign new_n14768_ = ~new_n2948_;
  assign new_n14769_ = ~new_n1992_;
  assign new_n14770_ = ~new_n2947_;
  assign new_n14771_ = ~new_n1985_;
  assign new_n14772_ = ~new_n2945_;
  assign new_n14773_ = ~new_n1984_;
  assign new_n14774_ = ~new_n1984_ | ~new_n14736_;
  assign new_n14775_ = ~new_n1980_;
  assign new_n14776_ = ~new_n2944_;
  assign new_n14777_ = ~new_n1981_;
  assign new_n14778_ = ~new_n14988_ | ~new_n14987_;
  assign new_n14779_ = ~new_n14767_ | ~new_n15003_;
  assign new_n14780_ = ~new_n14753_ | ~new_n15014_;
  assign new_n14781_ = ~new_n14743_ | ~new_n15025_;
  assign new_n14782_ = ~new_n2004_;
  assign new_n14783_ = ~new_n15082_ | ~new_n15081_;
  assign new_n14784_ = ~new_n15096_ | ~new_n15095_;
  assign new_n14785_ = ~new_n15101_ | ~new_n15100_;
  assign new_n14786_ = ~new_n15117_ | ~new_n15116_;
  assign new_n14787_ = ~new_n15122_ | ~new_n15121_;
  assign new_n14788_ = ~new_n15127_ | ~new_n15126_;
  assign new_n14789_ = ~new_n15132_ | ~new_n15131_;
  assign new_n14790_ = ~new_n15137_ | ~new_n15136_;
  assign new_n14791_ = ~new_n15153_ | ~new_n15152_;
  assign new_n14792_ = ~new_n15158_ | ~new_n15157_;
  assign new_n14793_ = ~new_n15041_ | ~new_n15040_;
  assign new_n14794_ = ~new_n15050_ | ~new_n15049_;
  assign new_n14795_ = ~new_n15057_ | ~new_n15056_;
  assign new_n14796_ = ~new_n15061_ | ~new_n15060_;
  assign new_n14797_ = ~new_n15070_ | ~new_n15069_;
  assign new_n14798_ = ~new_n15091_ | ~new_n15090_;
  assign new_n14799_ = ~new_n15108_ | ~new_n15107_;
  assign new_n14800_ = ~new_n15112_ | ~new_n15111_;
  assign new_n14801_ = ~new_n15144_ | ~new_n15143_;
  assign new_n14802_ = ~new_n15148_ | ~new_n15147_;
  assign new_n14803_ = ~new_n15165_ | ~new_n15164_;
  assign new_n14804_ = new_n14884_ & new_n14872_;
  assign new_n14805_ = new_n14887_ & new_n14888_;
  assign new_n14806_ = new_n14900_ & new_n14874_;
  assign new_n14807_ = new_n14903_ & new_n14904_;
  assign new_n14808_ = new_n14729_ & new_n15043_ & new_n15042_;
  assign new_n14809_ = new_n15046_ & new_n14874_;
  assign new_n14810_ = new_n14919_ & new_n14696_;
  assign new_n14811_ = new_n15053_ & new_n14873_;
  assign new_n14812_ = new_n14718_ & new_n15063_ & new_n15062_;
  assign new_n14813_ = new_n15066_ & new_n14872_;
  assign new_n14814_ = new_n14906_ & new_n14697_;
  assign new_n14815_ = new_n14951_ & new_n14869_;
  assign new_n14816_ = new_n14977_ & new_n14870_;
  assign new_n14817_ = new_n14993_ & new_n14994_;
  assign new_n14818_ = new_n14996_ & new_n15075_;
  assign new_n14819_ = new_n14997_ & new_n14994_ & new_n14993_;
  assign new_n14820_ = ~new_n15079_ | ~new_n15078_;
  assign new_n14821_ = new_n14774_ & new_n15084_ & new_n15083_;
  assign new_n14822_ = new_n15087_ & new_n14871_;
  assign new_n14823_ = ~new_n15093_ | ~new_n15092_;
  assign new_n14824_ = ~new_n15098_ | ~new_n15097_;
  assign new_n14825_ = new_n15104_ & new_n14870_;
  assign new_n14826_ = ~new_n15114_ | ~new_n15113_;
  assign new_n14827_ = ~new_n15119_ | ~new_n15118_;
  assign new_n14828_ = ~new_n15124_ | ~new_n15123_;
  assign new_n14829_ = ~new_n15129_ | ~new_n15128_;
  assign new_n14830_ = ~new_n15134_ | ~new_n15133_;
  assign new_n14831_ = new_n15140_ & new_n14869_;
  assign new_n14832_ = ~new_n15150_ | ~new_n15149_;
  assign new_n14833_ = ~new_n15155_ | ~new_n15154_;
  assign new_n14834_ = new_n15031_ & new_n14698_;
  assign new_n14835_ = new_n15161_ & new_n14868_;
  assign new_n14836_ = new_n15039_ & new_n15038_;
  assign new_n14837_ = ~new_n14807_ | ~new_n14901_;
  assign new_n14838_ = new_n15048_ & new_n15047_;
  assign new_n14839_ = new_n15055_ & new_n15054_;
  assign new_n14840_ = new_n15059_ & new_n15058_;
  assign new_n14841_ = ~new_n14805_ | ~new_n14885_;
  assign new_n14842_ = new_n15068_ & new_n15067_;
  assign new_n14843_ = ~new_n2955_;
  assign new_n14844_ = ~new_n1982_;
  assign new_n14845_ = new_n15077_ & new_n15076_;
  assign new_n14846_ = ~new_n14817_ | ~new_n14991_;
  assign new_n14847_ = new_n15089_ & new_n15088_;
  assign new_n14848_ = ~new_n14984_ | ~new_n14983_;
  assign new_n14849_ = ~new_n14980_ | ~new_n14979_;
  assign new_n14850_ = new_n15106_ & new_n15105_;
  assign new_n14851_ = new_n15110_ & new_n15109_;
  assign new_n14852_ = ~new_n14970_ | ~new_n14969_;
  assign new_n14853_ = ~new_n14966_ | ~new_n14965_;
  assign new_n14854_ = ~new_n2388_;
  assign new_n14855_ = ~new_n14962_ | ~new_n14961_;
  assign new_n14856_ = ~new_n2439_;
  assign new_n14857_ = ~new_n14954_ | ~new_n14953_;
  assign new_n14858_ = new_n15142_ & new_n15141_;
  assign new_n14859_ = new_n15146_ & new_n15145_;
  assign new_n14860_ = ~new_n14944_ | ~new_n14943_;
  assign new_n14861_ = ~new_n14940_ | ~new_n14939_;
  assign new_n14862_ = ~new_n14936_ | ~new_n14935_;
  assign new_n14863_ = new_n15163_ & new_n15162_;
  assign new_n14864_ = ~new_n14818_ | ~new_n14846_;
  assign new_n14865_ = ~new_n14774_;
  assign new_n14866_ = ~new_n14718_;
  assign new_n14867_ = ~new_n14729_;
  assign new_n14868_ = ~new_n2415_ | ~new_n14742_;
  assign new_n14869_ = ~new_n2430_ | ~new_n14751_;
  assign new_n14870_ = ~new_n2950_ | ~new_n14765_;
  assign new_n14871_ = ~new_n2946_ | ~new_n14773_;
  assign new_n14872_ = ~new_n2391_ | ~new_n14717_;
  assign new_n14873_ = ~new_n2400_ | ~new_n14724_;
  assign new_n14874_ = ~new_n2406_ | ~new_n14728_;
  assign new_n14875_ = ~new_n14753_;
  assign new_n14876_ = ~new_n14767_;
  assign new_n14877_ = ~new_n14726_;
  assign new_n14878_ = ~new_n14743_;
  assign new_n14879_ = ~new_n14714_;
  assign new_n14880_ = ~new_n14879_ | ~new_n14715_;
  assign new_n14881_ = ~new_n14880_ | ~new_n14854_;
  assign new_n14882_ = ~new_n2005_ | ~new_n14714_;
  assign new_n14883_ = ~new_n14735_;
  assign new_n14884_ = ~new_n2394_ | ~new_n14719_;
  assign new_n14885_ = ~new_n14804_ | ~new_n14735_;
  assign new_n14886_ = ~new_n14719_ | ~new_n14718_;
  assign new_n14887_ = ~new_n14886_ | ~new_n14716_;
  assign new_n14888_ = ~new_n1991_ | ~new_n14866_;
  assign new_n14889_ = ~new_n14841_;
  assign new_n14890_ = ~new_n2403_ | ~new_n14723_;
  assign new_n14891_ = ~new_n1998_ | ~new_n14720_;
  assign new_n14892_ = ~new_n1994_ | ~new_n14721_;
  assign new_n14893_ = ~new_n14877_ | ~new_n14695_;
  assign new_n14894_ = ~new_n14696_ | ~new_n14893_;
  assign new_n14895_ = ~new_n2397_ | ~new_n14725_;
  assign new_n14896_ = ~new_n2403_ | ~new_n14723_;
  assign new_n14897_ = ~new_n14695_ | ~new_n14895_ | ~new_n14841_;
  assign new_n14898_ = ~new_n14896_ | ~new_n14894_;
  assign new_n14899_ = ~new_n14733_;
  assign new_n14900_ = ~new_n2409_ | ~new_n14730_;
  assign new_n14901_ = ~new_n14806_ | ~new_n14733_;
  assign new_n14902_ = ~new_n14730_ | ~new_n14729_;
  assign new_n14903_ = ~new_n14902_ | ~new_n14727_;
  assign new_n14904_ = ~new_n2011_ | ~new_n14867_;
  assign new_n14905_ = ~new_n14837_;
  assign new_n14906_ = ~new_n2412_ | ~new_n14732_;
  assign new_n14907_ = ~new_n14906_ | ~new_n14743_;
  assign new_n14908_ = ~new_n14899_ | ~new_n14729_;
  assign new_n14909_ = ~new_n14809_ | ~new_n14908_;
  assign new_n14910_ = ~new_n14733_ | ~new_n14874_;
  assign new_n14911_ = ~new_n14808_ | ~new_n14910_;
  assign new_n14912_ = ~new_n14729_ | ~new_n14874_;
  assign new_n14913_ = ~new_n14895_ | ~new_n14841_;
  assign new_n14914_ = ~new_n14734_;
  assign new_n14915_ = ~new_n1994_ | ~new_n14721_;
  assign new_n14916_ = ~new_n14914_ | ~new_n14915_;
  assign new_n14917_ = ~new_n14811_ | ~new_n14916_;
  assign new_n14918_ = ~new_n14734_ | ~new_n14873_;
  assign new_n14919_ = ~new_n2403_ | ~new_n14723_;
  assign new_n14920_ = ~new_n14810_ | ~new_n14918_;
  assign new_n14921_ = ~new_n1994_ | ~new_n14721_;
  assign new_n14922_ = ~new_n14873_ | ~new_n14921_;
  assign new_n14923_ = ~new_n14895_ | ~new_n14726_;
  assign new_n14924_ = ~new_n14883_ | ~new_n14718_;
  assign new_n14925_ = ~new_n14813_ | ~new_n14924_;
  assign new_n14926_ = ~new_n14735_ | ~new_n14872_;
  assign new_n14927_ = ~new_n14812_ | ~new_n14926_;
  assign new_n14928_ = ~new_n14718_ | ~new_n14872_;
  assign new_n14929_ = ~new_n2418_ | ~new_n14741_;
  assign new_n14930_ = ~new_n1990_ | ~new_n14739_;
  assign new_n14931_ = ~new_n1989_ | ~new_n14740_;
  assign new_n14932_ = ~new_n14878_ | ~new_n14697_;
  assign new_n14933_ = ~new_n14698_ | ~new_n14932_;
  assign new_n14934_ = ~new_n2418_ | ~new_n14741_;
  assign new_n14935_ = ~new_n14814_ | ~new_n14837_;
  assign new_n14936_ = ~new_n14934_ | ~new_n14933_;
  assign new_n14937_ = ~new_n14862_;
  assign new_n14938_ = ~new_n2421_ | ~new_n14745_;
  assign new_n14939_ = ~new_n14938_ | ~new_n14862_;
  assign new_n14940_ = ~new_n1999_ | ~new_n14744_;
  assign new_n14941_ = ~new_n14861_;
  assign new_n14942_ = ~new_n2424_ | ~new_n14747_;
  assign new_n14943_ = ~new_n14942_ | ~new_n14861_;
  assign new_n14944_ = ~new_n2007_ | ~new_n14746_;
  assign new_n14945_ = ~new_n14860_;
  assign new_n14946_ = ~new_n2433_ | ~new_n14750_;
  assign new_n14947_ = ~new_n2000_ | ~new_n14748_;
  assign new_n14948_ = ~new_n2001_ | ~new_n14738_;
  assign new_n14949_ = ~new_n14875_ | ~new_n14869_;
  assign new_n14950_ = ~new_n14699_ | ~new_n14949_;
  assign new_n14951_ = ~new_n2427_ | ~new_n14752_;
  assign new_n14952_ = ~new_n2433_ | ~new_n14750_;
  assign new_n14953_ = ~new_n14946_ | ~new_n14860_ | ~new_n14815_;
  assign new_n14954_ = ~new_n14952_ | ~new_n14950_;
  assign new_n14955_ = ~new_n14857_;
  assign new_n14956_ = ~new_n2436_ | ~new_n14755_;
  assign new_n14957_ = ~new_n14956_ | ~new_n14857_;
  assign new_n14958_ = ~new_n1996_ | ~new_n14754_;
  assign new_n14959_ = ~new_n14756_;
  assign new_n14960_ = ~new_n14959_ | ~new_n14757_;
  assign new_n14961_ = ~new_n14960_ | ~new_n14856_;
  assign new_n14962_ = ~new_n2009_ | ~new_n14756_;
  assign new_n14963_ = ~new_n14855_;
  assign new_n14964_ = ~new_n2441_ | ~new_n14759_;
  assign new_n14965_ = ~new_n14964_ | ~new_n14855_;
  assign new_n14966_ = ~new_n2008_ | ~new_n14758_;
  assign new_n14967_ = ~new_n14853_;
  assign new_n14968_ = ~new_n2952_ | ~new_n14761_;
  assign new_n14969_ = ~new_n14968_ | ~new_n14853_;
  assign new_n14970_ = ~new_n2003_ | ~new_n14760_;
  assign new_n14971_ = ~new_n14852_;
  assign new_n14972_ = ~new_n2949_ | ~new_n14764_;
  assign new_n14973_ = ~new_n1993_ | ~new_n14762_;
  assign new_n14974_ = ~new_n1988_ | ~new_n14737_;
  assign new_n14975_ = ~new_n14876_ | ~new_n14870_;
  assign new_n14976_ = ~new_n14700_ | ~new_n14975_;
  assign new_n14977_ = ~new_n2951_ | ~new_n14766_;
  assign new_n14978_ = ~new_n2949_ | ~new_n14764_;
  assign new_n14979_ = ~new_n14972_ | ~new_n14852_ | ~new_n14816_;
  assign new_n14980_ = ~new_n14978_ | ~new_n14976_;
  assign new_n14981_ = ~new_n14849_;
  assign new_n14982_ = ~new_n2948_ | ~new_n14769_;
  assign new_n14983_ = ~new_n14982_ | ~new_n14849_;
  assign new_n14984_ = ~new_n1992_ | ~new_n14768_;
  assign new_n14985_ = ~new_n14848_;
  assign new_n14986_ = ~new_n2947_ | ~new_n14771_;
  assign new_n14987_ = ~new_n14986_ | ~new_n14848_;
  assign new_n14988_ = ~new_n1985_ | ~new_n14770_;
  assign new_n14989_ = ~new_n14778_;
  assign new_n14990_ = ~new_n2945_ | ~new_n14775_;
  assign new_n14991_ = ~new_n14990_ | ~new_n14778_ | ~new_n14871_;
  assign new_n14992_ = ~new_n14775_ | ~new_n14774_;
  assign new_n14993_ = ~new_n14992_ | ~new_n14772_;
  assign new_n14994_ = ~new_n1980_ | ~new_n14865_;
  assign new_n14995_ = ~new_n14846_;
  assign new_n14996_ = ~new_n2944_ | ~new_n14777_;
  assign new_n14997_ = ~new_n1981_ | ~new_n14776_;
  assign new_n14998_ = ~new_n14989_ | ~new_n14774_;
  assign new_n14999_ = ~new_n14822_ | ~new_n14998_;
  assign new_n15000_ = ~new_n14778_ | ~new_n14871_;
  assign new_n15001_ = ~new_n14821_ | ~new_n15000_;
  assign new_n15002_ = ~new_n14774_ | ~new_n14871_;
  assign new_n15003_ = ~new_n14977_ | ~new_n14852_;
  assign new_n15004_ = ~new_n14779_;
  assign new_n15005_ = ~new_n1988_ | ~new_n14737_;
  assign new_n15006_ = ~new_n15004_ | ~new_n15005_;
  assign new_n15007_ = ~new_n14825_ | ~new_n15006_;
  assign new_n15008_ = ~new_n14779_ | ~new_n14870_;
  assign new_n15009_ = ~new_n2949_ | ~new_n14764_;
  assign new_n15010_ = ~new_n14700_ | ~new_n15009_ | ~new_n15008_;
  assign new_n15011_ = ~new_n1988_ | ~new_n14737_;
  assign new_n15012_ = ~new_n14870_ | ~new_n15011_;
  assign new_n15013_ = ~new_n14977_ | ~new_n14767_;
  assign new_n15014_ = ~new_n14951_ | ~new_n14860_;
  assign new_n15015_ = ~new_n14780_;
  assign new_n15016_ = ~new_n2001_ | ~new_n14738_;
  assign new_n15017_ = ~new_n15015_ | ~new_n15016_;
  assign new_n15018_ = ~new_n14831_ | ~new_n15017_;
  assign new_n15019_ = ~new_n14780_ | ~new_n14869_;
  assign new_n15020_ = ~new_n2433_ | ~new_n14750_;
  assign new_n15021_ = ~new_n14699_ | ~new_n15020_ | ~new_n15019_;
  assign new_n15022_ = ~new_n2001_ | ~new_n14738_;
  assign new_n15023_ = ~new_n14869_ | ~new_n15022_;
  assign new_n15024_ = ~new_n14951_ | ~new_n14753_;
  assign new_n15025_ = ~new_n14906_ | ~new_n14837_;
  assign new_n15026_ = ~new_n14781_;
  assign new_n15027_ = ~new_n1989_ | ~new_n14740_;
  assign new_n15028_ = ~new_n15026_ | ~new_n15027_;
  assign new_n15029_ = ~new_n14835_ | ~new_n15028_;
  assign new_n15030_ = ~new_n14781_ | ~new_n14868_;
  assign new_n15031_ = ~new_n2418_ | ~new_n14741_;
  assign new_n15032_ = ~new_n14834_ | ~new_n15030_;
  assign new_n15033_ = ~new_n1989_ | ~new_n14740_;
  assign new_n15034_ = ~new_n14868_ | ~new_n15033_;
  assign new_n15035_ = ~new_n2004_ | ~new_n14713_;
  assign new_n15036_ = ~new_n14990_ | ~new_n14778_ | ~new_n14871_;
  assign new_n15037_ = ~new_n14819_ | ~new_n14701_ | ~new_n15036_;
  assign new_n15038_ = ~new_n2412_ | ~new_n14732_;
  assign new_n15039_ = ~new_n2010_ | ~new_n14731_;
  assign new_n15040_ = ~new_n14907_ | ~new_n14837_;
  assign new_n15041_ = ~new_n14905_ | ~new_n14836_;
  assign new_n15042_ = ~new_n2409_ | ~new_n14730_;
  assign new_n15043_ = ~new_n2011_ | ~new_n14727_;
  assign new_n15044_ = ~new_n2409_ | ~new_n14730_;
  assign new_n15045_ = ~new_n2011_ | ~new_n14727_;
  assign new_n15046_ = ~new_n15045_ | ~new_n15044_;
  assign new_n15047_ = ~new_n2406_ | ~new_n14728_;
  assign new_n15048_ = ~new_n1997_ | ~new_n14711_;
  assign new_n15049_ = ~new_n14912_ | ~new_n14733_;
  assign new_n15050_ = ~new_n14838_ | ~new_n14899_;
  assign new_n15051_ = ~new_n2403_ | ~new_n14723_;
  assign new_n15052_ = ~new_n1998_ | ~new_n14720_;
  assign new_n15053_ = ~new_n15052_ | ~new_n15051_;
  assign new_n15054_ = ~new_n2400_ | ~new_n14724_;
  assign new_n15055_ = ~new_n1994_ | ~new_n14721_;
  assign new_n15056_ = ~new_n14922_ | ~new_n14734_;
  assign new_n15057_ = ~new_n14839_ | ~new_n14914_;
  assign new_n15058_ = ~new_n2397_ | ~new_n14725_;
  assign new_n15059_ = ~new_n1987_ | ~new_n14722_;
  assign new_n15060_ = ~new_n14923_ | ~new_n14841_;
  assign new_n15061_ = ~new_n14889_ | ~new_n14840_;
  assign new_n15062_ = ~new_n2394_ | ~new_n14719_;
  assign new_n15063_ = ~new_n1991_ | ~new_n14716_;
  assign new_n15064_ = ~new_n2394_ | ~new_n14719_;
  assign new_n15065_ = ~new_n1991_ | ~new_n14716_;
  assign new_n15066_ = ~new_n15065_ | ~new_n15064_;
  assign new_n15067_ = ~new_n2391_ | ~new_n14717_;
  assign new_n15068_ = ~new_n1995_ | ~new_n14712_;
  assign new_n15069_ = ~new_n14928_ | ~new_n14735_;
  assign new_n15070_ = ~new_n14842_ | ~new_n14883_;
  assign new_n15071_ = ~new_n2955_ | ~new_n14844_;
  assign new_n15072_ = ~new_n1982_ | ~new_n14843_;
  assign new_n15073_ = ~new_n2955_ | ~new_n14844_;
  assign new_n15074_ = ~new_n1982_ | ~new_n14843_;
  assign new_n15075_ = ~new_n15074_ | ~new_n15073_;
  assign new_n15076_ = ~new_n14776_ | ~new_n1981_ | ~new_n15075_;
  assign new_n15077_ = ~new_n2944_ | ~new_n14701_ | ~new_n14777_;
  assign new_n15078_ = ~new_n2944_ | ~new_n14777_;
  assign new_n15079_ = ~new_n1981_ | ~new_n14776_;
  assign new_n15080_ = ~new_n14820_;
  assign new_n15081_ = ~new_n14995_ | ~new_n15080_;
  assign new_n15082_ = ~new_n14820_ | ~new_n14846_;
  assign new_n15083_ = ~new_n2945_ | ~new_n14775_;
  assign new_n15084_ = ~new_n1980_ | ~new_n14772_;
  assign new_n15085_ = ~new_n2945_ | ~new_n14775_;
  assign new_n15086_ = ~new_n1980_ | ~new_n14772_;
  assign new_n15087_ = ~new_n15086_ | ~new_n15085_;
  assign new_n15088_ = ~new_n2946_ | ~new_n14773_;
  assign new_n15089_ = ~new_n1984_ | ~new_n14736_;
  assign new_n15090_ = ~new_n15002_ | ~new_n14778_;
  assign new_n15091_ = ~new_n14847_ | ~new_n14989_;
  assign new_n15092_ = ~new_n2947_ | ~new_n14771_;
  assign new_n15093_ = ~new_n1985_ | ~new_n14770_;
  assign new_n15094_ = ~new_n14823_;
  assign new_n15095_ = ~new_n14985_ | ~new_n15094_;
  assign new_n15096_ = ~new_n14823_ | ~new_n14848_;
  assign new_n15097_ = ~new_n2948_ | ~new_n14769_;
  assign new_n15098_ = ~new_n1992_ | ~new_n14768_;
  assign new_n15099_ = ~new_n14824_;
  assign new_n15100_ = ~new_n14981_ | ~new_n15099_;
  assign new_n15101_ = ~new_n14824_ | ~new_n14849_;
  assign new_n15102_ = ~new_n2949_ | ~new_n14764_;
  assign new_n15103_ = ~new_n1993_ | ~new_n14762_;
  assign new_n15104_ = ~new_n15103_ | ~new_n15102_;
  assign new_n15105_ = ~new_n2950_ | ~new_n14765_;
  assign new_n15106_ = ~new_n1988_ | ~new_n14737_;
  assign new_n15107_ = ~new_n15012_ | ~new_n14779_;
  assign new_n15108_ = ~new_n14850_ | ~new_n15004_;
  assign new_n15109_ = ~new_n2951_ | ~new_n14766_;
  assign new_n15110_ = ~new_n2002_ | ~new_n14763_;
  assign new_n15111_ = ~new_n15013_ | ~new_n14852_;
  assign new_n15112_ = ~new_n14971_ | ~new_n14851_;
  assign new_n15113_ = ~new_n2952_ | ~new_n14761_;
  assign new_n15114_ = ~new_n2003_ | ~new_n14760_;
  assign new_n15115_ = ~new_n14826_;
  assign new_n15116_ = ~new_n14967_ | ~new_n15115_;
  assign new_n15117_ = ~new_n14826_ | ~new_n14853_;
  assign new_n15118_ = ~new_n2388_ | ~new_n14715_;
  assign new_n15119_ = ~new_n2005_ | ~new_n14854_;
  assign new_n15120_ = ~new_n14827_;
  assign new_n15121_ = ~new_n15120_ | ~new_n14879_;
  assign new_n15122_ = ~new_n14827_ | ~new_n14714_;
  assign new_n15123_ = ~new_n2441_ | ~new_n14759_;
  assign new_n15124_ = ~new_n2008_ | ~new_n14758_;
  assign new_n15125_ = ~new_n14828_;
  assign new_n15126_ = ~new_n14963_ | ~new_n15125_;
  assign new_n15127_ = ~new_n14828_ | ~new_n14855_;
  assign new_n15128_ = ~new_n2439_ | ~new_n14757_;
  assign new_n15129_ = ~new_n2009_ | ~new_n14856_;
  assign new_n15130_ = ~new_n14829_;
  assign new_n15131_ = ~new_n15130_ | ~new_n14959_;
  assign new_n15132_ = ~new_n14829_ | ~new_n14756_;
  assign new_n15133_ = ~new_n2436_ | ~new_n14755_;
  assign new_n15134_ = ~new_n1996_ | ~new_n14754_;
  assign new_n15135_ = ~new_n14830_;
  assign new_n15136_ = ~new_n14955_ | ~new_n15135_;
  assign new_n15137_ = ~new_n14830_ | ~new_n14857_;
  assign new_n15138_ = ~new_n2433_ | ~new_n14750_;
  assign new_n15139_ = ~new_n2000_ | ~new_n14748_;
  assign new_n15140_ = ~new_n15139_ | ~new_n15138_;
  assign new_n15141_ = ~new_n2430_ | ~new_n14751_;
  assign new_n15142_ = ~new_n2001_ | ~new_n14738_;
  assign new_n15143_ = ~new_n15023_ | ~new_n14780_;
  assign new_n15144_ = ~new_n14858_ | ~new_n15015_;
  assign new_n15145_ = ~new_n2427_ | ~new_n14752_;
  assign new_n15146_ = ~new_n2006_ | ~new_n14749_;
  assign new_n15147_ = ~new_n15024_ | ~new_n14860_;
  assign new_n15148_ = ~new_n14945_ | ~new_n14859_;
  assign new_n15149_ = ~new_n2424_ | ~new_n14747_;
  assign new_n15150_ = ~new_n2007_ | ~new_n14746_;
  assign new_n15151_ = ~new_n14832_;
  assign new_n15152_ = ~new_n14941_ | ~new_n15151_;
  assign new_n15153_ = ~new_n14832_ | ~new_n14861_;
  assign new_n15154_ = ~new_n2421_ | ~new_n14745_;
  assign new_n15155_ = ~new_n1999_ | ~new_n14744_;
  assign new_n15156_ = ~new_n14833_;
  assign new_n15157_ = ~new_n14937_ | ~new_n15156_;
  assign new_n15158_ = ~new_n14833_ | ~new_n14862_;
  assign new_n15159_ = ~new_n2418_ | ~new_n14741_;
  assign new_n15160_ = ~new_n1990_ | ~new_n14739_;
  assign new_n15161_ = ~new_n15160_ | ~new_n15159_;
  assign new_n15162_ = ~new_n2415_ | ~new_n14742_;
  assign new_n15163_ = ~new_n1989_ | ~new_n14740_;
  assign new_n15164_ = ~new_n15034_ | ~new_n14781_;
  assign new_n15165_ = ~new_n14863_ | ~new_n15026_;
  assign new_n15166_ = new_n15168_ & new_n15351_;
  assign new_n15167_ = new_n15349_ & new_n15350_ & new_n15260_;
  assign new_n15168_ = new_n15355_ & new_n15354_;
  assign new_n15169_ = ~new_n15167_ | ~new_n15352_;
  assign new_n15170_ = ~new_n2015_;
  assign new_n15171_ = ~new_n2014_;
  assign new_n15172_ = ~new_n2048_;
  assign new_n15173_ = ~new_n2047_;
  assign new_n15174_ = ~new_n2079_;
  assign new_n15175_ = ~new_n2044_;
  assign new_n15176_ = ~new_n2076_;
  assign new_n15177_ = ~new_n2075_;
  assign new_n15178_ = ~new_n2043_;
  assign new_n15179_ = ~new_n2042_;
  assign new_n15180_ = ~new_n2074_;
  assign new_n15181_ = ~new_n2073_;
  assign new_n15182_ = ~new_n2041_;
  assign new_n15183_ = ~new_n2040_;
  assign new_n15184_ = ~new_n2072_;
  assign new_n15185_ = ~new_n2071_;
  assign new_n15186_ = ~new_n2039_;
  assign new_n15187_ = ~new_n2038_;
  assign new_n15188_ = ~new_n2070_;
  assign new_n15189_ = ~new_n2069_;
  assign new_n15190_ = ~new_n2037_;
  assign new_n15191_ = ~new_n2036_;
  assign new_n15192_ = ~new_n2068_;
  assign new_n15193_ = ~new_n2067_;
  assign new_n15194_ = ~new_n2035_;
  assign new_n15195_ = ~new_n2034_;
  assign new_n15196_ = ~new_n2066_;
  assign new_n15197_ = ~new_n2065_;
  assign new_n15198_ = ~new_n2033_;
  assign new_n15199_ = ~new_n2032_;
  assign new_n15200_ = ~new_n2064_;
  assign new_n15201_ = ~new_n2063_;
  assign new_n15202_ = ~new_n2031_;
  assign new_n15203_ = ~new_n2030_;
  assign new_n15204_ = ~new_n2062_;
  assign new_n15205_ = ~new_n2061_;
  assign new_n15206_ = ~new_n2029_;
  assign new_n15207_ = ~new_n2028_;
  assign new_n15208_ = ~new_n2060_;
  assign new_n15209_ = ~new_n2059_;
  assign new_n15210_ = ~new_n2027_;
  assign new_n15211_ = ~new_n2026_;
  assign new_n15212_ = ~new_n2058_;
  assign new_n15213_ = ~new_n2057_;
  assign new_n15214_ = ~new_n2025_;
  assign new_n15215_ = ~new_n2024_;
  assign new_n15216_ = ~new_n2056_;
  assign new_n15217_ = ~new_n2055_;
  assign new_n15218_ = ~new_n2023_;
  assign new_n15219_ = ~new_n2022_;
  assign new_n15220_ = ~new_n2054_;
  assign new_n15221_ = ~new_n2053_;
  assign new_n15222_ = ~new_n2021_;
  assign new_n15223_ = ~new_n2020_;
  assign new_n15224_ = ~new_n2052_;
  assign new_n15225_ = ~new_n2051_;
  assign new_n15226_ = ~new_n2019_;
  assign new_n15227_ = ~new_n2018_;
  assign new_n15228_ = ~new_n2050_;
  assign new_n15229_ = ~new_n2016_;
  assign new_n15230_ = new_n15267_ & new_n15268_;
  assign new_n15231_ = new_n15270_ & new_n15271_;
  assign new_n15232_ = new_n15273_ & new_n15274_;
  assign new_n15233_ = new_n15276_ & new_n15277_;
  assign new_n15234_ = new_n15279_ & new_n15280_;
  assign new_n15235_ = new_n15282_ & new_n15283_;
  assign new_n15236_ = new_n15285_ & new_n15286_;
  assign new_n15237_ = new_n15288_ & new_n15289_;
  assign new_n15238_ = new_n15291_ & new_n15292_;
  assign new_n15239_ = new_n15294_ & new_n15295_;
  assign new_n15240_ = new_n15297_ & new_n15298_;
  assign new_n15241_ = new_n15300_ & new_n15301_;
  assign new_n15242_ = new_n15303_ & new_n15304_;
  assign new_n15243_ = new_n15306_ & new_n15307_;
  assign new_n15244_ = new_n15309_ & new_n15310_;
  assign new_n15245_ = new_n15312_ & new_n15313_;
  assign new_n15246_ = new_n15315_ & new_n15316_;
  assign new_n15247_ = new_n15318_ & new_n15319_;
  assign new_n15248_ = new_n15321_ & new_n15322_;
  assign new_n15249_ = new_n15324_ & new_n15325_;
  assign new_n15250_ = new_n15327_ & new_n15328_;
  assign new_n15251_ = new_n15330_ & new_n15331_;
  assign new_n15252_ = new_n15333_ & new_n15334_;
  assign new_n15253_ = new_n15336_ & new_n15337_;
  assign new_n15254_ = new_n15339_ & new_n15340_;
  assign new_n15255_ = new_n15342_ & new_n15343_;
  assign new_n15256_ = new_n15346_ & new_n15261_;
  assign new_n15257_ = new_n15346_ & new_n2017_;
  assign new_n15258_ = new_n15347_ & new_n15348_;
  assign new_n15259_ = ~new_n2046_;
  assign new_n15260_ = new_n15357_ & new_n15356_;
  assign new_n15261_ = ~new_n2049_;
  assign new_n15262_ = ~new_n2077_ | ~new_n2078_;
  assign new_n15263_ = ~new_n2045_ | ~new_n15262_;
  assign new_n15264_ = new_n2077_ | new_n2078_;
  assign new_n15265_ = ~new_n2044_ | ~new_n15176_;
  assign new_n15266_ = ~new_n15263_ | ~new_n15264_ | ~new_n15265_;
  assign new_n15267_ = ~new_n2076_ | ~new_n15175_;
  assign new_n15268_ = ~new_n2075_ | ~new_n15178_;
  assign new_n15269_ = ~new_n15230_ | ~new_n15266_;
  assign new_n15270_ = ~new_n2043_ | ~new_n15177_;
  assign new_n15271_ = ~new_n2042_ | ~new_n15180_;
  assign new_n15272_ = ~new_n15231_ | ~new_n15269_;
  assign new_n15273_ = ~new_n2074_ | ~new_n15179_;
  assign new_n15274_ = ~new_n2073_ | ~new_n15182_;
  assign new_n15275_ = ~new_n15232_ | ~new_n15272_;
  assign new_n15276_ = ~new_n2041_ | ~new_n15181_;
  assign new_n15277_ = ~new_n2040_ | ~new_n15184_;
  assign new_n15278_ = ~new_n15233_ | ~new_n15275_;
  assign new_n15279_ = ~new_n2072_ | ~new_n15183_;
  assign new_n15280_ = ~new_n2071_ | ~new_n15186_;
  assign new_n15281_ = ~new_n15234_ | ~new_n15278_;
  assign new_n15282_ = ~new_n2039_ | ~new_n15185_;
  assign new_n15283_ = ~new_n2038_ | ~new_n15188_;
  assign new_n15284_ = ~new_n15235_ | ~new_n15281_;
  assign new_n15285_ = ~new_n2070_ | ~new_n15187_;
  assign new_n15286_ = ~new_n2069_ | ~new_n15190_;
  assign new_n15287_ = ~new_n15236_ | ~new_n15284_;
  assign new_n15288_ = ~new_n2037_ | ~new_n15189_;
  assign new_n15289_ = ~new_n2036_ | ~new_n15192_;
  assign new_n15290_ = ~new_n15237_ | ~new_n15287_;
  assign new_n15291_ = ~new_n2068_ | ~new_n15191_;
  assign new_n15292_ = ~new_n2067_ | ~new_n15194_;
  assign new_n15293_ = ~new_n15238_ | ~new_n15290_;
  assign new_n15294_ = ~new_n2035_ | ~new_n15193_;
  assign new_n15295_ = ~new_n2034_ | ~new_n15196_;
  assign new_n15296_ = ~new_n15239_ | ~new_n15293_;
  assign new_n15297_ = ~new_n2066_ | ~new_n15195_;
  assign new_n15298_ = ~new_n2065_ | ~new_n15198_;
  assign new_n15299_ = ~new_n15240_ | ~new_n15296_;
  assign new_n15300_ = ~new_n2033_ | ~new_n15197_;
  assign new_n15301_ = ~new_n2032_ | ~new_n15200_;
  assign new_n15302_ = ~new_n15241_ | ~new_n15299_;
  assign new_n15303_ = ~new_n2064_ | ~new_n15199_;
  assign new_n15304_ = ~new_n2063_ | ~new_n15202_;
  assign new_n15305_ = ~new_n15242_ | ~new_n15302_;
  assign new_n15306_ = ~new_n2031_ | ~new_n15201_;
  assign new_n15307_ = ~new_n2030_ | ~new_n15204_;
  assign new_n15308_ = ~new_n15243_ | ~new_n15305_;
  assign new_n15309_ = ~new_n2062_ | ~new_n15203_;
  assign new_n15310_ = ~new_n2061_ | ~new_n15206_;
  assign new_n15311_ = ~new_n15244_ | ~new_n15308_;
  assign new_n15312_ = ~new_n2029_ | ~new_n15205_;
  assign new_n15313_ = ~new_n2028_ | ~new_n15208_;
  assign new_n15314_ = ~new_n15245_ | ~new_n15311_;
  assign new_n15315_ = ~new_n2060_ | ~new_n15207_;
  assign new_n15316_ = ~new_n2059_ | ~new_n15210_;
  assign new_n15317_ = ~new_n15246_ | ~new_n15314_;
  assign new_n15318_ = ~new_n2027_ | ~new_n15209_;
  assign new_n15319_ = ~new_n2026_ | ~new_n15212_;
  assign new_n15320_ = ~new_n15247_ | ~new_n15317_;
  assign new_n15321_ = ~new_n2058_ | ~new_n15211_;
  assign new_n15322_ = ~new_n2057_ | ~new_n15214_;
  assign new_n15323_ = ~new_n15248_ | ~new_n15320_;
  assign new_n15324_ = ~new_n2025_ | ~new_n15213_;
  assign new_n15325_ = ~new_n2024_ | ~new_n15216_;
  assign new_n15326_ = ~new_n15249_ | ~new_n15323_;
  assign new_n15327_ = ~new_n2056_ | ~new_n15215_;
  assign new_n15328_ = ~new_n2055_ | ~new_n15218_;
  assign new_n15329_ = ~new_n15250_ | ~new_n15326_;
  assign new_n15330_ = ~new_n2023_ | ~new_n15217_;
  assign new_n15331_ = ~new_n2022_ | ~new_n15220_;
  assign new_n15332_ = ~new_n15251_ | ~new_n15329_;
  assign new_n15333_ = ~new_n2054_ | ~new_n15219_;
  assign new_n15334_ = ~new_n2053_ | ~new_n15222_;
  assign new_n15335_ = ~new_n15252_ | ~new_n15332_;
  assign new_n15336_ = ~new_n2021_ | ~new_n15221_;
  assign new_n15337_ = ~new_n2020_ | ~new_n15224_;
  assign new_n15338_ = ~new_n15253_ | ~new_n15335_;
  assign new_n15339_ = ~new_n2052_ | ~new_n15223_;
  assign new_n15340_ = ~new_n2051_ | ~new_n15226_;
  assign new_n15341_ = ~new_n15254_ | ~new_n15338_;
  assign new_n15342_ = ~new_n2019_ | ~new_n15225_;
  assign new_n15343_ = ~new_n2018_ | ~new_n15228_;
  assign new_n15344_ = ~new_n15255_ | ~new_n15341_;
  assign new_n15345_ = ~new_n15256_ | ~new_n15344_;
  assign new_n15346_ = ~new_n2050_ | ~new_n15227_;
  assign new_n15347_ = ~new_n2017_ | ~new_n15261_;
  assign new_n15348_ = ~new_n2016_ | ~new_n15172_;
  assign new_n15349_ = ~new_n15351_ | ~new_n15229_ | ~new_n2048_ | ~new_n15168_;
  assign new_n15350_ = ~new_n2047_ | ~new_n15168_ | ~new_n15170_;
  assign new_n15351_ = ~new_n2015_ | ~new_n15173_;
  assign new_n15352_ = ~new_n15353_ | ~new_n15345_ | ~new_n15258_ | ~new_n15166_;
  assign new_n15353_ = ~new_n15257_ | ~new_n15344_;
  assign new_n15354_ = ~new_n2014_ | ~new_n15259_;
  assign new_n15355_ = ~new_n2046_ | ~new_n15171_;
  assign new_n15356_ = ~new_n15259_ | ~new_n2079_ | ~new_n2014_;
  assign new_n15357_ = ~new_n2046_ | ~new_n15174_ | ~new_n15171_;
  assign new_n15358_ = new_n1986_ & new_n15359_;
  assign new_n15359_ = ~new_n1983_;
  assign new_n15360_ = new_n15538_ & new_n15555_;
  assign new_n15361_ = new_n15557_ & new_n15556_;
  assign new_n15362_ = new_n15533_ & new_n15594_;
  assign new_n15363_ = new_n15596_ & new_n15595_;
  assign new_n15364_ = new_n15613_ & new_n15612_;
  assign new_n15365_ = new_n15639_ & new_n15638_;
  assign new_n15366_ = new_n15737_ & new_n15736_;
  assign new_n15367_ = ~new_n15694_ | ~new_n15697_;
  assign new_n15368_ = ~new_n15683_ | ~new_n15686_;
  assign new_n15369_ = ~new_n15672_ | ~new_n15675_;
  assign new_n15370_ = ~new_n15664_ | ~new_n15666_;
  assign new_n15371_ = ~new_n15702_ | ~new_n15510_ | ~new_n15529_;
  assign new_n15372_ = ~new_n15590_ | ~new_n15592_;
  assign new_n15373_ = ~new_n15582_ | ~new_n15585_;
  assign new_n15374_ = ~new_n15574_ | ~new_n15576_;
  assign new_n15375_ = ~new_n15379_ | ~new_n15700_;
  assign new_n15376_ = ~new_n2406_;
  assign new_n15377_ = ~new_n2391_;
  assign new_n15378_ = ~new_n2383_;
  assign new_n15379_ = ~new_n2383_ | ~new_n15447_;
  assign new_n15380_ = ~new_n2005_;
  assign new_n15381_ = ~new_n2394_;
  assign new_n15382_ = ~new_n1995_;
  assign new_n15383_ = ~new_n1995_ | ~new_n15377_;
  assign new_n15384_ = ~new_n1991_;
  assign new_n15385_ = ~new_n2403_;
  assign new_n15386_ = ~new_n2400_;
  assign new_n15387_ = ~new_n2397_;
  assign new_n15388_ = ~new_n1998_;
  assign new_n15389_ = ~new_n1994_;
  assign new_n15390_ = ~new_n1987_;
  assign new_n15391_ = ~new_n1987_ | ~new_n15387_;
  assign new_n15392_ = ~new_n2409_;
  assign new_n15393_ = ~new_n1997_;
  assign new_n15394_ = ~new_n1997_ | ~new_n15376_;
  assign new_n15395_ = ~new_n2011_;
  assign new_n15396_ = ~new_n2412_;
  assign new_n15397_ = ~new_n2010_;
  assign new_n15398_ = ~new_n15563_ | ~new_n15562_;
  assign new_n15399_ = ~new_n15391_ | ~new_n15578_;
  assign new_n15400_ = ~new_n15547_ | ~new_n15546_;
  assign new_n15401_ = ~new_n2946_;
  assign new_n15402_ = ~new_n2950_;
  assign new_n15403_ = ~new_n2430_;
  assign new_n15404_ = ~new_n2418_;
  assign new_n15405_ = ~new_n2415_;
  assign new_n15406_ = ~new_n1990_;
  assign new_n15407_ = ~new_n1989_;
  assign new_n15408_ = ~new_n2010_ | ~new_n15396_;
  assign new_n15409_ = ~new_n2421_;
  assign new_n15410_ = ~new_n1999_;
  assign new_n15411_ = ~new_n2424_;
  assign new_n15412_ = ~new_n2007_;
  assign new_n15413_ = ~new_n2433_;
  assign new_n15414_ = ~new_n2427_;
  assign new_n15415_ = ~new_n2000_;
  assign new_n15416_ = ~new_n2001_;
  assign new_n15417_ = ~new_n2006_;
  assign new_n15418_ = ~new_n2006_ | ~new_n15414_;
  assign new_n15419_ = ~new_n2436_;
  assign new_n15420_ = ~new_n1996_;
  assign new_n15421_ = ~new_n15623_ | ~new_n15622_;
  assign new_n15422_ = ~new_n2009_;
  assign new_n15423_ = ~new_n2441_;
  assign new_n15424_ = ~new_n2008_;
  assign new_n15425_ = ~new_n2952_;
  assign new_n15426_ = ~new_n2003_;
  assign new_n15427_ = ~new_n2949_;
  assign new_n15428_ = ~new_n2951_;
  assign new_n15429_ = ~new_n1993_;
  assign new_n15430_ = ~new_n1988_;
  assign new_n15431_ = ~new_n2002_;
  assign new_n15432_ = ~new_n2002_ | ~new_n15428_;
  assign new_n15433_ = ~new_n2948_;
  assign new_n15434_ = ~new_n1992_;
  assign new_n15435_ = ~new_n2947_;
  assign new_n15436_ = ~new_n1985_;
  assign new_n15437_ = ~new_n2945_;
  assign new_n15438_ = ~new_n1984_;
  assign new_n15439_ = ~new_n1984_ | ~new_n15401_;
  assign new_n15440_ = ~new_n1980_;
  assign new_n15441_ = ~new_n2944_;
  assign new_n15442_ = ~new_n1981_;
  assign new_n15443_ = ~new_n15653_ | ~new_n15652_;
  assign new_n15444_ = ~new_n15432_ | ~new_n15668_;
  assign new_n15445_ = ~new_n15418_ | ~new_n15679_;
  assign new_n15446_ = ~new_n15408_ | ~new_n15690_;
  assign new_n15447_ = ~new_n2004_;
  assign new_n15448_ = ~new_n15747_ | ~new_n15746_;
  assign new_n15449_ = ~new_n15761_ | ~new_n15760_;
  assign new_n15450_ = ~new_n15766_ | ~new_n15765_;
  assign new_n15451_ = ~new_n15782_ | ~new_n15781_;
  assign new_n15452_ = ~new_n15787_ | ~new_n15786_;
  assign new_n15453_ = ~new_n15792_ | ~new_n15791_;
  assign new_n15454_ = ~new_n15797_ | ~new_n15796_;
  assign new_n15455_ = ~new_n15802_ | ~new_n15801_;
  assign new_n15456_ = ~new_n15818_ | ~new_n15817_;
  assign new_n15457_ = ~new_n15823_ | ~new_n15822_;
  assign new_n15458_ = ~new_n15706_ | ~new_n15705_;
  assign new_n15459_ = ~new_n15715_ | ~new_n15714_;
  assign new_n15460_ = ~new_n15722_ | ~new_n15721_;
  assign new_n15461_ = ~new_n15726_ | ~new_n15725_;
  assign new_n15462_ = ~new_n15735_ | ~new_n15734_;
  assign new_n15463_ = ~new_n15756_ | ~new_n15755_;
  assign new_n15464_ = ~new_n15773_ | ~new_n15772_;
  assign new_n15465_ = ~new_n15777_ | ~new_n15776_;
  assign new_n15466_ = ~new_n15809_ | ~new_n15808_;
  assign new_n15467_ = ~new_n15813_ | ~new_n15812_;
  assign new_n15468_ = ~new_n15830_ | ~new_n15829_;
  assign new_n15469_ = new_n15549_ & new_n15537_;
  assign new_n15470_ = new_n15552_ & new_n15553_;
  assign new_n15471_ = new_n15565_ & new_n15539_;
  assign new_n15472_ = new_n15568_ & new_n15569_;
  assign new_n15473_ = new_n15394_ & new_n15708_ & new_n15707_;
  assign new_n15474_ = new_n15711_ & new_n15539_;
  assign new_n15475_ = new_n15584_ & new_n15361_;
  assign new_n15476_ = new_n15718_ & new_n15538_;
  assign new_n15477_ = new_n15383_ & new_n15728_ & new_n15727_;
  assign new_n15478_ = new_n15731_ & new_n15537_;
  assign new_n15479_ = new_n15571_ & new_n15362_;
  assign new_n15480_ = new_n15616_ & new_n15534_;
  assign new_n15481_ = new_n15642_ & new_n15535_;
  assign new_n15482_ = new_n15658_ & new_n15659_;
  assign new_n15483_ = new_n15661_ & new_n15740_;
  assign new_n15484_ = new_n15662_ & new_n15659_ & new_n15658_;
  assign new_n15485_ = ~new_n15744_ | ~new_n15743_;
  assign new_n15486_ = new_n15439_ & new_n15749_ & new_n15748_;
  assign new_n15487_ = new_n15752_ & new_n15536_;
  assign new_n15488_ = ~new_n15758_ | ~new_n15757_;
  assign new_n15489_ = ~new_n15763_ | ~new_n15762_;
  assign new_n15490_ = new_n15769_ & new_n15535_;
  assign new_n15491_ = ~new_n15779_ | ~new_n15778_;
  assign new_n15492_ = ~new_n15784_ | ~new_n15783_;
  assign new_n15493_ = ~new_n15789_ | ~new_n15788_;
  assign new_n15494_ = ~new_n15794_ | ~new_n15793_;
  assign new_n15495_ = ~new_n15799_ | ~new_n15798_;
  assign new_n15496_ = new_n15805_ & new_n15534_;
  assign new_n15497_ = ~new_n15815_ | ~new_n15814_;
  assign new_n15498_ = ~new_n15820_ | ~new_n15819_;
  assign new_n15499_ = new_n15696_ & new_n15363_;
  assign new_n15500_ = new_n15826_ & new_n15533_;
  assign new_n15501_ = new_n15704_ & new_n15703_;
  assign new_n15502_ = ~new_n15472_ | ~new_n15566_;
  assign new_n15503_ = new_n15713_ & new_n15712_;
  assign new_n15504_ = new_n15720_ & new_n15719_;
  assign new_n15505_ = new_n15724_ & new_n15723_;
  assign new_n15506_ = ~new_n15470_ | ~new_n15550_;
  assign new_n15507_ = new_n15733_ & new_n15732_;
  assign new_n15508_ = ~new_n2955_;
  assign new_n15509_ = ~new_n1982_;
  assign new_n15510_ = new_n15742_ & new_n15741_;
  assign new_n15511_ = ~new_n15482_ | ~new_n15656_;
  assign new_n15512_ = new_n15754_ & new_n15753_;
  assign new_n15513_ = ~new_n15649_ | ~new_n15648_;
  assign new_n15514_ = ~new_n15645_ | ~new_n15644_;
  assign new_n15515_ = new_n15771_ & new_n15770_;
  assign new_n15516_ = new_n15775_ & new_n15774_;
  assign new_n15517_ = ~new_n15635_ | ~new_n15634_;
  assign new_n15518_ = ~new_n15631_ | ~new_n15630_;
  assign new_n15519_ = ~new_n2388_;
  assign new_n15520_ = ~new_n15627_ | ~new_n15626_;
  assign new_n15521_ = ~new_n2439_;
  assign new_n15522_ = ~new_n15619_ | ~new_n15618_;
  assign new_n15523_ = new_n15807_ & new_n15806_;
  assign new_n15524_ = new_n15811_ & new_n15810_;
  assign new_n15525_ = ~new_n15609_ | ~new_n15608_;
  assign new_n15526_ = ~new_n15605_ | ~new_n15604_;
  assign new_n15527_ = ~new_n15601_ | ~new_n15600_;
  assign new_n15528_ = new_n15828_ & new_n15827_;
  assign new_n15529_ = ~new_n15483_ | ~new_n15511_;
  assign new_n15530_ = ~new_n15439_;
  assign new_n15531_ = ~new_n15383_;
  assign new_n15532_ = ~new_n15394_;
  assign new_n15533_ = ~new_n2415_ | ~new_n15407_;
  assign new_n15534_ = ~new_n2430_ | ~new_n15416_;
  assign new_n15535_ = ~new_n2950_ | ~new_n15430_;
  assign new_n15536_ = ~new_n2946_ | ~new_n15438_;
  assign new_n15537_ = ~new_n2391_ | ~new_n15382_;
  assign new_n15538_ = ~new_n2400_ | ~new_n15389_;
  assign new_n15539_ = ~new_n2406_ | ~new_n15393_;
  assign new_n15540_ = ~new_n15418_;
  assign new_n15541_ = ~new_n15432_;
  assign new_n15542_ = ~new_n15391_;
  assign new_n15543_ = ~new_n15408_;
  assign new_n15544_ = ~new_n15379_;
  assign new_n15545_ = ~new_n15544_ | ~new_n15380_;
  assign new_n15546_ = ~new_n15545_ | ~new_n15519_;
  assign new_n15547_ = ~new_n2005_ | ~new_n15379_;
  assign new_n15548_ = ~new_n15400_;
  assign new_n15549_ = ~new_n2394_ | ~new_n15384_;
  assign new_n15550_ = ~new_n15469_ | ~new_n15400_;
  assign new_n15551_ = ~new_n15384_ | ~new_n15383_;
  assign new_n15552_ = ~new_n15551_ | ~new_n15381_;
  assign new_n15553_ = ~new_n1991_ | ~new_n15531_;
  assign new_n15554_ = ~new_n15506_;
  assign new_n15555_ = ~new_n2403_ | ~new_n15388_;
  assign new_n15556_ = ~new_n1998_ | ~new_n15385_;
  assign new_n15557_ = ~new_n1994_ | ~new_n15386_;
  assign new_n15558_ = ~new_n15542_ | ~new_n15360_;
  assign new_n15559_ = ~new_n15361_ | ~new_n15558_;
  assign new_n15560_ = ~new_n2397_ | ~new_n15390_;
  assign new_n15561_ = ~new_n2403_ | ~new_n15388_;
  assign new_n15562_ = ~new_n15360_ | ~new_n15560_ | ~new_n15506_;
  assign new_n15563_ = ~new_n15561_ | ~new_n15559_;
  assign new_n15564_ = ~new_n15398_;
  assign new_n15565_ = ~new_n2409_ | ~new_n15395_;
  assign new_n15566_ = ~new_n15471_ | ~new_n15398_;
  assign new_n15567_ = ~new_n15395_ | ~new_n15394_;
  assign new_n15568_ = ~new_n15567_ | ~new_n15392_;
  assign new_n15569_ = ~new_n2011_ | ~new_n15532_;
  assign new_n15570_ = ~new_n15502_;
  assign new_n15571_ = ~new_n2412_ | ~new_n15397_;
  assign new_n15572_ = ~new_n15571_ | ~new_n15408_;
  assign new_n15573_ = ~new_n15564_ | ~new_n15394_;
  assign new_n15574_ = ~new_n15474_ | ~new_n15573_;
  assign new_n15575_ = ~new_n15398_ | ~new_n15539_;
  assign new_n15576_ = ~new_n15473_ | ~new_n15575_;
  assign new_n15577_ = ~new_n15394_ | ~new_n15539_;
  assign new_n15578_ = ~new_n15560_ | ~new_n15506_;
  assign new_n15579_ = ~new_n15399_;
  assign new_n15580_ = ~new_n1994_ | ~new_n15386_;
  assign new_n15581_ = ~new_n15579_ | ~new_n15580_;
  assign new_n15582_ = ~new_n15476_ | ~new_n15581_;
  assign new_n15583_ = ~new_n15399_ | ~new_n15538_;
  assign new_n15584_ = ~new_n2403_ | ~new_n15388_;
  assign new_n15585_ = ~new_n15475_ | ~new_n15583_;
  assign new_n15586_ = ~new_n1994_ | ~new_n15386_;
  assign new_n15587_ = ~new_n15538_ | ~new_n15586_;
  assign new_n15588_ = ~new_n15560_ | ~new_n15391_;
  assign new_n15589_ = ~new_n15548_ | ~new_n15383_;
  assign new_n15590_ = ~new_n15478_ | ~new_n15589_;
  assign new_n15591_ = ~new_n15400_ | ~new_n15537_;
  assign new_n15592_ = ~new_n15477_ | ~new_n15591_;
  assign new_n15593_ = ~new_n15383_ | ~new_n15537_;
  assign new_n15594_ = ~new_n2418_ | ~new_n15406_;
  assign new_n15595_ = ~new_n1990_ | ~new_n15404_;
  assign new_n15596_ = ~new_n1989_ | ~new_n15405_;
  assign new_n15597_ = ~new_n15543_ | ~new_n15362_;
  assign new_n15598_ = ~new_n15363_ | ~new_n15597_;
  assign new_n15599_ = ~new_n2418_ | ~new_n15406_;
  assign new_n15600_ = ~new_n15479_ | ~new_n15502_;
  assign new_n15601_ = ~new_n15599_ | ~new_n15598_;
  assign new_n15602_ = ~new_n15527_;
  assign new_n15603_ = ~new_n2421_ | ~new_n15410_;
  assign new_n15604_ = ~new_n15603_ | ~new_n15527_;
  assign new_n15605_ = ~new_n1999_ | ~new_n15409_;
  assign new_n15606_ = ~new_n15526_;
  assign new_n15607_ = ~new_n2424_ | ~new_n15412_;
  assign new_n15608_ = ~new_n15607_ | ~new_n15526_;
  assign new_n15609_ = ~new_n2007_ | ~new_n15411_;
  assign new_n15610_ = ~new_n15525_;
  assign new_n15611_ = ~new_n2433_ | ~new_n15415_;
  assign new_n15612_ = ~new_n2000_ | ~new_n15413_;
  assign new_n15613_ = ~new_n2001_ | ~new_n15403_;
  assign new_n15614_ = ~new_n15540_ | ~new_n15534_;
  assign new_n15615_ = ~new_n15364_ | ~new_n15614_;
  assign new_n15616_ = ~new_n2427_ | ~new_n15417_;
  assign new_n15617_ = ~new_n2433_ | ~new_n15415_;
  assign new_n15618_ = ~new_n15611_ | ~new_n15525_ | ~new_n15480_;
  assign new_n15619_ = ~new_n15617_ | ~new_n15615_;
  assign new_n15620_ = ~new_n15522_;
  assign new_n15621_ = ~new_n2436_ | ~new_n15420_;
  assign new_n15622_ = ~new_n15621_ | ~new_n15522_;
  assign new_n15623_ = ~new_n1996_ | ~new_n15419_;
  assign new_n15624_ = ~new_n15421_;
  assign new_n15625_ = ~new_n15624_ | ~new_n15422_;
  assign new_n15626_ = ~new_n15625_ | ~new_n15521_;
  assign new_n15627_ = ~new_n2009_ | ~new_n15421_;
  assign new_n15628_ = ~new_n15520_;
  assign new_n15629_ = ~new_n2441_ | ~new_n15424_;
  assign new_n15630_ = ~new_n15629_ | ~new_n15520_;
  assign new_n15631_ = ~new_n2008_ | ~new_n15423_;
  assign new_n15632_ = ~new_n15518_;
  assign new_n15633_ = ~new_n2952_ | ~new_n15426_;
  assign new_n15634_ = ~new_n15633_ | ~new_n15518_;
  assign new_n15635_ = ~new_n2003_ | ~new_n15425_;
  assign new_n15636_ = ~new_n15517_;
  assign new_n15637_ = ~new_n2949_ | ~new_n15429_;
  assign new_n15638_ = ~new_n1993_ | ~new_n15427_;
  assign new_n15639_ = ~new_n1988_ | ~new_n15402_;
  assign new_n15640_ = ~new_n15541_ | ~new_n15535_;
  assign new_n15641_ = ~new_n15365_ | ~new_n15640_;
  assign new_n15642_ = ~new_n2951_ | ~new_n15431_;
  assign new_n15643_ = ~new_n2949_ | ~new_n15429_;
  assign new_n15644_ = ~new_n15637_ | ~new_n15517_ | ~new_n15481_;
  assign new_n15645_ = ~new_n15643_ | ~new_n15641_;
  assign new_n15646_ = ~new_n15514_;
  assign new_n15647_ = ~new_n2948_ | ~new_n15434_;
  assign new_n15648_ = ~new_n15647_ | ~new_n15514_;
  assign new_n15649_ = ~new_n1992_ | ~new_n15433_;
  assign new_n15650_ = ~new_n15513_;
  assign new_n15651_ = ~new_n2947_ | ~new_n15436_;
  assign new_n15652_ = ~new_n15651_ | ~new_n15513_;
  assign new_n15653_ = ~new_n1985_ | ~new_n15435_;
  assign new_n15654_ = ~new_n15443_;
  assign new_n15655_ = ~new_n2945_ | ~new_n15440_;
  assign new_n15656_ = ~new_n15655_ | ~new_n15443_ | ~new_n15536_;
  assign new_n15657_ = ~new_n15440_ | ~new_n15439_;
  assign new_n15658_ = ~new_n15657_ | ~new_n15437_;
  assign new_n15659_ = ~new_n1980_ | ~new_n15530_;
  assign new_n15660_ = ~new_n15511_;
  assign new_n15661_ = ~new_n2944_ | ~new_n15442_;
  assign new_n15662_ = ~new_n1981_ | ~new_n15441_;
  assign new_n15663_ = ~new_n15654_ | ~new_n15439_;
  assign new_n15664_ = ~new_n15487_ | ~new_n15663_;
  assign new_n15665_ = ~new_n15443_ | ~new_n15536_;
  assign new_n15666_ = ~new_n15486_ | ~new_n15665_;
  assign new_n15667_ = ~new_n15439_ | ~new_n15536_;
  assign new_n15668_ = ~new_n15642_ | ~new_n15517_;
  assign new_n15669_ = ~new_n15444_;
  assign new_n15670_ = ~new_n1988_ | ~new_n15402_;
  assign new_n15671_ = ~new_n15669_ | ~new_n15670_;
  assign new_n15672_ = ~new_n15490_ | ~new_n15671_;
  assign new_n15673_ = ~new_n15444_ | ~new_n15535_;
  assign new_n15674_ = ~new_n2949_ | ~new_n15429_;
  assign new_n15675_ = ~new_n15365_ | ~new_n15674_ | ~new_n15673_;
  assign new_n15676_ = ~new_n1988_ | ~new_n15402_;
  assign new_n15677_ = ~new_n15535_ | ~new_n15676_;
  assign new_n15678_ = ~new_n15642_ | ~new_n15432_;
  assign new_n15679_ = ~new_n15616_ | ~new_n15525_;
  assign new_n15680_ = ~new_n15445_;
  assign new_n15681_ = ~new_n2001_ | ~new_n15403_;
  assign new_n15682_ = ~new_n15680_ | ~new_n15681_;
  assign new_n15683_ = ~new_n15496_ | ~new_n15682_;
  assign new_n15684_ = ~new_n15445_ | ~new_n15534_;
  assign new_n15685_ = ~new_n2433_ | ~new_n15415_;
  assign new_n15686_ = ~new_n15364_ | ~new_n15685_ | ~new_n15684_;
  assign new_n15687_ = ~new_n2001_ | ~new_n15403_;
  assign new_n15688_ = ~new_n15534_ | ~new_n15687_;
  assign new_n15689_ = ~new_n15616_ | ~new_n15418_;
  assign new_n15690_ = ~new_n15571_ | ~new_n15502_;
  assign new_n15691_ = ~new_n15446_;
  assign new_n15692_ = ~new_n1989_ | ~new_n15405_;
  assign new_n15693_ = ~new_n15691_ | ~new_n15692_;
  assign new_n15694_ = ~new_n15500_ | ~new_n15693_;
  assign new_n15695_ = ~new_n15446_ | ~new_n15533_;
  assign new_n15696_ = ~new_n2418_ | ~new_n15406_;
  assign new_n15697_ = ~new_n15499_ | ~new_n15695_;
  assign new_n15698_ = ~new_n1989_ | ~new_n15405_;
  assign new_n15699_ = ~new_n15533_ | ~new_n15698_;
  assign new_n15700_ = ~new_n2004_ | ~new_n15378_;
  assign new_n15701_ = ~new_n15655_ | ~new_n15443_ | ~new_n15536_;
  assign new_n15702_ = ~new_n15484_ | ~new_n15366_ | ~new_n15701_;
  assign new_n15703_ = ~new_n2412_ | ~new_n15397_;
  assign new_n15704_ = ~new_n2010_ | ~new_n15396_;
  assign new_n15705_ = ~new_n15572_ | ~new_n15502_;
  assign new_n15706_ = ~new_n15570_ | ~new_n15501_;
  assign new_n15707_ = ~new_n2409_ | ~new_n15395_;
  assign new_n15708_ = ~new_n2011_ | ~new_n15392_;
  assign new_n15709_ = ~new_n2409_ | ~new_n15395_;
  assign new_n15710_ = ~new_n2011_ | ~new_n15392_;
  assign new_n15711_ = ~new_n15710_ | ~new_n15709_;
  assign new_n15712_ = ~new_n2406_ | ~new_n15393_;
  assign new_n15713_ = ~new_n1997_ | ~new_n15376_;
  assign new_n15714_ = ~new_n15577_ | ~new_n15398_;
  assign new_n15715_ = ~new_n15503_ | ~new_n15564_;
  assign new_n15716_ = ~new_n2403_ | ~new_n15388_;
  assign new_n15717_ = ~new_n1998_ | ~new_n15385_;
  assign new_n15718_ = ~new_n15717_ | ~new_n15716_;
  assign new_n15719_ = ~new_n2400_ | ~new_n15389_;
  assign new_n15720_ = ~new_n1994_ | ~new_n15386_;
  assign new_n15721_ = ~new_n15587_ | ~new_n15399_;
  assign new_n15722_ = ~new_n15504_ | ~new_n15579_;
  assign new_n15723_ = ~new_n2397_ | ~new_n15390_;
  assign new_n15724_ = ~new_n1987_ | ~new_n15387_;
  assign new_n15725_ = ~new_n15588_ | ~new_n15506_;
  assign new_n15726_ = ~new_n15554_ | ~new_n15505_;
  assign new_n15727_ = ~new_n2394_ | ~new_n15384_;
  assign new_n15728_ = ~new_n1991_ | ~new_n15381_;
  assign new_n15729_ = ~new_n2394_ | ~new_n15384_;
  assign new_n15730_ = ~new_n1991_ | ~new_n15381_;
  assign new_n15731_ = ~new_n15730_ | ~new_n15729_;
  assign new_n15732_ = ~new_n2391_ | ~new_n15382_;
  assign new_n15733_ = ~new_n1995_ | ~new_n15377_;
  assign new_n15734_ = ~new_n15593_ | ~new_n15400_;
  assign new_n15735_ = ~new_n15507_ | ~new_n15548_;
  assign new_n15736_ = ~new_n2955_ | ~new_n15509_;
  assign new_n15737_ = ~new_n1982_ | ~new_n15508_;
  assign new_n15738_ = ~new_n2955_ | ~new_n15509_;
  assign new_n15739_ = ~new_n1982_ | ~new_n15508_;
  assign new_n15740_ = ~new_n15739_ | ~new_n15738_;
  assign new_n15741_ = ~new_n15441_ | ~new_n1981_ | ~new_n15740_;
  assign new_n15742_ = ~new_n2944_ | ~new_n15366_ | ~new_n15442_;
  assign new_n15743_ = ~new_n2944_ | ~new_n15442_;
  assign new_n15744_ = ~new_n1981_ | ~new_n15441_;
  assign new_n15745_ = ~new_n15485_;
  assign new_n15746_ = ~new_n15660_ | ~new_n15745_;
  assign new_n15747_ = ~new_n15485_ | ~new_n15511_;
  assign new_n15748_ = ~new_n2945_ | ~new_n15440_;
  assign new_n15749_ = ~new_n1980_ | ~new_n15437_;
  assign new_n15750_ = ~new_n2945_ | ~new_n15440_;
  assign new_n15751_ = ~new_n1980_ | ~new_n15437_;
  assign new_n15752_ = ~new_n15751_ | ~new_n15750_;
  assign new_n15753_ = ~new_n2946_ | ~new_n15438_;
  assign new_n15754_ = ~new_n1984_ | ~new_n15401_;
  assign new_n15755_ = ~new_n15667_ | ~new_n15443_;
  assign new_n15756_ = ~new_n15512_ | ~new_n15654_;
  assign new_n15757_ = ~new_n2947_ | ~new_n15436_;
  assign new_n15758_ = ~new_n1985_ | ~new_n15435_;
  assign new_n15759_ = ~new_n15488_;
  assign new_n15760_ = ~new_n15650_ | ~new_n15759_;
  assign new_n15761_ = ~new_n15488_ | ~new_n15513_;
  assign new_n15762_ = ~new_n2948_ | ~new_n15434_;
  assign new_n15763_ = ~new_n1992_ | ~new_n15433_;
  assign new_n15764_ = ~new_n15489_;
  assign new_n15765_ = ~new_n15646_ | ~new_n15764_;
  assign new_n15766_ = ~new_n15489_ | ~new_n15514_;
  assign new_n15767_ = ~new_n2949_ | ~new_n15429_;
  assign new_n15768_ = ~new_n1993_ | ~new_n15427_;
  assign new_n15769_ = ~new_n15768_ | ~new_n15767_;
  assign new_n15770_ = ~new_n2950_ | ~new_n15430_;
  assign new_n15771_ = ~new_n1988_ | ~new_n15402_;
  assign new_n15772_ = ~new_n15677_ | ~new_n15444_;
  assign new_n15773_ = ~new_n15515_ | ~new_n15669_;
  assign new_n15774_ = ~new_n2951_ | ~new_n15431_;
  assign new_n15775_ = ~new_n2002_ | ~new_n15428_;
  assign new_n15776_ = ~new_n15678_ | ~new_n15517_;
  assign new_n15777_ = ~new_n15636_ | ~new_n15516_;
  assign new_n15778_ = ~new_n2952_ | ~new_n15426_;
  assign new_n15779_ = ~new_n2003_ | ~new_n15425_;
  assign new_n15780_ = ~new_n15491_;
  assign new_n15781_ = ~new_n15632_ | ~new_n15780_;
  assign new_n15782_ = ~new_n15491_ | ~new_n15518_;
  assign new_n15783_ = ~new_n2388_ | ~new_n15380_;
  assign new_n15784_ = ~new_n2005_ | ~new_n15519_;
  assign new_n15785_ = ~new_n15492_;
  assign new_n15786_ = ~new_n15785_ | ~new_n15544_;
  assign new_n15787_ = ~new_n15492_ | ~new_n15379_;
  assign new_n15788_ = ~new_n2441_ | ~new_n15424_;
  assign new_n15789_ = ~new_n2008_ | ~new_n15423_;
  assign new_n15790_ = ~new_n15493_;
  assign new_n15791_ = ~new_n15628_ | ~new_n15790_;
  assign new_n15792_ = ~new_n15493_ | ~new_n15520_;
  assign new_n15793_ = ~new_n2439_ | ~new_n15422_;
  assign new_n15794_ = ~new_n2009_ | ~new_n15521_;
  assign new_n15795_ = ~new_n15494_;
  assign new_n15796_ = ~new_n15795_ | ~new_n15624_;
  assign new_n15797_ = ~new_n15494_ | ~new_n15421_;
  assign new_n15798_ = ~new_n2436_ | ~new_n15420_;
  assign new_n15799_ = ~new_n1996_ | ~new_n15419_;
  assign new_n15800_ = ~new_n15495_;
  assign new_n15801_ = ~new_n15620_ | ~new_n15800_;
  assign new_n15802_ = ~new_n15495_ | ~new_n15522_;
  assign new_n15803_ = ~new_n2433_ | ~new_n15415_;
  assign new_n15804_ = ~new_n2000_ | ~new_n15413_;
  assign new_n15805_ = ~new_n15804_ | ~new_n15803_;
  assign new_n15806_ = ~new_n2430_ | ~new_n15416_;
  assign new_n15807_ = ~new_n2001_ | ~new_n15403_;
  assign new_n15808_ = ~new_n15688_ | ~new_n15445_;
  assign new_n15809_ = ~new_n15523_ | ~new_n15680_;
  assign new_n15810_ = ~new_n2427_ | ~new_n15417_;
  assign new_n15811_ = ~new_n2006_ | ~new_n15414_;
  assign new_n15812_ = ~new_n15689_ | ~new_n15525_;
  assign new_n15813_ = ~new_n15610_ | ~new_n15524_;
  assign new_n15814_ = ~new_n2424_ | ~new_n15412_;
  assign new_n15815_ = ~new_n2007_ | ~new_n15411_;
  assign new_n15816_ = ~new_n15497_;
  assign new_n15817_ = ~new_n15606_ | ~new_n15816_;
  assign new_n15818_ = ~new_n15497_ | ~new_n15526_;
  assign new_n15819_ = ~new_n2421_ | ~new_n15410_;
  assign new_n15820_ = ~new_n1999_ | ~new_n15409_;
  assign new_n15821_ = ~new_n15498_;
  assign new_n15822_ = ~new_n15602_ | ~new_n15821_;
  assign new_n15823_ = ~new_n15498_ | ~new_n15527_;
  assign new_n15824_ = ~new_n2418_ | ~new_n15406_;
  assign new_n15825_ = ~new_n1990_ | ~new_n15404_;
  assign new_n15826_ = ~new_n15825_ | ~new_n15824_;
  assign new_n15827_ = ~new_n2415_ | ~new_n15407_;
  assign new_n15828_ = ~new_n1989_ | ~new_n15405_;
  assign new_n15829_ = ~new_n15699_ | ~new_n15446_;
  assign new_n15830_ = ~new_n15528_ | ~new_n15691_;
  assign new_n15831_ = new_n16029_ & new_n16028_;
  assign new_n15832_ = new_n16044_ & new_n16043_;
  assign new_n15833_ = new_n16078_ & new_n16077_;
  assign new_n15834_ = new_n16096_ & new_n16095_;
  assign new_n15835_ = new_n16108_ & new_n16107_;
  assign new_n15836_ = new_n16166_ & new_n16163_;
  assign new_n15837_ = new_n16157_ & new_n16154_;
  assign new_n15838_ = new_n16150_ & new_n16147_;
  assign new_n15839_ = new_n16141_ & new_n16138_;
  assign new_n15840_ = new_n16067_ & new_n16064_;
  assign new_n15841_ = new_n16060_ & new_n16057_;
  assign new_n15842_ = ~new_n2138_;
  assign new_n15843_ = ~new_n2102_;
  assign new_n15844_ = ~new_n2102_ | ~new_n15886_;
  assign new_n15845_ = ~new_n2101_;
  assign new_n15846_ = ~new_n2106_;
  assign new_n15847_ = ~new_n2106_ | ~new_n15888_;
  assign new_n15848_ = ~new_n2105_;
  assign new_n15849_ = ~new_n2108_;
  assign new_n15850_ = ~new_n2107_;
  assign new_n15851_ = ~new_n15937_ | ~new_n16033_;
  assign new_n15852_ = ~new_n2104_;
  assign new_n15853_ = ~new_n2103_;
  assign new_n15854_ = ~new_n2100_;
  assign new_n15855_ = ~new_n2099_;
  assign new_n15856_ = ~new_n16053_ | ~new_n16052_;
  assign new_n15857_ = ~new_n16041_ | ~new_n16040_;
  assign new_n15858_ = ~new_n16026_ | ~new_n16025_;
  assign new_n15859_ = ~new_n2081_;
  assign new_n15860_ = ~new_n2082_;
  assign new_n15861_ = ~new_n2083_;
  assign new_n15862_ = ~new_n2084_;
  assign new_n15863_ = ~new_n2087_;
  assign new_n15864_ = ~new_n2092_;
  assign new_n15865_ = ~new_n2092_ | ~new_n15900_;
  assign new_n15866_ = ~new_n2091_;
  assign new_n15867_ = ~new_n2098_;
  assign new_n15868_ = ~new_n2096_;
  assign new_n15869_ = ~new_n2097_;
  assign new_n15870_ = ~new_n2097_ | ~new_n15903_;
  assign new_n15871_ = ~new_n2095_;
  assign new_n15872_ = ~new_n2094_;
  assign new_n15873_ = ~new_n2093_;
  assign new_n15874_ = ~new_n2090_;
  assign new_n15875_ = ~new_n2089_;
  assign new_n15876_ = ~new_n2089_ | ~new_n15909_;
  assign new_n15877_ = ~new_n2088_;
  assign new_n15878_ = ~new_n2086_;
  assign new_n15879_ = ~new_n2085_;
  assign new_n15880_ = ~new_n2082_ | ~new_n15897_;
  assign new_n15881_ = ~new_n16019_ | ~new_n16134_;
  assign new_n15882_ = ~new_n15876_ | ~new_n16143_;
  assign new_n15883_ = ~new_n16093_ | ~new_n16092_;
  assign new_n15884_ = ~new_n15870_ | ~new_n16159_;
  assign new_n15885_ = ~new_n16186_ | ~new_n16185_;
  assign new_n15886_ = ~new_n16215_ | ~new_n16214_;
  assign new_n15887_ = ~new_n16212_ | ~new_n16211_;
  assign new_n15888_ = ~new_n16203_ | ~new_n16202_;
  assign new_n15889_ = ~new_n16200_ | ~new_n16199_;
  assign new_n15890_ = ~new_n16194_ | ~new_n16193_;
  assign new_n15891_ = ~new_n16197_ | ~new_n16196_;
  assign new_n15892_ = ~new_n16206_ | ~new_n16205_;
  assign new_n15893_ = ~new_n16209_ | ~new_n16208_;
  assign new_n15894_ = ~new_n16218_ | ~new_n16217_;
  assign new_n15895_ = ~new_n16258_ | ~new_n16257_;
  assign new_n15896_ = ~new_n16261_ | ~new_n16260_;
  assign new_n15897_ = ~new_n16264_ | ~new_n16263_;
  assign new_n15898_ = ~new_n16267_ | ~new_n16266_;
  assign new_n15899_ = ~new_n16270_ | ~new_n16269_;
  assign new_n15900_ = ~new_n16300_ | ~new_n16299_;
  assign new_n15901_ = ~new_n16297_ | ~new_n16296_;
  assign new_n15902_ = ~new_n16279_ | ~new_n16278_;
  assign new_n15903_ = ~new_n16288_ | ~new_n16287_;
  assign new_n15904_ = ~new_n16282_ | ~new_n16281_;
  assign new_n15905_ = ~new_n16285_ | ~new_n16284_;
  assign new_n15906_ = ~new_n16291_ | ~new_n16290_;
  assign new_n15907_ = ~new_n16294_ | ~new_n16293_;
  assign new_n15908_ = ~new_n16303_ | ~new_n16302_;
  assign new_n15909_ = ~new_n16276_ | ~new_n16275_;
  assign new_n15910_ = ~new_n16273_ | ~new_n16272_;
  assign new_n15911_ = ~new_n16306_ | ~new_n16305_;
  assign new_n15912_ = ~new_n16309_ | ~new_n16308_;
  assign new_n15913_ = ~new_n16315_ | ~new_n16314_;
  assign new_n15914_ = ~new_n16422_ | ~new_n16421_;
  assign new_n15915_ = ~new_n16221_ | ~new_n16220_;
  assign new_n15916_ = ~new_n16228_ | ~new_n16227_;
  assign new_n15917_ = ~new_n16235_ | ~new_n16234_;
  assign new_n15918_ = ~new_n16242_ | ~new_n16241_;
  assign new_n15919_ = ~new_n16249_ | ~new_n16248_;
  assign new_n15920_ = ~new_n16256_ | ~new_n16255_;
  assign new_n15921_ = ~new_n16318_ | ~new_n16317_;
  assign new_n15922_ = ~new_n16325_ | ~new_n16324_;
  assign new_n15923_ = ~new_n16332_ | ~new_n16331_;
  assign new_n15924_ = ~new_n16337_ | ~new_n16336_;
  assign new_n15925_ = ~new_n16344_ | ~new_n16343_;
  assign new_n15926_ = ~new_n16351_ | ~new_n16350_;
  assign new_n15927_ = ~new_n16358_ | ~new_n16357_;
  assign new_n15928_ = ~new_n16365_ | ~new_n16364_;
  assign new_n15929_ = ~new_n16370_ | ~new_n16369_;
  assign new_n15930_ = ~new_n16377_ | ~new_n16376_;
  assign new_n15931_ = ~new_n16384_ | ~new_n16383_;
  assign new_n15932_ = ~new_n16391_ | ~new_n16390_;
  assign new_n15933_ = ~new_n16398_ | ~new_n16397_;
  assign new_n15934_ = ~new_n16405_ | ~new_n16404_;
  assign new_n15935_ = ~new_n16410_ | ~new_n16409_;
  assign new_n15936_ = ~new_n16417_ | ~new_n16416_;
  assign new_n15937_ = new_n16032_ & new_n16031_;
  assign new_n15938_ = new_n16048_ & new_n16047_;
  assign new_n15939_ = new_n15844_ & new_n16230_ & new_n16229_;
  assign new_n15940_ = new_n16059_ & new_n15832_;
  assign new_n15941_ = new_n15847_ & new_n16251_ & new_n16250_;
  assign new_n15942_ = new_n16066_ & new_n15831_;
  assign new_n15943_ = new_n16082_ & new_n15833_;
  assign new_n15944_ = new_n16080_ & new_n16014_;
  assign new_n15945_ = new_n16100_ & new_n16099_;
  assign new_n15946_ = new_n16184_ & new_n15880_;
  assign new_n15947_ = new_n16133_ & new_n16128_;
  assign new_n15948_ = new_n16181_ & new_n16132_;
  assign new_n15949_ = ~new_n16312_ | ~new_n16311_;
  assign new_n15950_ = new_n16016_ & new_n16327_ & new_n16326_;
  assign new_n15951_ = new_n16015_ & new_n16353_ & new_n16352_;
  assign new_n15952_ = new_n15865_ & new_n16379_ & new_n16378_;
  assign new_n15953_ = new_n16156_ & new_n15834_;
  assign new_n15954_ = new_n16014_ & new_n16400_ & new_n16399_;
  assign new_n15955_ = new_n16165_ & new_n15833_;
  assign new_n15956_ = ~new_n16419_ | ~new_n16418_;
  assign new_n15957_ = ~new_n2128_;
  assign new_n15958_ = new_n16189_ & new_n16188_;
  assign new_n15959_ = ~new_n2137_;
  assign new_n15960_ = ~new_n2136_;
  assign new_n15961_ = ~new_n2134_;
  assign new_n15962_ = ~new_n2135_;
  assign new_n15963_ = ~new_n2133_;
  assign new_n15964_ = ~new_n2132_;
  assign new_n15965_ = ~new_n2130_;
  assign new_n15966_ = ~new_n2131_;
  assign new_n15967_ = ~new_n2129_;
  assign new_n15968_ = new_n16223_ & new_n16222_;
  assign new_n15969_ = ~new_n15938_ | ~new_n16049_;
  assign new_n15970_ = new_n16237_ & new_n16236_;
  assign new_n15971_ = ~new_n16037_ | ~new_n16036_;
  assign new_n15972_ = new_n16244_ & new_n16243_;
  assign new_n15973_ = ~new_n2110_;
  assign new_n15974_ = ~new_n2112_;
  assign new_n15975_ = ~new_n2111_;
  assign new_n15976_ = ~new_n2113_;
  assign new_n15977_ = ~new_n2116_;
  assign new_n15978_ = ~new_n2117_;
  assign new_n15979_ = ~new_n2118_;
  assign new_n15980_ = ~new_n2127_;
  assign new_n15981_ = ~new_n2124_;
  assign new_n15982_ = ~new_n2125_;
  assign new_n15983_ = ~new_n2126_;
  assign new_n15984_ = ~new_n2123_;
  assign new_n15985_ = ~new_n2122_;
  assign new_n15986_ = ~new_n2120_;
  assign new_n15987_ = ~new_n2121_;
  assign new_n15988_ = ~new_n2119_;
  assign new_n15989_ = ~new_n2115_;
  assign new_n15990_ = ~new_n2114_;
  assign new_n15991_ = ~new_n2080_;
  assign new_n15992_ = ~new_n2109_;
  assign new_n15993_ = new_n16320_ & new_n16319_;
  assign new_n15994_ = ~new_n15880_ | ~new_n16178_ | ~new_n16129_;
  assign new_n15995_ = ~new_n16123_ | ~new_n16122_;
  assign new_n15996_ = new_n16339_ & new_n16338_;
  assign new_n15997_ = ~new_n16119_ | ~new_n16118_;
  assign new_n15998_ = new_n16346_ & new_n16345_;
  assign new_n15999_ = ~new_n16115_ | ~new_n16114_ | ~new_n16110_;
  assign new_n16000_ = new_n16360_ & new_n16359_;
  assign new_n16001_ = ~new_n16022_ | ~new_n16021_;
  assign new_n16002_ = ~new_n16105_ | ~new_n16104_;
  assign new_n16003_ = new_n16372_ & new_n16371_;
  assign new_n16004_ = ~new_n15945_ | ~new_n16101_;
  assign new_n16005_ = new_n16386_ & new_n16385_;
  assign new_n16006_ = ~new_n16089_ | ~new_n16088_;
  assign new_n16007_ = new_n16393_ & new_n16392_;
  assign new_n16008_ = ~new_n16085_ | ~new_n16084_;
  assign new_n16009_ = ~new_n16075_ | ~new_n16074_;
  assign new_n16010_ = new_n16412_ & new_n16411_;
  assign new_n16011_ = ~new_n16071_ | ~new_n16070_;
  assign new_n16012_ = ~new_n16180_ | ~new_n16179_;
  assign new_n16013_ = ~new_n15847_;
  assign new_n16014_ = ~new_n2096_ | ~new_n15905_;
  assign new_n16015_ = ~new_n2088_ | ~new_n15910_;
  assign new_n16016_ = ~new_n2083_ | ~new_n15896_;
  assign new_n16017_ = ~new_n15870_;
  assign new_n16018_ = ~new_n15876_;
  assign new_n16019_ = ~new_n2084_ | ~new_n15898_;
  assign new_n16020_ = new_n2138_ | new_n2108_;
  assign new_n16021_ = ~new_n15890_ | ~new_n16020_;
  assign new_n16022_ = ~new_n2108_ | ~new_n2138_;
  assign new_n16023_ = ~new_n16001_;
  assign new_n16024_ = ~new_n16198_ | ~new_n15850_;
  assign new_n16025_ = ~new_n16024_ | ~new_n16001_;
  assign new_n16026_ = ~new_n2107_ | ~new_n15891_;
  assign new_n16027_ = ~new_n15858_;
  assign new_n16028_ = ~new_n16201_ | ~new_n15848_;
  assign new_n16029_ = ~new_n16204_ | ~new_n15846_;
  assign new_n16030_ = ~new_n15848_ | ~new_n15847_;
  assign new_n16031_ = ~new_n15889_ | ~new_n16030_;
  assign new_n16032_ = ~new_n2105_ | ~new_n16013_;
  assign new_n16033_ = ~new_n15831_ | ~new_n15858_;
  assign new_n16034_ = ~new_n15851_;
  assign new_n16035_ = ~new_n16034_ | ~new_n15852_;
  assign new_n16036_ = ~new_n15892_ | ~new_n16035_;
  assign new_n16037_ = ~new_n2104_ | ~new_n15851_;
  assign new_n16038_ = ~new_n15971_;
  assign new_n16039_ = ~new_n16210_ | ~new_n15853_;
  assign new_n16040_ = ~new_n16039_ | ~new_n15971_;
  assign new_n16041_ = ~new_n2103_ | ~new_n15893_;
  assign new_n16042_ = ~new_n15857_;
  assign new_n16043_ = ~new_n16213_ | ~new_n15845_;
  assign new_n16044_ = ~new_n16216_ | ~new_n15843_;
  assign new_n16045_ = ~new_n15844_;
  assign new_n16046_ = ~new_n15845_ | ~new_n15844_;
  assign new_n16047_ = ~new_n15887_ | ~new_n16046_;
  assign new_n16048_ = ~new_n2101_ | ~new_n16045_;
  assign new_n16049_ = ~new_n15832_ | ~new_n15857_;
  assign new_n16050_ = ~new_n15969_;
  assign new_n16051_ = ~new_n16219_ | ~new_n15854_;
  assign new_n16052_ = ~new_n16051_ | ~new_n15969_;
  assign new_n16053_ = ~new_n2100_ | ~new_n15894_;
  assign new_n16054_ = ~new_n15856_;
  assign new_n16055_ = ~new_n16216_ | ~new_n15843_;
  assign new_n16056_ = ~new_n16055_ | ~new_n15857_;
  assign new_n16057_ = ~new_n15939_ | ~new_n16056_;
  assign new_n16058_ = ~new_n16042_ | ~new_n15844_;
  assign new_n16059_ = ~new_n2101_ | ~new_n15887_;
  assign new_n16060_ = ~new_n15940_ | ~new_n16058_;
  assign new_n16061_ = ~new_n16216_ | ~new_n15843_;
  assign new_n16062_ = ~new_n16204_ | ~new_n15846_;
  assign new_n16063_ = ~new_n16062_ | ~new_n15858_;
  assign new_n16064_ = ~new_n15941_ | ~new_n16063_;
  assign new_n16065_ = ~new_n16027_ | ~new_n15847_;
  assign new_n16066_ = ~new_n2105_ | ~new_n15889_;
  assign new_n16067_ = ~new_n15942_ | ~new_n16065_;
  assign new_n16068_ = ~new_n16204_ | ~new_n15846_;
  assign new_n16069_ = ~new_n16054_ | ~new_n15855_;
  assign new_n16070_ = ~new_n15885_ | ~new_n16069_;
  assign new_n16071_ = ~new_n2099_ | ~new_n15856_;
  assign new_n16072_ = ~new_n16011_;
  assign new_n16073_ = ~new_n16280_ | ~new_n15867_;
  assign new_n16074_ = ~new_n16073_ | ~new_n16011_;
  assign new_n16075_ = ~new_n2098_ | ~new_n15902_;
  assign new_n16076_ = ~new_n16009_;
  assign new_n16077_ = ~new_n16283_ | ~new_n15871_;
  assign new_n16078_ = ~new_n16286_ | ~new_n15868_;
  assign new_n16079_ = ~new_n16017_ | ~new_n15833_;
  assign new_n16080_ = ~new_n2095_ | ~new_n15904_;
  assign new_n16081_ = ~new_n15944_ | ~new_n16079_;
  assign new_n16082_ = ~new_n16289_ | ~new_n15869_;
  assign new_n16083_ = ~new_n16283_ | ~new_n15871_;
  assign new_n16084_ = ~new_n15943_ | ~new_n16009_;
  assign new_n16085_ = ~new_n16083_ | ~new_n16081_;
  assign new_n16086_ = ~new_n16008_;
  assign new_n16087_ = ~new_n16292_ | ~new_n15872_;
  assign new_n16088_ = ~new_n16087_ | ~new_n16008_;
  assign new_n16089_ = ~new_n2094_ | ~new_n15906_;
  assign new_n16090_ = ~new_n16006_;
  assign new_n16091_ = ~new_n16295_ | ~new_n15873_;
  assign new_n16092_ = ~new_n16091_ | ~new_n16006_;
  assign new_n16093_ = ~new_n2093_ | ~new_n15907_;
  assign new_n16094_ = ~new_n15883_;
  assign new_n16095_ = ~new_n16298_ | ~new_n15866_;
  assign new_n16096_ = ~new_n16301_ | ~new_n15864_;
  assign new_n16097_ = ~new_n15865_;
  assign new_n16098_ = ~new_n15866_ | ~new_n15865_;
  assign new_n16099_ = ~new_n15901_ | ~new_n16098_;
  assign new_n16100_ = ~new_n2091_ | ~new_n16097_;
  assign new_n16101_ = ~new_n15834_ | ~new_n15883_;
  assign new_n16102_ = ~new_n16004_;
  assign new_n16103_ = ~new_n16304_ | ~new_n15874_;
  assign new_n16104_ = ~new_n16103_ | ~new_n16004_;
  assign new_n16105_ = ~new_n2090_ | ~new_n15908_;
  assign new_n16106_ = ~new_n16002_;
  assign new_n16107_ = ~new_n16271_ | ~new_n15863_;
  assign new_n16108_ = ~new_n16274_ | ~new_n15877_;
  assign new_n16109_ = ~new_n16018_ | ~new_n15835_;
  assign new_n16110_ = ~new_n2087_ | ~new_n15899_;
  assign new_n16111_ = ~new_n16015_ | ~new_n16109_;
  assign new_n16112_ = ~new_n16277_ | ~new_n15875_;
  assign new_n16113_ = ~new_n16271_ | ~new_n15863_;
  assign new_n16114_ = ~new_n15835_ | ~new_n16112_ | ~new_n16002_;
  assign new_n16115_ = ~new_n16113_ | ~new_n16111_;
  assign new_n16116_ = ~new_n15999_;
  assign new_n16117_ = ~new_n16307_ | ~new_n15878_;
  assign new_n16118_ = ~new_n16117_ | ~new_n15999_;
  assign new_n16119_ = ~new_n2086_ | ~new_n15911_;
  assign new_n16120_ = ~new_n15997_;
  assign new_n16121_ = ~new_n16310_ | ~new_n15879_;
  assign new_n16122_ = ~new_n16121_ | ~new_n15997_;
  assign new_n16123_ = ~new_n2085_ | ~new_n15912_;
  assign new_n16124_ = ~new_n15995_;
  assign new_n16125_ = ~new_n16262_ | ~new_n15861_;
  assign new_n16126_ = ~new_n16019_ | ~new_n16016_;
  assign new_n16127_ = ~new_n15880_;
  assign new_n16128_ = ~new_n16268_ | ~new_n15862_;
  assign new_n16129_ = ~new_n16012_ | ~new_n15995_ | ~new_n16128_;
  assign new_n16130_ = ~new_n15994_;
  assign new_n16131_ = ~new_n16259_ | ~new_n15859_;
  assign new_n16132_ = ~new_n2081_ | ~new_n15895_;
  assign new_n16133_ = ~new_n16259_ | ~new_n15859_;
  assign new_n16134_ = ~new_n16128_ | ~new_n15995_;
  assign new_n16135_ = ~new_n15881_;
  assign new_n16136_ = ~new_n16262_ | ~new_n15861_;
  assign new_n16137_ = ~new_n16136_ | ~new_n15881_;
  assign new_n16138_ = ~new_n15950_ | ~new_n16137_;
  assign new_n16139_ = ~new_n16135_ | ~new_n16016_;
  assign new_n16140_ = ~new_n2082_ | ~new_n15897_;
  assign new_n16141_ = ~new_n16012_ | ~new_n16139_ | ~new_n16140_;
  assign new_n16142_ = ~new_n16262_ | ~new_n15861_;
  assign new_n16143_ = ~new_n16112_ | ~new_n16002_;
  assign new_n16144_ = ~new_n15882_;
  assign new_n16145_ = ~new_n16274_ | ~new_n15877_;
  assign new_n16146_ = ~new_n16145_ | ~new_n15882_;
  assign new_n16147_ = ~new_n15951_ | ~new_n16146_;
  assign new_n16148_ = ~new_n16144_ | ~new_n16015_;
  assign new_n16149_ = ~new_n2087_ | ~new_n15899_;
  assign new_n16150_ = ~new_n15835_ | ~new_n16149_ | ~new_n16148_;
  assign new_n16151_ = ~new_n16274_ | ~new_n15877_;
  assign new_n16152_ = ~new_n16301_ | ~new_n15864_;
  assign new_n16153_ = ~new_n16152_ | ~new_n15883_;
  assign new_n16154_ = ~new_n15952_ | ~new_n16153_;
  assign new_n16155_ = ~new_n16094_ | ~new_n15865_;
  assign new_n16156_ = ~new_n2091_ | ~new_n15901_;
  assign new_n16157_ = ~new_n15953_ | ~new_n16155_;
  assign new_n16158_ = ~new_n16301_ | ~new_n15864_;
  assign new_n16159_ = ~new_n16082_ | ~new_n16009_;
  assign new_n16160_ = ~new_n15884_;
  assign new_n16161_ = ~new_n16286_ | ~new_n15868_;
  assign new_n16162_ = ~new_n16161_ | ~new_n15884_;
  assign new_n16163_ = ~new_n15954_ | ~new_n16162_;
  assign new_n16164_ = ~new_n16160_ | ~new_n16014_;
  assign new_n16165_ = ~new_n2095_ | ~new_n15904_;
  assign new_n16166_ = ~new_n15955_ | ~new_n16164_;
  assign new_n16167_ = ~new_n16286_ | ~new_n15868_;
  assign new_n16168_ = ~new_n16061_ | ~new_n15844_;
  assign new_n16169_ = ~new_n16068_ | ~new_n15847_;
  assign new_n16170_ = ~new_n16142_ | ~new_n16016_;
  assign new_n16171_ = ~new_n16128_ | ~new_n16019_;
  assign new_n16172_ = ~new_n16151_ | ~new_n16015_;
  assign new_n16173_ = ~new_n16112_ | ~new_n15876_;
  assign new_n16174_ = ~new_n16158_ | ~new_n15865_;
  assign new_n16175_ = ~new_n16167_ | ~new_n16014_;
  assign new_n16176_ = ~new_n16082_ | ~new_n15870_;
  assign new_n16177_ = ~new_n15946_ | ~new_n16178_ | ~new_n16129_;
  assign new_n16178_ = ~new_n16126_ | ~new_n16012_;
  assign new_n16179_ = ~new_n15897_ | ~new_n16125_;
  assign new_n16180_ = ~new_n2082_ | ~new_n16125_;
  assign new_n16181_ = ~new_n16133_ | ~new_n16126_ | ~new_n16012_;
  assign new_n16182_ = ~new_n15947_ | ~new_n15995_ | ~new_n16012_;
  assign new_n16183_ = ~new_n16127_ | ~new_n16133_;
  assign new_n16184_ = ~new_n2081_ | ~new_n15895_;
  assign new_n16185_ = ~new_n2138_ | ~new_n15957_;
  assign new_n16186_ = ~new_n2128_ | ~new_n15842_;
  assign new_n16187_ = ~new_n15885_;
  assign new_n16188_ = ~new_n16187_ | ~new_n2099_;
  assign new_n16189_ = ~new_n15885_ | ~new_n15855_;
  assign new_n16190_ = ~new_n16187_ | ~new_n2099_;
  assign new_n16191_ = ~new_n15885_ | ~new_n15855_;
  assign new_n16192_ = ~new_n16191_ | ~new_n16190_;
  assign new_n16193_ = ~new_n2138_ | ~new_n15959_;
  assign new_n16194_ = ~new_n2137_ | ~new_n15842_;
  assign new_n16195_ = ~new_n15890_;
  assign new_n16196_ = ~new_n2138_ | ~new_n15960_;
  assign new_n16197_ = ~new_n2136_ | ~new_n15842_;
  assign new_n16198_ = ~new_n15891_;
  assign new_n16199_ = ~new_n2138_ | ~new_n15961_;
  assign new_n16200_ = ~new_n2134_ | ~new_n15842_;
  assign new_n16201_ = ~new_n15889_;
  assign new_n16202_ = ~new_n2138_ | ~new_n15962_;
  assign new_n16203_ = ~new_n2135_ | ~new_n15842_;
  assign new_n16204_ = ~new_n15888_;
  assign new_n16205_ = ~new_n2138_ | ~new_n15963_;
  assign new_n16206_ = ~new_n2133_ | ~new_n15842_;
  assign new_n16207_ = ~new_n15892_;
  assign new_n16208_ = ~new_n2138_ | ~new_n15964_;
  assign new_n16209_ = ~new_n2132_ | ~new_n15842_;
  assign new_n16210_ = ~new_n15893_;
  assign new_n16211_ = ~new_n2138_ | ~new_n15965_;
  assign new_n16212_ = ~new_n2130_ | ~new_n15842_;
  assign new_n16213_ = ~new_n15887_;
  assign new_n16214_ = ~new_n2138_ | ~new_n15966_;
  assign new_n16215_ = ~new_n2131_ | ~new_n15842_;
  assign new_n16216_ = ~new_n15886_;
  assign new_n16217_ = ~new_n2138_ | ~new_n15967_;
  assign new_n16218_ = ~new_n2129_ | ~new_n15842_;
  assign new_n16219_ = ~new_n15894_;
  assign new_n16220_ = ~new_n15958_ | ~new_n15856_;
  assign new_n16221_ = ~new_n16192_ | ~new_n16054_;
  assign new_n16222_ = ~new_n16219_ | ~new_n2100_;
  assign new_n16223_ = ~new_n15894_ | ~new_n15854_;
  assign new_n16224_ = ~new_n16219_ | ~new_n2100_;
  assign new_n16225_ = ~new_n15894_ | ~new_n15854_;
  assign new_n16226_ = ~new_n16225_ | ~new_n16224_;
  assign new_n16227_ = ~new_n15968_ | ~new_n15969_;
  assign new_n16228_ = ~new_n16050_ | ~new_n16226_;
  assign new_n16229_ = ~new_n16213_ | ~new_n2101_;
  assign new_n16230_ = ~new_n15887_ | ~new_n15845_;
  assign new_n16231_ = ~new_n16216_ | ~new_n2102_;
  assign new_n16232_ = ~new_n15886_ | ~new_n15843_;
  assign new_n16233_ = ~new_n16232_ | ~new_n16231_;
  assign new_n16234_ = ~new_n16168_ | ~new_n15857_;
  assign new_n16235_ = ~new_n16233_ | ~new_n16042_;
  assign new_n16236_ = ~new_n16210_ | ~new_n2103_;
  assign new_n16237_ = ~new_n15893_ | ~new_n15853_;
  assign new_n16238_ = ~new_n16210_ | ~new_n2103_;
  assign new_n16239_ = ~new_n15893_ | ~new_n15853_;
  assign new_n16240_ = ~new_n16239_ | ~new_n16238_;
  assign new_n16241_ = ~new_n15970_ | ~new_n15971_;
  assign new_n16242_ = ~new_n16038_ | ~new_n16240_;
  assign new_n16243_ = ~new_n16207_ | ~new_n2104_;
  assign new_n16244_ = ~new_n15892_ | ~new_n15852_;
  assign new_n16245_ = ~new_n16207_ | ~new_n2104_;
  assign new_n16246_ = ~new_n15892_ | ~new_n15852_;
  assign new_n16247_ = ~new_n16246_ | ~new_n16245_;
  assign new_n16248_ = ~new_n15972_ | ~new_n15851_;
  assign new_n16249_ = ~new_n16247_ | ~new_n16034_;
  assign new_n16250_ = ~new_n16201_ | ~new_n2105_;
  assign new_n16251_ = ~new_n15889_ | ~new_n15848_;
  assign new_n16252_ = ~new_n16204_ | ~new_n2106_;
  assign new_n16253_ = ~new_n15888_ | ~new_n15846_;
  assign new_n16254_ = ~new_n16253_ | ~new_n16252_;
  assign new_n16255_ = ~new_n16169_ | ~new_n15858_;
  assign new_n16256_ = ~new_n16254_ | ~new_n16027_;
  assign new_n16257_ = ~new_n2138_ | ~new_n15973_;
  assign new_n16258_ = ~new_n2110_ | ~new_n15842_;
  assign new_n16259_ = ~new_n15895_;
  assign new_n16260_ = ~new_n2138_ | ~new_n15974_;
  assign new_n16261_ = ~new_n2112_ | ~new_n15842_;
  assign new_n16262_ = ~new_n15896_;
  assign new_n16263_ = ~new_n2138_ | ~new_n15975_;
  assign new_n16264_ = ~new_n2111_ | ~new_n15842_;
  assign new_n16265_ = ~new_n15897_;
  assign new_n16266_ = ~new_n2138_ | ~new_n15976_;
  assign new_n16267_ = ~new_n2113_ | ~new_n15842_;
  assign new_n16268_ = ~new_n15898_;
  assign new_n16269_ = ~new_n2138_ | ~new_n15977_;
  assign new_n16270_ = ~new_n2116_ | ~new_n15842_;
  assign new_n16271_ = ~new_n15899_;
  assign new_n16272_ = ~new_n2138_ | ~new_n15978_;
  assign new_n16273_ = ~new_n2117_ | ~new_n15842_;
  assign new_n16274_ = ~new_n15910_;
  assign new_n16275_ = ~new_n2138_ | ~new_n15979_;
  assign new_n16276_ = ~new_n2118_ | ~new_n15842_;
  assign new_n16277_ = ~new_n15909_;
  assign new_n16278_ = ~new_n2138_ | ~new_n15980_;
  assign new_n16279_ = ~new_n2127_ | ~new_n15842_;
  assign new_n16280_ = ~new_n15902_;
  assign new_n16281_ = ~new_n2138_ | ~new_n15981_;
  assign new_n16282_ = ~new_n2124_ | ~new_n15842_;
  assign new_n16283_ = ~new_n15904_;
  assign new_n16284_ = ~new_n2138_ | ~new_n15982_;
  assign new_n16285_ = ~new_n2125_ | ~new_n15842_;
  assign new_n16286_ = ~new_n15905_;
  assign new_n16287_ = ~new_n2138_ | ~new_n15983_;
  assign new_n16288_ = ~new_n2126_ | ~new_n15842_;
  assign new_n16289_ = ~new_n15903_;
  assign new_n16290_ = ~new_n2138_ | ~new_n15984_;
  assign new_n16291_ = ~new_n2123_ | ~new_n15842_;
  assign new_n16292_ = ~new_n15906_;
  assign new_n16293_ = ~new_n2138_ | ~new_n15985_;
  assign new_n16294_ = ~new_n2122_ | ~new_n15842_;
  assign new_n16295_ = ~new_n15907_;
  assign new_n16296_ = ~new_n2138_ | ~new_n15986_;
  assign new_n16297_ = ~new_n2120_ | ~new_n15842_;
  assign new_n16298_ = ~new_n15901_;
  assign new_n16299_ = ~new_n2138_ | ~new_n15987_;
  assign new_n16300_ = ~new_n2121_ | ~new_n15842_;
  assign new_n16301_ = ~new_n15900_;
  assign new_n16302_ = ~new_n2138_ | ~new_n15988_;
  assign new_n16303_ = ~new_n2119_ | ~new_n15842_;
  assign new_n16304_ = ~new_n15908_;
  assign new_n16305_ = ~new_n2138_ | ~new_n15989_;
  assign new_n16306_ = ~new_n2115_ | ~new_n15842_;
  assign new_n16307_ = ~new_n15911_;
  assign new_n16308_ = ~new_n2138_ | ~new_n15990_;
  assign new_n16309_ = ~new_n2114_ | ~new_n15842_;
  assign new_n16310_ = ~new_n15912_;
  assign new_n16311_ = ~new_n2138_ | ~new_n15991_;
  assign new_n16312_ = ~new_n2080_ | ~new_n15842_;
  assign new_n16313_ = ~new_n15949_;
  assign new_n16314_ = ~new_n2109_ | ~new_n16313_;
  assign new_n16315_ = ~new_n15949_ | ~new_n15992_;
  assign new_n16316_ = ~new_n15913_;
  assign new_n16317_ = ~new_n16316_ | ~new_n16177_ | ~new_n16131_;
  assign new_n16318_ = ~new_n16182_ | ~new_n15913_ | ~new_n15948_ | ~new_n16183_;
  assign new_n16319_ = ~new_n16259_ | ~new_n2081_;
  assign new_n16320_ = ~new_n15895_ | ~new_n15859_;
  assign new_n16321_ = ~new_n16259_ | ~new_n2081_;
  assign new_n16322_ = ~new_n15895_ | ~new_n15859_;
  assign new_n16323_ = ~new_n16322_ | ~new_n16321_;
  assign new_n16324_ = ~new_n15993_ | ~new_n15994_;
  assign new_n16325_ = ~new_n16130_ | ~new_n16323_;
  assign new_n16326_ = ~new_n16265_ | ~new_n2082_;
  assign new_n16327_ = ~new_n15897_ | ~new_n15860_;
  assign new_n16328_ = ~new_n16262_ | ~new_n2083_;
  assign new_n16329_ = ~new_n15896_ | ~new_n15861_;
  assign new_n16330_ = ~new_n16329_ | ~new_n16328_;
  assign new_n16331_ = ~new_n16170_ | ~new_n15881_;
  assign new_n16332_ = ~new_n16330_ | ~new_n16135_;
  assign new_n16333_ = ~new_n16268_ | ~new_n2084_;
  assign new_n16334_ = ~new_n15898_ | ~new_n15862_;
  assign new_n16335_ = ~new_n16334_ | ~new_n16333_;
  assign new_n16336_ = ~new_n16171_ | ~new_n15995_;
  assign new_n16337_ = ~new_n16124_ | ~new_n16335_;
  assign new_n16338_ = ~new_n16310_ | ~new_n2085_;
  assign new_n16339_ = ~new_n15912_ | ~new_n15879_;
  assign new_n16340_ = ~new_n16310_ | ~new_n2085_;
  assign new_n16341_ = ~new_n15912_ | ~new_n15879_;
  assign new_n16342_ = ~new_n16341_ | ~new_n16340_;
  assign new_n16343_ = ~new_n15996_ | ~new_n15997_;
  assign new_n16344_ = ~new_n16120_ | ~new_n16342_;
  assign new_n16345_ = ~new_n16307_ | ~new_n2086_;
  assign new_n16346_ = ~new_n15911_ | ~new_n15878_;
  assign new_n16347_ = ~new_n16307_ | ~new_n2086_;
  assign new_n16348_ = ~new_n15911_ | ~new_n15878_;
  assign new_n16349_ = ~new_n16348_ | ~new_n16347_;
  assign new_n16350_ = ~new_n15998_ | ~new_n15999_;
  assign new_n16351_ = ~new_n16116_ | ~new_n16349_;
  assign new_n16352_ = ~new_n16271_ | ~new_n2087_;
  assign new_n16353_ = ~new_n15899_ | ~new_n15863_;
  assign new_n16354_ = ~new_n16274_ | ~new_n2088_;
  assign new_n16355_ = ~new_n15910_ | ~new_n15877_;
  assign new_n16356_ = ~new_n16355_ | ~new_n16354_;
  assign new_n16357_ = ~new_n16172_ | ~new_n15882_;
  assign new_n16358_ = ~new_n16356_ | ~new_n16144_;
  assign new_n16359_ = ~new_n16198_ | ~new_n2107_;
  assign new_n16360_ = ~new_n15891_ | ~new_n15850_;
  assign new_n16361_ = ~new_n16198_ | ~new_n2107_;
  assign new_n16362_ = ~new_n15891_ | ~new_n15850_;
  assign new_n16363_ = ~new_n16362_ | ~new_n16361_;
  assign new_n16364_ = ~new_n16000_ | ~new_n16001_;
  assign new_n16365_ = ~new_n16023_ | ~new_n16363_;
  assign new_n16366_ = ~new_n16277_ | ~new_n2089_;
  assign new_n16367_ = ~new_n15909_ | ~new_n15875_;
  assign new_n16368_ = ~new_n16367_ | ~new_n16366_;
  assign new_n16369_ = ~new_n16173_ | ~new_n16002_;
  assign new_n16370_ = ~new_n16106_ | ~new_n16368_;
  assign new_n16371_ = ~new_n16304_ | ~new_n2090_;
  assign new_n16372_ = ~new_n15908_ | ~new_n15874_;
  assign new_n16373_ = ~new_n16304_ | ~new_n2090_;
  assign new_n16374_ = ~new_n15908_ | ~new_n15874_;
  assign new_n16375_ = ~new_n16374_ | ~new_n16373_;
  assign new_n16376_ = ~new_n16003_ | ~new_n16004_;
  assign new_n16377_ = ~new_n16102_ | ~new_n16375_;
  assign new_n16378_ = ~new_n16298_ | ~new_n2091_;
  assign new_n16379_ = ~new_n15901_ | ~new_n15866_;
  assign new_n16380_ = ~new_n16301_ | ~new_n2092_;
  assign new_n16381_ = ~new_n15900_ | ~new_n15864_;
  assign new_n16382_ = ~new_n16381_ | ~new_n16380_;
  assign new_n16383_ = ~new_n16174_ | ~new_n15883_;
  assign new_n16384_ = ~new_n16382_ | ~new_n16094_;
  assign new_n16385_ = ~new_n16295_ | ~new_n2093_;
  assign new_n16386_ = ~new_n15907_ | ~new_n15873_;
  assign new_n16387_ = ~new_n16295_ | ~new_n2093_;
  assign new_n16388_ = ~new_n15907_ | ~new_n15873_;
  assign new_n16389_ = ~new_n16388_ | ~new_n16387_;
  assign new_n16390_ = ~new_n16005_ | ~new_n16006_;
  assign new_n16391_ = ~new_n16090_ | ~new_n16389_;
  assign new_n16392_ = ~new_n16292_ | ~new_n2094_;
  assign new_n16393_ = ~new_n15906_ | ~new_n15872_;
  assign new_n16394_ = ~new_n16292_ | ~new_n2094_;
  assign new_n16395_ = ~new_n15906_ | ~new_n15872_;
  assign new_n16396_ = ~new_n16395_ | ~new_n16394_;
  assign new_n16397_ = ~new_n16007_ | ~new_n16008_;
  assign new_n16398_ = ~new_n16086_ | ~new_n16396_;
  assign new_n16399_ = ~new_n16283_ | ~new_n2095_;
  assign new_n16400_ = ~new_n15904_ | ~new_n15871_;
  assign new_n16401_ = ~new_n16286_ | ~new_n2096_;
  assign new_n16402_ = ~new_n15905_ | ~new_n15868_;
  assign new_n16403_ = ~new_n16402_ | ~new_n16401_;
  assign new_n16404_ = ~new_n16175_ | ~new_n15884_;
  assign new_n16405_ = ~new_n16403_ | ~new_n16160_;
  assign new_n16406_ = ~new_n16289_ | ~new_n2097_;
  assign new_n16407_ = ~new_n15903_ | ~new_n15869_;
  assign new_n16408_ = ~new_n16407_ | ~new_n16406_;
  assign new_n16409_ = ~new_n16176_ | ~new_n16009_;
  assign new_n16410_ = ~new_n16076_ | ~new_n16408_;
  assign new_n16411_ = ~new_n16280_ | ~new_n2098_;
  assign new_n16412_ = ~new_n15902_ | ~new_n15867_;
  assign new_n16413_ = ~new_n16280_ | ~new_n2098_;
  assign new_n16414_ = ~new_n15902_ | ~new_n15867_;
  assign new_n16415_ = ~new_n16414_ | ~new_n16413_;
  assign new_n16416_ = ~new_n16010_ | ~new_n16011_;
  assign new_n16417_ = ~new_n16072_ | ~new_n16415_;
  assign new_n16418_ = ~new_n2108_ | ~new_n15842_;
  assign new_n16419_ = ~new_n2138_ | ~new_n15849_;
  assign new_n16420_ = ~new_n15956_;
  assign new_n16421_ = ~new_n15890_ | ~new_n16420_;
  assign new_n16422_ = ~new_n15956_ | ~new_n16195_;
  assign new_n16423_ = new_n16601_ & new_n16618_;
  assign new_n16424_ = new_n16620_ & new_n16619_;
  assign new_n16425_ = new_n16596_ & new_n16657_;
  assign new_n16426_ = new_n16659_ & new_n16658_;
  assign new_n16427_ = new_n16676_ & new_n16675_;
  assign new_n16428_ = new_n16702_ & new_n16701_;
  assign new_n16429_ = new_n16800_ & new_n16799_;
  assign new_n16430_ = ~new_n16757_ | ~new_n16760_;
  assign new_n16431_ = ~new_n16746_ | ~new_n16749_;
  assign new_n16432_ = ~new_n16735_ | ~new_n16738_;
  assign new_n16433_ = ~new_n16727_ | ~new_n16729_;
  assign new_n16434_ = ~new_n16765_ | ~new_n16573_ | ~new_n16592_;
  assign new_n16435_ = ~new_n16653_ | ~new_n16655_;
  assign new_n16436_ = ~new_n16645_ | ~new_n16648_;
  assign new_n16437_ = ~new_n16637_ | ~new_n16639_;
  assign new_n16438_ = ~new_n16442_ | ~new_n16763_;
  assign new_n16439_ = ~new_n2406_;
  assign new_n16440_ = ~new_n2391_;
  assign new_n16441_ = ~new_n2383_;
  assign new_n16442_ = ~new_n2383_ | ~new_n16510_;
  assign new_n16443_ = ~new_n2005_;
  assign new_n16444_ = ~new_n2394_;
  assign new_n16445_ = ~new_n1995_;
  assign new_n16446_ = ~new_n1995_ | ~new_n16440_;
  assign new_n16447_ = ~new_n1991_;
  assign new_n16448_ = ~new_n2403_;
  assign new_n16449_ = ~new_n2400_;
  assign new_n16450_ = ~new_n2397_;
  assign new_n16451_ = ~new_n1998_;
  assign new_n16452_ = ~new_n1994_;
  assign new_n16453_ = ~new_n1987_;
  assign new_n16454_ = ~new_n1987_ | ~new_n16450_;
  assign new_n16455_ = ~new_n2409_;
  assign new_n16456_ = ~new_n1997_;
  assign new_n16457_ = ~new_n1997_ | ~new_n16439_;
  assign new_n16458_ = ~new_n2011_;
  assign new_n16459_ = ~new_n2412_;
  assign new_n16460_ = ~new_n2010_;
  assign new_n16461_ = ~new_n16626_ | ~new_n16625_;
  assign new_n16462_ = ~new_n16454_ | ~new_n16641_;
  assign new_n16463_ = ~new_n16610_ | ~new_n16609_;
  assign new_n16464_ = ~new_n2946_;
  assign new_n16465_ = ~new_n2950_;
  assign new_n16466_ = ~new_n2430_;
  assign new_n16467_ = ~new_n2418_;
  assign new_n16468_ = ~new_n2415_;
  assign new_n16469_ = ~new_n1990_;
  assign new_n16470_ = ~new_n1989_;
  assign new_n16471_ = ~new_n2010_ | ~new_n16459_;
  assign new_n16472_ = ~new_n2421_;
  assign new_n16473_ = ~new_n1999_;
  assign new_n16474_ = ~new_n2424_;
  assign new_n16475_ = ~new_n2007_;
  assign new_n16476_ = ~new_n2433_;
  assign new_n16477_ = ~new_n2427_;
  assign new_n16478_ = ~new_n2000_;
  assign new_n16479_ = ~new_n2001_;
  assign new_n16480_ = ~new_n2006_;
  assign new_n16481_ = ~new_n2006_ | ~new_n16477_;
  assign new_n16482_ = ~new_n2436_;
  assign new_n16483_ = ~new_n1996_;
  assign new_n16484_ = ~new_n16686_ | ~new_n16685_;
  assign new_n16485_ = ~new_n2009_;
  assign new_n16486_ = ~new_n2441_;
  assign new_n16487_ = ~new_n2008_;
  assign new_n16488_ = ~new_n2952_;
  assign new_n16489_ = ~new_n2003_;
  assign new_n16490_ = ~new_n2949_;
  assign new_n16491_ = ~new_n2951_;
  assign new_n16492_ = ~new_n1993_;
  assign new_n16493_ = ~new_n1988_;
  assign new_n16494_ = ~new_n2002_;
  assign new_n16495_ = ~new_n2002_ | ~new_n16491_;
  assign new_n16496_ = ~new_n2948_;
  assign new_n16497_ = ~new_n1992_;
  assign new_n16498_ = ~new_n2947_;
  assign new_n16499_ = ~new_n1985_;
  assign new_n16500_ = ~new_n2945_;
  assign new_n16501_ = ~new_n1984_;
  assign new_n16502_ = ~new_n1984_ | ~new_n16464_;
  assign new_n16503_ = ~new_n1980_;
  assign new_n16504_ = ~new_n2944_;
  assign new_n16505_ = ~new_n1981_;
  assign new_n16506_ = ~new_n16716_ | ~new_n16715_;
  assign new_n16507_ = ~new_n16495_ | ~new_n16731_;
  assign new_n16508_ = ~new_n16481_ | ~new_n16742_;
  assign new_n16509_ = ~new_n16471_ | ~new_n16753_;
  assign new_n16510_ = ~new_n2004_;
  assign new_n16511_ = ~new_n16810_ | ~new_n16809_;
  assign new_n16512_ = ~new_n16824_ | ~new_n16823_;
  assign new_n16513_ = ~new_n16829_ | ~new_n16828_;
  assign new_n16514_ = ~new_n16845_ | ~new_n16844_;
  assign new_n16515_ = ~new_n16850_ | ~new_n16849_;
  assign new_n16516_ = ~new_n16855_ | ~new_n16854_;
  assign new_n16517_ = ~new_n16860_ | ~new_n16859_;
  assign new_n16518_ = ~new_n16865_ | ~new_n16864_;
  assign new_n16519_ = ~new_n16881_ | ~new_n16880_;
  assign new_n16520_ = ~new_n16886_ | ~new_n16885_;
  assign new_n16521_ = ~new_n16769_ | ~new_n16768_;
  assign new_n16522_ = ~new_n16778_ | ~new_n16777_;
  assign new_n16523_ = ~new_n16785_ | ~new_n16784_;
  assign new_n16524_ = ~new_n16789_ | ~new_n16788_;
  assign new_n16525_ = ~new_n16798_ | ~new_n16797_;
  assign new_n16526_ = ~new_n16819_ | ~new_n16818_;
  assign new_n16527_ = ~new_n16836_ | ~new_n16835_;
  assign new_n16528_ = ~new_n16840_ | ~new_n16839_;
  assign new_n16529_ = ~new_n16872_ | ~new_n16871_;
  assign new_n16530_ = ~new_n16876_ | ~new_n16875_;
  assign new_n16531_ = ~new_n16893_ | ~new_n16892_;
  assign new_n16532_ = new_n16612_ & new_n16600_;
  assign new_n16533_ = new_n16615_ & new_n16616_;
  assign new_n16534_ = new_n16628_ & new_n16602_;
  assign new_n16535_ = new_n16631_ & new_n16632_;
  assign new_n16536_ = new_n16457_ & new_n16771_ & new_n16770_;
  assign new_n16537_ = new_n16774_ & new_n16602_;
  assign new_n16538_ = new_n16647_ & new_n16424_;
  assign new_n16539_ = new_n16781_ & new_n16601_;
  assign new_n16540_ = new_n16446_ & new_n16791_ & new_n16790_;
  assign new_n16541_ = new_n16794_ & new_n16600_;
  assign new_n16542_ = new_n16634_ & new_n16425_;
  assign new_n16543_ = new_n16679_ & new_n16597_;
  assign new_n16544_ = new_n16705_ & new_n16598_;
  assign new_n16545_ = new_n16721_ & new_n16722_;
  assign new_n16546_ = new_n16724_ & new_n16803_;
  assign new_n16547_ = new_n16725_ & new_n16722_ & new_n16721_;
  assign new_n16548_ = ~new_n16807_ | ~new_n16806_;
  assign new_n16549_ = new_n16502_ & new_n16812_ & new_n16811_;
  assign new_n16550_ = new_n16815_ & new_n16599_;
  assign new_n16551_ = ~new_n16821_ | ~new_n16820_;
  assign new_n16552_ = ~new_n16826_ | ~new_n16825_;
  assign new_n16553_ = new_n16832_ & new_n16598_;
  assign new_n16554_ = ~new_n16842_ | ~new_n16841_;
  assign new_n16555_ = ~new_n16847_ | ~new_n16846_;
  assign new_n16556_ = ~new_n16852_ | ~new_n16851_;
  assign new_n16557_ = ~new_n16857_ | ~new_n16856_;
  assign new_n16558_ = ~new_n16862_ | ~new_n16861_;
  assign new_n16559_ = new_n16868_ & new_n16597_;
  assign new_n16560_ = ~new_n16878_ | ~new_n16877_;
  assign new_n16561_ = ~new_n16883_ | ~new_n16882_;
  assign new_n16562_ = new_n16759_ & new_n16426_;
  assign new_n16563_ = new_n16889_ & new_n16596_;
  assign new_n16564_ = new_n16767_ & new_n16766_;
  assign new_n16565_ = ~new_n16535_ | ~new_n16629_;
  assign new_n16566_ = new_n16776_ & new_n16775_;
  assign new_n16567_ = new_n16783_ & new_n16782_;
  assign new_n16568_ = new_n16787_ & new_n16786_;
  assign new_n16569_ = ~new_n16533_ | ~new_n16613_;
  assign new_n16570_ = new_n16796_ & new_n16795_;
  assign new_n16571_ = ~new_n2955_;
  assign new_n16572_ = ~new_n1982_;
  assign new_n16573_ = new_n16805_ & new_n16804_;
  assign new_n16574_ = ~new_n16545_ | ~new_n16719_;
  assign new_n16575_ = new_n16817_ & new_n16816_;
  assign new_n16576_ = ~new_n16712_ | ~new_n16711_;
  assign new_n16577_ = ~new_n16708_ | ~new_n16707_;
  assign new_n16578_ = new_n16834_ & new_n16833_;
  assign new_n16579_ = new_n16838_ & new_n16837_;
  assign new_n16580_ = ~new_n16698_ | ~new_n16697_;
  assign new_n16581_ = ~new_n16694_ | ~new_n16693_;
  assign new_n16582_ = ~new_n2388_;
  assign new_n16583_ = ~new_n16690_ | ~new_n16689_;
  assign new_n16584_ = ~new_n2439_;
  assign new_n16585_ = ~new_n16682_ | ~new_n16681_;
  assign new_n16586_ = new_n16870_ & new_n16869_;
  assign new_n16587_ = new_n16874_ & new_n16873_;
  assign new_n16588_ = ~new_n16672_ | ~new_n16671_;
  assign new_n16589_ = ~new_n16668_ | ~new_n16667_;
  assign new_n16590_ = ~new_n16664_ | ~new_n16663_;
  assign new_n16591_ = new_n16891_ & new_n16890_;
  assign new_n16592_ = ~new_n16546_ | ~new_n16574_;
  assign new_n16593_ = ~new_n16502_;
  assign new_n16594_ = ~new_n16446_;
  assign new_n16595_ = ~new_n16457_;
  assign new_n16596_ = ~new_n2415_ | ~new_n16470_;
  assign new_n16597_ = ~new_n2430_ | ~new_n16479_;
  assign new_n16598_ = ~new_n2950_ | ~new_n16493_;
  assign new_n16599_ = ~new_n2946_ | ~new_n16501_;
  assign new_n16600_ = ~new_n2391_ | ~new_n16445_;
  assign new_n16601_ = ~new_n2400_ | ~new_n16452_;
  assign new_n16602_ = ~new_n2406_ | ~new_n16456_;
  assign new_n16603_ = ~new_n16481_;
  assign new_n16604_ = ~new_n16495_;
  assign new_n16605_ = ~new_n16454_;
  assign new_n16606_ = ~new_n16471_;
  assign new_n16607_ = ~new_n16442_;
  assign new_n16608_ = ~new_n16607_ | ~new_n16443_;
  assign new_n16609_ = ~new_n16608_ | ~new_n16582_;
  assign new_n16610_ = ~new_n2005_ | ~new_n16442_;
  assign new_n16611_ = ~new_n16463_;
  assign new_n16612_ = ~new_n2394_ | ~new_n16447_;
  assign new_n16613_ = ~new_n16532_ | ~new_n16463_;
  assign new_n16614_ = ~new_n16447_ | ~new_n16446_;
  assign new_n16615_ = ~new_n16614_ | ~new_n16444_;
  assign new_n16616_ = ~new_n1991_ | ~new_n16594_;
  assign new_n16617_ = ~new_n16569_;
  assign new_n16618_ = ~new_n2403_ | ~new_n16451_;
  assign new_n16619_ = ~new_n1998_ | ~new_n16448_;
  assign new_n16620_ = ~new_n1994_ | ~new_n16449_;
  assign new_n16621_ = ~new_n16605_ | ~new_n16423_;
  assign new_n16622_ = ~new_n16424_ | ~new_n16621_;
  assign new_n16623_ = ~new_n2397_ | ~new_n16453_;
  assign new_n16624_ = ~new_n2403_ | ~new_n16451_;
  assign new_n16625_ = ~new_n16423_ | ~new_n16623_ | ~new_n16569_;
  assign new_n16626_ = ~new_n16624_ | ~new_n16622_;
  assign new_n16627_ = ~new_n16461_;
  assign new_n16628_ = ~new_n2409_ | ~new_n16458_;
  assign new_n16629_ = ~new_n16534_ | ~new_n16461_;
  assign new_n16630_ = ~new_n16458_ | ~new_n16457_;
  assign new_n16631_ = ~new_n16630_ | ~new_n16455_;
  assign new_n16632_ = ~new_n2011_ | ~new_n16595_;
  assign new_n16633_ = ~new_n16565_;
  assign new_n16634_ = ~new_n2412_ | ~new_n16460_;
  assign new_n16635_ = ~new_n16634_ | ~new_n16471_;
  assign new_n16636_ = ~new_n16627_ | ~new_n16457_;
  assign new_n16637_ = ~new_n16537_ | ~new_n16636_;
  assign new_n16638_ = ~new_n16461_ | ~new_n16602_;
  assign new_n16639_ = ~new_n16536_ | ~new_n16638_;
  assign new_n16640_ = ~new_n16457_ | ~new_n16602_;
  assign new_n16641_ = ~new_n16623_ | ~new_n16569_;
  assign new_n16642_ = ~new_n16462_;
  assign new_n16643_ = ~new_n1994_ | ~new_n16449_;
  assign new_n16644_ = ~new_n16642_ | ~new_n16643_;
  assign new_n16645_ = ~new_n16539_ | ~new_n16644_;
  assign new_n16646_ = ~new_n16462_ | ~new_n16601_;
  assign new_n16647_ = ~new_n2403_ | ~new_n16451_;
  assign new_n16648_ = ~new_n16538_ | ~new_n16646_;
  assign new_n16649_ = ~new_n1994_ | ~new_n16449_;
  assign new_n16650_ = ~new_n16601_ | ~new_n16649_;
  assign new_n16651_ = ~new_n16623_ | ~new_n16454_;
  assign new_n16652_ = ~new_n16611_ | ~new_n16446_;
  assign new_n16653_ = ~new_n16541_ | ~new_n16652_;
  assign new_n16654_ = ~new_n16463_ | ~new_n16600_;
  assign new_n16655_ = ~new_n16540_ | ~new_n16654_;
  assign new_n16656_ = ~new_n16446_ | ~new_n16600_;
  assign new_n16657_ = ~new_n2418_ | ~new_n16469_;
  assign new_n16658_ = ~new_n1990_ | ~new_n16467_;
  assign new_n16659_ = ~new_n1989_ | ~new_n16468_;
  assign new_n16660_ = ~new_n16606_ | ~new_n16425_;
  assign new_n16661_ = ~new_n16426_ | ~new_n16660_;
  assign new_n16662_ = ~new_n2418_ | ~new_n16469_;
  assign new_n16663_ = ~new_n16542_ | ~new_n16565_;
  assign new_n16664_ = ~new_n16662_ | ~new_n16661_;
  assign new_n16665_ = ~new_n16590_;
  assign new_n16666_ = ~new_n2421_ | ~new_n16473_;
  assign new_n16667_ = ~new_n16666_ | ~new_n16590_;
  assign new_n16668_ = ~new_n1999_ | ~new_n16472_;
  assign new_n16669_ = ~new_n16589_;
  assign new_n16670_ = ~new_n2424_ | ~new_n16475_;
  assign new_n16671_ = ~new_n16670_ | ~new_n16589_;
  assign new_n16672_ = ~new_n2007_ | ~new_n16474_;
  assign new_n16673_ = ~new_n16588_;
  assign new_n16674_ = ~new_n2433_ | ~new_n16478_;
  assign new_n16675_ = ~new_n2000_ | ~new_n16476_;
  assign new_n16676_ = ~new_n2001_ | ~new_n16466_;
  assign new_n16677_ = ~new_n16603_ | ~new_n16597_;
  assign new_n16678_ = ~new_n16427_ | ~new_n16677_;
  assign new_n16679_ = ~new_n2427_ | ~new_n16480_;
  assign new_n16680_ = ~new_n2433_ | ~new_n16478_;
  assign new_n16681_ = ~new_n16674_ | ~new_n16588_ | ~new_n16543_;
  assign new_n16682_ = ~new_n16680_ | ~new_n16678_;
  assign new_n16683_ = ~new_n16585_;
  assign new_n16684_ = ~new_n2436_ | ~new_n16483_;
  assign new_n16685_ = ~new_n16684_ | ~new_n16585_;
  assign new_n16686_ = ~new_n1996_ | ~new_n16482_;
  assign new_n16687_ = ~new_n16484_;
  assign new_n16688_ = ~new_n16687_ | ~new_n16485_;
  assign new_n16689_ = ~new_n16688_ | ~new_n16584_;
  assign new_n16690_ = ~new_n2009_ | ~new_n16484_;
  assign new_n16691_ = ~new_n16583_;
  assign new_n16692_ = ~new_n2441_ | ~new_n16487_;
  assign new_n16693_ = ~new_n16692_ | ~new_n16583_;
  assign new_n16694_ = ~new_n2008_ | ~new_n16486_;
  assign new_n16695_ = ~new_n16581_;
  assign new_n16696_ = ~new_n2952_ | ~new_n16489_;
  assign new_n16697_ = ~new_n16696_ | ~new_n16581_;
  assign new_n16698_ = ~new_n2003_ | ~new_n16488_;
  assign new_n16699_ = ~new_n16580_;
  assign new_n16700_ = ~new_n2949_ | ~new_n16492_;
  assign new_n16701_ = ~new_n1993_ | ~new_n16490_;
  assign new_n16702_ = ~new_n1988_ | ~new_n16465_;
  assign new_n16703_ = ~new_n16604_ | ~new_n16598_;
  assign new_n16704_ = ~new_n16428_ | ~new_n16703_;
  assign new_n16705_ = ~new_n2951_ | ~new_n16494_;
  assign new_n16706_ = ~new_n2949_ | ~new_n16492_;
  assign new_n16707_ = ~new_n16700_ | ~new_n16580_ | ~new_n16544_;
  assign new_n16708_ = ~new_n16706_ | ~new_n16704_;
  assign new_n16709_ = ~new_n16577_;
  assign new_n16710_ = ~new_n2948_ | ~new_n16497_;
  assign new_n16711_ = ~new_n16710_ | ~new_n16577_;
  assign new_n16712_ = ~new_n1992_ | ~new_n16496_;
  assign new_n16713_ = ~new_n16576_;
  assign new_n16714_ = ~new_n2947_ | ~new_n16499_;
  assign new_n16715_ = ~new_n16714_ | ~new_n16576_;
  assign new_n16716_ = ~new_n1985_ | ~new_n16498_;
  assign new_n16717_ = ~new_n16506_;
  assign new_n16718_ = ~new_n2945_ | ~new_n16503_;
  assign new_n16719_ = ~new_n16718_ | ~new_n16506_ | ~new_n16599_;
  assign new_n16720_ = ~new_n16503_ | ~new_n16502_;
  assign new_n16721_ = ~new_n16720_ | ~new_n16500_;
  assign new_n16722_ = ~new_n1980_ | ~new_n16593_;
  assign new_n16723_ = ~new_n16574_;
  assign new_n16724_ = ~new_n2944_ | ~new_n16505_;
  assign new_n16725_ = ~new_n1981_ | ~new_n16504_;
  assign new_n16726_ = ~new_n16717_ | ~new_n16502_;
  assign new_n16727_ = ~new_n16550_ | ~new_n16726_;
  assign new_n16728_ = ~new_n16506_ | ~new_n16599_;
  assign new_n16729_ = ~new_n16549_ | ~new_n16728_;
  assign new_n16730_ = ~new_n16502_ | ~new_n16599_;
  assign new_n16731_ = ~new_n16705_ | ~new_n16580_;
  assign new_n16732_ = ~new_n16507_;
  assign new_n16733_ = ~new_n1988_ | ~new_n16465_;
  assign new_n16734_ = ~new_n16732_ | ~new_n16733_;
  assign new_n16735_ = ~new_n16553_ | ~new_n16734_;
  assign new_n16736_ = ~new_n16507_ | ~new_n16598_;
  assign new_n16737_ = ~new_n2949_ | ~new_n16492_;
  assign new_n16738_ = ~new_n16428_ | ~new_n16737_ | ~new_n16736_;
  assign new_n16739_ = ~new_n1988_ | ~new_n16465_;
  assign new_n16740_ = ~new_n16598_ | ~new_n16739_;
  assign new_n16741_ = ~new_n16705_ | ~new_n16495_;
  assign new_n16742_ = ~new_n16679_ | ~new_n16588_;
  assign new_n16743_ = ~new_n16508_;
  assign new_n16744_ = ~new_n2001_ | ~new_n16466_;
  assign new_n16745_ = ~new_n16743_ | ~new_n16744_;
  assign new_n16746_ = ~new_n16559_ | ~new_n16745_;
  assign new_n16747_ = ~new_n16508_ | ~new_n16597_;
  assign new_n16748_ = ~new_n2433_ | ~new_n16478_;
  assign new_n16749_ = ~new_n16427_ | ~new_n16748_ | ~new_n16747_;
  assign new_n16750_ = ~new_n2001_ | ~new_n16466_;
  assign new_n16751_ = ~new_n16597_ | ~new_n16750_;
  assign new_n16752_ = ~new_n16679_ | ~new_n16481_;
  assign new_n16753_ = ~new_n16634_ | ~new_n16565_;
  assign new_n16754_ = ~new_n16509_;
  assign new_n16755_ = ~new_n1989_ | ~new_n16468_;
  assign new_n16756_ = ~new_n16754_ | ~new_n16755_;
  assign new_n16757_ = ~new_n16563_ | ~new_n16756_;
  assign new_n16758_ = ~new_n16509_ | ~new_n16596_;
  assign new_n16759_ = ~new_n2418_ | ~new_n16469_;
  assign new_n16760_ = ~new_n16562_ | ~new_n16758_;
  assign new_n16761_ = ~new_n1989_ | ~new_n16468_;
  assign new_n16762_ = ~new_n16596_ | ~new_n16761_;
  assign new_n16763_ = ~new_n2004_ | ~new_n16441_;
  assign new_n16764_ = ~new_n16718_ | ~new_n16506_ | ~new_n16599_;
  assign new_n16765_ = ~new_n16547_ | ~new_n16429_ | ~new_n16764_;
  assign new_n16766_ = ~new_n2412_ | ~new_n16460_;
  assign new_n16767_ = ~new_n2010_ | ~new_n16459_;
  assign new_n16768_ = ~new_n16635_ | ~new_n16565_;
  assign new_n16769_ = ~new_n16633_ | ~new_n16564_;
  assign new_n16770_ = ~new_n2409_ | ~new_n16458_;
  assign new_n16771_ = ~new_n2011_ | ~new_n16455_;
  assign new_n16772_ = ~new_n2409_ | ~new_n16458_;
  assign new_n16773_ = ~new_n2011_ | ~new_n16455_;
  assign new_n16774_ = ~new_n16773_ | ~new_n16772_;
  assign new_n16775_ = ~new_n2406_ | ~new_n16456_;
  assign new_n16776_ = ~new_n1997_ | ~new_n16439_;
  assign new_n16777_ = ~new_n16640_ | ~new_n16461_;
  assign new_n16778_ = ~new_n16566_ | ~new_n16627_;
  assign new_n16779_ = ~new_n2403_ | ~new_n16451_;
  assign new_n16780_ = ~new_n1998_ | ~new_n16448_;
  assign new_n16781_ = ~new_n16780_ | ~new_n16779_;
  assign new_n16782_ = ~new_n2400_ | ~new_n16452_;
  assign new_n16783_ = ~new_n1994_ | ~new_n16449_;
  assign new_n16784_ = ~new_n16650_ | ~new_n16462_;
  assign new_n16785_ = ~new_n16567_ | ~new_n16642_;
  assign new_n16786_ = ~new_n2397_ | ~new_n16453_;
  assign new_n16787_ = ~new_n1987_ | ~new_n16450_;
  assign new_n16788_ = ~new_n16651_ | ~new_n16569_;
  assign new_n16789_ = ~new_n16617_ | ~new_n16568_;
  assign new_n16790_ = ~new_n2394_ | ~new_n16447_;
  assign new_n16791_ = ~new_n1991_ | ~new_n16444_;
  assign new_n16792_ = ~new_n2394_ | ~new_n16447_;
  assign new_n16793_ = ~new_n1991_ | ~new_n16444_;
  assign new_n16794_ = ~new_n16793_ | ~new_n16792_;
  assign new_n16795_ = ~new_n2391_ | ~new_n16445_;
  assign new_n16796_ = ~new_n1995_ | ~new_n16440_;
  assign new_n16797_ = ~new_n16656_ | ~new_n16463_;
  assign new_n16798_ = ~new_n16570_ | ~new_n16611_;
  assign new_n16799_ = ~new_n2955_ | ~new_n16572_;
  assign new_n16800_ = ~new_n1982_ | ~new_n16571_;
  assign new_n16801_ = ~new_n2955_ | ~new_n16572_;
  assign new_n16802_ = ~new_n1982_ | ~new_n16571_;
  assign new_n16803_ = ~new_n16802_ | ~new_n16801_;
  assign new_n16804_ = ~new_n16504_ | ~new_n1981_ | ~new_n16803_;
  assign new_n16805_ = ~new_n2944_ | ~new_n16429_ | ~new_n16505_;
  assign new_n16806_ = ~new_n2944_ | ~new_n16505_;
  assign new_n16807_ = ~new_n1981_ | ~new_n16504_;
  assign new_n16808_ = ~new_n16548_;
  assign new_n16809_ = ~new_n16723_ | ~new_n16808_;
  assign new_n16810_ = ~new_n16548_ | ~new_n16574_;
  assign new_n16811_ = ~new_n2945_ | ~new_n16503_;
  assign new_n16812_ = ~new_n1980_ | ~new_n16500_;
  assign new_n16813_ = ~new_n2945_ | ~new_n16503_;
  assign new_n16814_ = ~new_n1980_ | ~new_n16500_;
  assign new_n16815_ = ~new_n16814_ | ~new_n16813_;
  assign new_n16816_ = ~new_n2946_ | ~new_n16501_;
  assign new_n16817_ = ~new_n1984_ | ~new_n16464_;
  assign new_n16818_ = ~new_n16730_ | ~new_n16506_;
  assign new_n16819_ = ~new_n16575_ | ~new_n16717_;
  assign new_n16820_ = ~new_n2947_ | ~new_n16499_;
  assign new_n16821_ = ~new_n1985_ | ~new_n16498_;
  assign new_n16822_ = ~new_n16551_;
  assign new_n16823_ = ~new_n16713_ | ~new_n16822_;
  assign new_n16824_ = ~new_n16551_ | ~new_n16576_;
  assign new_n16825_ = ~new_n2948_ | ~new_n16497_;
  assign new_n16826_ = ~new_n1992_ | ~new_n16496_;
  assign new_n16827_ = ~new_n16552_;
  assign new_n16828_ = ~new_n16709_ | ~new_n16827_;
  assign new_n16829_ = ~new_n16552_ | ~new_n16577_;
  assign new_n16830_ = ~new_n2949_ | ~new_n16492_;
  assign new_n16831_ = ~new_n1993_ | ~new_n16490_;
  assign new_n16832_ = ~new_n16831_ | ~new_n16830_;
  assign new_n16833_ = ~new_n2950_ | ~new_n16493_;
  assign new_n16834_ = ~new_n1988_ | ~new_n16465_;
  assign new_n16835_ = ~new_n16740_ | ~new_n16507_;
  assign new_n16836_ = ~new_n16578_ | ~new_n16732_;
  assign new_n16837_ = ~new_n2951_ | ~new_n16494_;
  assign new_n16838_ = ~new_n2002_ | ~new_n16491_;
  assign new_n16839_ = ~new_n16741_ | ~new_n16580_;
  assign new_n16840_ = ~new_n16699_ | ~new_n16579_;
  assign new_n16841_ = ~new_n2952_ | ~new_n16489_;
  assign new_n16842_ = ~new_n2003_ | ~new_n16488_;
  assign new_n16843_ = ~new_n16554_;
  assign new_n16844_ = ~new_n16695_ | ~new_n16843_;
  assign new_n16845_ = ~new_n16554_ | ~new_n16581_;
  assign new_n16846_ = ~new_n2388_ | ~new_n16443_;
  assign new_n16847_ = ~new_n2005_ | ~new_n16582_;
  assign new_n16848_ = ~new_n16555_;
  assign new_n16849_ = ~new_n16848_ | ~new_n16607_;
  assign new_n16850_ = ~new_n16555_ | ~new_n16442_;
  assign new_n16851_ = ~new_n2441_ | ~new_n16487_;
  assign new_n16852_ = ~new_n2008_ | ~new_n16486_;
  assign new_n16853_ = ~new_n16556_;
  assign new_n16854_ = ~new_n16691_ | ~new_n16853_;
  assign new_n16855_ = ~new_n16556_ | ~new_n16583_;
  assign new_n16856_ = ~new_n2439_ | ~new_n16485_;
  assign new_n16857_ = ~new_n2009_ | ~new_n16584_;
  assign new_n16858_ = ~new_n16557_;
  assign new_n16859_ = ~new_n16858_ | ~new_n16687_;
  assign new_n16860_ = ~new_n16557_ | ~new_n16484_;
  assign new_n16861_ = ~new_n2436_ | ~new_n16483_;
  assign new_n16862_ = ~new_n1996_ | ~new_n16482_;
  assign new_n16863_ = ~new_n16558_;
  assign new_n16864_ = ~new_n16683_ | ~new_n16863_;
  assign new_n16865_ = ~new_n16558_ | ~new_n16585_;
  assign new_n16866_ = ~new_n2433_ | ~new_n16478_;
  assign new_n16867_ = ~new_n2000_ | ~new_n16476_;
  assign new_n16868_ = ~new_n16867_ | ~new_n16866_;
  assign new_n16869_ = ~new_n2430_ | ~new_n16479_;
  assign new_n16870_ = ~new_n2001_ | ~new_n16466_;
  assign new_n16871_ = ~new_n16751_ | ~new_n16508_;
  assign new_n16872_ = ~new_n16586_ | ~new_n16743_;
  assign new_n16873_ = ~new_n2427_ | ~new_n16480_;
  assign new_n16874_ = ~new_n2006_ | ~new_n16477_;
  assign new_n16875_ = ~new_n16752_ | ~new_n16588_;
  assign new_n16876_ = ~new_n16673_ | ~new_n16587_;
  assign new_n16877_ = ~new_n2424_ | ~new_n16475_;
  assign new_n16878_ = ~new_n2007_ | ~new_n16474_;
  assign new_n16879_ = ~new_n16560_;
  assign new_n16880_ = ~new_n16669_ | ~new_n16879_;
  assign new_n16881_ = ~new_n16560_ | ~new_n16589_;
  assign new_n16882_ = ~new_n2421_ | ~new_n16473_;
  assign new_n16883_ = ~new_n1999_ | ~new_n16472_;
  assign new_n16884_ = ~new_n16561_;
  assign new_n16885_ = ~new_n16665_ | ~new_n16884_;
  assign new_n16886_ = ~new_n16561_ | ~new_n16590_;
  assign new_n16887_ = ~new_n2418_ | ~new_n16469_;
  assign new_n16888_ = ~new_n1990_ | ~new_n16467_;
  assign new_n16889_ = ~new_n16888_ | ~new_n16887_;
  assign new_n16890_ = ~new_n2415_ | ~new_n16470_;
  assign new_n16891_ = ~new_n1989_ | ~new_n16468_;
  assign new_n16892_ = ~new_n16762_ | ~new_n16509_;
  assign new_n16893_ = ~new_n16591_ | ~new_n16754_;
  assign new_n16894_ = new_n17072_ & new_n17089_;
  assign new_n16895_ = new_n17091_ & new_n17090_;
  assign new_n16896_ = new_n17067_ & new_n17128_;
  assign new_n16897_ = new_n17130_ & new_n17129_;
  assign new_n16898_ = new_n17147_ & new_n17146_;
  assign new_n16899_ = new_n17173_ & new_n17172_;
  assign new_n16900_ = new_n17271_ & new_n17270_;
  assign new_n16901_ = ~new_n17228_ | ~new_n17231_;
  assign new_n16902_ = ~new_n17217_ | ~new_n17220_;
  assign new_n16903_ = ~new_n17206_ | ~new_n17209_;
  assign new_n16904_ = ~new_n17198_ | ~new_n17200_;
  assign new_n16905_ = ~new_n17236_ | ~new_n17044_ | ~new_n17063_;
  assign new_n16906_ = ~new_n17124_ | ~new_n17126_;
  assign new_n16907_ = ~new_n17116_ | ~new_n17119_;
  assign new_n16908_ = ~new_n17108_ | ~new_n17110_;
  assign new_n16909_ = ~new_n16913_ | ~new_n17234_;
  assign new_n16910_ = ~new_n2406_;
  assign new_n16911_ = ~new_n2391_;
  assign new_n16912_ = ~new_n2383_;
  assign new_n16913_ = ~new_n2383_ | ~new_n16981_;
  assign new_n16914_ = ~new_n2005_;
  assign new_n16915_ = ~new_n2394_;
  assign new_n16916_ = ~new_n1995_;
  assign new_n16917_ = ~new_n1995_ | ~new_n16911_;
  assign new_n16918_ = ~new_n1991_;
  assign new_n16919_ = ~new_n2403_;
  assign new_n16920_ = ~new_n2400_;
  assign new_n16921_ = ~new_n2397_;
  assign new_n16922_ = ~new_n1998_;
  assign new_n16923_ = ~new_n1994_;
  assign new_n16924_ = ~new_n1987_;
  assign new_n16925_ = ~new_n1987_ | ~new_n16921_;
  assign new_n16926_ = ~new_n2409_;
  assign new_n16927_ = ~new_n1997_;
  assign new_n16928_ = ~new_n1997_ | ~new_n16910_;
  assign new_n16929_ = ~new_n2011_;
  assign new_n16930_ = ~new_n2412_;
  assign new_n16931_ = ~new_n2010_;
  assign new_n16932_ = ~new_n17097_ | ~new_n17096_;
  assign new_n16933_ = ~new_n16925_ | ~new_n17112_;
  assign new_n16934_ = ~new_n17081_ | ~new_n17080_;
  assign new_n16935_ = ~new_n2946_;
  assign new_n16936_ = ~new_n2950_;
  assign new_n16937_ = ~new_n2430_;
  assign new_n16938_ = ~new_n2418_;
  assign new_n16939_ = ~new_n2415_;
  assign new_n16940_ = ~new_n1990_;
  assign new_n16941_ = ~new_n1989_;
  assign new_n16942_ = ~new_n2010_ | ~new_n16930_;
  assign new_n16943_ = ~new_n2421_;
  assign new_n16944_ = ~new_n1999_;
  assign new_n16945_ = ~new_n2424_;
  assign new_n16946_ = ~new_n2007_;
  assign new_n16947_ = ~new_n2433_;
  assign new_n16948_ = ~new_n2427_;
  assign new_n16949_ = ~new_n2000_;
  assign new_n16950_ = ~new_n2001_;
  assign new_n16951_ = ~new_n2006_;
  assign new_n16952_ = ~new_n2006_ | ~new_n16948_;
  assign new_n16953_ = ~new_n2436_;
  assign new_n16954_ = ~new_n1996_;
  assign new_n16955_ = ~new_n17157_ | ~new_n17156_;
  assign new_n16956_ = ~new_n2009_;
  assign new_n16957_ = ~new_n2441_;
  assign new_n16958_ = ~new_n2008_;
  assign new_n16959_ = ~new_n2952_;
  assign new_n16960_ = ~new_n2003_;
  assign new_n16961_ = ~new_n2949_;
  assign new_n16962_ = ~new_n2951_;
  assign new_n16963_ = ~new_n1993_;
  assign new_n16964_ = ~new_n1988_;
  assign new_n16965_ = ~new_n2002_;
  assign new_n16966_ = ~new_n2002_ | ~new_n16962_;
  assign new_n16967_ = ~new_n2948_;
  assign new_n16968_ = ~new_n1992_;
  assign new_n16969_ = ~new_n2947_;
  assign new_n16970_ = ~new_n1985_;
  assign new_n16971_ = ~new_n2945_;
  assign new_n16972_ = ~new_n1984_;
  assign new_n16973_ = ~new_n1984_ | ~new_n16935_;
  assign new_n16974_ = ~new_n1980_;
  assign new_n16975_ = ~new_n2944_;
  assign new_n16976_ = ~new_n1981_;
  assign new_n16977_ = ~new_n17187_ | ~new_n17186_;
  assign new_n16978_ = ~new_n16966_ | ~new_n17202_;
  assign new_n16979_ = ~new_n16952_ | ~new_n17213_;
  assign new_n16980_ = ~new_n16942_ | ~new_n17224_;
  assign new_n16981_ = ~new_n2004_;
  assign new_n16982_ = ~new_n17281_ | ~new_n17280_;
  assign new_n16983_ = ~new_n17295_ | ~new_n17294_;
  assign new_n16984_ = ~new_n17300_ | ~new_n17299_;
  assign new_n16985_ = ~new_n17316_ | ~new_n17315_;
  assign new_n16986_ = ~new_n17321_ | ~new_n17320_;
  assign new_n16987_ = ~new_n17326_ | ~new_n17325_;
  assign new_n16988_ = ~new_n17331_ | ~new_n17330_;
  assign new_n16989_ = ~new_n17336_ | ~new_n17335_;
  assign new_n16990_ = ~new_n17352_ | ~new_n17351_;
  assign new_n16991_ = ~new_n17357_ | ~new_n17356_;
  assign new_n16992_ = ~new_n17240_ | ~new_n17239_;
  assign new_n16993_ = ~new_n17249_ | ~new_n17248_;
  assign new_n16994_ = ~new_n17256_ | ~new_n17255_;
  assign new_n16995_ = ~new_n17260_ | ~new_n17259_;
  assign new_n16996_ = ~new_n17269_ | ~new_n17268_;
  assign new_n16997_ = ~new_n17290_ | ~new_n17289_;
  assign new_n16998_ = ~new_n17307_ | ~new_n17306_;
  assign new_n16999_ = ~new_n17311_ | ~new_n17310_;
  assign new_n17000_ = ~new_n17343_ | ~new_n17342_;
  assign new_n17001_ = ~new_n17347_ | ~new_n17346_;
  assign new_n17002_ = ~new_n17364_ | ~new_n17363_;
  assign new_n17003_ = new_n17083_ & new_n17071_;
  assign new_n17004_ = new_n17086_ & new_n17087_;
  assign new_n17005_ = new_n17099_ & new_n17073_;
  assign new_n17006_ = new_n17102_ & new_n17103_;
  assign new_n17007_ = new_n16928_ & new_n17242_ & new_n17241_;
  assign new_n17008_ = new_n17245_ & new_n17073_;
  assign new_n17009_ = new_n17118_ & new_n16895_;
  assign new_n17010_ = new_n17252_ & new_n17072_;
  assign new_n17011_ = new_n16917_ & new_n17262_ & new_n17261_;
  assign new_n17012_ = new_n17265_ & new_n17071_;
  assign new_n17013_ = new_n17105_ & new_n16896_;
  assign new_n17014_ = new_n17150_ & new_n17068_;
  assign new_n17015_ = new_n17176_ & new_n17069_;
  assign new_n17016_ = new_n17192_ & new_n17193_;
  assign new_n17017_ = new_n17195_ & new_n17274_;
  assign new_n17018_ = new_n17196_ & new_n17193_ & new_n17192_;
  assign new_n17019_ = ~new_n17278_ | ~new_n17277_;
  assign new_n17020_ = new_n16973_ & new_n17283_ & new_n17282_;
  assign new_n17021_ = new_n17286_ & new_n17070_;
  assign new_n17022_ = ~new_n17292_ | ~new_n17291_;
  assign new_n17023_ = ~new_n17297_ | ~new_n17296_;
  assign new_n17024_ = new_n17303_ & new_n17069_;
  assign new_n17025_ = ~new_n17313_ | ~new_n17312_;
  assign new_n17026_ = ~new_n17318_ | ~new_n17317_;
  assign new_n17027_ = ~new_n17323_ | ~new_n17322_;
  assign new_n17028_ = ~new_n17328_ | ~new_n17327_;
  assign new_n17029_ = ~new_n17333_ | ~new_n17332_;
  assign new_n17030_ = new_n17339_ & new_n17068_;
  assign new_n17031_ = ~new_n17349_ | ~new_n17348_;
  assign new_n17032_ = ~new_n17354_ | ~new_n17353_;
  assign new_n17033_ = new_n17230_ & new_n16897_;
  assign new_n17034_ = new_n17360_ & new_n17067_;
  assign new_n17035_ = new_n17238_ & new_n17237_;
  assign new_n17036_ = ~new_n17006_ | ~new_n17100_;
  assign new_n17037_ = new_n17247_ & new_n17246_;
  assign new_n17038_ = new_n17254_ & new_n17253_;
  assign new_n17039_ = new_n17258_ & new_n17257_;
  assign new_n17040_ = ~new_n17004_ | ~new_n17084_;
  assign new_n17041_ = new_n17267_ & new_n17266_;
  assign new_n17042_ = ~new_n2955_;
  assign new_n17043_ = ~new_n1982_;
  assign new_n17044_ = new_n17276_ & new_n17275_;
  assign new_n17045_ = ~new_n17016_ | ~new_n17190_;
  assign new_n17046_ = new_n17288_ & new_n17287_;
  assign new_n17047_ = ~new_n17183_ | ~new_n17182_;
  assign new_n17048_ = ~new_n17179_ | ~new_n17178_;
  assign new_n17049_ = new_n17305_ & new_n17304_;
  assign new_n17050_ = new_n17309_ & new_n17308_;
  assign new_n17051_ = ~new_n17169_ | ~new_n17168_;
  assign new_n17052_ = ~new_n17165_ | ~new_n17164_;
  assign new_n17053_ = ~new_n2388_;
  assign new_n17054_ = ~new_n17161_ | ~new_n17160_;
  assign new_n17055_ = ~new_n2439_;
  assign new_n17056_ = ~new_n17153_ | ~new_n17152_;
  assign new_n17057_ = new_n17341_ & new_n17340_;
  assign new_n17058_ = new_n17345_ & new_n17344_;
  assign new_n17059_ = ~new_n17143_ | ~new_n17142_;
  assign new_n17060_ = ~new_n17139_ | ~new_n17138_;
  assign new_n17061_ = ~new_n17135_ | ~new_n17134_;
  assign new_n17062_ = new_n17362_ & new_n17361_;
  assign new_n17063_ = ~new_n17017_ | ~new_n17045_;
  assign new_n17064_ = ~new_n16973_;
  assign new_n17065_ = ~new_n16917_;
  assign new_n17066_ = ~new_n16928_;
  assign new_n17067_ = ~new_n2415_ | ~new_n16941_;
  assign new_n17068_ = ~new_n2430_ | ~new_n16950_;
  assign new_n17069_ = ~new_n2950_ | ~new_n16964_;
  assign new_n17070_ = ~new_n2946_ | ~new_n16972_;
  assign new_n17071_ = ~new_n2391_ | ~new_n16916_;
  assign new_n17072_ = ~new_n2400_ | ~new_n16923_;
  assign new_n17073_ = ~new_n2406_ | ~new_n16927_;
  assign new_n17074_ = ~new_n16952_;
  assign new_n17075_ = ~new_n16966_;
  assign new_n17076_ = ~new_n16925_;
  assign new_n17077_ = ~new_n16942_;
  assign new_n17078_ = ~new_n16913_;
  assign new_n17079_ = ~new_n17078_ | ~new_n16914_;
  assign new_n17080_ = ~new_n17079_ | ~new_n17053_;
  assign new_n17081_ = ~new_n2005_ | ~new_n16913_;
  assign new_n17082_ = ~new_n16934_;
  assign new_n17083_ = ~new_n2394_ | ~new_n16918_;
  assign new_n17084_ = ~new_n17003_ | ~new_n16934_;
  assign new_n17085_ = ~new_n16918_ | ~new_n16917_;
  assign new_n17086_ = ~new_n17085_ | ~new_n16915_;
  assign new_n17087_ = ~new_n1991_ | ~new_n17065_;
  assign new_n17088_ = ~new_n17040_;
  assign new_n17089_ = ~new_n2403_ | ~new_n16922_;
  assign new_n17090_ = ~new_n1998_ | ~new_n16919_;
  assign new_n17091_ = ~new_n1994_ | ~new_n16920_;
  assign new_n17092_ = ~new_n17076_ | ~new_n16894_;
  assign new_n17093_ = ~new_n16895_ | ~new_n17092_;
  assign new_n17094_ = ~new_n2397_ | ~new_n16924_;
  assign new_n17095_ = ~new_n2403_ | ~new_n16922_;
  assign new_n17096_ = ~new_n16894_ | ~new_n17094_ | ~new_n17040_;
  assign new_n17097_ = ~new_n17095_ | ~new_n17093_;
  assign new_n17098_ = ~new_n16932_;
  assign new_n17099_ = ~new_n2409_ | ~new_n16929_;
  assign new_n17100_ = ~new_n17005_ | ~new_n16932_;
  assign new_n17101_ = ~new_n16929_ | ~new_n16928_;
  assign new_n17102_ = ~new_n17101_ | ~new_n16926_;
  assign new_n17103_ = ~new_n2011_ | ~new_n17066_;
  assign new_n17104_ = ~new_n17036_;
  assign new_n17105_ = ~new_n2412_ | ~new_n16931_;
  assign new_n17106_ = ~new_n17105_ | ~new_n16942_;
  assign new_n17107_ = ~new_n17098_ | ~new_n16928_;
  assign new_n17108_ = ~new_n17008_ | ~new_n17107_;
  assign new_n17109_ = ~new_n16932_ | ~new_n17073_;
  assign new_n17110_ = ~new_n17007_ | ~new_n17109_;
  assign new_n17111_ = ~new_n16928_ | ~new_n17073_;
  assign new_n17112_ = ~new_n17094_ | ~new_n17040_;
  assign new_n17113_ = ~new_n16933_;
  assign new_n17114_ = ~new_n1994_ | ~new_n16920_;
  assign new_n17115_ = ~new_n17113_ | ~new_n17114_;
  assign new_n17116_ = ~new_n17010_ | ~new_n17115_;
  assign new_n17117_ = ~new_n16933_ | ~new_n17072_;
  assign new_n17118_ = ~new_n2403_ | ~new_n16922_;
  assign new_n17119_ = ~new_n17009_ | ~new_n17117_;
  assign new_n17120_ = ~new_n1994_ | ~new_n16920_;
  assign new_n17121_ = ~new_n17072_ | ~new_n17120_;
  assign new_n17122_ = ~new_n17094_ | ~new_n16925_;
  assign new_n17123_ = ~new_n17082_ | ~new_n16917_;
  assign new_n17124_ = ~new_n17012_ | ~new_n17123_;
  assign new_n17125_ = ~new_n16934_ | ~new_n17071_;
  assign new_n17126_ = ~new_n17011_ | ~new_n17125_;
  assign new_n17127_ = ~new_n16917_ | ~new_n17071_;
  assign new_n17128_ = ~new_n2418_ | ~new_n16940_;
  assign new_n17129_ = ~new_n1990_ | ~new_n16938_;
  assign new_n17130_ = ~new_n1989_ | ~new_n16939_;
  assign new_n17131_ = ~new_n17077_ | ~new_n16896_;
  assign new_n17132_ = ~new_n16897_ | ~new_n17131_;
  assign new_n17133_ = ~new_n2418_ | ~new_n16940_;
  assign new_n17134_ = ~new_n17013_ | ~new_n17036_;
  assign new_n17135_ = ~new_n17133_ | ~new_n17132_;
  assign new_n17136_ = ~new_n17061_;
  assign new_n17137_ = ~new_n2421_ | ~new_n16944_;
  assign new_n17138_ = ~new_n17137_ | ~new_n17061_;
  assign new_n17139_ = ~new_n1999_ | ~new_n16943_;
  assign new_n17140_ = ~new_n17060_;
  assign new_n17141_ = ~new_n2424_ | ~new_n16946_;
  assign new_n17142_ = ~new_n17141_ | ~new_n17060_;
  assign new_n17143_ = ~new_n2007_ | ~new_n16945_;
  assign new_n17144_ = ~new_n17059_;
  assign new_n17145_ = ~new_n2433_ | ~new_n16949_;
  assign new_n17146_ = ~new_n2000_ | ~new_n16947_;
  assign new_n17147_ = ~new_n2001_ | ~new_n16937_;
  assign new_n17148_ = ~new_n17074_ | ~new_n17068_;
  assign new_n17149_ = ~new_n16898_ | ~new_n17148_;
  assign new_n17150_ = ~new_n2427_ | ~new_n16951_;
  assign new_n17151_ = ~new_n2433_ | ~new_n16949_;
  assign new_n17152_ = ~new_n17145_ | ~new_n17059_ | ~new_n17014_;
  assign new_n17153_ = ~new_n17151_ | ~new_n17149_;
  assign new_n17154_ = ~new_n17056_;
  assign new_n17155_ = ~new_n2436_ | ~new_n16954_;
  assign new_n17156_ = ~new_n17155_ | ~new_n17056_;
  assign new_n17157_ = ~new_n1996_ | ~new_n16953_;
  assign new_n17158_ = ~new_n16955_;
  assign new_n17159_ = ~new_n17158_ | ~new_n16956_;
  assign new_n17160_ = ~new_n17159_ | ~new_n17055_;
  assign new_n17161_ = ~new_n2009_ | ~new_n16955_;
  assign new_n17162_ = ~new_n17054_;
  assign new_n17163_ = ~new_n2441_ | ~new_n16958_;
  assign new_n17164_ = ~new_n17163_ | ~new_n17054_;
  assign new_n17165_ = ~new_n2008_ | ~new_n16957_;
  assign new_n17166_ = ~new_n17052_;
  assign new_n17167_ = ~new_n2952_ | ~new_n16960_;
  assign new_n17168_ = ~new_n17167_ | ~new_n17052_;
  assign new_n17169_ = ~new_n2003_ | ~new_n16959_;
  assign new_n17170_ = ~new_n17051_;
  assign new_n17171_ = ~new_n2949_ | ~new_n16963_;
  assign new_n17172_ = ~new_n1993_ | ~new_n16961_;
  assign new_n17173_ = ~new_n1988_ | ~new_n16936_;
  assign new_n17174_ = ~new_n17075_ | ~new_n17069_;
  assign new_n17175_ = ~new_n16899_ | ~new_n17174_;
  assign new_n17176_ = ~new_n2951_ | ~new_n16965_;
  assign new_n17177_ = ~new_n2949_ | ~new_n16963_;
  assign new_n17178_ = ~new_n17171_ | ~new_n17051_ | ~new_n17015_;
  assign new_n17179_ = ~new_n17177_ | ~new_n17175_;
  assign new_n17180_ = ~new_n17048_;
  assign new_n17181_ = ~new_n2948_ | ~new_n16968_;
  assign new_n17182_ = ~new_n17181_ | ~new_n17048_;
  assign new_n17183_ = ~new_n1992_ | ~new_n16967_;
  assign new_n17184_ = ~new_n17047_;
  assign new_n17185_ = ~new_n2947_ | ~new_n16970_;
  assign new_n17186_ = ~new_n17185_ | ~new_n17047_;
  assign new_n17187_ = ~new_n1985_ | ~new_n16969_;
  assign new_n17188_ = ~new_n16977_;
  assign new_n17189_ = ~new_n2945_ | ~new_n16974_;
  assign new_n17190_ = ~new_n17189_ | ~new_n16977_ | ~new_n17070_;
  assign new_n17191_ = ~new_n16974_ | ~new_n16973_;
  assign new_n17192_ = ~new_n17191_ | ~new_n16971_;
  assign new_n17193_ = ~new_n1980_ | ~new_n17064_;
  assign new_n17194_ = ~new_n17045_;
  assign new_n17195_ = ~new_n2944_ | ~new_n16976_;
  assign new_n17196_ = ~new_n1981_ | ~new_n16975_;
  assign new_n17197_ = ~new_n17188_ | ~new_n16973_;
  assign new_n17198_ = ~new_n17021_ | ~new_n17197_;
  assign new_n17199_ = ~new_n16977_ | ~new_n17070_;
  assign new_n17200_ = ~new_n17020_ | ~new_n17199_;
  assign new_n17201_ = ~new_n16973_ | ~new_n17070_;
  assign new_n17202_ = ~new_n17176_ | ~new_n17051_;
  assign new_n17203_ = ~new_n16978_;
  assign new_n17204_ = ~new_n1988_ | ~new_n16936_;
  assign new_n17205_ = ~new_n17203_ | ~new_n17204_;
  assign new_n17206_ = ~new_n17024_ | ~new_n17205_;
  assign new_n17207_ = ~new_n16978_ | ~new_n17069_;
  assign new_n17208_ = ~new_n2949_ | ~new_n16963_;
  assign new_n17209_ = ~new_n16899_ | ~new_n17208_ | ~new_n17207_;
  assign new_n17210_ = ~new_n1988_ | ~new_n16936_;
  assign new_n17211_ = ~new_n17069_ | ~new_n17210_;
  assign new_n17212_ = ~new_n17176_ | ~new_n16966_;
  assign new_n17213_ = ~new_n17150_ | ~new_n17059_;
  assign new_n17214_ = ~new_n16979_;
  assign new_n17215_ = ~new_n2001_ | ~new_n16937_;
  assign new_n17216_ = ~new_n17214_ | ~new_n17215_;
  assign new_n17217_ = ~new_n17030_ | ~new_n17216_;
  assign new_n17218_ = ~new_n16979_ | ~new_n17068_;
  assign new_n17219_ = ~new_n2433_ | ~new_n16949_;
  assign new_n17220_ = ~new_n16898_ | ~new_n17219_ | ~new_n17218_;
  assign new_n17221_ = ~new_n2001_ | ~new_n16937_;
  assign new_n17222_ = ~new_n17068_ | ~new_n17221_;
  assign new_n17223_ = ~new_n17150_ | ~new_n16952_;
  assign new_n17224_ = ~new_n17105_ | ~new_n17036_;
  assign new_n17225_ = ~new_n16980_;
  assign new_n17226_ = ~new_n1989_ | ~new_n16939_;
  assign new_n17227_ = ~new_n17225_ | ~new_n17226_;
  assign new_n17228_ = ~new_n17034_ | ~new_n17227_;
  assign new_n17229_ = ~new_n16980_ | ~new_n17067_;
  assign new_n17230_ = ~new_n2418_ | ~new_n16940_;
  assign new_n17231_ = ~new_n17033_ | ~new_n17229_;
  assign new_n17232_ = ~new_n1989_ | ~new_n16939_;
  assign new_n17233_ = ~new_n17067_ | ~new_n17232_;
  assign new_n17234_ = ~new_n2004_ | ~new_n16912_;
  assign new_n17235_ = ~new_n17189_ | ~new_n16977_ | ~new_n17070_;
  assign new_n17236_ = ~new_n17018_ | ~new_n16900_ | ~new_n17235_;
  assign new_n17237_ = ~new_n2412_ | ~new_n16931_;
  assign new_n17238_ = ~new_n2010_ | ~new_n16930_;
  assign new_n17239_ = ~new_n17106_ | ~new_n17036_;
  assign new_n17240_ = ~new_n17104_ | ~new_n17035_;
  assign new_n17241_ = ~new_n2409_ | ~new_n16929_;
  assign new_n17242_ = ~new_n2011_ | ~new_n16926_;
  assign new_n17243_ = ~new_n2409_ | ~new_n16929_;
  assign new_n17244_ = ~new_n2011_ | ~new_n16926_;
  assign new_n17245_ = ~new_n17244_ | ~new_n17243_;
  assign new_n17246_ = ~new_n2406_ | ~new_n16927_;
  assign new_n17247_ = ~new_n1997_ | ~new_n16910_;
  assign new_n17248_ = ~new_n17111_ | ~new_n16932_;
  assign new_n17249_ = ~new_n17037_ | ~new_n17098_;
  assign new_n17250_ = ~new_n2403_ | ~new_n16922_;
  assign new_n17251_ = ~new_n1998_ | ~new_n16919_;
  assign new_n17252_ = ~new_n17251_ | ~new_n17250_;
  assign new_n17253_ = ~new_n2400_ | ~new_n16923_;
  assign new_n17254_ = ~new_n1994_ | ~new_n16920_;
  assign new_n17255_ = ~new_n17121_ | ~new_n16933_;
  assign new_n17256_ = ~new_n17038_ | ~new_n17113_;
  assign new_n17257_ = ~new_n2397_ | ~new_n16924_;
  assign new_n17258_ = ~new_n1987_ | ~new_n16921_;
  assign new_n17259_ = ~new_n17122_ | ~new_n17040_;
  assign new_n17260_ = ~new_n17088_ | ~new_n17039_;
  assign new_n17261_ = ~new_n2394_ | ~new_n16918_;
  assign new_n17262_ = ~new_n1991_ | ~new_n16915_;
  assign new_n17263_ = ~new_n2394_ | ~new_n16918_;
  assign new_n17264_ = ~new_n1991_ | ~new_n16915_;
  assign new_n17265_ = ~new_n17264_ | ~new_n17263_;
  assign new_n17266_ = ~new_n2391_ | ~new_n16916_;
  assign new_n17267_ = ~new_n1995_ | ~new_n16911_;
  assign new_n17268_ = ~new_n17127_ | ~new_n16934_;
  assign new_n17269_ = ~new_n17041_ | ~new_n17082_;
  assign new_n17270_ = ~new_n2955_ | ~new_n17043_;
  assign new_n17271_ = ~new_n1982_ | ~new_n17042_;
  assign new_n17272_ = ~new_n2955_ | ~new_n17043_;
  assign new_n17273_ = ~new_n1982_ | ~new_n17042_;
  assign new_n17274_ = ~new_n17273_ | ~new_n17272_;
  assign new_n17275_ = ~new_n16975_ | ~new_n1981_ | ~new_n17274_;
  assign new_n17276_ = ~new_n2944_ | ~new_n16900_ | ~new_n16976_;
  assign new_n17277_ = ~new_n2944_ | ~new_n16976_;
  assign new_n17278_ = ~new_n1981_ | ~new_n16975_;
  assign new_n17279_ = ~new_n17019_;
  assign new_n17280_ = ~new_n17194_ | ~new_n17279_;
  assign new_n17281_ = ~new_n17019_ | ~new_n17045_;
  assign new_n17282_ = ~new_n2945_ | ~new_n16974_;
  assign new_n17283_ = ~new_n1980_ | ~new_n16971_;
  assign new_n17284_ = ~new_n2945_ | ~new_n16974_;
  assign new_n17285_ = ~new_n1980_ | ~new_n16971_;
  assign new_n17286_ = ~new_n17285_ | ~new_n17284_;
  assign new_n17287_ = ~new_n2946_ | ~new_n16972_;
  assign new_n17288_ = ~new_n1984_ | ~new_n16935_;
  assign new_n17289_ = ~new_n17201_ | ~new_n16977_;
  assign new_n17290_ = ~new_n17046_ | ~new_n17188_;
  assign new_n17291_ = ~new_n2947_ | ~new_n16970_;
  assign new_n17292_ = ~new_n1985_ | ~new_n16969_;
  assign new_n17293_ = ~new_n17022_;
  assign new_n17294_ = ~new_n17184_ | ~new_n17293_;
  assign new_n17295_ = ~new_n17022_ | ~new_n17047_;
  assign new_n17296_ = ~new_n2948_ | ~new_n16968_;
  assign new_n17297_ = ~new_n1992_ | ~new_n16967_;
  assign new_n17298_ = ~new_n17023_;
  assign new_n17299_ = ~new_n17180_ | ~new_n17298_;
  assign new_n17300_ = ~new_n17023_ | ~new_n17048_;
  assign new_n17301_ = ~new_n2949_ | ~new_n16963_;
  assign new_n17302_ = ~new_n1993_ | ~new_n16961_;
  assign new_n17303_ = ~new_n17302_ | ~new_n17301_;
  assign new_n17304_ = ~new_n2950_ | ~new_n16964_;
  assign new_n17305_ = ~new_n1988_ | ~new_n16936_;
  assign new_n17306_ = ~new_n17211_ | ~new_n16978_;
  assign new_n17307_ = ~new_n17049_ | ~new_n17203_;
  assign new_n17308_ = ~new_n2951_ | ~new_n16965_;
  assign new_n17309_ = ~new_n2002_ | ~new_n16962_;
  assign new_n17310_ = ~new_n17212_ | ~new_n17051_;
  assign new_n17311_ = ~new_n17170_ | ~new_n17050_;
  assign new_n17312_ = ~new_n2952_ | ~new_n16960_;
  assign new_n17313_ = ~new_n2003_ | ~new_n16959_;
  assign new_n17314_ = ~new_n17025_;
  assign new_n17315_ = ~new_n17166_ | ~new_n17314_;
  assign new_n17316_ = ~new_n17025_ | ~new_n17052_;
  assign new_n17317_ = ~new_n2388_ | ~new_n16914_;
  assign new_n17318_ = ~new_n2005_ | ~new_n17053_;
  assign new_n17319_ = ~new_n17026_;
  assign new_n17320_ = ~new_n17319_ | ~new_n17078_;
  assign new_n17321_ = ~new_n17026_ | ~new_n16913_;
  assign new_n17322_ = ~new_n2441_ | ~new_n16958_;
  assign new_n17323_ = ~new_n2008_ | ~new_n16957_;
  assign new_n17324_ = ~new_n17027_;
  assign new_n17325_ = ~new_n17162_ | ~new_n17324_;
  assign new_n17326_ = ~new_n17027_ | ~new_n17054_;
  assign new_n17327_ = ~new_n2439_ | ~new_n16956_;
  assign new_n17328_ = ~new_n2009_ | ~new_n17055_;
  assign new_n17329_ = ~new_n17028_;
  assign new_n17330_ = ~new_n17329_ | ~new_n17158_;
  assign new_n17331_ = ~new_n17028_ | ~new_n16955_;
  assign new_n17332_ = ~new_n2436_ | ~new_n16954_;
  assign new_n17333_ = ~new_n1996_ | ~new_n16953_;
  assign new_n17334_ = ~new_n17029_;
  assign new_n17335_ = ~new_n17154_ | ~new_n17334_;
  assign new_n17336_ = ~new_n17029_ | ~new_n17056_;
  assign new_n17337_ = ~new_n2433_ | ~new_n16949_;
  assign new_n17338_ = ~new_n2000_ | ~new_n16947_;
  assign new_n17339_ = ~new_n17338_ | ~new_n17337_;
  assign new_n17340_ = ~new_n2430_ | ~new_n16950_;
  assign new_n17341_ = ~new_n2001_ | ~new_n16937_;
  assign new_n17342_ = ~new_n17222_ | ~new_n16979_;
  assign new_n17343_ = ~new_n17057_ | ~new_n17214_;
  assign new_n17344_ = ~new_n2427_ | ~new_n16951_;
  assign new_n17345_ = ~new_n2006_ | ~new_n16948_;
  assign new_n17346_ = ~new_n17223_ | ~new_n17059_;
  assign new_n17347_ = ~new_n17144_ | ~new_n17058_;
  assign new_n17348_ = ~new_n2424_ | ~new_n16946_;
  assign new_n17349_ = ~new_n2007_ | ~new_n16945_;
  assign new_n17350_ = ~new_n17031_;
  assign new_n17351_ = ~new_n17140_ | ~new_n17350_;
  assign new_n17352_ = ~new_n17031_ | ~new_n17060_;
  assign new_n17353_ = ~new_n2421_ | ~new_n16944_;
  assign new_n17354_ = ~new_n1999_ | ~new_n16943_;
  assign new_n17355_ = ~new_n17032_;
  assign new_n17356_ = ~new_n17136_ | ~new_n17355_;
  assign new_n17357_ = ~new_n17032_ | ~new_n17061_;
  assign new_n17358_ = ~new_n2418_ | ~new_n16940_;
  assign new_n17359_ = ~new_n1990_ | ~new_n16938_;
  assign new_n17360_ = ~new_n17359_ | ~new_n17358_;
  assign new_n17361_ = ~new_n2415_ | ~new_n16941_;
  assign new_n17362_ = ~new_n1989_ | ~new_n16939_;
  assign new_n17363_ = ~new_n17233_ | ~new_n16980_;
  assign new_n17364_ = ~new_n17062_ | ~new_n17225_;
  assign new_n17365_ = new_n17537_ & new_n17536_;
  assign new_n17366_ = new_n17538_ & new_n17539_;
  assign new_n17367_ = new_n17555_ & new_n17554_;
  assign new_n17368_ = new_n17595_ & new_n17594_;
  assign new_n17369_ = new_n17604_ & new_n17603_;
  assign new_n17370_ = new_n17622_ & new_n17621_;
  assign new_n17371_ = new_n17630_ & new_n17629_;
  assign new_n17372_ = new_n17709_ & new_n17706_;
  assign new_n17373_ = new_n17702_ & new_n17699_;
  assign new_n17374_ = new_n17693_ & new_n17690_;
  assign new_n17375_ = new_n17684_ & new_n17681_;
  assign new_n17376_ = new_n17678_ & new_n17676_;
  assign new_n17377_ = new_n17671_ & new_n17668_;
  assign new_n17378_ = new_n17593_ & new_n17590_;
  assign new_n17379_ = new_n17585_ & new_n17582_;
  assign new_n17380_ = new_n17571_ & new_n17568_;
  assign new_n17381_ = ~new_n2403_;
  assign new_n17382_ = ~new_n1998_;
  assign new_n17383_ = ~new_n1997_;
  assign new_n17384_ = ~new_n1998_ | ~new_n2403_;
  assign new_n17385_ = ~new_n2406_;
  assign new_n17386_ = ~new_n2397_;
  assign new_n17387_ = ~new_n1987_;
  assign new_n17388_ = ~new_n1994_;
  assign new_n17389_ = ~new_n2391_;
  assign new_n17390_ = ~new_n1995_;
  assign new_n17391_ = ~new_n2383_;
  assign new_n17392_ = ~new_n2004_;
  assign new_n17393_ = ~new_n2004_ | ~new_n2383_;
  assign new_n17394_ = ~new_n2394_;
  assign new_n17395_ = ~new_n1991_;
  assign new_n17396_ = ~new_n1987_ | ~new_n2397_;
  assign new_n17397_ = ~new_n2400_;
  assign new_n17398_ = ~new_n2409_;
  assign new_n17399_ = ~new_n2011_;
  assign new_n17400_ = ~new_n2010_;
  assign new_n17401_ = ~new_n2412_;
  assign new_n17402_ = ~new_n17423_ | ~new_n17563_;
  assign new_n17403_ = ~new_n17479_ | ~new_n17551_;
  assign new_n17404_ = ~new_n17540_ | ~new_n17541_;
  assign new_n17405_ = ~new_n2388_ | ~new_n2005_;
  assign new_n17406_ = ~new_n17483_ | ~new_n17577_;
  assign new_n17407_ = ~new_n17574_ | ~new_n17573_;
  assign new_n17408_ = ~new_n2945_;
  assign new_n17409_ = ~new_n1980_;
  assign new_n17410_ = ~new_n1984_;
  assign new_n17411_ = ~new_n2946_;
  assign new_n17412_ = ~new_n2947_;
  assign new_n17413_ = ~new_n1985_;
  assign new_n17414_ = ~new_n2948_;
  assign new_n17415_ = ~new_n1992_;
  assign new_n17416_ = ~new_n2951_;
  assign new_n17417_ = ~new_n2002_;
  assign new_n17418_ = ~new_n2433_;
  assign new_n17419_ = ~new_n2000_;
  assign new_n17420_ = ~new_n1996_;
  assign new_n17421_ = ~new_n2000_ | ~new_n2433_;
  assign new_n17422_ = ~new_n2436_;
  assign new_n17423_ = ~new_n2011_ | ~new_n2409_;
  assign new_n17424_ = ~new_n2415_;
  assign new_n17425_ = ~new_n1989_;
  assign new_n17426_ = ~new_n2421_;
  assign new_n17427_ = ~new_n1999_;
  assign new_n17428_ = ~new_n2418_;
  assign new_n17429_ = ~new_n1990_;
  assign new_n17430_ = ~new_n1990_ | ~new_n2418_;
  assign new_n17431_ = ~new_n2424_;
  assign new_n17432_ = ~new_n2007_;
  assign new_n17433_ = ~new_n2427_;
  assign new_n17434_ = ~new_n2006_;
  assign new_n17435_ = ~new_n2430_;
  assign new_n17436_ = ~new_n2001_;
  assign new_n17437_ = ~new_n2439_;
  assign new_n17438_ = ~new_n2009_;
  assign new_n17439_ = ~new_n2009_ | ~new_n2439_;
  assign new_n17440_ = ~new_n2441_;
  assign new_n17441_ = ~new_n2008_;
  assign new_n17442_ = ~new_n2008_ | ~new_n2441_;
  assign new_n17443_ = ~new_n2952_;
  assign new_n17444_ = ~new_n2950_;
  assign new_n17445_ = ~new_n1988_;
  assign new_n17446_ = ~new_n2949_;
  assign new_n17447_ = ~new_n1993_;
  assign new_n17448_ = ~new_n2946_ | ~new_n1984_;
  assign new_n17449_ = ~new_n1981_;
  assign new_n17450_ = ~new_n2944_;
  assign new_n17451_ = ~new_n17664_ | ~new_n17534_;
  assign new_n17452_ = ~new_n2003_;
  assign new_n17453_ = ~new_n17439_ | ~new_n17673_;
  assign new_n17454_ = ~new_n17619_ | ~new_n17618_;
  assign new_n17455_ = ~new_n17430_ | ~new_n17695_;
  assign new_n17456_ = ~new_n17815_ | ~new_n17814_;
  assign new_n17457_ = ~new_n17862_ | ~new_n17861_;
  assign new_n17458_ = ~new_n17733_ | ~new_n17732_;
  assign new_n17459_ = ~new_n17738_ | ~new_n17737_;
  assign new_n17460_ = ~new_n17745_ | ~new_n17744_;
  assign new_n17461_ = ~new_n17752_ | ~new_n17751_;
  assign new_n17462_ = ~new_n17757_ | ~new_n17756_;
  assign new_n17463_ = ~new_n17766_ | ~new_n17765_;
  assign new_n17464_ = ~new_n17773_ | ~new_n17772_;
  assign new_n17465_ = ~new_n17780_ | ~new_n17779_;
  assign new_n17466_ = ~new_n17787_ | ~new_n17786_;
  assign new_n17467_ = ~new_n17792_ | ~new_n17791_;
  assign new_n17468_ = ~new_n17799_ | ~new_n17798_;
  assign new_n17469_ = ~new_n17806_ | ~new_n17805_;
  assign new_n17470_ = ~new_n17820_ | ~new_n17819_;
  assign new_n17471_ = ~new_n17825_ | ~new_n17824_;
  assign new_n17472_ = ~new_n17832_ | ~new_n17831_;
  assign new_n17473_ = ~new_n17839_ | ~new_n17838_;
  assign new_n17474_ = ~new_n17846_ | ~new_n17845_;
  assign new_n17475_ = ~new_n17853_ | ~new_n17852_;
  assign new_n17476_ = ~new_n17858_ | ~new_n17857_;
  assign new_n17477_ = new_n2391_ & new_n1995_;
  assign new_n17478_ = new_n17547_ & new_n17545_;
  assign new_n17479_ = new_n17552_ & new_n17550_;
  assign new_n17480_ = new_n17559_ & new_n17558_;
  assign new_n17481_ = new_n17384_ & new_n17740_ & new_n17739_;
  assign new_n17482_ = new_n17570_ & new_n17367_;
  assign new_n17483_ = new_n17578_ & new_n17576_;
  assign new_n17484_ = new_n17396_ & new_n17747_ & new_n17746_;
  assign new_n17485_ = new_n17584_ & new_n17365_;
  assign new_n17486_ = new_n17592_ & new_n17539_;
  assign new_n17487_ = new_n17562_ & new_n17368_;
  assign new_n17488_ = new_n17597_ & new_n17529_;
  assign new_n17489_ = new_n17606_ & new_n17530_;
  assign new_n17490_ = new_n17626_ & new_n17625_;
  assign new_n17491_ = new_n17371_ & new_n17640_;
  assign new_n17492_ = new_n17643_ & new_n17638_;
  assign new_n17493_ = new_n17659_ & new_n17656_;
  assign new_n17494_ = new_n17726_ & new_n17660_;
  assign new_n17495_ = new_n17517_ & new_n17636_;
  assign new_n17496_ = new_n17421_ & new_n17827_ & new_n17826_;
  assign new_n17497_ = new_n17530_ & new_n17848_ & new_n17847_;
  assign new_n17498_ = new_n17701_ & new_n17369_;
  assign new_n17499_ = new_n17529_ & new_n17860_ & new_n17859_;
  assign new_n17500_ = new_n17708_ & new_n17368_;
  assign new_n17501_ = ~new_n17480_ | ~new_n17560_;
  assign new_n17502_ = ~new_n17575_ | ~new_n17587_;
  assign new_n17503_ = ~new_n1982_;
  assign new_n17504_ = ~new_n2955_;
  assign new_n17505_ = new_n17761_ & new_n17760_;
  assign new_n17506_ = ~new_n17722_ | ~new_n17662_ | ~new_n17527_;
  assign new_n17507_ = new_n17768_ & new_n17767_;
  assign new_n17508_ = ~new_n17494_ | ~new_n17728_ | ~new_n17727_;
  assign new_n17509_ = new_n17775_ & new_n17774_;
  assign new_n17510_ = ~new_n17448_ | ~new_n17723_ | ~new_n17657_;
  assign new_n17511_ = new_n17782_ & new_n17781_;
  assign new_n17512_ = ~new_n17651_ | ~new_n17650_;
  assign new_n17513_ = new_n17794_ & new_n17793_;
  assign new_n17514_ = ~new_n17647_ | ~new_n17646_;
  assign new_n17515_ = new_n17801_ & new_n17800_;
  assign new_n17516_ = ~new_n17492_ | ~new_n17642_;
  assign new_n17517_ = new_n17808_ & new_n17807_;
  assign new_n17518_ = new_n17813_ & new_n17812_;
  assign new_n17519_ = ~new_n17405_ | ~new_n17685_;
  assign new_n17520_ = ~new_n17490_ | ~new_n17627_;
  assign new_n17521_ = new_n17834_ & new_n17833_;
  assign new_n17522_ = ~new_n17615_ | ~new_n17614_;
  assign new_n17523_ = new_n17841_ & new_n17840_;
  assign new_n17524_ = ~new_n17611_ | ~new_n17610_;
  assign new_n17525_ = ~new_n17601_ | ~new_n17600_;
  assign new_n17526_ = ~new_n17725_ | ~new_n17724_;
  assign new_n17527_ = ~new_n1981_ | ~new_n17508_;
  assign new_n17528_ = ~new_n17396_;
  assign new_n17529_ = ~new_n2412_ | ~new_n2010_;
  assign new_n17530_ = ~new_n1999_ | ~new_n2421_;
  assign new_n17531_ = ~new_n1985_ | ~new_n2947_;
  assign new_n17532_ = ~new_n17430_;
  assign new_n17533_ = ~new_n17439_;
  assign new_n17534_ = ~new_n1992_ | ~new_n2948_;
  assign new_n17535_ = ~new_n17423_;
  assign new_n17536_ = new_n1994_ | new_n2400_;
  assign new_n17537_ = new_n1987_ | new_n2397_;
  assign new_n17538_ = new_n2394_ | new_n1991_;
  assign new_n17539_ = new_n2391_ | new_n1995_;
  assign new_n17540_ = ~new_n17393_;
  assign new_n17541_ = new_n2388_ | new_n2005_;
  assign new_n17542_ = ~new_n17404_;
  assign new_n17543_ = ~new_n17405_;
  assign new_n17544_ = ~new_n17404_ | ~new_n17405_;
  assign new_n17545_ = ~new_n17477_ | ~new_n17538_;
  assign new_n17546_ = ~new_n17366_ | ~new_n17544_;
  assign new_n17547_ = ~new_n1991_ | ~new_n2394_;
  assign new_n17548_ = ~new_n17478_ | ~new_n17546_;
  assign new_n17549_ = ~new_n17397_ | ~new_n17396_;
  assign new_n17550_ = ~new_n1994_ | ~new_n17549_;
  assign new_n17551_ = ~new_n17365_ | ~new_n17548_;
  assign new_n17552_ = ~new_n2400_ | ~new_n17528_;
  assign new_n17553_ = ~new_n17403_;
  assign new_n17554_ = new_n1997_ | new_n2406_;
  assign new_n17555_ = new_n1998_ | new_n2403_;
  assign new_n17556_ = ~new_n17384_;
  assign new_n17557_ = ~new_n17385_ | ~new_n17384_;
  assign new_n17558_ = ~new_n1997_ | ~new_n17557_;
  assign new_n17559_ = ~new_n2406_ | ~new_n17556_;
  assign new_n17560_ = ~new_n17367_ | ~new_n17403_;
  assign new_n17561_ = ~new_n17501_;
  assign new_n17562_ = new_n2409_ | new_n2011_;
  assign new_n17563_ = ~new_n17562_ | ~new_n17501_;
  assign new_n17564_ = ~new_n17402_;
  assign new_n17565_ = new_n2010_ | new_n2412_;
  assign new_n17566_ = new_n2403_ | new_n1998_;
  assign new_n17567_ = ~new_n17566_ | ~new_n17403_;
  assign new_n17568_ = ~new_n17481_ | ~new_n17567_;
  assign new_n17569_ = ~new_n17553_ | ~new_n17384_;
  assign new_n17570_ = ~new_n2406_ | ~new_n1997_;
  assign new_n17571_ = ~new_n17482_ | ~new_n17569_;
  assign new_n17572_ = new_n1998_ | new_n2403_;
  assign new_n17573_ = ~new_n17543_ | ~new_n17539_;
  assign new_n17574_ = ~new_n1995_ | ~new_n2391_;
  assign new_n17575_ = ~new_n17407_;
  assign new_n17576_ = ~new_n17542_ | ~new_n17366_;
  assign new_n17577_ = ~new_n17407_ | ~new_n17538_;
  assign new_n17578_ = ~new_n1991_ | ~new_n2394_;
  assign new_n17579_ = ~new_n17406_;
  assign new_n17580_ = new_n2397_ | new_n1987_;
  assign new_n17581_ = ~new_n17580_ | ~new_n17406_;
  assign new_n17582_ = ~new_n17484_ | ~new_n17581_;
  assign new_n17583_ = ~new_n17579_ | ~new_n17396_;
  assign new_n17584_ = ~new_n2400_ | ~new_n1994_;
  assign new_n17585_ = ~new_n17485_ | ~new_n17583_;
  assign new_n17586_ = new_n1987_ | new_n2397_;
  assign new_n17587_ = ~new_n17542_ | ~new_n17539_;
  assign new_n17588_ = ~new_n17502_;
  assign new_n17589_ = ~new_n1991_ | ~new_n2394_;
  assign new_n17590_ = ~new_n17758_ | ~new_n17404_ | ~new_n17405_ | ~new_n17759_;
  assign new_n17591_ = ~new_n17405_ | ~new_n17404_;
  assign new_n17592_ = ~new_n1995_ | ~new_n2391_;
  assign new_n17593_ = ~new_n17486_ | ~new_n17591_;
  assign new_n17594_ = new_n2010_ | new_n2412_;
  assign new_n17595_ = new_n1989_ | new_n2415_;
  assign new_n17596_ = ~new_n17535_ | ~new_n17368_;
  assign new_n17597_ = ~new_n1989_ | ~new_n2415_;
  assign new_n17598_ = ~new_n17488_ | ~new_n17596_;
  assign new_n17599_ = new_n2415_ | new_n1989_;
  assign new_n17600_ = ~new_n17487_ | ~new_n17501_;
  assign new_n17601_ = ~new_n17599_ | ~new_n17598_;
  assign new_n17602_ = ~new_n17525_;
  assign new_n17603_ = new_n2007_ | new_n2424_;
  assign new_n17604_ = new_n1999_ | new_n2421_;
  assign new_n17605_ = ~new_n17532_ | ~new_n17369_;
  assign new_n17606_ = ~new_n2007_ | ~new_n2424_;
  assign new_n17607_ = ~new_n17489_ | ~new_n17605_;
  assign new_n17608_ = new_n2418_ | new_n1990_;
  assign new_n17609_ = new_n2424_ | new_n2007_;
  assign new_n17610_ = ~new_n17369_ | ~new_n17608_ | ~new_n17525_;
  assign new_n17611_ = ~new_n17609_ | ~new_n17607_;
  assign new_n17612_ = ~new_n17524_;
  assign new_n17613_ = new_n2427_ | new_n2006_;
  assign new_n17614_ = ~new_n17613_ | ~new_n17524_;
  assign new_n17615_ = ~new_n2006_ | ~new_n2427_;
  assign new_n17616_ = ~new_n17522_;
  assign new_n17617_ = new_n2430_ | new_n2001_;
  assign new_n17618_ = ~new_n17617_ | ~new_n17522_;
  assign new_n17619_ = ~new_n2001_ | ~new_n2430_;
  assign new_n17620_ = ~new_n17454_;
  assign new_n17621_ = new_n1996_ | new_n2436_;
  assign new_n17622_ = new_n2000_ | new_n2433_;
  assign new_n17623_ = ~new_n17421_;
  assign new_n17624_ = ~new_n17422_ | ~new_n17421_;
  assign new_n17625_ = ~new_n1996_ | ~new_n17624_;
  assign new_n17626_ = ~new_n2436_ | ~new_n17623_;
  assign new_n17627_ = ~new_n17370_ | ~new_n17454_;
  assign new_n17628_ = ~new_n17520_;
  assign new_n17629_ = new_n2003_ | new_n2952_;
  assign new_n17630_ = new_n2008_ | new_n2441_;
  assign new_n17631_ = new_n2002_ | new_n2951_;
  assign new_n17632_ = ~new_n17442_;
  assign new_n17633_ = ~new_n2952_ | ~new_n17632_;
  assign new_n17634_ = ~new_n17633_ | ~new_n17452_;
  assign new_n17635_ = ~new_n17442_ | ~new_n17443_;
  assign new_n17636_ = ~new_n17635_ | ~new_n17634_;
  assign new_n17637_ = ~new_n17533_ | ~new_n17371_;
  assign new_n17638_ = ~new_n2002_ | ~new_n2951_;
  assign new_n17639_ = ~new_n17636_ | ~new_n17637_;
  assign new_n17640_ = new_n2439_ | new_n2009_;
  assign new_n17641_ = new_n2951_ | new_n2002_;
  assign new_n17642_ = ~new_n17491_ | ~new_n17631_ | ~new_n17520_;
  assign new_n17643_ = ~new_n17641_ | ~new_n17639_;
  assign new_n17644_ = ~new_n17516_;
  assign new_n17645_ = new_n2950_ | new_n1988_;
  assign new_n17646_ = ~new_n17645_ | ~new_n17516_;
  assign new_n17647_ = ~new_n1988_ | ~new_n2950_;
  assign new_n17648_ = ~new_n17514_;
  assign new_n17649_ = new_n2949_ | new_n1993_;
  assign new_n17650_ = ~new_n17649_ | ~new_n17514_;
  assign new_n17651_ = ~new_n1993_ | ~new_n2949_;
  assign new_n17652_ = ~new_n17512_;
  assign new_n17653_ = new_n1985_ | new_n2947_;
  assign new_n17654_ = ~new_n17534_ | ~new_n17531_;
  assign new_n17655_ = ~new_n17448_;
  assign new_n17656_ = new_n2948_ | new_n1992_;
  assign new_n17657_ = ~new_n17526_ | ~new_n17512_ | ~new_n17656_;
  assign new_n17658_ = ~new_n17510_;
  assign new_n17659_ = new_n2945_ | new_n1980_;
  assign new_n17660_ = ~new_n1980_ | ~new_n2945_;
  assign new_n17661_ = ~new_n17508_;
  assign new_n17662_ = ~new_n2944_ | ~new_n17508_;
  assign new_n17663_ = ~new_n17506_;
  assign new_n17664_ = ~new_n17656_ | ~new_n17512_;
  assign new_n17665_ = ~new_n17451_;
  assign new_n17666_ = new_n2947_ | new_n1985_;
  assign new_n17667_ = ~new_n17666_ | ~new_n17451_;
  assign new_n17668_ = ~new_n17511_ | ~new_n17667_ | ~new_n17531_;
  assign new_n17669_ = ~new_n17665_ | ~new_n17531_;
  assign new_n17670_ = ~new_n2946_ | ~new_n1984_;
  assign new_n17671_ = ~new_n17526_ | ~new_n17669_ | ~new_n17670_;
  assign new_n17672_ = new_n1985_ | new_n2947_;
  assign new_n17673_ = ~new_n17640_ | ~new_n17520_;
  assign new_n17674_ = ~new_n17453_;
  assign new_n17675_ = ~new_n17371_ | ~new_n17453_;
  assign new_n17676_ = ~new_n17495_ | ~new_n17675_;
  assign new_n17677_ = ~new_n17675_ | ~new_n17636_;
  assign new_n17678_ = ~new_n17811_ | ~new_n17677_;
  assign new_n17679_ = new_n2441_ | new_n2008_;
  assign new_n17680_ = ~new_n17679_ | ~new_n17453_;
  assign new_n17681_ = ~new_n17518_ | ~new_n17680_ | ~new_n17442_;
  assign new_n17682_ = ~new_n17674_ | ~new_n17442_;
  assign new_n17683_ = ~new_n2003_ | ~new_n2952_;
  assign new_n17684_ = ~new_n17371_ | ~new_n17683_ | ~new_n17682_;
  assign new_n17685_ = new_n2388_ | new_n2005_;
  assign new_n17686_ = ~new_n17519_;
  assign new_n17687_ = new_n2008_ | new_n2441_;
  assign new_n17688_ = new_n2433_ | new_n2000_;
  assign new_n17689_ = ~new_n17688_ | ~new_n17454_;
  assign new_n17690_ = ~new_n17496_ | ~new_n17689_;
  assign new_n17691_ = ~new_n17620_ | ~new_n17421_;
  assign new_n17692_ = ~new_n2436_ | ~new_n1996_;
  assign new_n17693_ = ~new_n17370_ | ~new_n17692_ | ~new_n17691_;
  assign new_n17694_ = new_n2000_ | new_n2433_;
  assign new_n17695_ = ~new_n17608_ | ~new_n17525_;
  assign new_n17696_ = ~new_n17455_;
  assign new_n17697_ = new_n2421_ | new_n1999_;
  assign new_n17698_ = ~new_n17697_ | ~new_n17455_;
  assign new_n17699_ = ~new_n17497_ | ~new_n17698_;
  assign new_n17700_ = ~new_n17696_ | ~new_n17530_;
  assign new_n17701_ = ~new_n2007_ | ~new_n2424_;
  assign new_n17702_ = ~new_n17498_ | ~new_n17700_;
  assign new_n17703_ = new_n1999_ | new_n2421_;
  assign new_n17704_ = new_n2412_ | new_n2010_;
  assign new_n17705_ = ~new_n17704_ | ~new_n17402_;
  assign new_n17706_ = ~new_n17499_ | ~new_n17705_;
  assign new_n17707_ = ~new_n17564_ | ~new_n17529_;
  assign new_n17708_ = ~new_n1989_ | ~new_n2415_;
  assign new_n17709_ = ~new_n17500_ | ~new_n17707_;
  assign new_n17710_ = ~new_n17565_ | ~new_n17529_;
  assign new_n17711_ = ~new_n17562_ | ~new_n17423_;
  assign new_n17712_ = ~new_n17572_ | ~new_n17384_;
  assign new_n17713_ = ~new_n17586_ | ~new_n17396_;
  assign new_n17714_ = ~new_n17589_ | ~new_n17538_;
  assign new_n17715_ = ~new_n17672_ | ~new_n17531_;
  assign new_n17716_ = ~new_n17656_ | ~new_n17534_;
  assign new_n17717_ = ~new_n17687_ | ~new_n17442_;
  assign new_n17718_ = ~new_n17640_ | ~new_n17439_;
  assign new_n17719_ = ~new_n17694_ | ~new_n17421_;
  assign new_n17720_ = ~new_n17703_ | ~new_n17530_;
  assign new_n17721_ = ~new_n17608_ | ~new_n17430_;
  assign new_n17722_ = ~new_n2944_ | ~new_n1981_;
  assign new_n17723_ = ~new_n17654_ | ~new_n17526_;
  assign new_n17724_ = ~new_n1984_ | ~new_n17653_;
  assign new_n17725_ = ~new_n2946_ | ~new_n17653_;
  assign new_n17726_ = ~new_n17659_ | ~new_n17654_ | ~new_n17526_;
  assign new_n17727_ = ~new_n17493_ | ~new_n17512_ | ~new_n17526_;
  assign new_n17728_ = ~new_n17655_ | ~new_n17659_;
  assign new_n17729_ = ~new_n2010_ | ~new_n17401_;
  assign new_n17730_ = ~new_n2412_ | ~new_n17400_;
  assign new_n17731_ = ~new_n17730_ | ~new_n17729_;
  assign new_n17732_ = ~new_n17710_ | ~new_n17402_;
  assign new_n17733_ = ~new_n17731_ | ~new_n17564_;
  assign new_n17734_ = ~new_n2011_ | ~new_n17398_;
  assign new_n17735_ = ~new_n2409_ | ~new_n17399_;
  assign new_n17736_ = ~new_n17735_ | ~new_n17734_;
  assign new_n17737_ = ~new_n17711_ | ~new_n17501_;
  assign new_n17738_ = ~new_n17561_ | ~new_n17736_;
  assign new_n17739_ = ~new_n1997_ | ~new_n17385_;
  assign new_n17740_ = ~new_n2406_ | ~new_n17383_;
  assign new_n17741_ = ~new_n1998_ | ~new_n17381_;
  assign new_n17742_ = ~new_n2403_ | ~new_n17382_;
  assign new_n17743_ = ~new_n17742_ | ~new_n17741_;
  assign new_n17744_ = ~new_n17712_ | ~new_n17403_;
  assign new_n17745_ = ~new_n17743_ | ~new_n17553_;
  assign new_n17746_ = ~new_n1994_ | ~new_n17397_;
  assign new_n17747_ = ~new_n2400_ | ~new_n17388_;
  assign new_n17748_ = ~new_n1987_ | ~new_n17386_;
  assign new_n17749_ = ~new_n2397_ | ~new_n17387_;
  assign new_n17750_ = ~new_n17749_ | ~new_n17748_;
  assign new_n17751_ = ~new_n17713_ | ~new_n17406_;
  assign new_n17752_ = ~new_n17750_ | ~new_n17579_;
  assign new_n17753_ = ~new_n1991_ | ~new_n17394_;
  assign new_n17754_ = ~new_n2394_ | ~new_n17395_;
  assign new_n17755_ = ~new_n17754_ | ~new_n17753_;
  assign new_n17756_ = ~new_n17714_ | ~new_n17502_;
  assign new_n17757_ = ~new_n17588_ | ~new_n17755_;
  assign new_n17758_ = ~new_n1995_ | ~new_n17389_;
  assign new_n17759_ = ~new_n2391_ | ~new_n17390_;
  assign new_n17760_ = ~new_n1982_ | ~new_n17504_;
  assign new_n17761_ = ~new_n2955_ | ~new_n17503_;
  assign new_n17762_ = ~new_n1982_ | ~new_n17504_;
  assign new_n17763_ = ~new_n2955_ | ~new_n17503_;
  assign new_n17764_ = ~new_n17763_ | ~new_n17762_;
  assign new_n17765_ = ~new_n17505_ | ~new_n17506_;
  assign new_n17766_ = ~new_n17663_ | ~new_n17764_;
  assign new_n17767_ = ~new_n1981_ | ~new_n17450_;
  assign new_n17768_ = ~new_n2944_ | ~new_n17449_;
  assign new_n17769_ = ~new_n1981_ | ~new_n17450_;
  assign new_n17770_ = ~new_n2944_ | ~new_n17449_;
  assign new_n17771_ = ~new_n17770_ | ~new_n17769_;
  assign new_n17772_ = ~new_n17507_ | ~new_n17508_;
  assign new_n17773_ = ~new_n17661_ | ~new_n17771_;
  assign new_n17774_ = ~new_n1980_ | ~new_n17408_;
  assign new_n17775_ = ~new_n2945_ | ~new_n17409_;
  assign new_n17776_ = ~new_n1980_ | ~new_n17408_;
  assign new_n17777_ = ~new_n2945_ | ~new_n17409_;
  assign new_n17778_ = ~new_n17777_ | ~new_n17776_;
  assign new_n17779_ = ~new_n17509_ | ~new_n17510_;
  assign new_n17780_ = ~new_n17658_ | ~new_n17778_;
  assign new_n17781_ = ~new_n1984_ | ~new_n17411_;
  assign new_n17782_ = ~new_n2946_ | ~new_n17410_;
  assign new_n17783_ = ~new_n1985_ | ~new_n17412_;
  assign new_n17784_ = ~new_n2947_ | ~new_n17413_;
  assign new_n17785_ = ~new_n17784_ | ~new_n17783_;
  assign new_n17786_ = ~new_n17715_ | ~new_n17451_;
  assign new_n17787_ = ~new_n17785_ | ~new_n17665_;
  assign new_n17788_ = ~new_n1992_ | ~new_n17414_;
  assign new_n17789_ = ~new_n2948_ | ~new_n17415_;
  assign new_n17790_ = ~new_n17789_ | ~new_n17788_;
  assign new_n17791_ = ~new_n17716_ | ~new_n17512_;
  assign new_n17792_ = ~new_n17652_ | ~new_n17790_;
  assign new_n17793_ = ~new_n1993_ | ~new_n17446_;
  assign new_n17794_ = ~new_n2949_ | ~new_n17447_;
  assign new_n17795_ = ~new_n1993_ | ~new_n17446_;
  assign new_n17796_ = ~new_n2949_ | ~new_n17447_;
  assign new_n17797_ = ~new_n17796_ | ~new_n17795_;
  assign new_n17798_ = ~new_n17513_ | ~new_n17514_;
  assign new_n17799_ = ~new_n17648_ | ~new_n17797_;
  assign new_n17800_ = ~new_n1988_ | ~new_n17444_;
  assign new_n17801_ = ~new_n2950_ | ~new_n17445_;
  assign new_n17802_ = ~new_n1988_ | ~new_n17444_;
  assign new_n17803_ = ~new_n2950_ | ~new_n17445_;
  assign new_n17804_ = ~new_n17803_ | ~new_n17802_;
  assign new_n17805_ = ~new_n17515_ | ~new_n17516_;
  assign new_n17806_ = ~new_n17644_ | ~new_n17804_;
  assign new_n17807_ = ~new_n2002_ | ~new_n17416_;
  assign new_n17808_ = ~new_n2951_ | ~new_n17417_;
  assign new_n17809_ = ~new_n2002_ | ~new_n17416_;
  assign new_n17810_ = ~new_n2951_ | ~new_n17417_;
  assign new_n17811_ = ~new_n17810_ | ~new_n17809_;
  assign new_n17812_ = ~new_n2003_ | ~new_n17443_;
  assign new_n17813_ = ~new_n2952_ | ~new_n17452_;
  assign new_n17814_ = ~new_n17540_ | ~new_n17519_;
  assign new_n17815_ = ~new_n17686_ | ~new_n17393_;
  assign new_n17816_ = ~new_n2008_ | ~new_n17440_;
  assign new_n17817_ = ~new_n2441_ | ~new_n17441_;
  assign new_n17818_ = ~new_n17817_ | ~new_n17816_;
  assign new_n17819_ = ~new_n17717_ | ~new_n17453_;
  assign new_n17820_ = ~new_n17818_ | ~new_n17674_;
  assign new_n17821_ = ~new_n2009_ | ~new_n17437_;
  assign new_n17822_ = ~new_n2439_ | ~new_n17438_;
  assign new_n17823_ = ~new_n17822_ | ~new_n17821_;
  assign new_n17824_ = ~new_n17718_ | ~new_n17520_;
  assign new_n17825_ = ~new_n17628_ | ~new_n17823_;
  assign new_n17826_ = ~new_n1996_ | ~new_n17422_;
  assign new_n17827_ = ~new_n2436_ | ~new_n17420_;
  assign new_n17828_ = ~new_n2000_ | ~new_n17418_;
  assign new_n17829_ = ~new_n2433_ | ~new_n17419_;
  assign new_n17830_ = ~new_n17829_ | ~new_n17828_;
  assign new_n17831_ = ~new_n17719_ | ~new_n17454_;
  assign new_n17832_ = ~new_n17830_ | ~new_n17620_;
  assign new_n17833_ = ~new_n2001_ | ~new_n17435_;
  assign new_n17834_ = ~new_n2430_ | ~new_n17436_;
  assign new_n17835_ = ~new_n2001_ | ~new_n17435_;
  assign new_n17836_ = ~new_n2430_ | ~new_n17436_;
  assign new_n17837_ = ~new_n17836_ | ~new_n17835_;
  assign new_n17838_ = ~new_n17521_ | ~new_n17522_;
  assign new_n17839_ = ~new_n17616_ | ~new_n17837_;
  assign new_n17840_ = ~new_n2006_ | ~new_n17433_;
  assign new_n17841_ = ~new_n2427_ | ~new_n17434_;
  assign new_n17842_ = ~new_n2006_ | ~new_n17433_;
  assign new_n17843_ = ~new_n2427_ | ~new_n17434_;
  assign new_n17844_ = ~new_n17843_ | ~new_n17842_;
  assign new_n17845_ = ~new_n17523_ | ~new_n17524_;
  assign new_n17846_ = ~new_n17612_ | ~new_n17844_;
  assign new_n17847_ = ~new_n2007_ | ~new_n17431_;
  assign new_n17848_ = ~new_n2424_ | ~new_n17432_;
  assign new_n17849_ = ~new_n1999_ | ~new_n17426_;
  assign new_n17850_ = ~new_n2421_ | ~new_n17427_;
  assign new_n17851_ = ~new_n17850_ | ~new_n17849_;
  assign new_n17852_ = ~new_n17720_ | ~new_n17455_;
  assign new_n17853_ = ~new_n17851_ | ~new_n17696_;
  assign new_n17854_ = ~new_n1990_ | ~new_n17428_;
  assign new_n17855_ = ~new_n2418_ | ~new_n17429_;
  assign new_n17856_ = ~new_n17855_ | ~new_n17854_;
  assign new_n17857_ = ~new_n17721_ | ~new_n17525_;
  assign new_n17858_ = ~new_n17602_ | ~new_n17856_;
  assign new_n17859_ = ~new_n1989_ | ~new_n17424_;
  assign new_n17860_ = ~new_n2415_ | ~new_n17425_;
  assign new_n17861_ = ~new_n2004_ | ~new_n17391_;
  assign new_n17862_ = ~new_n2383_ | ~new_n17392_;
  assign new_n17863_ = new_n18035_ & new_n18034_;
  assign new_n17864_ = new_n18036_ & new_n18037_;
  assign new_n17865_ = new_n18053_ & new_n18052_;
  assign new_n17866_ = new_n18093_ & new_n18092_;
  assign new_n17867_ = new_n18102_ & new_n18101_;
  assign new_n17868_ = new_n18120_ & new_n18119_;
  assign new_n17869_ = new_n18128_ & new_n18127_;
  assign new_n17870_ = new_n18207_ & new_n18204_;
  assign new_n17871_ = new_n18200_ & new_n18197_;
  assign new_n17872_ = new_n18191_ & new_n18188_;
  assign new_n17873_ = new_n18182_ & new_n18179_;
  assign new_n17874_ = new_n18176_ & new_n18174_;
  assign new_n17875_ = new_n18169_ & new_n18166_;
  assign new_n17876_ = new_n18091_ & new_n18088_;
  assign new_n17877_ = new_n18083_ & new_n18080_;
  assign new_n17878_ = new_n18069_ & new_n18066_;
  assign new_n17879_ = ~new_n2403_;
  assign new_n17880_ = ~new_n1998_;
  assign new_n17881_ = ~new_n1997_;
  assign new_n17882_ = ~new_n1998_ | ~new_n2403_;
  assign new_n17883_ = ~new_n2406_;
  assign new_n17884_ = ~new_n2397_;
  assign new_n17885_ = ~new_n1987_;
  assign new_n17886_ = ~new_n1994_;
  assign new_n17887_ = ~new_n2391_;
  assign new_n17888_ = ~new_n1995_;
  assign new_n17889_ = ~new_n2383_;
  assign new_n17890_ = ~new_n2004_;
  assign new_n17891_ = ~new_n2004_ | ~new_n2383_;
  assign new_n17892_ = ~new_n2394_;
  assign new_n17893_ = ~new_n1991_;
  assign new_n17894_ = ~new_n1987_ | ~new_n2397_;
  assign new_n17895_ = ~new_n2400_;
  assign new_n17896_ = ~new_n2409_;
  assign new_n17897_ = ~new_n2011_;
  assign new_n17898_ = ~new_n2010_;
  assign new_n17899_ = ~new_n2412_;
  assign new_n17900_ = ~new_n17921_ | ~new_n18061_;
  assign new_n17901_ = ~new_n17977_ | ~new_n18049_;
  assign new_n17902_ = ~new_n18038_ | ~new_n18039_;
  assign new_n17903_ = ~new_n2388_ | ~new_n2005_;
  assign new_n17904_ = ~new_n17981_ | ~new_n18075_;
  assign new_n17905_ = ~new_n18072_ | ~new_n18071_;
  assign new_n17906_ = ~new_n2945_;
  assign new_n17907_ = ~new_n1980_;
  assign new_n17908_ = ~new_n1984_;
  assign new_n17909_ = ~new_n2946_;
  assign new_n17910_ = ~new_n2947_;
  assign new_n17911_ = ~new_n1985_;
  assign new_n17912_ = ~new_n2948_;
  assign new_n17913_ = ~new_n1992_;
  assign new_n17914_ = ~new_n2951_;
  assign new_n17915_ = ~new_n2002_;
  assign new_n17916_ = ~new_n2433_;
  assign new_n17917_ = ~new_n2000_;
  assign new_n17918_ = ~new_n1996_;
  assign new_n17919_ = ~new_n2000_ | ~new_n2433_;
  assign new_n17920_ = ~new_n2436_;
  assign new_n17921_ = ~new_n2011_ | ~new_n2409_;
  assign new_n17922_ = ~new_n2415_;
  assign new_n17923_ = ~new_n1989_;
  assign new_n17924_ = ~new_n2421_;
  assign new_n17925_ = ~new_n1999_;
  assign new_n17926_ = ~new_n2418_;
  assign new_n17927_ = ~new_n1990_;
  assign new_n17928_ = ~new_n1990_ | ~new_n2418_;
  assign new_n17929_ = ~new_n2424_;
  assign new_n17930_ = ~new_n2007_;
  assign new_n17931_ = ~new_n2427_;
  assign new_n17932_ = ~new_n2006_;
  assign new_n17933_ = ~new_n2430_;
  assign new_n17934_ = ~new_n2001_;
  assign new_n17935_ = ~new_n2439_;
  assign new_n17936_ = ~new_n2009_;
  assign new_n17937_ = ~new_n2009_ | ~new_n2439_;
  assign new_n17938_ = ~new_n2441_;
  assign new_n17939_ = ~new_n2008_;
  assign new_n17940_ = ~new_n2008_ | ~new_n2441_;
  assign new_n17941_ = ~new_n2952_;
  assign new_n17942_ = ~new_n2950_;
  assign new_n17943_ = ~new_n1988_;
  assign new_n17944_ = ~new_n2949_;
  assign new_n17945_ = ~new_n1993_;
  assign new_n17946_ = ~new_n2946_ | ~new_n1984_;
  assign new_n17947_ = ~new_n1981_;
  assign new_n17948_ = ~new_n2944_;
  assign new_n17949_ = ~new_n18162_ | ~new_n18032_;
  assign new_n17950_ = ~new_n2003_;
  assign new_n17951_ = ~new_n17937_ | ~new_n18171_;
  assign new_n17952_ = ~new_n18117_ | ~new_n18116_;
  assign new_n17953_ = ~new_n17928_ | ~new_n18193_;
  assign new_n17954_ = ~new_n18313_ | ~new_n18312_;
  assign new_n17955_ = ~new_n18360_ | ~new_n18359_;
  assign new_n17956_ = ~new_n18231_ | ~new_n18230_;
  assign new_n17957_ = ~new_n18236_ | ~new_n18235_;
  assign new_n17958_ = ~new_n18243_ | ~new_n18242_;
  assign new_n17959_ = ~new_n18250_ | ~new_n18249_;
  assign new_n17960_ = ~new_n18255_ | ~new_n18254_;
  assign new_n17961_ = ~new_n18264_ | ~new_n18263_;
  assign new_n17962_ = ~new_n18271_ | ~new_n18270_;
  assign new_n17963_ = ~new_n18278_ | ~new_n18277_;
  assign new_n17964_ = ~new_n18285_ | ~new_n18284_;
  assign new_n17965_ = ~new_n18290_ | ~new_n18289_;
  assign new_n17966_ = ~new_n18297_ | ~new_n18296_;
  assign new_n17967_ = ~new_n18304_ | ~new_n18303_;
  assign new_n17968_ = ~new_n18318_ | ~new_n18317_;
  assign new_n17969_ = ~new_n18323_ | ~new_n18322_;
  assign new_n17970_ = ~new_n18330_ | ~new_n18329_;
  assign new_n17971_ = ~new_n18337_ | ~new_n18336_;
  assign new_n17972_ = ~new_n18344_ | ~new_n18343_;
  assign new_n17973_ = ~new_n18351_ | ~new_n18350_;
  assign new_n17974_ = ~new_n18356_ | ~new_n18355_;
  assign new_n17975_ = new_n2391_ & new_n1995_;
  assign new_n17976_ = new_n18045_ & new_n18043_;
  assign new_n17977_ = new_n18050_ & new_n18048_;
  assign new_n17978_ = new_n18057_ & new_n18056_;
  assign new_n17979_ = new_n17882_ & new_n18238_ & new_n18237_;
  assign new_n17980_ = new_n18068_ & new_n17865_;
  assign new_n17981_ = new_n18076_ & new_n18074_;
  assign new_n17982_ = new_n17894_ & new_n18245_ & new_n18244_;
  assign new_n17983_ = new_n18082_ & new_n17863_;
  assign new_n17984_ = new_n18090_ & new_n18037_;
  assign new_n17985_ = new_n18060_ & new_n17866_;
  assign new_n17986_ = new_n18095_ & new_n18027_;
  assign new_n17987_ = new_n18104_ & new_n18028_;
  assign new_n17988_ = new_n18124_ & new_n18123_;
  assign new_n17989_ = new_n17869_ & new_n18138_;
  assign new_n17990_ = new_n18141_ & new_n18136_;
  assign new_n17991_ = new_n18157_ & new_n18154_;
  assign new_n17992_ = new_n18224_ & new_n18158_;
  assign new_n17993_ = new_n18015_ & new_n18134_;
  assign new_n17994_ = new_n17919_ & new_n18325_ & new_n18324_;
  assign new_n17995_ = new_n18028_ & new_n18346_ & new_n18345_;
  assign new_n17996_ = new_n18199_ & new_n17867_;
  assign new_n17997_ = new_n18027_ & new_n18358_ & new_n18357_;
  assign new_n17998_ = new_n18206_ & new_n17866_;
  assign new_n17999_ = ~new_n17978_ | ~new_n18058_;
  assign new_n18000_ = ~new_n18073_ | ~new_n18085_;
  assign new_n18001_ = ~new_n1982_;
  assign new_n18002_ = ~new_n2955_;
  assign new_n18003_ = new_n18259_ & new_n18258_;
  assign new_n18004_ = ~new_n18220_ | ~new_n18160_ | ~new_n18025_;
  assign new_n18005_ = new_n18266_ & new_n18265_;
  assign new_n18006_ = ~new_n17992_ | ~new_n18226_ | ~new_n18225_;
  assign new_n18007_ = new_n18273_ & new_n18272_;
  assign new_n18008_ = ~new_n17946_ | ~new_n18221_ | ~new_n18155_;
  assign new_n18009_ = new_n18280_ & new_n18279_;
  assign new_n18010_ = ~new_n18149_ | ~new_n18148_;
  assign new_n18011_ = new_n18292_ & new_n18291_;
  assign new_n18012_ = ~new_n18145_ | ~new_n18144_;
  assign new_n18013_ = new_n18299_ & new_n18298_;
  assign new_n18014_ = ~new_n17990_ | ~new_n18140_;
  assign new_n18015_ = new_n18306_ & new_n18305_;
  assign new_n18016_ = new_n18311_ & new_n18310_;
  assign new_n18017_ = ~new_n17903_ | ~new_n18183_;
  assign new_n18018_ = ~new_n17988_ | ~new_n18125_;
  assign new_n18019_ = new_n18332_ & new_n18331_;
  assign new_n18020_ = ~new_n18113_ | ~new_n18112_;
  assign new_n18021_ = new_n18339_ & new_n18338_;
  assign new_n18022_ = ~new_n18109_ | ~new_n18108_;
  assign new_n18023_ = ~new_n18099_ | ~new_n18098_;
  assign new_n18024_ = ~new_n18223_ | ~new_n18222_;
  assign new_n18025_ = ~new_n1981_ | ~new_n18006_;
  assign new_n18026_ = ~new_n17894_;
  assign new_n18027_ = ~new_n2412_ | ~new_n2010_;
  assign new_n18028_ = ~new_n1999_ | ~new_n2421_;
  assign new_n18029_ = ~new_n1985_ | ~new_n2947_;
  assign new_n18030_ = ~new_n17928_;
  assign new_n18031_ = ~new_n17937_;
  assign new_n18032_ = ~new_n1992_ | ~new_n2948_;
  assign new_n18033_ = ~new_n17921_;
  assign new_n18034_ = new_n1994_ | new_n2400_;
  assign new_n18035_ = new_n1987_ | new_n2397_;
  assign new_n18036_ = new_n2394_ | new_n1991_;
  assign new_n18037_ = new_n2391_ | new_n1995_;
  assign new_n18038_ = ~new_n17891_;
  assign new_n18039_ = new_n2388_ | new_n2005_;
  assign new_n18040_ = ~new_n17902_;
  assign new_n18041_ = ~new_n17903_;
  assign new_n18042_ = ~new_n17902_ | ~new_n17903_;
  assign new_n18043_ = ~new_n17975_ | ~new_n18036_;
  assign new_n18044_ = ~new_n17864_ | ~new_n18042_;
  assign new_n18045_ = ~new_n1991_ | ~new_n2394_;
  assign new_n18046_ = ~new_n17976_ | ~new_n18044_;
  assign new_n18047_ = ~new_n17895_ | ~new_n17894_;
  assign new_n18048_ = ~new_n1994_ | ~new_n18047_;
  assign new_n18049_ = ~new_n17863_ | ~new_n18046_;
  assign new_n18050_ = ~new_n2400_ | ~new_n18026_;
  assign new_n18051_ = ~new_n17901_;
  assign new_n18052_ = new_n1997_ | new_n2406_;
  assign new_n18053_ = new_n1998_ | new_n2403_;
  assign new_n18054_ = ~new_n17882_;
  assign new_n18055_ = ~new_n17883_ | ~new_n17882_;
  assign new_n18056_ = ~new_n1997_ | ~new_n18055_;
  assign new_n18057_ = ~new_n2406_ | ~new_n18054_;
  assign new_n18058_ = ~new_n17865_ | ~new_n17901_;
  assign new_n18059_ = ~new_n17999_;
  assign new_n18060_ = new_n2409_ | new_n2011_;
  assign new_n18061_ = ~new_n18060_ | ~new_n17999_;
  assign new_n18062_ = ~new_n17900_;
  assign new_n18063_ = new_n2010_ | new_n2412_;
  assign new_n18064_ = new_n2403_ | new_n1998_;
  assign new_n18065_ = ~new_n18064_ | ~new_n17901_;
  assign new_n18066_ = ~new_n17979_ | ~new_n18065_;
  assign new_n18067_ = ~new_n18051_ | ~new_n17882_;
  assign new_n18068_ = ~new_n2406_ | ~new_n1997_;
  assign new_n18069_ = ~new_n17980_ | ~new_n18067_;
  assign new_n18070_ = new_n1998_ | new_n2403_;
  assign new_n18071_ = ~new_n18041_ | ~new_n18037_;
  assign new_n18072_ = ~new_n1995_ | ~new_n2391_;
  assign new_n18073_ = ~new_n17905_;
  assign new_n18074_ = ~new_n18040_ | ~new_n17864_;
  assign new_n18075_ = ~new_n17905_ | ~new_n18036_;
  assign new_n18076_ = ~new_n1991_ | ~new_n2394_;
  assign new_n18077_ = ~new_n17904_;
  assign new_n18078_ = new_n2397_ | new_n1987_;
  assign new_n18079_ = ~new_n18078_ | ~new_n17904_;
  assign new_n18080_ = ~new_n17982_ | ~new_n18079_;
  assign new_n18081_ = ~new_n18077_ | ~new_n17894_;
  assign new_n18082_ = ~new_n2400_ | ~new_n1994_;
  assign new_n18083_ = ~new_n17983_ | ~new_n18081_;
  assign new_n18084_ = new_n1987_ | new_n2397_;
  assign new_n18085_ = ~new_n18040_ | ~new_n18037_;
  assign new_n18086_ = ~new_n18000_;
  assign new_n18087_ = ~new_n1991_ | ~new_n2394_;
  assign new_n18088_ = ~new_n18256_ | ~new_n17902_ | ~new_n17903_ | ~new_n18257_;
  assign new_n18089_ = ~new_n17903_ | ~new_n17902_;
  assign new_n18090_ = ~new_n1995_ | ~new_n2391_;
  assign new_n18091_ = ~new_n17984_ | ~new_n18089_;
  assign new_n18092_ = new_n2010_ | new_n2412_;
  assign new_n18093_ = new_n1989_ | new_n2415_;
  assign new_n18094_ = ~new_n18033_ | ~new_n17866_;
  assign new_n18095_ = ~new_n1989_ | ~new_n2415_;
  assign new_n18096_ = ~new_n17986_ | ~new_n18094_;
  assign new_n18097_ = new_n2415_ | new_n1989_;
  assign new_n18098_ = ~new_n17985_ | ~new_n17999_;
  assign new_n18099_ = ~new_n18097_ | ~new_n18096_;
  assign new_n18100_ = ~new_n18023_;
  assign new_n18101_ = new_n2007_ | new_n2424_;
  assign new_n18102_ = new_n1999_ | new_n2421_;
  assign new_n18103_ = ~new_n18030_ | ~new_n17867_;
  assign new_n18104_ = ~new_n2007_ | ~new_n2424_;
  assign new_n18105_ = ~new_n17987_ | ~new_n18103_;
  assign new_n18106_ = new_n2418_ | new_n1990_;
  assign new_n18107_ = new_n2424_ | new_n2007_;
  assign new_n18108_ = ~new_n17867_ | ~new_n18106_ | ~new_n18023_;
  assign new_n18109_ = ~new_n18107_ | ~new_n18105_;
  assign new_n18110_ = ~new_n18022_;
  assign new_n18111_ = new_n2427_ | new_n2006_;
  assign new_n18112_ = ~new_n18111_ | ~new_n18022_;
  assign new_n18113_ = ~new_n2006_ | ~new_n2427_;
  assign new_n18114_ = ~new_n18020_;
  assign new_n18115_ = new_n2430_ | new_n2001_;
  assign new_n18116_ = ~new_n18115_ | ~new_n18020_;
  assign new_n18117_ = ~new_n2001_ | ~new_n2430_;
  assign new_n18118_ = ~new_n17952_;
  assign new_n18119_ = new_n1996_ | new_n2436_;
  assign new_n18120_ = new_n2000_ | new_n2433_;
  assign new_n18121_ = ~new_n17919_;
  assign new_n18122_ = ~new_n17920_ | ~new_n17919_;
  assign new_n18123_ = ~new_n1996_ | ~new_n18122_;
  assign new_n18124_ = ~new_n2436_ | ~new_n18121_;
  assign new_n18125_ = ~new_n17868_ | ~new_n17952_;
  assign new_n18126_ = ~new_n18018_;
  assign new_n18127_ = new_n2003_ | new_n2952_;
  assign new_n18128_ = new_n2008_ | new_n2441_;
  assign new_n18129_ = new_n2002_ | new_n2951_;
  assign new_n18130_ = ~new_n17940_;
  assign new_n18131_ = ~new_n2952_ | ~new_n18130_;
  assign new_n18132_ = ~new_n18131_ | ~new_n17950_;
  assign new_n18133_ = ~new_n17940_ | ~new_n17941_;
  assign new_n18134_ = ~new_n18133_ | ~new_n18132_;
  assign new_n18135_ = ~new_n18031_ | ~new_n17869_;
  assign new_n18136_ = ~new_n2002_ | ~new_n2951_;
  assign new_n18137_ = ~new_n18134_ | ~new_n18135_;
  assign new_n18138_ = new_n2439_ | new_n2009_;
  assign new_n18139_ = new_n2951_ | new_n2002_;
  assign new_n18140_ = ~new_n17989_ | ~new_n18129_ | ~new_n18018_;
  assign new_n18141_ = ~new_n18139_ | ~new_n18137_;
  assign new_n18142_ = ~new_n18014_;
  assign new_n18143_ = new_n2950_ | new_n1988_;
  assign new_n18144_ = ~new_n18143_ | ~new_n18014_;
  assign new_n18145_ = ~new_n1988_ | ~new_n2950_;
  assign new_n18146_ = ~new_n18012_;
  assign new_n18147_ = new_n2949_ | new_n1993_;
  assign new_n18148_ = ~new_n18147_ | ~new_n18012_;
  assign new_n18149_ = ~new_n1993_ | ~new_n2949_;
  assign new_n18150_ = ~new_n18010_;
  assign new_n18151_ = new_n1985_ | new_n2947_;
  assign new_n18152_ = ~new_n18032_ | ~new_n18029_;
  assign new_n18153_ = ~new_n17946_;
  assign new_n18154_ = new_n2948_ | new_n1992_;
  assign new_n18155_ = ~new_n18024_ | ~new_n18010_ | ~new_n18154_;
  assign new_n18156_ = ~new_n18008_;
  assign new_n18157_ = new_n2945_ | new_n1980_;
  assign new_n18158_ = ~new_n1980_ | ~new_n2945_;
  assign new_n18159_ = ~new_n18006_;
  assign new_n18160_ = ~new_n2944_ | ~new_n18006_;
  assign new_n18161_ = ~new_n18004_;
  assign new_n18162_ = ~new_n18154_ | ~new_n18010_;
  assign new_n18163_ = ~new_n17949_;
  assign new_n18164_ = new_n2947_ | new_n1985_;
  assign new_n18165_ = ~new_n18164_ | ~new_n17949_;
  assign new_n18166_ = ~new_n18009_ | ~new_n18165_ | ~new_n18029_;
  assign new_n18167_ = ~new_n18163_ | ~new_n18029_;
  assign new_n18168_ = ~new_n2946_ | ~new_n1984_;
  assign new_n18169_ = ~new_n18024_ | ~new_n18167_ | ~new_n18168_;
  assign new_n18170_ = new_n1985_ | new_n2947_;
  assign new_n18171_ = ~new_n18138_ | ~new_n18018_;
  assign new_n18172_ = ~new_n17951_;
  assign new_n18173_ = ~new_n17869_ | ~new_n17951_;
  assign new_n18174_ = ~new_n17993_ | ~new_n18173_;
  assign new_n18175_ = ~new_n18173_ | ~new_n18134_;
  assign new_n18176_ = ~new_n18309_ | ~new_n18175_;
  assign new_n18177_ = new_n2441_ | new_n2008_;
  assign new_n18178_ = ~new_n18177_ | ~new_n17951_;
  assign new_n18179_ = ~new_n18016_ | ~new_n18178_ | ~new_n17940_;
  assign new_n18180_ = ~new_n18172_ | ~new_n17940_;
  assign new_n18181_ = ~new_n2003_ | ~new_n2952_;
  assign new_n18182_ = ~new_n17869_ | ~new_n18181_ | ~new_n18180_;
  assign new_n18183_ = new_n2388_ | new_n2005_;
  assign new_n18184_ = ~new_n18017_;
  assign new_n18185_ = new_n2008_ | new_n2441_;
  assign new_n18186_ = new_n2433_ | new_n2000_;
  assign new_n18187_ = ~new_n18186_ | ~new_n17952_;
  assign new_n18188_ = ~new_n17994_ | ~new_n18187_;
  assign new_n18189_ = ~new_n18118_ | ~new_n17919_;
  assign new_n18190_ = ~new_n2436_ | ~new_n1996_;
  assign new_n18191_ = ~new_n17868_ | ~new_n18190_ | ~new_n18189_;
  assign new_n18192_ = new_n2000_ | new_n2433_;
  assign new_n18193_ = ~new_n18106_ | ~new_n18023_;
  assign new_n18194_ = ~new_n17953_;
  assign new_n18195_ = new_n2421_ | new_n1999_;
  assign new_n18196_ = ~new_n18195_ | ~new_n17953_;
  assign new_n18197_ = ~new_n17995_ | ~new_n18196_;
  assign new_n18198_ = ~new_n18194_ | ~new_n18028_;
  assign new_n18199_ = ~new_n2007_ | ~new_n2424_;
  assign new_n18200_ = ~new_n17996_ | ~new_n18198_;
  assign new_n18201_ = new_n1999_ | new_n2421_;
  assign new_n18202_ = new_n2412_ | new_n2010_;
  assign new_n18203_ = ~new_n18202_ | ~new_n17900_;
  assign new_n18204_ = ~new_n17997_ | ~new_n18203_;
  assign new_n18205_ = ~new_n18062_ | ~new_n18027_;
  assign new_n18206_ = ~new_n1989_ | ~new_n2415_;
  assign new_n18207_ = ~new_n17998_ | ~new_n18205_;
  assign new_n18208_ = ~new_n18063_ | ~new_n18027_;
  assign new_n18209_ = ~new_n18060_ | ~new_n17921_;
  assign new_n18210_ = ~new_n18070_ | ~new_n17882_;
  assign new_n18211_ = ~new_n18084_ | ~new_n17894_;
  assign new_n18212_ = ~new_n18087_ | ~new_n18036_;
  assign new_n18213_ = ~new_n18170_ | ~new_n18029_;
  assign new_n18214_ = ~new_n18154_ | ~new_n18032_;
  assign new_n18215_ = ~new_n18185_ | ~new_n17940_;
  assign new_n18216_ = ~new_n18138_ | ~new_n17937_;
  assign new_n18217_ = ~new_n18192_ | ~new_n17919_;
  assign new_n18218_ = ~new_n18201_ | ~new_n18028_;
  assign new_n18219_ = ~new_n18106_ | ~new_n17928_;
  assign new_n18220_ = ~new_n2944_ | ~new_n1981_;
  assign new_n18221_ = ~new_n18152_ | ~new_n18024_;
  assign new_n18222_ = ~new_n1984_ | ~new_n18151_;
  assign new_n18223_ = ~new_n2946_ | ~new_n18151_;
  assign new_n18224_ = ~new_n18157_ | ~new_n18152_ | ~new_n18024_;
  assign new_n18225_ = ~new_n17991_ | ~new_n18010_ | ~new_n18024_;
  assign new_n18226_ = ~new_n18153_ | ~new_n18157_;
  assign new_n18227_ = ~new_n2010_ | ~new_n17899_;
  assign new_n18228_ = ~new_n2412_ | ~new_n17898_;
  assign new_n18229_ = ~new_n18228_ | ~new_n18227_;
  assign new_n18230_ = ~new_n18208_ | ~new_n17900_;
  assign new_n18231_ = ~new_n18229_ | ~new_n18062_;
  assign new_n18232_ = ~new_n2011_ | ~new_n17896_;
  assign new_n18233_ = ~new_n2409_ | ~new_n17897_;
  assign new_n18234_ = ~new_n18233_ | ~new_n18232_;
  assign new_n18235_ = ~new_n18209_ | ~new_n17999_;
  assign new_n18236_ = ~new_n18059_ | ~new_n18234_;
  assign new_n18237_ = ~new_n1997_ | ~new_n17883_;
  assign new_n18238_ = ~new_n2406_ | ~new_n17881_;
  assign new_n18239_ = ~new_n1998_ | ~new_n17879_;
  assign new_n18240_ = ~new_n2403_ | ~new_n17880_;
  assign new_n18241_ = ~new_n18240_ | ~new_n18239_;
  assign new_n18242_ = ~new_n18210_ | ~new_n17901_;
  assign new_n18243_ = ~new_n18241_ | ~new_n18051_;
  assign new_n18244_ = ~new_n1994_ | ~new_n17895_;
  assign new_n18245_ = ~new_n2400_ | ~new_n17886_;
  assign new_n18246_ = ~new_n1987_ | ~new_n17884_;
  assign new_n18247_ = ~new_n2397_ | ~new_n17885_;
  assign new_n18248_ = ~new_n18247_ | ~new_n18246_;
  assign new_n18249_ = ~new_n18211_ | ~new_n17904_;
  assign new_n18250_ = ~new_n18248_ | ~new_n18077_;
  assign new_n18251_ = ~new_n1991_ | ~new_n17892_;
  assign new_n18252_ = ~new_n2394_ | ~new_n17893_;
  assign new_n18253_ = ~new_n18252_ | ~new_n18251_;
  assign new_n18254_ = ~new_n18212_ | ~new_n18000_;
  assign new_n18255_ = ~new_n18086_ | ~new_n18253_;
  assign new_n18256_ = ~new_n1995_ | ~new_n17887_;
  assign new_n18257_ = ~new_n2391_ | ~new_n17888_;
  assign new_n18258_ = ~new_n1982_ | ~new_n18002_;
  assign new_n18259_ = ~new_n2955_ | ~new_n18001_;
  assign new_n18260_ = ~new_n1982_ | ~new_n18002_;
  assign new_n18261_ = ~new_n2955_ | ~new_n18001_;
  assign new_n18262_ = ~new_n18261_ | ~new_n18260_;
  assign new_n18263_ = ~new_n18003_ | ~new_n18004_;
  assign new_n18264_ = ~new_n18161_ | ~new_n18262_;
  assign new_n18265_ = ~new_n1981_ | ~new_n17948_;
  assign new_n18266_ = ~new_n2944_ | ~new_n17947_;
  assign new_n18267_ = ~new_n1981_ | ~new_n17948_;
  assign new_n18268_ = ~new_n2944_ | ~new_n17947_;
  assign new_n18269_ = ~new_n18268_ | ~new_n18267_;
  assign new_n18270_ = ~new_n18005_ | ~new_n18006_;
  assign new_n18271_ = ~new_n18159_ | ~new_n18269_;
  assign new_n18272_ = ~new_n1980_ | ~new_n17906_;
  assign new_n18273_ = ~new_n2945_ | ~new_n17907_;
  assign new_n18274_ = ~new_n1980_ | ~new_n17906_;
  assign new_n18275_ = ~new_n2945_ | ~new_n17907_;
  assign new_n18276_ = ~new_n18275_ | ~new_n18274_;
  assign new_n18277_ = ~new_n18007_ | ~new_n18008_;
  assign new_n18278_ = ~new_n18156_ | ~new_n18276_;
  assign new_n18279_ = ~new_n1984_ | ~new_n17909_;
  assign new_n18280_ = ~new_n2946_ | ~new_n17908_;
  assign new_n18281_ = ~new_n1985_ | ~new_n17910_;
  assign new_n18282_ = ~new_n2947_ | ~new_n17911_;
  assign new_n18283_ = ~new_n18282_ | ~new_n18281_;
  assign new_n18284_ = ~new_n18213_ | ~new_n17949_;
  assign new_n18285_ = ~new_n18283_ | ~new_n18163_;
  assign new_n18286_ = ~new_n1992_ | ~new_n17912_;
  assign new_n18287_ = ~new_n2948_ | ~new_n17913_;
  assign new_n18288_ = ~new_n18287_ | ~new_n18286_;
  assign new_n18289_ = ~new_n18214_ | ~new_n18010_;
  assign new_n18290_ = ~new_n18150_ | ~new_n18288_;
  assign new_n18291_ = ~new_n1993_ | ~new_n17944_;
  assign new_n18292_ = ~new_n2949_ | ~new_n17945_;
  assign new_n18293_ = ~new_n1993_ | ~new_n17944_;
  assign new_n18294_ = ~new_n2949_ | ~new_n17945_;
  assign new_n18295_ = ~new_n18294_ | ~new_n18293_;
  assign new_n18296_ = ~new_n18011_ | ~new_n18012_;
  assign new_n18297_ = ~new_n18146_ | ~new_n18295_;
  assign new_n18298_ = ~new_n1988_ | ~new_n17942_;
  assign new_n18299_ = ~new_n2950_ | ~new_n17943_;
  assign new_n18300_ = ~new_n1988_ | ~new_n17942_;
  assign new_n18301_ = ~new_n2950_ | ~new_n17943_;
  assign new_n18302_ = ~new_n18301_ | ~new_n18300_;
  assign new_n18303_ = ~new_n18013_ | ~new_n18014_;
  assign new_n18304_ = ~new_n18142_ | ~new_n18302_;
  assign new_n18305_ = ~new_n2002_ | ~new_n17914_;
  assign new_n18306_ = ~new_n2951_ | ~new_n17915_;
  assign new_n18307_ = ~new_n2002_ | ~new_n17914_;
  assign new_n18308_ = ~new_n2951_ | ~new_n17915_;
  assign new_n18309_ = ~new_n18308_ | ~new_n18307_;
  assign new_n18310_ = ~new_n2003_ | ~new_n17941_;
  assign new_n18311_ = ~new_n2952_ | ~new_n17950_;
  assign new_n18312_ = ~new_n18038_ | ~new_n18017_;
  assign new_n18313_ = ~new_n18184_ | ~new_n17891_;
  assign new_n18314_ = ~new_n2008_ | ~new_n17938_;
  assign new_n18315_ = ~new_n2441_ | ~new_n17939_;
  assign new_n18316_ = ~new_n18315_ | ~new_n18314_;
  assign new_n18317_ = ~new_n18215_ | ~new_n17951_;
  assign new_n18318_ = ~new_n18316_ | ~new_n18172_;
  assign new_n18319_ = ~new_n2009_ | ~new_n17935_;
  assign new_n18320_ = ~new_n2439_ | ~new_n17936_;
  assign new_n18321_ = ~new_n18320_ | ~new_n18319_;
  assign new_n18322_ = ~new_n18216_ | ~new_n18018_;
  assign new_n18323_ = ~new_n18126_ | ~new_n18321_;
  assign new_n18324_ = ~new_n1996_ | ~new_n17920_;
  assign new_n18325_ = ~new_n2436_ | ~new_n17918_;
  assign new_n18326_ = ~new_n2000_ | ~new_n17916_;
  assign new_n18327_ = ~new_n2433_ | ~new_n17917_;
  assign new_n18328_ = ~new_n18327_ | ~new_n18326_;
  assign new_n18329_ = ~new_n18217_ | ~new_n17952_;
  assign new_n18330_ = ~new_n18328_ | ~new_n18118_;
  assign new_n18331_ = ~new_n2001_ | ~new_n17933_;
  assign new_n18332_ = ~new_n2430_ | ~new_n17934_;
  assign new_n18333_ = ~new_n2001_ | ~new_n17933_;
  assign new_n18334_ = ~new_n2430_ | ~new_n17934_;
  assign new_n18335_ = ~new_n18334_ | ~new_n18333_;
  assign new_n18336_ = ~new_n18019_ | ~new_n18020_;
  assign new_n18337_ = ~new_n18114_ | ~new_n18335_;
  assign new_n18338_ = ~new_n2006_ | ~new_n17931_;
  assign new_n18339_ = ~new_n2427_ | ~new_n17932_;
  assign new_n18340_ = ~new_n2006_ | ~new_n17931_;
  assign new_n18341_ = ~new_n2427_ | ~new_n17932_;
  assign new_n18342_ = ~new_n18341_ | ~new_n18340_;
  assign new_n18343_ = ~new_n18021_ | ~new_n18022_;
  assign new_n18344_ = ~new_n18110_ | ~new_n18342_;
  assign new_n18345_ = ~new_n2007_ | ~new_n17929_;
  assign new_n18346_ = ~new_n2424_ | ~new_n17930_;
  assign new_n18347_ = ~new_n1999_ | ~new_n17924_;
  assign new_n18348_ = ~new_n2421_ | ~new_n17925_;
  assign new_n18349_ = ~new_n18348_ | ~new_n18347_;
  assign new_n18350_ = ~new_n18218_ | ~new_n17953_;
  assign new_n18351_ = ~new_n18349_ | ~new_n18194_;
  assign new_n18352_ = ~new_n1990_ | ~new_n17926_;
  assign new_n18353_ = ~new_n2418_ | ~new_n17927_;
  assign new_n18354_ = ~new_n18353_ | ~new_n18352_;
  assign new_n18355_ = ~new_n18219_ | ~new_n18023_;
  assign new_n18356_ = ~new_n18100_ | ~new_n18354_;
  assign new_n18357_ = ~new_n1989_ | ~new_n17922_;
  assign new_n18358_ = ~new_n2415_ | ~new_n17923_;
  assign new_n18359_ = ~new_n2004_ | ~new_n17889_;
  assign new_n18360_ = ~new_n2383_ | ~new_n17890_;
  assign new_n18361_ = new_n18533_ & new_n18532_;
  assign new_n18362_ = new_n18534_ & new_n18535_;
  assign new_n18363_ = new_n18551_ & new_n18550_;
  assign new_n18364_ = new_n18591_ & new_n18590_;
  assign new_n18365_ = new_n18600_ & new_n18599_;
  assign new_n18366_ = new_n18618_ & new_n18617_;
  assign new_n18367_ = new_n18626_ & new_n18625_;
  assign new_n18368_ = new_n18705_ & new_n18702_;
  assign new_n18369_ = new_n18698_ & new_n18695_;
  assign new_n18370_ = new_n18689_ & new_n18686_;
  assign new_n18371_ = new_n18680_ & new_n18677_;
  assign new_n18372_ = new_n18674_ & new_n18672_;
  assign new_n18373_ = new_n18667_ & new_n18664_;
  assign new_n18374_ = new_n18589_ & new_n18586_;
  assign new_n18375_ = new_n18581_ & new_n18578_;
  assign new_n18376_ = new_n18567_ & new_n18564_;
  assign new_n18377_ = ~new_n2403_;
  assign new_n18378_ = ~new_n1998_;
  assign new_n18379_ = ~new_n1997_;
  assign new_n18380_ = ~new_n1998_ | ~new_n2403_;
  assign new_n18381_ = ~new_n2406_;
  assign new_n18382_ = ~new_n2397_;
  assign new_n18383_ = ~new_n1987_;
  assign new_n18384_ = ~new_n1994_;
  assign new_n18385_ = ~new_n2391_;
  assign new_n18386_ = ~new_n1995_;
  assign new_n18387_ = ~new_n2383_;
  assign new_n18388_ = ~new_n2004_;
  assign new_n18389_ = ~new_n2004_ | ~new_n2383_;
  assign new_n18390_ = ~new_n2394_;
  assign new_n18391_ = ~new_n1991_;
  assign new_n18392_ = ~new_n1987_ | ~new_n2397_;
  assign new_n18393_ = ~new_n2400_;
  assign new_n18394_ = ~new_n2409_;
  assign new_n18395_ = ~new_n2011_;
  assign new_n18396_ = ~new_n2010_;
  assign new_n18397_ = ~new_n2412_;
  assign new_n18398_ = ~new_n18419_ | ~new_n18559_;
  assign new_n18399_ = ~new_n18475_ | ~new_n18547_;
  assign new_n18400_ = ~new_n18536_ | ~new_n18537_;
  assign new_n18401_ = ~new_n2388_ | ~new_n2005_;
  assign new_n18402_ = ~new_n18479_ | ~new_n18573_;
  assign new_n18403_ = ~new_n18570_ | ~new_n18569_;
  assign new_n18404_ = ~new_n2945_;
  assign new_n18405_ = ~new_n1980_;
  assign new_n18406_ = ~new_n1984_;
  assign new_n18407_ = ~new_n2946_;
  assign new_n18408_ = ~new_n2947_;
  assign new_n18409_ = ~new_n1985_;
  assign new_n18410_ = ~new_n2948_;
  assign new_n18411_ = ~new_n1992_;
  assign new_n18412_ = ~new_n2951_;
  assign new_n18413_ = ~new_n2002_;
  assign new_n18414_ = ~new_n2433_;
  assign new_n18415_ = ~new_n2000_;
  assign new_n18416_ = ~new_n1996_;
  assign new_n18417_ = ~new_n2000_ | ~new_n2433_;
  assign new_n18418_ = ~new_n2436_;
  assign new_n18419_ = ~new_n2011_ | ~new_n2409_;
  assign new_n18420_ = ~new_n2415_;
  assign new_n18421_ = ~new_n1989_;
  assign new_n18422_ = ~new_n2421_;
  assign new_n18423_ = ~new_n1999_;
  assign new_n18424_ = ~new_n2418_;
  assign new_n18425_ = ~new_n1990_;
  assign new_n18426_ = ~new_n1990_ | ~new_n2418_;
  assign new_n18427_ = ~new_n2424_;
  assign new_n18428_ = ~new_n2007_;
  assign new_n18429_ = ~new_n2427_;
  assign new_n18430_ = ~new_n2006_;
  assign new_n18431_ = ~new_n2430_;
  assign new_n18432_ = ~new_n2001_;
  assign new_n18433_ = ~new_n2439_;
  assign new_n18434_ = ~new_n2009_;
  assign new_n18435_ = ~new_n2009_ | ~new_n2439_;
  assign new_n18436_ = ~new_n2441_;
  assign new_n18437_ = ~new_n2008_;
  assign new_n18438_ = ~new_n2008_ | ~new_n2441_;
  assign new_n18439_ = ~new_n2952_;
  assign new_n18440_ = ~new_n2950_;
  assign new_n18441_ = ~new_n1988_;
  assign new_n18442_ = ~new_n2949_;
  assign new_n18443_ = ~new_n1993_;
  assign new_n18444_ = ~new_n2946_ | ~new_n1984_;
  assign new_n18445_ = ~new_n1981_;
  assign new_n18446_ = ~new_n2944_;
  assign new_n18447_ = ~new_n18660_ | ~new_n18530_;
  assign new_n18448_ = ~new_n2003_;
  assign new_n18449_ = ~new_n18435_ | ~new_n18669_;
  assign new_n18450_ = ~new_n18615_ | ~new_n18614_;
  assign new_n18451_ = ~new_n18426_ | ~new_n18691_;
  assign new_n18452_ = ~new_n18811_ | ~new_n18810_;
  assign new_n18453_ = ~new_n18858_ | ~new_n18857_;
  assign new_n18454_ = ~new_n18729_ | ~new_n18728_;
  assign new_n18455_ = ~new_n18734_ | ~new_n18733_;
  assign new_n18456_ = ~new_n18741_ | ~new_n18740_;
  assign new_n18457_ = ~new_n18748_ | ~new_n18747_;
  assign new_n18458_ = ~new_n18753_ | ~new_n18752_;
  assign new_n18459_ = ~new_n18762_ | ~new_n18761_;
  assign new_n18460_ = ~new_n18769_ | ~new_n18768_;
  assign new_n18461_ = ~new_n18776_ | ~new_n18775_;
  assign new_n18462_ = ~new_n18783_ | ~new_n18782_;
  assign new_n18463_ = ~new_n18788_ | ~new_n18787_;
  assign new_n18464_ = ~new_n18795_ | ~new_n18794_;
  assign new_n18465_ = ~new_n18802_ | ~new_n18801_;
  assign new_n18466_ = ~new_n18816_ | ~new_n18815_;
  assign new_n18467_ = ~new_n18821_ | ~new_n18820_;
  assign new_n18468_ = ~new_n18828_ | ~new_n18827_;
  assign new_n18469_ = ~new_n18835_ | ~new_n18834_;
  assign new_n18470_ = ~new_n18842_ | ~new_n18841_;
  assign new_n18471_ = ~new_n18849_ | ~new_n18848_;
  assign new_n18472_ = ~new_n18854_ | ~new_n18853_;
  assign new_n18473_ = new_n2391_ & new_n1995_;
  assign new_n18474_ = new_n18543_ & new_n18541_;
  assign new_n18475_ = new_n18548_ & new_n18546_;
  assign new_n18476_ = new_n18555_ & new_n18554_;
  assign new_n18477_ = new_n18380_ & new_n18736_ & new_n18735_;
  assign new_n18478_ = new_n18566_ & new_n18363_;
  assign new_n18479_ = new_n18574_ & new_n18572_;
  assign new_n18480_ = new_n18392_ & new_n18743_ & new_n18742_;
  assign new_n18481_ = new_n18580_ & new_n18361_;
  assign new_n18482_ = new_n18588_ & new_n18535_;
  assign new_n18483_ = new_n18558_ & new_n18364_;
  assign new_n18484_ = new_n18593_ & new_n18525_;
  assign new_n18485_ = new_n18602_ & new_n18526_;
  assign new_n18486_ = new_n18622_ & new_n18621_;
  assign new_n18487_ = new_n18367_ & new_n18636_;
  assign new_n18488_ = new_n18639_ & new_n18634_;
  assign new_n18489_ = new_n18655_ & new_n18652_;
  assign new_n18490_ = new_n18722_ & new_n18656_;
  assign new_n18491_ = new_n18513_ & new_n18632_;
  assign new_n18492_ = new_n18417_ & new_n18823_ & new_n18822_;
  assign new_n18493_ = new_n18526_ & new_n18844_ & new_n18843_;
  assign new_n18494_ = new_n18697_ & new_n18365_;
  assign new_n18495_ = new_n18525_ & new_n18856_ & new_n18855_;
  assign new_n18496_ = new_n18704_ & new_n18364_;
  assign new_n18497_ = ~new_n18476_ | ~new_n18556_;
  assign new_n18498_ = ~new_n18571_ | ~new_n18583_;
  assign new_n18499_ = ~new_n1982_;
  assign new_n18500_ = ~new_n2955_;
  assign new_n18501_ = new_n18757_ & new_n18756_;
  assign new_n18502_ = ~new_n18718_ | ~new_n18658_ | ~new_n18523_;
  assign new_n18503_ = new_n18764_ & new_n18763_;
  assign new_n18504_ = ~new_n18490_ | ~new_n18724_ | ~new_n18723_;
  assign new_n18505_ = new_n18771_ & new_n18770_;
  assign new_n18506_ = ~new_n18444_ | ~new_n18719_ | ~new_n18653_;
  assign new_n18507_ = new_n18778_ & new_n18777_;
  assign new_n18508_ = ~new_n18647_ | ~new_n18646_;
  assign new_n18509_ = new_n18790_ & new_n18789_;
  assign new_n18510_ = ~new_n18643_ | ~new_n18642_;
  assign new_n18511_ = new_n18797_ & new_n18796_;
  assign new_n18512_ = ~new_n18488_ | ~new_n18638_;
  assign new_n18513_ = new_n18804_ & new_n18803_;
  assign new_n18514_ = new_n18809_ & new_n18808_;
  assign new_n18515_ = ~new_n18401_ | ~new_n18681_;
  assign new_n18516_ = ~new_n18486_ | ~new_n18623_;
  assign new_n18517_ = new_n18830_ & new_n18829_;
  assign new_n18518_ = ~new_n18611_ | ~new_n18610_;
  assign new_n18519_ = new_n18837_ & new_n18836_;
  assign new_n18520_ = ~new_n18607_ | ~new_n18606_;
  assign new_n18521_ = ~new_n18597_ | ~new_n18596_;
  assign new_n18522_ = ~new_n18721_ | ~new_n18720_;
  assign new_n18523_ = ~new_n1981_ | ~new_n18504_;
  assign new_n18524_ = ~new_n18392_;
  assign new_n18525_ = ~new_n2412_ | ~new_n2010_;
  assign new_n18526_ = ~new_n1999_ | ~new_n2421_;
  assign new_n18527_ = ~new_n1985_ | ~new_n2947_;
  assign new_n18528_ = ~new_n18426_;
  assign new_n18529_ = ~new_n18435_;
  assign new_n18530_ = ~new_n1992_ | ~new_n2948_;
  assign new_n18531_ = ~new_n18419_;
  assign new_n18532_ = new_n1994_ | new_n2400_;
  assign new_n18533_ = new_n1987_ | new_n2397_;
  assign new_n18534_ = new_n2394_ | new_n1991_;
  assign new_n18535_ = new_n2391_ | new_n1995_;
  assign new_n18536_ = ~new_n18389_;
  assign new_n18537_ = new_n2388_ | new_n2005_;
  assign new_n18538_ = ~new_n18400_;
  assign new_n18539_ = ~new_n18401_;
  assign new_n18540_ = ~new_n18400_ | ~new_n18401_;
  assign new_n18541_ = ~new_n18473_ | ~new_n18534_;
  assign new_n18542_ = ~new_n18362_ | ~new_n18540_;
  assign new_n18543_ = ~new_n1991_ | ~new_n2394_;
  assign new_n18544_ = ~new_n18474_ | ~new_n18542_;
  assign new_n18545_ = ~new_n18393_ | ~new_n18392_;
  assign new_n18546_ = ~new_n1994_ | ~new_n18545_;
  assign new_n18547_ = ~new_n18361_ | ~new_n18544_;
  assign new_n18548_ = ~new_n2400_ | ~new_n18524_;
  assign new_n18549_ = ~new_n18399_;
  assign new_n18550_ = new_n1997_ | new_n2406_;
  assign new_n18551_ = new_n1998_ | new_n2403_;
  assign new_n18552_ = ~new_n18380_;
  assign new_n18553_ = ~new_n18381_ | ~new_n18380_;
  assign new_n18554_ = ~new_n1997_ | ~new_n18553_;
  assign new_n18555_ = ~new_n2406_ | ~new_n18552_;
  assign new_n18556_ = ~new_n18363_ | ~new_n18399_;
  assign new_n18557_ = ~new_n18497_;
  assign new_n18558_ = new_n2409_ | new_n2011_;
  assign new_n18559_ = ~new_n18558_ | ~new_n18497_;
  assign new_n18560_ = ~new_n18398_;
  assign new_n18561_ = new_n2010_ | new_n2412_;
  assign new_n18562_ = new_n2403_ | new_n1998_;
  assign new_n18563_ = ~new_n18562_ | ~new_n18399_;
  assign new_n18564_ = ~new_n18477_ | ~new_n18563_;
  assign new_n18565_ = ~new_n18549_ | ~new_n18380_;
  assign new_n18566_ = ~new_n2406_ | ~new_n1997_;
  assign new_n18567_ = ~new_n18478_ | ~new_n18565_;
  assign new_n18568_ = new_n1998_ | new_n2403_;
  assign new_n18569_ = ~new_n18539_ | ~new_n18535_;
  assign new_n18570_ = ~new_n1995_ | ~new_n2391_;
  assign new_n18571_ = ~new_n18403_;
  assign new_n18572_ = ~new_n18538_ | ~new_n18362_;
  assign new_n18573_ = ~new_n18403_ | ~new_n18534_;
  assign new_n18574_ = ~new_n1991_ | ~new_n2394_;
  assign new_n18575_ = ~new_n18402_;
  assign new_n18576_ = new_n2397_ | new_n1987_;
  assign new_n18577_ = ~new_n18576_ | ~new_n18402_;
  assign new_n18578_ = ~new_n18480_ | ~new_n18577_;
  assign new_n18579_ = ~new_n18575_ | ~new_n18392_;
  assign new_n18580_ = ~new_n2400_ | ~new_n1994_;
  assign new_n18581_ = ~new_n18481_ | ~new_n18579_;
  assign new_n18582_ = new_n1987_ | new_n2397_;
  assign new_n18583_ = ~new_n18538_ | ~new_n18535_;
  assign new_n18584_ = ~new_n18498_;
  assign new_n18585_ = ~new_n1991_ | ~new_n2394_;
  assign new_n18586_ = ~new_n18754_ | ~new_n18400_ | ~new_n18401_ | ~new_n18755_;
  assign new_n18587_ = ~new_n18401_ | ~new_n18400_;
  assign new_n18588_ = ~new_n1995_ | ~new_n2391_;
  assign new_n18589_ = ~new_n18482_ | ~new_n18587_;
  assign new_n18590_ = new_n2010_ | new_n2412_;
  assign new_n18591_ = new_n1989_ | new_n2415_;
  assign new_n18592_ = ~new_n18531_ | ~new_n18364_;
  assign new_n18593_ = ~new_n1989_ | ~new_n2415_;
  assign new_n18594_ = ~new_n18484_ | ~new_n18592_;
  assign new_n18595_ = new_n2415_ | new_n1989_;
  assign new_n18596_ = ~new_n18483_ | ~new_n18497_;
  assign new_n18597_ = ~new_n18595_ | ~new_n18594_;
  assign new_n18598_ = ~new_n18521_;
  assign new_n18599_ = new_n2007_ | new_n2424_;
  assign new_n18600_ = new_n1999_ | new_n2421_;
  assign new_n18601_ = ~new_n18528_ | ~new_n18365_;
  assign new_n18602_ = ~new_n2007_ | ~new_n2424_;
  assign new_n18603_ = ~new_n18485_ | ~new_n18601_;
  assign new_n18604_ = new_n2418_ | new_n1990_;
  assign new_n18605_ = new_n2424_ | new_n2007_;
  assign new_n18606_ = ~new_n18365_ | ~new_n18604_ | ~new_n18521_;
  assign new_n18607_ = ~new_n18605_ | ~new_n18603_;
  assign new_n18608_ = ~new_n18520_;
  assign new_n18609_ = new_n2427_ | new_n2006_;
  assign new_n18610_ = ~new_n18609_ | ~new_n18520_;
  assign new_n18611_ = ~new_n2006_ | ~new_n2427_;
  assign new_n18612_ = ~new_n18518_;
  assign new_n18613_ = new_n2430_ | new_n2001_;
  assign new_n18614_ = ~new_n18613_ | ~new_n18518_;
  assign new_n18615_ = ~new_n2001_ | ~new_n2430_;
  assign new_n18616_ = ~new_n18450_;
  assign new_n18617_ = new_n1996_ | new_n2436_;
  assign new_n18618_ = new_n2000_ | new_n2433_;
  assign new_n18619_ = ~new_n18417_;
  assign new_n18620_ = ~new_n18418_ | ~new_n18417_;
  assign new_n18621_ = ~new_n1996_ | ~new_n18620_;
  assign new_n18622_ = ~new_n2436_ | ~new_n18619_;
  assign new_n18623_ = ~new_n18366_ | ~new_n18450_;
  assign new_n18624_ = ~new_n18516_;
  assign new_n18625_ = new_n2003_ | new_n2952_;
  assign new_n18626_ = new_n2008_ | new_n2441_;
  assign new_n18627_ = new_n2002_ | new_n2951_;
  assign new_n18628_ = ~new_n18438_;
  assign new_n18629_ = ~new_n2952_ | ~new_n18628_;
  assign new_n18630_ = ~new_n18629_ | ~new_n18448_;
  assign new_n18631_ = ~new_n18438_ | ~new_n18439_;
  assign new_n18632_ = ~new_n18631_ | ~new_n18630_;
  assign new_n18633_ = ~new_n18529_ | ~new_n18367_;
  assign new_n18634_ = ~new_n2002_ | ~new_n2951_;
  assign new_n18635_ = ~new_n18632_ | ~new_n18633_;
  assign new_n18636_ = new_n2439_ | new_n2009_;
  assign new_n18637_ = new_n2951_ | new_n2002_;
  assign new_n18638_ = ~new_n18487_ | ~new_n18627_ | ~new_n18516_;
  assign new_n18639_ = ~new_n18637_ | ~new_n18635_;
  assign new_n18640_ = ~new_n18512_;
  assign new_n18641_ = new_n2950_ | new_n1988_;
  assign new_n18642_ = ~new_n18641_ | ~new_n18512_;
  assign new_n18643_ = ~new_n1988_ | ~new_n2950_;
  assign new_n18644_ = ~new_n18510_;
  assign new_n18645_ = new_n2949_ | new_n1993_;
  assign new_n18646_ = ~new_n18645_ | ~new_n18510_;
  assign new_n18647_ = ~new_n1993_ | ~new_n2949_;
  assign new_n18648_ = ~new_n18508_;
  assign new_n18649_ = new_n1985_ | new_n2947_;
  assign new_n18650_ = ~new_n18530_ | ~new_n18527_;
  assign new_n18651_ = ~new_n18444_;
  assign new_n18652_ = new_n2948_ | new_n1992_;
  assign new_n18653_ = ~new_n18522_ | ~new_n18508_ | ~new_n18652_;
  assign new_n18654_ = ~new_n18506_;
  assign new_n18655_ = new_n2945_ | new_n1980_;
  assign new_n18656_ = ~new_n1980_ | ~new_n2945_;
  assign new_n18657_ = ~new_n18504_;
  assign new_n18658_ = ~new_n2944_ | ~new_n18504_;
  assign new_n18659_ = ~new_n18502_;
  assign new_n18660_ = ~new_n18652_ | ~new_n18508_;
  assign new_n18661_ = ~new_n18447_;
  assign new_n18662_ = new_n2947_ | new_n1985_;
  assign new_n18663_ = ~new_n18662_ | ~new_n18447_;
  assign new_n18664_ = ~new_n18507_ | ~new_n18663_ | ~new_n18527_;
  assign new_n18665_ = ~new_n18661_ | ~new_n18527_;
  assign new_n18666_ = ~new_n2946_ | ~new_n1984_;
  assign new_n18667_ = ~new_n18522_ | ~new_n18665_ | ~new_n18666_;
  assign new_n18668_ = new_n1985_ | new_n2947_;
  assign new_n18669_ = ~new_n18636_ | ~new_n18516_;
  assign new_n18670_ = ~new_n18449_;
  assign new_n18671_ = ~new_n18367_ | ~new_n18449_;
  assign new_n18672_ = ~new_n18491_ | ~new_n18671_;
  assign new_n18673_ = ~new_n18671_ | ~new_n18632_;
  assign new_n18674_ = ~new_n18807_ | ~new_n18673_;
  assign new_n18675_ = new_n2441_ | new_n2008_;
  assign new_n18676_ = ~new_n18675_ | ~new_n18449_;
  assign new_n18677_ = ~new_n18514_ | ~new_n18676_ | ~new_n18438_;
  assign new_n18678_ = ~new_n18670_ | ~new_n18438_;
  assign new_n18679_ = ~new_n2003_ | ~new_n2952_;
  assign new_n18680_ = ~new_n18367_ | ~new_n18679_ | ~new_n18678_;
  assign new_n18681_ = new_n2388_ | new_n2005_;
  assign new_n18682_ = ~new_n18515_;
  assign new_n18683_ = new_n2008_ | new_n2441_;
  assign new_n18684_ = new_n2433_ | new_n2000_;
  assign new_n18685_ = ~new_n18684_ | ~new_n18450_;
  assign new_n18686_ = ~new_n18492_ | ~new_n18685_;
  assign new_n18687_ = ~new_n18616_ | ~new_n18417_;
  assign new_n18688_ = ~new_n2436_ | ~new_n1996_;
  assign new_n18689_ = ~new_n18366_ | ~new_n18688_ | ~new_n18687_;
  assign new_n18690_ = new_n2000_ | new_n2433_;
  assign new_n18691_ = ~new_n18604_ | ~new_n18521_;
  assign new_n18692_ = ~new_n18451_;
  assign new_n18693_ = new_n2421_ | new_n1999_;
  assign new_n18694_ = ~new_n18693_ | ~new_n18451_;
  assign new_n18695_ = ~new_n18493_ | ~new_n18694_;
  assign new_n18696_ = ~new_n18692_ | ~new_n18526_;
  assign new_n18697_ = ~new_n2007_ | ~new_n2424_;
  assign new_n18698_ = ~new_n18494_ | ~new_n18696_;
  assign new_n18699_ = new_n1999_ | new_n2421_;
  assign new_n18700_ = new_n2412_ | new_n2010_;
  assign new_n18701_ = ~new_n18700_ | ~new_n18398_;
  assign new_n18702_ = ~new_n18495_ | ~new_n18701_;
  assign new_n18703_ = ~new_n18560_ | ~new_n18525_;
  assign new_n18704_ = ~new_n1989_ | ~new_n2415_;
  assign new_n18705_ = ~new_n18496_ | ~new_n18703_;
  assign new_n18706_ = ~new_n18561_ | ~new_n18525_;
  assign new_n18707_ = ~new_n18558_ | ~new_n18419_;
  assign new_n18708_ = ~new_n18568_ | ~new_n18380_;
  assign new_n18709_ = ~new_n18582_ | ~new_n18392_;
  assign new_n18710_ = ~new_n18585_ | ~new_n18534_;
  assign new_n18711_ = ~new_n18668_ | ~new_n18527_;
  assign new_n18712_ = ~new_n18652_ | ~new_n18530_;
  assign new_n18713_ = ~new_n18683_ | ~new_n18438_;
  assign new_n18714_ = ~new_n18636_ | ~new_n18435_;
  assign new_n18715_ = ~new_n18690_ | ~new_n18417_;
  assign new_n18716_ = ~new_n18699_ | ~new_n18526_;
  assign new_n18717_ = ~new_n18604_ | ~new_n18426_;
  assign new_n18718_ = ~new_n2944_ | ~new_n1981_;
  assign new_n18719_ = ~new_n18650_ | ~new_n18522_;
  assign new_n18720_ = ~new_n1984_ | ~new_n18649_;
  assign new_n18721_ = ~new_n2946_ | ~new_n18649_;
  assign new_n18722_ = ~new_n18655_ | ~new_n18650_ | ~new_n18522_;
  assign new_n18723_ = ~new_n18489_ | ~new_n18508_ | ~new_n18522_;
  assign new_n18724_ = ~new_n18651_ | ~new_n18655_;
  assign new_n18725_ = ~new_n2010_ | ~new_n18397_;
  assign new_n18726_ = ~new_n2412_ | ~new_n18396_;
  assign new_n18727_ = ~new_n18726_ | ~new_n18725_;
  assign new_n18728_ = ~new_n18706_ | ~new_n18398_;
  assign new_n18729_ = ~new_n18727_ | ~new_n18560_;
  assign new_n18730_ = ~new_n2011_ | ~new_n18394_;
  assign new_n18731_ = ~new_n2409_ | ~new_n18395_;
  assign new_n18732_ = ~new_n18731_ | ~new_n18730_;
  assign new_n18733_ = ~new_n18707_ | ~new_n18497_;
  assign new_n18734_ = ~new_n18557_ | ~new_n18732_;
  assign new_n18735_ = ~new_n1997_ | ~new_n18381_;
  assign new_n18736_ = ~new_n2406_ | ~new_n18379_;
  assign new_n18737_ = ~new_n1998_ | ~new_n18377_;
  assign new_n18738_ = ~new_n2403_ | ~new_n18378_;
  assign new_n18739_ = ~new_n18738_ | ~new_n18737_;
  assign new_n18740_ = ~new_n18708_ | ~new_n18399_;
  assign new_n18741_ = ~new_n18739_ | ~new_n18549_;
  assign new_n18742_ = ~new_n1994_ | ~new_n18393_;
  assign new_n18743_ = ~new_n2400_ | ~new_n18384_;
  assign new_n18744_ = ~new_n1987_ | ~new_n18382_;
  assign new_n18745_ = ~new_n2397_ | ~new_n18383_;
  assign new_n18746_ = ~new_n18745_ | ~new_n18744_;
  assign new_n18747_ = ~new_n18709_ | ~new_n18402_;
  assign new_n18748_ = ~new_n18746_ | ~new_n18575_;
  assign new_n18749_ = ~new_n1991_ | ~new_n18390_;
  assign new_n18750_ = ~new_n2394_ | ~new_n18391_;
  assign new_n18751_ = ~new_n18750_ | ~new_n18749_;
  assign new_n18752_ = ~new_n18710_ | ~new_n18498_;
  assign new_n18753_ = ~new_n18584_ | ~new_n18751_;
  assign new_n18754_ = ~new_n1995_ | ~new_n18385_;
  assign new_n18755_ = ~new_n2391_ | ~new_n18386_;
  assign new_n18756_ = ~new_n1982_ | ~new_n18500_;
  assign new_n18757_ = ~new_n2955_ | ~new_n18499_;
  assign new_n18758_ = ~new_n1982_ | ~new_n18500_;
  assign new_n18759_ = ~new_n2955_ | ~new_n18499_;
  assign new_n18760_ = ~new_n18759_ | ~new_n18758_;
  assign new_n18761_ = ~new_n18501_ | ~new_n18502_;
  assign new_n18762_ = ~new_n18659_ | ~new_n18760_;
  assign new_n18763_ = ~new_n1981_ | ~new_n18446_;
  assign new_n18764_ = ~new_n2944_ | ~new_n18445_;
  assign new_n18765_ = ~new_n1981_ | ~new_n18446_;
  assign new_n18766_ = ~new_n2944_ | ~new_n18445_;
  assign new_n18767_ = ~new_n18766_ | ~new_n18765_;
  assign new_n18768_ = ~new_n18503_ | ~new_n18504_;
  assign new_n18769_ = ~new_n18657_ | ~new_n18767_;
  assign new_n18770_ = ~new_n1980_ | ~new_n18404_;
  assign new_n18771_ = ~new_n2945_ | ~new_n18405_;
  assign new_n18772_ = ~new_n1980_ | ~new_n18404_;
  assign new_n18773_ = ~new_n2945_ | ~new_n18405_;
  assign new_n18774_ = ~new_n18773_ | ~new_n18772_;
  assign new_n18775_ = ~new_n18505_ | ~new_n18506_;
  assign new_n18776_ = ~new_n18654_ | ~new_n18774_;
  assign new_n18777_ = ~new_n1984_ | ~new_n18407_;
  assign new_n18778_ = ~new_n2946_ | ~new_n18406_;
  assign new_n18779_ = ~new_n1985_ | ~new_n18408_;
  assign new_n18780_ = ~new_n2947_ | ~new_n18409_;
  assign new_n18781_ = ~new_n18780_ | ~new_n18779_;
  assign new_n18782_ = ~new_n18711_ | ~new_n18447_;
  assign new_n18783_ = ~new_n18781_ | ~new_n18661_;
  assign new_n18784_ = ~new_n1992_ | ~new_n18410_;
  assign new_n18785_ = ~new_n2948_ | ~new_n18411_;
  assign new_n18786_ = ~new_n18785_ | ~new_n18784_;
  assign new_n18787_ = ~new_n18712_ | ~new_n18508_;
  assign new_n18788_ = ~new_n18648_ | ~new_n18786_;
  assign new_n18789_ = ~new_n1993_ | ~new_n18442_;
  assign new_n18790_ = ~new_n2949_ | ~new_n18443_;
  assign new_n18791_ = ~new_n1993_ | ~new_n18442_;
  assign new_n18792_ = ~new_n2949_ | ~new_n18443_;
  assign new_n18793_ = ~new_n18792_ | ~new_n18791_;
  assign new_n18794_ = ~new_n18509_ | ~new_n18510_;
  assign new_n18795_ = ~new_n18644_ | ~new_n18793_;
  assign new_n18796_ = ~new_n1988_ | ~new_n18440_;
  assign new_n18797_ = ~new_n2950_ | ~new_n18441_;
  assign new_n18798_ = ~new_n1988_ | ~new_n18440_;
  assign new_n18799_ = ~new_n2950_ | ~new_n18441_;
  assign new_n18800_ = ~new_n18799_ | ~new_n18798_;
  assign new_n18801_ = ~new_n18511_ | ~new_n18512_;
  assign new_n18802_ = ~new_n18640_ | ~new_n18800_;
  assign new_n18803_ = ~new_n2002_ | ~new_n18412_;
  assign new_n18804_ = ~new_n2951_ | ~new_n18413_;
  assign new_n18805_ = ~new_n2002_ | ~new_n18412_;
  assign new_n18806_ = ~new_n2951_ | ~new_n18413_;
  assign new_n18807_ = ~new_n18806_ | ~new_n18805_;
  assign new_n18808_ = ~new_n2003_ | ~new_n18439_;
  assign new_n18809_ = ~new_n2952_ | ~new_n18448_;
  assign new_n18810_ = ~new_n18536_ | ~new_n18515_;
  assign new_n18811_ = ~new_n18682_ | ~new_n18389_;
  assign new_n18812_ = ~new_n2008_ | ~new_n18436_;
  assign new_n18813_ = ~new_n2441_ | ~new_n18437_;
  assign new_n18814_ = ~new_n18813_ | ~new_n18812_;
  assign new_n18815_ = ~new_n18713_ | ~new_n18449_;
  assign new_n18816_ = ~new_n18814_ | ~new_n18670_;
  assign new_n18817_ = ~new_n2009_ | ~new_n18433_;
  assign new_n18818_ = ~new_n2439_ | ~new_n18434_;
  assign new_n18819_ = ~new_n18818_ | ~new_n18817_;
  assign new_n18820_ = ~new_n18714_ | ~new_n18516_;
  assign new_n18821_ = ~new_n18624_ | ~new_n18819_;
  assign new_n18822_ = ~new_n1996_ | ~new_n18418_;
  assign new_n18823_ = ~new_n2436_ | ~new_n18416_;
  assign new_n18824_ = ~new_n2000_ | ~new_n18414_;
  assign new_n18825_ = ~new_n2433_ | ~new_n18415_;
  assign new_n18826_ = ~new_n18825_ | ~new_n18824_;
  assign new_n18827_ = ~new_n18715_ | ~new_n18450_;
  assign new_n18828_ = ~new_n18826_ | ~new_n18616_;
  assign new_n18829_ = ~new_n2001_ | ~new_n18431_;
  assign new_n18830_ = ~new_n2430_ | ~new_n18432_;
  assign new_n18831_ = ~new_n2001_ | ~new_n18431_;
  assign new_n18832_ = ~new_n2430_ | ~new_n18432_;
  assign new_n18833_ = ~new_n18832_ | ~new_n18831_;
  assign new_n18834_ = ~new_n18517_ | ~new_n18518_;
  assign new_n18835_ = ~new_n18612_ | ~new_n18833_;
  assign new_n18836_ = ~new_n2006_ | ~new_n18429_;
  assign new_n18837_ = ~new_n2427_ | ~new_n18430_;
  assign new_n18838_ = ~new_n2006_ | ~new_n18429_;
  assign new_n18839_ = ~new_n2427_ | ~new_n18430_;
  assign new_n18840_ = ~new_n18839_ | ~new_n18838_;
  assign new_n18841_ = ~new_n18519_ | ~new_n18520_;
  assign new_n18842_ = ~new_n18608_ | ~new_n18840_;
  assign new_n18843_ = ~new_n2007_ | ~new_n18427_;
  assign new_n18844_ = ~new_n2424_ | ~new_n18428_;
  assign new_n18845_ = ~new_n1999_ | ~new_n18422_;
  assign new_n18846_ = ~new_n2421_ | ~new_n18423_;
  assign new_n18847_ = ~new_n18846_ | ~new_n18845_;
  assign new_n18848_ = ~new_n18716_ | ~new_n18451_;
  assign new_n18849_ = ~new_n18847_ | ~new_n18692_;
  assign new_n18850_ = ~new_n1990_ | ~new_n18424_;
  assign new_n18851_ = ~new_n2418_ | ~new_n18425_;
  assign new_n18852_ = ~new_n18851_ | ~new_n18850_;
  assign new_n18853_ = ~new_n18717_ | ~new_n18521_;
  assign new_n18854_ = ~new_n18598_ | ~new_n18852_;
  assign new_n18855_ = ~new_n1989_ | ~new_n18420_;
  assign new_n18856_ = ~new_n2415_ | ~new_n18421_;
  assign new_n18857_ = ~new_n2004_ | ~new_n18387_;
  assign new_n18858_ = ~new_n2383_ | ~new_n18388_;
  assign new_n18859_ = ~pi514;
  assign new_n18860_ = new_n18933_ & new_n18961_;
  assign new_n18861_ = ~pi505;
  assign new_n18862_ = ~pi502;
  assign new_n18863_ = ~pi502 | ~pi505 | ~pi514;
  assign new_n18864_ = ~pi519;
  assign new_n18865_ = ~pi493;
  assign new_n18866_ = ~new_n18930_ | ~new_n18940_;
  assign new_n18867_ = ~pi511;
  assign new_n18868_ = ~pi501;
  assign new_n18869_ = ~new_n18931_ | ~new_n18942_;
  assign new_n18870_ = ~pi496;
  assign new_n18871_ = ~pi515;
  assign new_n18872_ = ~new_n18932_ | ~new_n18944_;
  assign new_n18873_ = ~pi508;
  assign new_n18874_ = ~pi508 | ~new_n18946_;
  assign new_n18875_ = ~pi498;
  assign new_n18876_ = ~pi498 | ~new_n18947_;
  assign new_n18877_ = ~pi517;
  assign new_n18878_ = ~pi517 | ~new_n18948_;
  assign new_n18879_ = ~pi491;
  assign new_n18880_ = ~pi491 | ~new_n18949_;
  assign new_n18881_ = ~pi506;
  assign new_n18882_ = ~pi506 | ~new_n18950_;
  assign new_n18883_ = ~pi504;
  assign new_n18884_ = ~pi504 | ~new_n18951_;
  assign new_n18885_ = ~pi494;
  assign new_n18886_ = ~pi494 | ~new_n18952_;
  assign new_n18887_ = ~pi513;
  assign new_n18888_ = ~pi513 | ~new_n18953_;
  assign new_n18889_ = ~pi499;
  assign new_n18890_ = ~pi499 | ~new_n18954_;
  assign new_n18891_ = ~pi509;
  assign new_n18892_ = ~pi509 | ~new_n18955_;
  assign new_n18893_ = ~pi497;
  assign new_n18894_ = ~pi497 | ~new_n18956_;
  assign new_n18895_ = ~pi516;
  assign new_n18896_ = ~pi516 | ~new_n18957_;
  assign new_n18897_ = ~pi503;
  assign new_n18898_ = ~pi503 | ~new_n18958_;
  assign new_n18899_ = ~pi507;
  assign new_n18900_ = ~pi507 | ~new_n18959_;
  assign new_n18901_ = ~pi492;
  assign new_n18902_ = ~pi492 | ~new_n18960_;
  assign new_n18903_ = ~pi512;
  assign new_n18904_ = ~pi518;
  assign new_n18905_ = ~new_n18964_ | ~new_n18963_;
  assign new_n18906_ = ~new_n18966_ | ~new_n18965_;
  assign new_n18907_ = ~new_n18968_ | ~new_n18967_;
  assign new_n18908_ = ~new_n18970_ | ~new_n18969_;
  assign new_n18909_ = ~new_n18972_ | ~new_n18971_;
  assign new_n18910_ = ~new_n18974_ | ~new_n18973_;
  assign new_n18911_ = ~new_n18976_ | ~new_n18975_;
  assign new_n18912_ = ~new_n18978_ | ~new_n18977_;
  assign new_n18913_ = ~new_n18980_ | ~new_n18979_;
  assign new_n18914_ = ~new_n18982_ | ~new_n18981_;
  assign new_n18915_ = ~new_n18984_ | ~new_n18983_;
  assign new_n18916_ = ~new_n18986_ | ~new_n18985_;
  assign new_n18917_ = ~new_n18988_ | ~new_n18987_;
  assign new_n18918_ = ~new_n18990_ | ~new_n18989_;
  assign new_n18919_ = ~new_n18992_ | ~new_n18991_;
  assign new_n18920_ = ~new_n18994_ | ~new_n18993_;
  assign new_n18921_ = ~new_n18996_ | ~new_n18995_;
  assign new_n18922_ = ~new_n18998_ | ~new_n18997_;
  assign new_n18923_ = ~new_n19000_ | ~new_n18999_;
  assign new_n18924_ = ~new_n19002_ | ~new_n19001_;
  assign new_n18925_ = ~new_n19004_ | ~new_n19003_;
  assign new_n18926_ = ~new_n19006_ | ~new_n19005_;
  assign new_n18927_ = ~new_n19008_ | ~new_n19007_;
  assign new_n18928_ = ~new_n19010_ | ~new_n19009_;
  assign new_n18929_ = ~new_n19012_ | ~new_n19011_;
  assign new_n18930_ = pi519 & pi493;
  assign new_n18931_ = pi511 & pi501;
  assign new_n18932_ = pi496 & pi515;
  assign new_n18933_ = pi512 & pi518;
  assign new_n18934_ = ~pi511 | ~new_n18942_;
  assign new_n18935_ = ~pi493 | ~new_n18940_;
  assign new_n18936_ = ~pi502 | ~pi514;
  assign new_n18937_ = ~pi518 | ~new_n18961_;
  assign new_n18938_ = ~pi515 | ~new_n18944_;
  assign new_n18939_ = ~new_n18936_;
  assign new_n18940_ = ~new_n18863_;
  assign new_n18941_ = ~new_n18935_;
  assign new_n18942_ = ~new_n18866_;
  assign new_n18943_ = ~new_n18934_;
  assign new_n18944_ = ~new_n18869_;
  assign new_n18945_ = ~new_n18938_;
  assign new_n18946_ = ~new_n18872_;
  assign new_n18947_ = ~new_n18874_;
  assign new_n18948_ = ~new_n18876_;
  assign new_n18949_ = ~new_n18878_;
  assign new_n18950_ = ~new_n18880_;
  assign new_n18951_ = ~new_n18882_;
  assign new_n18952_ = ~new_n18884_;
  assign new_n18953_ = ~new_n18886_;
  assign new_n18954_ = ~new_n18888_;
  assign new_n18955_ = ~new_n18890_;
  assign new_n18956_ = ~new_n18892_;
  assign new_n18957_ = ~new_n18894_;
  assign new_n18958_ = ~new_n18896_;
  assign new_n18959_ = ~new_n18898_;
  assign new_n18960_ = ~new_n18900_;
  assign new_n18961_ = ~new_n18902_;
  assign new_n18962_ = ~new_n18937_;
  assign new_n18963_ = ~pi501 | ~new_n18934_;
  assign new_n18964_ = ~new_n18943_ | ~new_n18868_;
  assign new_n18965_ = ~pi511 | ~new_n18866_;
  assign new_n18966_ = ~new_n18942_ | ~new_n18867_;
  assign new_n18967_ = ~pi519 | ~new_n18935_;
  assign new_n18968_ = ~new_n18941_ | ~new_n18864_;
  assign new_n18969_ = ~pi493 | ~new_n18863_;
  assign new_n18970_ = ~new_n18940_ | ~new_n18865_;
  assign new_n18971_ = ~pi505 | ~new_n18936_;
  assign new_n18972_ = ~new_n18939_ | ~new_n18861_;
  assign new_n18973_ = ~pi502 | ~new_n18859_;
  assign new_n18974_ = ~pi514 | ~new_n18862_;
  assign new_n18975_ = ~pi512 | ~new_n18937_;
  assign new_n18976_ = ~new_n18962_ | ~new_n18903_;
  assign new_n18977_ = ~pi518 | ~new_n18902_;
  assign new_n18978_ = ~new_n18961_ | ~new_n18904_;
  assign new_n18979_ = ~pi492 | ~new_n18900_;
  assign new_n18980_ = ~new_n18960_ | ~new_n18901_;
  assign new_n18981_ = ~pi507 | ~new_n18898_;
  assign new_n18982_ = ~new_n18959_ | ~new_n18899_;
  assign new_n18983_ = ~pi503 | ~new_n18896_;
  assign new_n18984_ = ~new_n18958_ | ~new_n18897_;
  assign new_n18985_ = ~pi516 | ~new_n18894_;
  assign new_n18986_ = ~new_n18957_ | ~new_n18895_;
  assign new_n18987_ = ~pi497 | ~new_n18892_;
  assign new_n18988_ = ~new_n18956_ | ~new_n18893_;
  assign new_n18989_ = ~pi509 | ~new_n18890_;
  assign new_n18990_ = ~new_n18955_ | ~new_n18891_;
  assign new_n18991_ = ~pi499 | ~new_n18888_;
  assign new_n18992_ = ~new_n18954_ | ~new_n18889_;
  assign new_n18993_ = ~pi513 | ~new_n18886_;
  assign new_n18994_ = ~new_n18953_ | ~new_n18887_;
  assign new_n18995_ = ~pi494 | ~new_n18884_;
  assign new_n18996_ = ~new_n18952_ | ~new_n18885_;
  assign new_n18997_ = ~pi504 | ~new_n18882_;
  assign new_n18998_ = ~new_n18951_ | ~new_n18883_;
  assign new_n18999_ = ~pi506 | ~new_n18880_;
  assign new_n19000_ = ~new_n18950_ | ~new_n18881_;
  assign new_n19001_ = ~pi491 | ~new_n18878_;
  assign new_n19002_ = ~new_n18949_ | ~new_n18879_;
  assign new_n19003_ = ~pi517 | ~new_n18876_;
  assign new_n19004_ = ~new_n18948_ | ~new_n18877_;
  assign new_n19005_ = ~pi498 | ~new_n18874_;
  assign new_n19006_ = ~new_n18947_ | ~new_n18875_;
  assign new_n19007_ = ~pi508 | ~new_n18872_;
  assign new_n19008_ = ~new_n18946_ | ~new_n18873_;
  assign new_n19009_ = ~pi496 | ~new_n18938_;
  assign new_n19010_ = ~new_n18945_ | ~new_n18870_;
  assign new_n19011_ = ~pi515 | ~new_n18869_;
  assign new_n19012_ = ~new_n18944_ | ~new_n18871_;
  assign new_n19013_ = new_n19179_ & new_n19047_;
  assign new_n19014_ = new_n19177_ & new_n19147_;
  assign new_n19015_ = new_n19176_ & new_n19044_;
  assign new_n19016_ = new_n19175_ & new_n19045_;
  assign new_n19017_ = new_n19173_ & new_n19150_;
  assign new_n19018_ = new_n19172_ & new_n19037_;
  assign new_n19019_ = new_n19171_ & new_n19043_;
  assign new_n19020_ = new_n19169_ & new_n19039_;
  assign new_n19021_ = new_n19167_ & new_n19040_;
  assign new_n19022_ = new_n19166_ & new_n19116_;
  assign new_n19023_ = new_n19164_ & new_n19036_;
  assign new_n19024_ = new_n19162_ & new_n19030_;
  assign new_n19025_ = new_n19145_ & new_n19135_;
  assign new_n19026_ = new_n19144_ & new_n19032_;
  assign new_n19027_ = new_n19143_ & new_n19033_;
  assign new_n19028_ = new_n19141_ & new_n19138_;
  assign new_n19029_ = new_n19140_ & new_n19031_;
  assign new_n19030_ = pi280 | pi279 | pi278;
  assign new_n19031_ = ~new_n19051_ | ~new_n19052_ | ~new_n19181_;
  assign new_n19032_ = ~new_n19053_ | ~new_n19181_;
  assign new_n19033_ = ~new_n19054_ | ~new_n19136_;
  assign new_n19034_ = ~pi285;
  assign new_n19035_ = ~pi281;
  assign new_n19036_ = ~new_n19064_ | ~new_n19059_;
  assign new_n19037_ = ~new_n19097_ | ~new_n19095_ | ~new_n19096_ | ~new_n19098_;
  assign new_n19038_ = ~new_n19099_ | ~new_n19151_;
  assign new_n19039_ = ~new_n19100_ | ~new_n19154_;
  assign new_n19040_ = ~new_n19156_ | ~new_n19041_;
  assign new_n19041_ = ~pi302;
  assign new_n19042_ = ~new_n19154_ | ~new_n19122_;
  assign new_n19043_ = ~new_n19101_ | ~new_n19151_;
  assign new_n19044_ = ~new_n19102_ | ~new_n19139_;
  assign new_n19045_ = ~new_n19103_ | ~new_n19148_;
  assign new_n19046_ = ~pi293;
  assign new_n19047_ = ~new_n19104_ | ~new_n19139_;
  assign new_n19048_ = ~pi289;
  assign new_n19049_ = ~new_n19203_ | ~new_n19202_;
  assign new_n19050_ = ~new_n19187_ | ~new_n19186_;
  assign new_n19051_ = ~pi282 & ~pi284 & ~pi283 & ~pi281;
  assign new_n19052_ = ~pi285 & ~pi286;
  assign new_n19053_ = ~pi281 & ~pi282;
  assign new_n19054_ = ~pi283 & ~pi284;
  assign new_n19055_ = ~pi289 & ~pi291 & ~pi290 & ~pi288;
  assign new_n19056_ = ~pi293 & ~pi295 & ~pi294 & ~pi292;
  assign new_n19057_ = ~pi297 & ~pi278 & ~pi279 & ~pi296;
  assign new_n19058_ = ~pi299 & ~pi300 & ~pi298;
  assign new_n19059_ = new_n19057_ & new_n19055_ & new_n19056_ & new_n19058_;
  assign new_n19060_ = ~pi302 & ~pi304 & ~pi303 & ~pi301;
  assign new_n19061_ = ~pi306 & ~pi280 & ~pi307 & ~pi305;
  assign new_n19062_ = ~pi282 & ~pi284 & ~pi283 & ~pi281;
  assign new_n19063_ = ~pi286 & ~pi287 & ~pi285;
  assign new_n19064_ = new_n19062_ & new_n19060_ & new_n19061_ & new_n19063_;
  assign new_n19065_ = ~pi289 & ~pi291 & ~pi290 & ~pi288;
  assign new_n19066_ = ~pi293 & ~pi295 & ~pi294 & ~pi292;
  assign new_n19067_ = ~pi297 & ~pi278 & ~pi279 & ~pi296;
  assign new_n19068_ = ~pi299 & ~pi300 & ~pi298;
  assign new_n19069_ = new_n19067_ & new_n19065_ & new_n19066_ & new_n19068_;
  assign new_n19070_ = ~pi302 & ~pi304 & ~pi303 & ~pi301;
  assign new_n19071_ = ~pi306 & ~pi280 & ~pi305;
  assign new_n19072_ = ~pi282 & ~pi284 & ~pi283 & ~pi281;
  assign new_n19073_ = ~pi286 & ~pi287 & ~pi285;
  assign new_n19074_ = new_n19072_ & new_n19070_ & new_n19071_ & new_n19073_;
  assign new_n19075_ = ~pi289 & ~pi291 & ~pi290 & ~pi288;
  assign new_n19076_ = ~pi293 & ~pi294 & ~pi292;
  assign new_n19077_ = ~pi296 & ~pi279 & ~pi297 & ~pi295;
  assign new_n19078_ = ~pi298 & ~pi299 & ~pi278;
  assign new_n19079_ = new_n19077_ & new_n19075_ & new_n19076_ & new_n19078_;
  assign new_n19080_ = ~pi301 & ~pi303 & ~pi302 & ~pi300;
  assign new_n19081_ = ~pi305 & ~pi280 & ~pi304;
  assign new_n19082_ = ~pi282 & ~pi284 & ~pi283 & ~pi281;
  assign new_n19083_ = ~pi286 & ~pi287 & ~pi285;
  assign new_n19084_ = new_n19082_ & new_n19080_ & new_n19081_ & new_n19083_;
  assign new_n19085_ = ~pi289 & ~pi291 & ~pi290 & ~pi288;
  assign new_n19086_ = ~pi293 & ~pi294 & ~pi292;
  assign new_n19087_ = ~pi296 & ~pi279 & ~pi297 & ~pi295;
  assign new_n19088_ = ~pi298 & ~pi299 & ~pi278;
  assign new_n19089_ = new_n19087_ & new_n19085_ & new_n19086_ & new_n19088_;
  assign new_n19090_ = ~pi301 & ~pi303 & ~pi302 & ~pi300;
  assign new_n19091_ = ~pi280 & ~pi281 & ~pi304;
  assign new_n19092_ = ~pi283 & ~pi284 & ~pi282;
  assign new_n19093_ = ~pi286 & ~pi287 & ~pi285;
  assign new_n19094_ = new_n19092_ & new_n19090_ & new_n19091_ & new_n19093_;
  assign new_n19095_ = ~pi292 & ~pi291 & ~pi289 & ~pi288 & ~pi290;
  assign new_n19096_ = ~pi294 & ~pi278 & ~pi279 & ~pi293;
  assign new_n19097_ = ~pi281 & ~pi283 & ~pi282 & ~pi280;
  assign new_n19098_ = ~pi285 & ~pi287 & ~pi286 & ~pi284;
  assign new_n19099_ = ~pi296 & ~pi298 & ~pi297 & ~pi295;
  assign new_n19100_ = ~pi300 & ~pi301 & ~pi299;
  assign new_n19101_ = ~pi295 & ~pi296;
  assign new_n19102_ = ~pi289 & ~pi287 & ~pi290 & ~pi288;
  assign new_n19103_ = ~pi291 & ~pi292;
  assign new_n19104_ = ~pi288 & ~pi287;
  assign new_n19105_ = ~pi287;
  assign new_n19106_ = new_n19183_ & new_n19182_;
  assign new_n19107_ = ~pi283;
  assign new_n19108_ = new_n19185_ & new_n19184_;
  assign new_n19109_ = ~pi309;
  assign new_n19110_ = ~pi308;
  assign new_n19111_ = new_n19189_ & new_n19188_;
  assign new_n19112_ = ~pi306;
  assign new_n19113_ = ~new_n19084_ | ~new_n19079_;
  assign new_n19114_ = new_n19191_ & new_n19190_;
  assign new_n19115_ = ~pi305;
  assign new_n19116_ = ~new_n19094_ | ~new_n19089_;
  assign new_n19117_ = new_n19193_ & new_n19192_;
  assign new_n19118_ = ~pi303;
  assign new_n19119_ = new_n19195_ & new_n19194_;
  assign new_n19120_ = ~pi300;
  assign new_n19121_ = new_n19197_ & new_n19196_;
  assign new_n19122_ = ~pi299;
  assign new_n19123_ = new_n19199_ & new_n19198_;
  assign new_n19124_ = ~pi298;
  assign new_n19125_ = ~new_n19152_ | ~new_n19129_;
  assign new_n19126_ = new_n19201_ & new_n19200_;
  assign new_n19127_ = ~pi279;
  assign new_n19128_ = ~pi278;
  assign new_n19129_ = ~pi297;
  assign new_n19130_ = new_n19205_ & new_n19204_;
  assign new_n19131_ = ~pi295;
  assign new_n19132_ = new_n19207_ & new_n19206_;
  assign new_n19133_ = ~pi291;
  assign new_n19134_ = new_n19209_ & new_n19208_;
  assign new_n19135_ = ~new_n19181_ | ~new_n19035_;
  assign new_n19136_ = ~new_n19032_;
  assign new_n19137_ = ~new_n19033_;
  assign new_n19138_ = ~new_n19137_ | ~new_n19034_;
  assign new_n19139_ = ~new_n19031_;
  assign new_n19140_ = ~pi286 | ~new_n19138_;
  assign new_n19141_ = ~pi285 | ~new_n19033_;
  assign new_n19142_ = ~new_n19136_ | ~new_n19107_;
  assign new_n19143_ = ~pi284 | ~new_n19142_;
  assign new_n19144_ = ~pi282 | ~new_n19135_;
  assign new_n19145_ = ~pi281 | ~new_n19030_;
  assign new_n19146_ = ~new_n19047_;
  assign new_n19147_ = ~new_n19146_ | ~new_n19048_;
  assign new_n19148_ = ~new_n19044_;
  assign new_n19149_ = ~new_n19045_;
  assign new_n19150_ = ~new_n19149_ | ~new_n19046_;
  assign new_n19151_ = ~new_n19037_;
  assign new_n19152_ = ~new_n19043_;
  assign new_n19153_ = ~new_n19125_;
  assign new_n19154_ = ~new_n19038_;
  assign new_n19155_ = ~new_n19042_;
  assign new_n19156_ = ~new_n19039_;
  assign new_n19157_ = ~new_n19040_;
  assign new_n19158_ = ~new_n19116_;
  assign new_n19159_ = ~new_n19113_;
  assign new_n19160_ = ~new_n19036_;
  assign new_n19161_ = pi279 | pi278;
  assign new_n19162_ = ~pi280 | ~new_n19161_;
  assign new_n19163_ = ~new_n19074_ | ~new_n19069_;
  assign new_n19164_ = ~pi307 | ~new_n19163_;
  assign new_n19165_ = ~new_n19157_ | ~new_n19118_;
  assign new_n19166_ = ~pi304 | ~new_n19165_;
  assign new_n19167_ = ~pi302 | ~new_n19039_;
  assign new_n19168_ = ~new_n19155_ | ~new_n19120_;
  assign new_n19169_ = ~pi301 | ~new_n19168_;
  assign new_n19170_ = ~new_n19151_ | ~new_n19131_;
  assign new_n19171_ = ~pi296 | ~new_n19170_;
  assign new_n19172_ = ~pi294 | ~new_n19150_;
  assign new_n19173_ = ~pi293 | ~new_n19045_;
  assign new_n19174_ = ~new_n19148_ | ~new_n19133_;
  assign new_n19175_ = ~pi292 | ~new_n19174_;
  assign new_n19176_ = ~pi290 | ~new_n19147_;
  assign new_n19177_ = ~pi289 | ~new_n19047_;
  assign new_n19178_ = ~new_n19139_ | ~new_n19105_;
  assign new_n19179_ = ~pi288 | ~new_n19178_;
  assign new_n19180_ = ~new_n19160_ | ~new_n19110_;
  assign new_n19181_ = ~new_n19030_;
  assign new_n19182_ = ~pi287 | ~new_n19031_;
  assign new_n19183_ = ~new_n19139_ | ~new_n19105_;
  assign new_n19184_ = ~pi283 | ~new_n19032_;
  assign new_n19185_ = ~new_n19136_ | ~new_n19107_;
  assign new_n19186_ = ~new_n19180_ | ~new_n19109_;
  assign new_n19187_ = ~pi309 | ~new_n19160_ | ~new_n19110_;
  assign new_n19188_ = ~pi308 | ~new_n19036_;
  assign new_n19189_ = ~new_n19160_ | ~new_n19110_;
  assign new_n19190_ = ~pi306 | ~new_n19113_;
  assign new_n19191_ = ~new_n19159_ | ~new_n19112_;
  assign new_n19192_ = ~pi305 | ~new_n19116_;
  assign new_n19193_ = ~new_n19158_ | ~new_n19115_;
  assign new_n19194_ = ~pi303 | ~new_n19040_;
  assign new_n19195_ = ~new_n19157_ | ~new_n19118_;
  assign new_n19196_ = ~pi300 | ~new_n19042_;
  assign new_n19197_ = ~new_n19155_ | ~new_n19120_;
  assign new_n19198_ = ~pi299 | ~new_n19038_;
  assign new_n19199_ = ~new_n19154_ | ~new_n19122_;
  assign new_n19200_ = ~pi298 | ~new_n19125_;
  assign new_n19201_ = ~new_n19153_ | ~new_n19124_;
  assign new_n19202_ = ~pi279 | ~new_n19128_;
  assign new_n19203_ = ~pi278 | ~new_n19127_;
  assign new_n19204_ = ~pi297 | ~new_n19043_;
  assign new_n19205_ = ~new_n19152_ | ~new_n19129_;
  assign new_n19206_ = ~pi295 | ~new_n19037_;
  assign new_n19207_ = ~new_n19151_ | ~new_n19131_;
  assign new_n19208_ = ~pi291 | ~new_n19044_;
  assign new_n19209_ = ~new_n19148_ | ~new_n19133_;
  assign new_n19210_ = new_n5281_ & new_n19211_;
  assign new_n19211_ = ~new_n5278_;
  assign new_n19212_ = new_n19377_ & new_n19378_ & new_n19376_;
  assign new_n19213_ = new_n19291_ & new_n19290_;
  assign new_n19214_ = new_n19213_ & new_n19379_;
  assign new_n19215_ = new_n19389_ & new_n19388_;
  assign new_n19216_ = new_n19419_ & new_n19418_;
  assign new_n19217_ = new_n19375_ & new_n19220_ & new_n19288_;
  assign new_n19218_ = new_n19362_ & new_n19360_ & new_n19361_ & new_n19363_;
  assign new_n19219_ = new_n19381_ & new_n19379_ & new_n19380_ & new_n19382_;
  assign new_n19220_ = new_n19370_ & new_n19368_ & new_n19367_;
  assign new_n19221_ = new_n19212_ & new_n19223_ & new_n19371_ & new_n19289_ & new_n19217_;
  assign new_n19222_ = new_n19371_ & new_n19369_;
  assign new_n19223_ = new_n19431_ & new_n19430_;
  assign new_n19224_ = ~new_n19358_ | ~new_n19350_ | ~new_n19353_ | ~new_n19356_ | ~new_n19357_;
  assign new_n19225_ = ~new_n5310_;
  assign new_n19226_ = ~new_n5313_;
  assign new_n19227_ = ~new_n5311_;
  assign new_n19228_ = ~new_n5312_;
  assign new_n19229_ = ~new_n5346_;
  assign new_n19230_ = ~new_n5343_;
  assign new_n19231_ = ~new_n5309_;
  assign new_n19232_ = ~new_n5341_;
  assign new_n19233_ = ~new_n5325_;
  assign new_n19234_ = ~new_n5326_;
  assign new_n19235_ = ~new_n5328_;
  assign new_n19236_ = ~new_n5327_;
  assign new_n19237_ = ~new_n5329_;
  assign new_n19238_ = ~new_n5330_;
  assign new_n19239_ = ~new_n5331_;
  assign new_n19240_ = ~new_n5332_;
  assign new_n19241_ = ~new_n5335_;
  assign new_n19242_ = ~new_n5336_;
  assign new_n19243_ = ~new_n5334_;
  assign new_n19244_ = ~new_n5333_;
  assign new_n19245_ = ~new_n5324_;
  assign new_n19246_ = ~new_n5314_;
  assign new_n19247_ = ~new_n5322_;
  assign new_n19248_ = ~new_n5321_;
  assign new_n19249_ = ~new_n5323_;
  assign new_n19250_ = ~new_n5320_;
  assign new_n19251_ = ~new_n5319_;
  assign new_n19252_ = ~new_n5315_;
  assign new_n19253_ = ~new_n5317_;
  assign new_n19254_ = ~new_n5318_;
  assign new_n19255_ = ~new_n5316_;
  assign new_n19256_ = ~new_n5369_;
  assign new_n19257_ = ~new_n5337_;
  assign new_n19258_ = ~new_n5338_;
  assign new_n19259_ = ~new_n5339_;
  assign new_n19260_ = ~new_n5371_;
  assign new_n19261_ = ~new_n5347_;
  assign new_n19262_ = ~new_n5345_;
  assign new_n19263_ = ~new_n5344_;
  assign new_n19264_ = ~new_n5360_;
  assign new_n19265_ = ~new_n5361_;
  assign new_n19266_ = ~new_n5363_;
  assign new_n19267_ = ~new_n5348_;
  assign new_n19268_ = ~new_n5349_;
  assign new_n19269_ = ~new_n5351_;
  assign new_n19270_ = ~new_n5354_;
  assign new_n19271_ = ~new_n5355_;
  assign new_n19272_ = ~new_n5357_;
  assign new_n19273_ = ~new_n5366_;
  assign new_n19274_ = ~new_n5367_;
  assign new_n19275_ = ~new_n5353_;
  assign new_n19276_ = ~new_n5359_;
  assign new_n19277_ = ~new_n5365_;
  assign new_n19278_ = ~new_n5350_;
  assign new_n19279_ = ~new_n5352_;
  assign new_n19280_ = ~new_n5356_;
  assign new_n19281_ = ~new_n5358_;
  assign new_n19282_ = ~new_n5362_;
  assign new_n19283_ = ~new_n5364_;
  assign new_n19284_ = ~new_n5368_;
  assign new_n19285_ = ~new_n5370_;
  assign new_n19286_ = ~new_n5342_;
  assign new_n19287_ = new_n19223_ & new_n19372_;
  assign new_n19288_ = new_n19366_ & new_n19365_;
  assign new_n19289_ = new_n19369_ & new_n19364_;
  assign new_n19290_ = new_n19382_ & new_n19380_ & new_n19381_ & new_n19383_;
  assign new_n19291_ = new_n19386_ & new_n19385_ & new_n19384_;
  assign new_n19292_ = new_n19257_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19293_ = new_n5369_ & new_n19218_;
  assign new_n19294_ = new_n19392_ & new_n19379_;
  assign new_n19295_ = new_n19294_ & new_n19372_ & new_n19373_ & new_n19374_ & new_n19391_;
  assign new_n19296_ = new_n19297_ & new_n19213_ & new_n19393_;
  assign new_n19297_ = new_n19215_ & new_n19218_;
  assign new_n19298_ = new_n19372_ & new_n19373_ & new_n19259_;
  assign new_n19299_ = new_n19218_ & new_n5371_ & new_n19215_;
  assign new_n19300_ = new_n5347_ & new_n19252_;
  assign new_n19301_ = new_n19400_ & new_n19401_;
  assign new_n19302_ = new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19303_ = new_n19235_ & new_n19374_ & new_n19379_ & new_n19373_;
  assign new_n19304_ = new_n5360_ & new_n19382_ & new_n19380_;
  assign new_n19305_ = new_n19237_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19306_ = new_n19219_ & new_n5361_;
  assign new_n19307_ = new_n19239_ & new_n19374_ & new_n19383_ & new_n19373_;
  assign new_n19308_ = new_n19309_ & new_n19219_;
  assign new_n19309_ = new_n5363_ & new_n19384_;
  assign new_n19310_ = new_n19255_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19311_ = new_n19370_ & new_n19372_ & new_n19373_ & new_n19374_ & new_n19253_;
  assign new_n19312_ = new_n19251_ & new_n19374_ & new_n19375_ & new_n19373_;
  assign new_n19313_ = new_n5351_ & new_n19222_;
  assign new_n19314_ = new_n19247_ & new_n19374_ & new_n19377_ & new_n19373_;
  assign new_n19315_ = new_n5354_ & new_n19222_;
  assign new_n19316_ = new_n19249_ & new_n19374_ & new_n19376_ & new_n19373_;
  assign new_n19317_ = new_n19217_ & new_n19372_ & new_n19318_ & new_n19223_ & new_n19377_;
  assign new_n19318_ = new_n5355_ & new_n19222_;
  assign new_n19319_ = new_n19372_ & new_n19373_ & new_n19233_;
  assign new_n19320_ = new_n5357_ & new_n19374_;
  assign new_n19321_ = new_n19243_ & new_n19372_ & new_n19373_ & new_n19363_;
  assign new_n19322_ = new_n19362_ & new_n19372_ & new_n19373_ & new_n19363_ & new_n19241_;
  assign new_n19323_ = new_n19248_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19324_ = new_n5353_ & new_n19222_;
  assign new_n19325_ = new_n19236_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19326_ = new_n5359_ & new_n19380_ & new_n19379_;
  assign new_n19327_ = new_n19244_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19328_ = new_n19367_ & new_n19372_ & new_n19373_ & new_n19370_ & new_n19254_;
  assign new_n19329_ = new_n19375_ & new_n19374_;
  assign new_n19330_ = new_n19366_ & new_n19372_ & new_n19373_ & new_n19374_ & new_n19250_;
  assign new_n19331_ = new_n5352_ & new_n19222_;
  assign new_n19332_ = new_n19373_ & new_n19245_;
  assign new_n19333_ = new_n19332_ & new_n19223_ & new_n19374_;
  assign new_n19334_ = new_n19212_ & new_n5356_;
  assign new_n19335_ = new_n19234_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19336_ = new_n5358_ & new_n19379_;
  assign new_n19337_ = new_n19238_ & new_n19372_ & new_n19373_ & new_n19374_;
  assign new_n19338_ = new_n19339_ & new_n19219_;
  assign new_n19339_ = new_n5362_ & new_n19383_;
  assign new_n19340_ = new_n19240_ & new_n19374_ & new_n19383_ & new_n19373_;
  assign new_n19341_ = new_n19219_ & new_n19342_;
  assign new_n19342_ = new_n5364_ & new_n19385_ & new_n19384_;
  assign new_n19343_ = new_n19363_ & new_n19372_ & new_n19242_ & new_n19360_ & new_n19362_;
  assign new_n19344_ = new_n19214_ & new_n19373_ & new_n19374_ & new_n5368_;
  assign new_n19345_ = new_n19258_ & new_n19374_ & new_n19427_ & new_n19373_;
  assign new_n19346_ = new_n5370_ & new_n19218_;
  assign new_n19347_ = new_n19387_ & new_n19359_;
  assign new_n19348_ = new_n19398_ & new_n19394_;
  assign new_n19349_ = new_n19404_ & new_n19405_ & new_n19403_;
  assign new_n19350_ = new_n19349_ & new_n19348_ & new_n19347_;
  assign new_n19351_ = new_n19409_ & new_n19408_;
  assign new_n19352_ = new_n19411_ & new_n19410_;
  assign new_n19353_ = new_n19407_ & new_n19412_ & new_n19352_ & new_n19351_ & new_n19406_;
  assign new_n19354_ = new_n19416_ & new_n19415_;
  assign new_n19355_ = new_n19420_ & new_n19421_;
  assign new_n19356_ = new_n19414_ & new_n19417_ & new_n19355_ & new_n19354_ & new_n19413_;
  assign new_n19357_ = new_n19424_ & new_n19422_ & new_n19423_ & new_n19425_;
  assign new_n19358_ = new_n19428_ & new_n19216_ & new_n19426_;
  assign new_n19359_ = ~new_n19287_ | ~new_n19397_;
  assign new_n19360_ = ~new_n5335_ | ~new_n19274_;
  assign new_n19361_ = ~new_n5336_ | ~new_n19284_;
  assign new_n19362_ = ~new_n5334_ | ~new_n19273_;
  assign new_n19363_ = ~new_n5333_ | ~new_n19277_;
  assign new_n19364_ = ~new_n5324_ | ~new_n19280_;
  assign new_n19365_ = ~new_n5320_ | ~new_n19279_;
  assign new_n19366_ = ~new_n5319_ | ~new_n19269_;
  assign new_n19367_ = ~new_n5317_ | ~new_n19268_;
  assign new_n19368_ = ~new_n5318_ | ~new_n19278_;
  assign new_n19369_ = ~new_n5314_ | ~new_n19229_;
  assign new_n19370_ = ~new_n5316_ | ~new_n19267_;
  assign new_n19371_ = ~new_n5313_ | ~new_n19262_;
  assign new_n19372_ = ~new_n5310_ | ~new_n19286_;
  assign new_n19373_ = ~new_n5311_ | ~new_n19230_;
  assign new_n19374_ = ~new_n5312_ | ~new_n19263_;
  assign new_n19375_ = ~new_n5315_ | ~new_n19261_;
  assign new_n19376_ = ~new_n5322_ | ~new_n19270_;
  assign new_n19377_ = ~new_n5321_ | ~new_n19275_;
  assign new_n19378_ = ~new_n5323_ | ~new_n19271_;
  assign new_n19379_ = ~new_n5325_ | ~new_n19272_;
  assign new_n19380_ = ~new_n5326_ | ~new_n19281_;
  assign new_n19381_ = ~new_n5328_ | ~new_n19264_;
  assign new_n19382_ = ~new_n5327_ | ~new_n19276_;
  assign new_n19383_ = ~new_n5329_ | ~new_n19265_;
  assign new_n19384_ = ~new_n5330_ | ~new_n19282_;
  assign new_n19385_ = ~new_n5331_ | ~new_n19266_;
  assign new_n19386_ = ~new_n5332_ | ~new_n19283_;
  assign new_n19387_ = ~new_n19293_ | ~new_n19292_ | ~new_n19221_ | ~new_n19214_;
  assign new_n19388_ = ~new_n5337_ | ~new_n19256_;
  assign new_n19389_ = ~new_n5338_ | ~new_n19285_;
  assign new_n19390_ = ~new_n5372_ | ~new_n5373_;
  assign new_n19391_ = ~new_n5340_ | ~new_n19390_;
  assign new_n19392_ = ~new_n5339_ | ~new_n19260_;
  assign new_n19393_ = new_n5372_ | new_n5373_;
  assign new_n19394_ = ~new_n19295_ | ~new_n19221_ | ~new_n19296_;
  assign new_n19395_ = ~new_n19371_ | ~new_n19374_ | ~new_n5346_ | ~new_n19373_ | ~new_n19246_;
  assign new_n19396_ = ~new_n5343_ | ~new_n19227_;
  assign new_n19397_ = ~new_n19396_ | ~new_n19395_;
  assign new_n19398_ = ~new_n19214_ | ~new_n19298_ | ~new_n19221_ | ~new_n19374_ | ~new_n19299_;
  assign new_n19399_ = ~new_n19300_ | ~new_n19222_;
  assign new_n19400_ = ~new_n5345_ | ~new_n19226_;
  assign new_n19401_ = ~new_n5344_ | ~new_n19228_;
  assign new_n19402_ = ~new_n19301_ | ~new_n19399_;
  assign new_n19403_ = ~new_n19302_ | ~new_n19223_ | ~new_n19402_;
  assign new_n19404_ = ~new_n19221_ | ~new_n19303_ | ~new_n19372_ | ~new_n19304_;
  assign new_n19405_ = ~new_n19305_ | ~new_n19306_ | ~new_n19221_;
  assign new_n19406_ = ~new_n19308_ | ~new_n19307_ | ~new_n19372_ | ~new_n19221_;
  assign new_n19407_ = ~new_n5348_ | ~new_n19310_ | ~new_n19375_ | ~new_n19223_ | ~new_n19222_;
  assign new_n19408_ = ~new_n5349_ | ~new_n19311_ | ~new_n19375_ | ~new_n19223_ | ~new_n19222_;
  assign new_n19409_ = ~new_n19223_ | ~new_n19312_ | ~new_n19372_ | ~new_n19313_ | ~new_n19220_;
  assign new_n19410_ = ~new_n19223_ | ~new_n19314_ | ~new_n19372_ | ~new_n19315_ | ~new_n19217_;
  assign new_n19411_ = ~new_n19316_ | ~new_n19317_;
  assign new_n19412_ = ~new_n19319_ | ~new_n19320_ | ~new_n19221_;
  assign new_n19413_ = ~new_n5366_ | ~new_n19321_ | ~new_n19221_ | ~new_n19374_ | ~new_n19214_;
  assign new_n19414_ = ~new_n5367_ | ~new_n19322_ | ~new_n19221_ | ~new_n19374_ | ~new_n19214_;
  assign new_n19415_ = ~new_n19217_ | ~new_n19323_ | ~new_n19324_ | ~new_n19223_;
  assign new_n19416_ = ~new_n19325_ | ~new_n19326_ | ~new_n19221_;
  assign new_n19417_ = ~new_n5365_ | ~new_n19327_ | ~new_n19221_ | ~new_n19214_;
  assign new_n19418_ = ~new_n19429_ | ~new_n19433_ | ~new_n19432_;
  assign new_n19419_ = ~new_n19225_ | ~new_n19223_ | ~new_n5342_;
  assign new_n19420_ = ~new_n5350_ | ~new_n19328_ | ~new_n19329_ | ~new_n19223_ | ~new_n19222_;
  assign new_n19421_ = ~new_n19220_ | ~new_n19330_ | ~new_n19331_ | ~new_n19223_ | ~new_n19375_;
  assign new_n19422_ = ~new_n19217_ | ~new_n19333_ | ~new_n19372_ | ~new_n19222_ | ~new_n19334_;
  assign new_n19423_ = ~new_n19335_ | ~new_n19336_ | ~new_n19221_;
  assign new_n19424_ = ~new_n19337_ | ~new_n19221_ | ~new_n19338_;
  assign new_n19425_ = ~new_n19341_ | ~new_n19340_ | ~new_n19372_ | ~new_n19221_;
  assign new_n19426_ = ~new_n19343_ | ~new_n19221_ | ~new_n19344_;
  assign new_n19427_ = ~new_n5337_ | ~new_n19256_;
  assign new_n19428_ = ~new_n19214_ | ~new_n19345_ | ~new_n19372_ | ~new_n19221_ | ~new_n19346_;
  assign new_n19429_ = ~new_n5341_ | ~new_n5309_;
  assign new_n19430_ = ~new_n5309_ | ~new_n19232_;
  assign new_n19431_ = ~new_n5341_ | ~new_n19231_;
  assign new_n19432_ = new_n5374_ | new_n5341_;
  assign new_n19433_ = ~new_n5374_ | ~new_n19231_;
  assign new_n19434_ = ~new_n5281_;
  assign new_n19435_ = ~new_n5278_;
  assign new_n19436_ = new_n19438_ & new_n19437_;
  assign new_n19437_ = ~new_n5278_ | ~new_n19434_;
  assign new_n19438_ = ~new_n5281_ | ~new_n19435_;
  assign new_n19439_ = new_n19530_ & new_n19529_;
  assign new_n19440_ = new_n19531_ & new_n19532_;
  assign new_n19441_ = new_n19548_ & new_n19547_;
  assign new_n19442_ = new_n19590_ & new_n19589_;
  assign new_n19443_ = new_n19599_ & new_n19598_;
  assign new_n19444_ = new_n19617_ & new_n19616_;
  assign new_n19445_ = new_n19653_ & new_n19650_;
  assign new_n19446_ = new_n19646_ & new_n19643_;
  assign new_n19447_ = new_n19637_ & new_n19634_;
  assign new_n19448_ = new_n19631_ & new_n19627_;
  assign new_n19449_ = new_n19586_ & new_n19583_;
  assign new_n19450_ = new_n19578_ & new_n19575_;
  assign new_n19451_ = new_n19564_ & new_n19561_;
  assign new_n19452_ = ~pi380;
  assign new_n19453_ = ~new_n5666_;
  assign new_n19454_ = ~new_n5669_;
  assign new_n19455_ = ~new_n5666_ | ~pi380;
  assign new_n19456_ = ~pi381;
  assign new_n19457_ = ~pi378;
  assign new_n19458_ = ~new_n5660_;
  assign new_n19459_ = ~new_n5663_;
  assign new_n19460_ = ~pi376;
  assign new_n19461_ = ~new_n5654_;
  assign new_n19462_ = ~pi374;
  assign new_n19463_ = ~new_n5645_;
  assign new_n19464_ = ~new_n5645_ | ~pi374;
  assign new_n19465_ = ~pi377;
  assign new_n19466_ = ~new_n5657_;
  assign new_n19467_ = ~new_n5660_ | ~pi378;
  assign new_n19468_ = ~pi379;
  assign new_n19469_ = ~pi382;
  assign new_n19470_ = ~new_n5672_;
  assign new_n19471_ = ~new_n5675_;
  assign new_n19472_ = ~pi383;
  assign new_n19473_ = ~new_n19484_ | ~new_n19556_;
  assign new_n19474_ = ~new_n19544_ | ~new_n19545_ | ~new_n19543_;
  assign new_n19475_ = ~new_n19533_ | ~new_n19534_;
  assign new_n19476_ = ~pi375 | ~new_n5651_;
  assign new_n19477_ = ~new_n19570_ | ~new_n19571_ | ~new_n19569_;
  assign new_n19478_ = ~new_n19567_ | ~new_n19566_;
  assign new_n19479_ = ~pi390;
  assign new_n19480_ = ~new_n5696_;
  assign new_n19481_ = ~new_n5699_;
  assign new_n19482_ = ~new_n5696_ | ~pi390;
  assign new_n19483_ = ~pi391;
  assign new_n19484_ = ~new_n5672_ | ~pi382;
  assign new_n19485_ = ~pi384;
  assign new_n19486_ = ~new_n5678_;
  assign new_n19487_ = ~pi386;
  assign new_n19488_ = ~new_n5684_;
  assign new_n19489_ = ~pi385;
  assign new_n19490_ = ~new_n5681_;
  assign new_n19491_ = ~new_n5681_ | ~pi385;
  assign new_n19492_ = ~pi387;
  assign new_n19493_ = ~new_n5687_;
  assign new_n19494_ = ~pi388;
  assign new_n19495_ = ~new_n5690_;
  assign new_n19496_ = ~pi389;
  assign new_n19497_ = ~new_n5693_;
  assign new_n19498_ = ~pi392;
  assign new_n19499_ = ~new_n5702_;
  assign new_n19500_ = ~new_n19622_ | ~new_n19621_ | ~new_n19620_;
  assign new_n19501_ = ~new_n19614_ | ~new_n19613_;
  assign new_n19502_ = ~new_n19491_ | ~new_n19639_;
  assign new_n19503_ = ~new_n19694_ | ~new_n19693_;
  assign new_n19504_ = ~new_n19743_ | ~new_n19742_;
  assign new_n19505_ = ~new_n19666_ | ~new_n19665_;
  assign new_n19506_ = ~new_n19671_ | ~new_n19670_;
  assign new_n19507_ = ~new_n19678_ | ~new_n19677_;
  assign new_n19508_ = ~new_n19685_ | ~new_n19684_;
  assign new_n19509_ = ~new_n19690_ | ~new_n19689_;
  assign new_n19510_ = ~new_n19706_ | ~new_n19705_;
  assign new_n19511_ = ~new_n19713_ | ~new_n19712_;
  assign new_n19512_ = ~new_n19720_ | ~new_n19719_;
  assign new_n19513_ = ~new_n19727_ | ~new_n19726_;
  assign new_n19514_ = ~new_n19734_ | ~new_n19733_;
  assign new_n19515_ = ~new_n19739_ | ~new_n19738_;
  assign new_n19516_ = ~new_n19553_ | ~new_n19552_ | ~new_n19551_;
  assign new_n19517_ = ~new_n19568_ | ~new_n19580_;
  assign new_n19518_ = ~new_n19476_ | ~new_n19587_;
  assign new_n19519_ = ~new_n5644_;
  assign new_n19520_ = ~pi393;
  assign new_n19521_ = ~new_n19610_ | ~new_n19609_;
  assign new_n19522_ = ~new_n19606_ | ~new_n19605_;
  assign new_n19523_ = ~new_n19596_ | ~new_n19595_;
  assign new_n19524_ = ~new_n19467_;
  assign new_n19525_ = ~pi383 | ~new_n5675_;
  assign new_n19526_ = ~new_n5684_ | ~pi386;
  assign new_n19527_ = ~new_n19491_;
  assign new_n19528_ = ~new_n19484_;
  assign new_n19529_ = new_n5663_ | pi379;
  assign new_n19530_ = new_n5660_ | pi378;
  assign new_n19531_ = pi377 | new_n5657_;
  assign new_n19532_ = pi376 | new_n5654_;
  assign new_n19533_ = ~new_n19464_;
  assign new_n19534_ = pi375 | new_n5651_;
  assign new_n19535_ = ~new_n19475_;
  assign new_n19536_ = ~new_n19476_;
  assign new_n19537_ = ~new_n19475_ | ~new_n19476_;
  assign new_n19538_ = ~new_n19531_ | ~pi376 | ~new_n5654_;
  assign new_n19539_ = ~new_n19440_ | ~new_n19537_;
  assign new_n19540_ = ~new_n5657_ | ~pi377;
  assign new_n19541_ = ~new_n19539_ | ~new_n19540_ | ~new_n19538_;
  assign new_n19542_ = ~new_n19468_ | ~new_n19467_;
  assign new_n19543_ = ~new_n5663_ | ~new_n19542_;
  assign new_n19544_ = ~new_n19439_ | ~new_n19541_;
  assign new_n19545_ = ~pi379 | ~new_n19524_;
  assign new_n19546_ = ~new_n19474_;
  assign new_n19547_ = new_n5669_ | pi381;
  assign new_n19548_ = new_n5666_ | pi380;
  assign new_n19549_ = ~new_n19455_;
  assign new_n19550_ = ~new_n19456_ | ~new_n19455_;
  assign new_n19551_ = ~new_n5669_ | ~new_n19550_;
  assign new_n19552_ = ~pi381 | ~new_n19549_;
  assign new_n19553_ = ~new_n19441_ | ~new_n19474_;
  assign new_n19554_ = ~new_n19516_;
  assign new_n19555_ = pi382 | new_n5672_;
  assign new_n19556_ = ~new_n19555_ | ~new_n19516_;
  assign new_n19557_ = ~new_n19473_;
  assign new_n19558_ = new_n5675_ | pi383;
  assign new_n19559_ = pi380 | new_n5666_;
  assign new_n19560_ = ~new_n19559_ | ~new_n19474_;
  assign new_n19561_ = ~new_n19672_ | ~new_n19560_ | ~new_n19455_ | ~new_n19673_;
  assign new_n19562_ = ~new_n19546_ | ~new_n19455_;
  assign new_n19563_ = ~pi381 | ~new_n5669_;
  assign new_n19564_ = ~new_n19562_ | ~new_n19563_ | ~new_n19441_;
  assign new_n19565_ = new_n5666_ | pi380;
  assign new_n19566_ = ~new_n19536_ | ~new_n19532_;
  assign new_n19567_ = ~new_n5654_ | ~pi376;
  assign new_n19568_ = ~new_n19478_;
  assign new_n19569_ = ~new_n19535_ | ~new_n19440_;
  assign new_n19570_ = ~new_n19478_ | ~new_n19531_;
  assign new_n19571_ = ~new_n5657_ | ~pi377;
  assign new_n19572_ = ~new_n19477_;
  assign new_n19573_ = pi378 | new_n5660_;
  assign new_n19574_ = ~new_n19573_ | ~new_n19477_;
  assign new_n19575_ = ~new_n19679_ | ~new_n19574_ | ~new_n19467_ | ~new_n19680_;
  assign new_n19576_ = ~new_n19572_ | ~new_n19467_;
  assign new_n19577_ = ~pi379 | ~new_n5663_;
  assign new_n19578_ = ~new_n19576_ | ~new_n19577_ | ~new_n19439_;
  assign new_n19579_ = new_n5660_ | pi378;
  assign new_n19580_ = ~new_n19535_ | ~new_n19532_;
  assign new_n19581_ = ~new_n19517_;
  assign new_n19582_ = ~new_n5657_ | ~pi377;
  assign new_n19583_ = ~new_n19691_ | ~new_n19475_ | ~new_n19476_ | ~new_n19692_;
  assign new_n19584_ = ~new_n19476_ | ~new_n19475_;
  assign new_n19585_ = ~new_n5654_ | ~pi376;
  assign new_n19586_ = ~new_n19584_ | ~new_n19585_ | ~new_n19532_;
  assign new_n19587_ = pi375 | new_n5651_;
  assign new_n19588_ = ~new_n19518_;
  assign new_n19589_ = new_n5675_ | pi383;
  assign new_n19590_ = new_n5678_ | pi384;
  assign new_n19591_ = ~new_n19528_ | ~new_n19442_;
  assign new_n19592_ = ~new_n5678_ | ~pi384;
  assign new_n19593_ = ~new_n19591_ | ~new_n19592_ | ~new_n19525_;
  assign new_n19594_ = pi384 | new_n5678_;
  assign new_n19595_ = ~new_n19516_ | ~new_n19555_ | ~new_n19442_;
  assign new_n19596_ = ~new_n19594_ | ~new_n19593_;
  assign new_n19597_ = ~new_n19523_;
  assign new_n19598_ = new_n5687_ | pi387;
  assign new_n19599_ = new_n5684_ | pi386;
  assign new_n19600_ = ~new_n19527_ | ~new_n19443_;
  assign new_n19601_ = ~new_n5687_ | ~pi387;
  assign new_n19602_ = ~new_n19600_ | ~new_n19601_ | ~new_n19526_;
  assign new_n19603_ = pi385 | new_n5681_;
  assign new_n19604_ = pi387 | new_n5687_;
  assign new_n19605_ = ~new_n19523_ | ~new_n19603_ | ~new_n19443_;
  assign new_n19606_ = ~new_n19604_ | ~new_n19602_;
  assign new_n19607_ = ~new_n19522_;
  assign new_n19608_ = pi388 | new_n5690_;
  assign new_n19609_ = ~new_n19608_ | ~new_n19522_;
  assign new_n19610_ = ~new_n5690_ | ~pi388;
  assign new_n19611_ = ~new_n19521_;
  assign new_n19612_ = pi389 | new_n5693_;
  assign new_n19613_ = ~new_n19612_ | ~new_n19521_;
  assign new_n19614_ = ~new_n5693_ | ~pi389;
  assign new_n19615_ = ~new_n19501_;
  assign new_n19616_ = new_n5699_ | pi391;
  assign new_n19617_ = new_n5696_ | pi390;
  assign new_n19618_ = ~new_n19482_;
  assign new_n19619_ = ~new_n19483_ | ~new_n19482_;
  assign new_n19620_ = ~new_n5699_ | ~new_n19619_;
  assign new_n19621_ = ~pi391 | ~new_n19618_;
  assign new_n19622_ = ~new_n19444_ | ~new_n19501_;
  assign new_n19623_ = ~new_n19500_;
  assign new_n19624_ = pi392 | new_n5702_;
  assign new_n19625_ = ~new_n19624_ | ~new_n19500_;
  assign new_n19626_ = ~new_n5702_ | ~pi392;
  assign new_n19627_ = ~new_n19695_ | ~new_n19625_ | ~new_n19626_ | ~new_n19696_;
  assign new_n19628_ = ~new_n5702_ | ~pi392;
  assign new_n19629_ = ~new_n19623_ | ~new_n19628_;
  assign new_n19630_ = new_n5702_ | pi392;
  assign new_n19631_ = ~new_n19629_ | ~new_n19630_ | ~new_n19699_;
  assign new_n19632_ = pi390 | new_n5696_;
  assign new_n19633_ = ~new_n19632_ | ~new_n19501_;
  assign new_n19634_ = ~new_n19707_ | ~new_n19633_ | ~new_n19482_ | ~new_n19708_;
  assign new_n19635_ = ~new_n19615_ | ~new_n19482_;
  assign new_n19636_ = ~pi391 | ~new_n5699_;
  assign new_n19637_ = ~new_n19635_ | ~new_n19636_ | ~new_n19444_;
  assign new_n19638_ = new_n5696_ | pi390;
  assign new_n19639_ = ~new_n19603_ | ~new_n19523_;
  assign new_n19640_ = ~new_n19502_;
  assign new_n19641_ = pi386 | new_n5684_;
  assign new_n19642_ = ~new_n19641_ | ~new_n19502_;
  assign new_n19643_ = ~new_n19728_ | ~new_n19642_ | ~new_n19526_ | ~new_n19729_;
  assign new_n19644_ = ~new_n19640_ | ~new_n19526_;
  assign new_n19645_ = ~new_n5687_ | ~pi387;
  assign new_n19646_ = ~new_n19644_ | ~new_n19645_ | ~new_n19443_;
  assign new_n19647_ = new_n5684_ | pi386;
  assign new_n19648_ = pi383 | new_n5675_;
  assign new_n19649_ = ~new_n19648_ | ~new_n19473_;
  assign new_n19650_ = ~new_n19740_ | ~new_n19649_ | ~new_n19525_ | ~new_n19741_;
  assign new_n19651_ = ~new_n19557_ | ~new_n19525_;
  assign new_n19652_ = ~new_n5678_ | ~pi384;
  assign new_n19653_ = ~new_n19651_ | ~new_n19652_ | ~new_n19442_;
  assign new_n19654_ = ~new_n19558_ | ~new_n19525_;
  assign new_n19655_ = ~new_n19555_ | ~new_n19484_;
  assign new_n19656_ = ~new_n19565_ | ~new_n19455_;
  assign new_n19657_ = ~new_n19579_ | ~new_n19467_;
  assign new_n19658_ = ~new_n19582_ | ~new_n19531_;
  assign new_n19659_ = ~new_n19638_ | ~new_n19482_;
  assign new_n19660_ = ~new_n19647_ | ~new_n19526_;
  assign new_n19661_ = ~new_n19603_ | ~new_n19491_;
  assign new_n19662_ = ~new_n5675_ | ~new_n19472_;
  assign new_n19663_ = ~pi383 | ~new_n19471_;
  assign new_n19664_ = ~new_n19663_ | ~new_n19662_;
  assign new_n19665_ = ~new_n19654_ | ~new_n19473_;
  assign new_n19666_ = ~new_n19664_ | ~new_n19557_;
  assign new_n19667_ = ~new_n5672_ | ~new_n19469_;
  assign new_n19668_ = ~pi382 | ~new_n19470_;
  assign new_n19669_ = ~new_n19668_ | ~new_n19667_;
  assign new_n19670_ = ~new_n19655_ | ~new_n19516_;
  assign new_n19671_ = ~new_n19554_ | ~new_n19669_;
  assign new_n19672_ = ~new_n5669_ | ~new_n19456_;
  assign new_n19673_ = ~pi381 | ~new_n19454_;
  assign new_n19674_ = ~new_n5666_ | ~new_n19452_;
  assign new_n19675_ = ~pi380 | ~new_n19453_;
  assign new_n19676_ = ~new_n19675_ | ~new_n19674_;
  assign new_n19677_ = ~new_n19656_ | ~new_n19474_;
  assign new_n19678_ = ~new_n19676_ | ~new_n19546_;
  assign new_n19679_ = ~new_n5663_ | ~new_n19468_;
  assign new_n19680_ = ~pi379 | ~new_n19459_;
  assign new_n19681_ = ~new_n5660_ | ~new_n19457_;
  assign new_n19682_ = ~pi378 | ~new_n19458_;
  assign new_n19683_ = ~new_n19682_ | ~new_n19681_;
  assign new_n19684_ = ~new_n19657_ | ~new_n19477_;
  assign new_n19685_ = ~new_n19683_ | ~new_n19572_;
  assign new_n19686_ = ~new_n5657_ | ~new_n19465_;
  assign new_n19687_ = ~pi377 | ~new_n19466_;
  assign new_n19688_ = ~new_n19687_ | ~new_n19686_;
  assign new_n19689_ = ~new_n19658_ | ~new_n19517_;
  assign new_n19690_ = ~new_n19581_ | ~new_n19688_;
  assign new_n19691_ = ~new_n5654_ | ~new_n19460_;
  assign new_n19692_ = ~pi376 | ~new_n19461_;
  assign new_n19693_ = ~new_n19533_ | ~new_n19518_;
  assign new_n19694_ = ~new_n19588_ | ~new_n19464_;
  assign new_n19695_ = ~new_n5644_ | ~new_n19520_;
  assign new_n19696_ = ~pi393 | ~new_n19519_;
  assign new_n19697_ = ~new_n5644_ | ~new_n19520_;
  assign new_n19698_ = ~pi393 | ~new_n19519_;
  assign new_n19699_ = ~new_n19698_ | ~new_n19697_;
  assign new_n19700_ = ~new_n5702_ | ~new_n19498_;
  assign new_n19701_ = ~pi392 | ~new_n19499_;
  assign new_n19702_ = ~new_n5702_ | ~new_n19498_;
  assign new_n19703_ = ~pi392 | ~new_n19499_;
  assign new_n19704_ = ~new_n19703_ | ~new_n19702_;
  assign new_n19705_ = ~new_n19500_ | ~new_n19701_ | ~new_n19700_;
  assign new_n19706_ = ~new_n19704_ | ~new_n19623_;
  assign new_n19707_ = ~new_n5699_ | ~new_n19483_;
  assign new_n19708_ = ~pi391 | ~new_n19481_;
  assign new_n19709_ = ~new_n5696_ | ~new_n19479_;
  assign new_n19710_ = ~pi390 | ~new_n19480_;
  assign new_n19711_ = ~new_n19710_ | ~new_n19709_;
  assign new_n19712_ = ~new_n19659_ | ~new_n19501_;
  assign new_n19713_ = ~new_n19711_ | ~new_n19615_;
  assign new_n19714_ = ~new_n5693_ | ~new_n19496_;
  assign new_n19715_ = ~pi389 | ~new_n19497_;
  assign new_n19716_ = ~new_n5693_ | ~new_n19496_;
  assign new_n19717_ = ~pi389 | ~new_n19497_;
  assign new_n19718_ = ~new_n19717_ | ~new_n19716_;
  assign new_n19719_ = ~new_n19521_ | ~new_n19715_ | ~new_n19714_;
  assign new_n19720_ = ~new_n19611_ | ~new_n19718_;
  assign new_n19721_ = ~new_n5690_ | ~new_n19494_;
  assign new_n19722_ = ~pi388 | ~new_n19495_;
  assign new_n19723_ = ~new_n5690_ | ~new_n19494_;
  assign new_n19724_ = ~pi388 | ~new_n19495_;
  assign new_n19725_ = ~new_n19724_ | ~new_n19723_;
  assign new_n19726_ = ~new_n19522_ | ~new_n19722_ | ~new_n19721_;
  assign new_n19727_ = ~new_n19607_ | ~new_n19725_;
  assign new_n19728_ = ~new_n5687_ | ~new_n19492_;
  assign new_n19729_ = ~pi387 | ~new_n19493_;
  assign new_n19730_ = ~new_n5684_ | ~new_n19487_;
  assign new_n19731_ = ~pi386 | ~new_n19488_;
  assign new_n19732_ = ~new_n19731_ | ~new_n19730_;
  assign new_n19733_ = ~new_n19660_ | ~new_n19502_;
  assign new_n19734_ = ~new_n19732_ | ~new_n19640_;
  assign new_n19735_ = ~new_n5681_ | ~new_n19489_;
  assign new_n19736_ = ~pi385 | ~new_n19490_;
  assign new_n19737_ = ~new_n19736_ | ~new_n19735_;
  assign new_n19738_ = ~new_n19661_ | ~new_n19523_;
  assign new_n19739_ = ~new_n19597_ | ~new_n19737_;
  assign new_n19740_ = ~new_n5678_ | ~new_n19485_;
  assign new_n19741_ = ~pi384 | ~new_n19486_;
  assign new_n19742_ = ~new_n5645_ | ~new_n19462_;
  assign new_n19743_ = ~pi374 | ~new_n19463_;
  assign new_n19744_ = new_n19835_ & new_n19834_;
  assign new_n19745_ = new_n19836_ & new_n19837_;
  assign new_n19746_ = new_n19853_ & new_n19852_;
  assign new_n19747_ = new_n19895_ & new_n19894_;
  assign new_n19748_ = new_n19904_ & new_n19903_;
  assign new_n19749_ = new_n19922_ & new_n19921_;
  assign new_n19750_ = new_n19958_ & new_n19955_;
  assign new_n19751_ = new_n19951_ & new_n19948_;
  assign new_n19752_ = new_n19942_ & new_n19939_;
  assign new_n19753_ = new_n19936_ & new_n19932_;
  assign new_n19754_ = new_n19891_ & new_n19888_;
  assign new_n19755_ = new_n19883_ & new_n19880_;
  assign new_n19756_ = new_n19869_ & new_n19866_;
  assign new_n19757_ = ~pi412;
  assign new_n19758_ = ~new_n5666_;
  assign new_n19759_ = ~new_n5669_;
  assign new_n19760_ = ~new_n5666_ | ~pi412;
  assign new_n19761_ = ~pi413;
  assign new_n19762_ = ~pi410;
  assign new_n19763_ = ~new_n5660_;
  assign new_n19764_ = ~new_n5663_;
  assign new_n19765_ = ~pi408;
  assign new_n19766_ = ~new_n5654_;
  assign new_n19767_ = ~pi406;
  assign new_n19768_ = ~new_n5645_;
  assign new_n19769_ = ~new_n5645_ | ~pi406;
  assign new_n19770_ = ~pi409;
  assign new_n19771_ = ~new_n5657_;
  assign new_n19772_ = ~new_n5660_ | ~pi410;
  assign new_n19773_ = ~pi411;
  assign new_n19774_ = ~pi414;
  assign new_n19775_ = ~new_n5672_;
  assign new_n19776_ = ~new_n5675_;
  assign new_n19777_ = ~pi415;
  assign new_n19778_ = ~new_n19789_ | ~new_n19861_;
  assign new_n19779_ = ~new_n19849_ | ~new_n19850_ | ~new_n19848_;
  assign new_n19780_ = ~new_n19838_ | ~new_n19839_;
  assign new_n19781_ = ~pi407 | ~new_n5651_;
  assign new_n19782_ = ~new_n19875_ | ~new_n19876_ | ~new_n19874_;
  assign new_n19783_ = ~new_n19872_ | ~new_n19871_;
  assign new_n19784_ = ~pi422;
  assign new_n19785_ = ~new_n5696_;
  assign new_n19786_ = ~new_n5699_;
  assign new_n19787_ = ~new_n5696_ | ~pi422;
  assign new_n19788_ = ~pi423;
  assign new_n19789_ = ~new_n5672_ | ~pi414;
  assign new_n19790_ = ~pi416;
  assign new_n19791_ = ~new_n5678_;
  assign new_n19792_ = ~pi418;
  assign new_n19793_ = ~new_n5684_;
  assign new_n19794_ = ~pi417;
  assign new_n19795_ = ~new_n5681_;
  assign new_n19796_ = ~new_n5681_ | ~pi417;
  assign new_n19797_ = ~pi419;
  assign new_n19798_ = ~new_n5687_;
  assign new_n19799_ = ~pi420;
  assign new_n19800_ = ~new_n5690_;
  assign new_n19801_ = ~pi421;
  assign new_n19802_ = ~new_n5693_;
  assign new_n19803_ = ~pi424;
  assign new_n19804_ = ~new_n5702_;
  assign new_n19805_ = ~new_n19927_ | ~new_n19926_ | ~new_n19925_;
  assign new_n19806_ = ~new_n19919_ | ~new_n19918_;
  assign new_n19807_ = ~new_n19796_ | ~new_n19944_;
  assign new_n19808_ = ~new_n19999_ | ~new_n19998_;
  assign new_n19809_ = ~new_n20048_ | ~new_n20047_;
  assign new_n19810_ = ~new_n19971_ | ~new_n19970_;
  assign new_n19811_ = ~new_n19976_ | ~new_n19975_;
  assign new_n19812_ = ~new_n19983_ | ~new_n19982_;
  assign new_n19813_ = ~new_n19990_ | ~new_n19989_;
  assign new_n19814_ = ~new_n19995_ | ~new_n19994_;
  assign new_n19815_ = ~new_n20011_ | ~new_n20010_;
  assign new_n19816_ = ~new_n20018_ | ~new_n20017_;
  assign new_n19817_ = ~new_n20025_ | ~new_n20024_;
  assign new_n19818_ = ~new_n20032_ | ~new_n20031_;
  assign new_n19819_ = ~new_n20039_ | ~new_n20038_;
  assign new_n19820_ = ~new_n20044_ | ~new_n20043_;
  assign new_n19821_ = ~new_n19858_ | ~new_n19857_ | ~new_n19856_;
  assign new_n19822_ = ~new_n19873_ | ~new_n19885_;
  assign new_n19823_ = ~new_n19781_ | ~new_n19892_;
  assign new_n19824_ = ~new_n5644_;
  assign new_n19825_ = ~pi425;
  assign new_n19826_ = ~new_n19915_ | ~new_n19914_;
  assign new_n19827_ = ~new_n19911_ | ~new_n19910_;
  assign new_n19828_ = ~new_n19901_ | ~new_n19900_;
  assign new_n19829_ = ~new_n19772_;
  assign new_n19830_ = ~pi415 | ~new_n5675_;
  assign new_n19831_ = ~new_n5684_ | ~pi418;
  assign new_n19832_ = ~new_n19796_;
  assign new_n19833_ = ~new_n19789_;
  assign new_n19834_ = new_n5663_ | pi411;
  assign new_n19835_ = new_n5660_ | pi410;
  assign new_n19836_ = pi409 | new_n5657_;
  assign new_n19837_ = pi408 | new_n5654_;
  assign new_n19838_ = ~new_n19769_;
  assign new_n19839_ = pi407 | new_n5651_;
  assign new_n19840_ = ~new_n19780_;
  assign new_n19841_ = ~new_n19781_;
  assign new_n19842_ = ~new_n19780_ | ~new_n19781_;
  assign new_n19843_ = ~new_n19836_ | ~pi408 | ~new_n5654_;
  assign new_n19844_ = ~new_n19745_ | ~new_n19842_;
  assign new_n19845_ = ~new_n5657_ | ~pi409;
  assign new_n19846_ = ~new_n19844_ | ~new_n19845_ | ~new_n19843_;
  assign new_n19847_ = ~new_n19773_ | ~new_n19772_;
  assign new_n19848_ = ~new_n5663_ | ~new_n19847_;
  assign new_n19849_ = ~new_n19744_ | ~new_n19846_;
  assign new_n19850_ = ~pi411 | ~new_n19829_;
  assign new_n19851_ = ~new_n19779_;
  assign new_n19852_ = new_n5669_ | pi413;
  assign new_n19853_ = new_n5666_ | pi412;
  assign new_n19854_ = ~new_n19760_;
  assign new_n19855_ = ~new_n19761_ | ~new_n19760_;
  assign new_n19856_ = ~new_n5669_ | ~new_n19855_;
  assign new_n19857_ = ~pi413 | ~new_n19854_;
  assign new_n19858_ = ~new_n19746_ | ~new_n19779_;
  assign new_n19859_ = ~new_n19821_;
  assign new_n19860_ = pi414 | new_n5672_;
  assign new_n19861_ = ~new_n19860_ | ~new_n19821_;
  assign new_n19862_ = ~new_n19778_;
  assign new_n19863_ = new_n5675_ | pi415;
  assign new_n19864_ = pi412 | new_n5666_;
  assign new_n19865_ = ~new_n19864_ | ~new_n19779_;
  assign new_n19866_ = ~new_n19977_ | ~new_n19865_ | ~new_n19760_ | ~new_n19978_;
  assign new_n19867_ = ~new_n19851_ | ~new_n19760_;
  assign new_n19868_ = ~pi413 | ~new_n5669_;
  assign new_n19869_ = ~new_n19867_ | ~new_n19868_ | ~new_n19746_;
  assign new_n19870_ = new_n5666_ | pi412;
  assign new_n19871_ = ~new_n19841_ | ~new_n19837_;
  assign new_n19872_ = ~new_n5654_ | ~pi408;
  assign new_n19873_ = ~new_n19783_;
  assign new_n19874_ = ~new_n19840_ | ~new_n19745_;
  assign new_n19875_ = ~new_n19783_ | ~new_n19836_;
  assign new_n19876_ = ~new_n5657_ | ~pi409;
  assign new_n19877_ = ~new_n19782_;
  assign new_n19878_ = pi410 | new_n5660_;
  assign new_n19879_ = ~new_n19878_ | ~new_n19782_;
  assign new_n19880_ = ~new_n19984_ | ~new_n19879_ | ~new_n19772_ | ~new_n19985_;
  assign new_n19881_ = ~new_n19877_ | ~new_n19772_;
  assign new_n19882_ = ~pi411 | ~new_n5663_;
  assign new_n19883_ = ~new_n19881_ | ~new_n19882_ | ~new_n19744_;
  assign new_n19884_ = new_n5660_ | pi410;
  assign new_n19885_ = ~new_n19840_ | ~new_n19837_;
  assign new_n19886_ = ~new_n19822_;
  assign new_n19887_ = ~new_n5657_ | ~pi409;
  assign new_n19888_ = ~new_n19996_ | ~new_n19780_ | ~new_n19781_ | ~new_n19997_;
  assign new_n19889_ = ~new_n19781_ | ~new_n19780_;
  assign new_n19890_ = ~new_n5654_ | ~pi408;
  assign new_n19891_ = ~new_n19889_ | ~new_n19890_ | ~new_n19837_;
  assign new_n19892_ = pi407 | new_n5651_;
  assign new_n19893_ = ~new_n19823_;
  assign new_n19894_ = new_n5675_ | pi415;
  assign new_n19895_ = new_n5678_ | pi416;
  assign new_n19896_ = ~new_n19833_ | ~new_n19747_;
  assign new_n19897_ = ~new_n5678_ | ~pi416;
  assign new_n19898_ = ~new_n19896_ | ~new_n19897_ | ~new_n19830_;
  assign new_n19899_ = pi416 | new_n5678_;
  assign new_n19900_ = ~new_n19821_ | ~new_n19860_ | ~new_n19747_;
  assign new_n19901_ = ~new_n19899_ | ~new_n19898_;
  assign new_n19902_ = ~new_n19828_;
  assign new_n19903_ = new_n5687_ | pi419;
  assign new_n19904_ = new_n5684_ | pi418;
  assign new_n19905_ = ~new_n19832_ | ~new_n19748_;
  assign new_n19906_ = ~new_n5687_ | ~pi419;
  assign new_n19907_ = ~new_n19905_ | ~new_n19906_ | ~new_n19831_;
  assign new_n19908_ = pi417 | new_n5681_;
  assign new_n19909_ = pi419 | new_n5687_;
  assign new_n19910_ = ~new_n19828_ | ~new_n19908_ | ~new_n19748_;
  assign new_n19911_ = ~new_n19909_ | ~new_n19907_;
  assign new_n19912_ = ~new_n19827_;
  assign new_n19913_ = pi420 | new_n5690_;
  assign new_n19914_ = ~new_n19913_ | ~new_n19827_;
  assign new_n19915_ = ~new_n5690_ | ~pi420;
  assign new_n19916_ = ~new_n19826_;
  assign new_n19917_ = pi421 | new_n5693_;
  assign new_n19918_ = ~new_n19917_ | ~new_n19826_;
  assign new_n19919_ = ~new_n5693_ | ~pi421;
  assign new_n19920_ = ~new_n19806_;
  assign new_n19921_ = new_n5699_ | pi423;
  assign new_n19922_ = new_n5696_ | pi422;
  assign new_n19923_ = ~new_n19787_;
  assign new_n19924_ = ~new_n19788_ | ~new_n19787_;
  assign new_n19925_ = ~new_n5699_ | ~new_n19924_;
  assign new_n19926_ = ~pi423 | ~new_n19923_;
  assign new_n19927_ = ~new_n19749_ | ~new_n19806_;
  assign new_n19928_ = ~new_n19805_;
  assign new_n19929_ = pi424 | new_n5702_;
  assign new_n19930_ = ~new_n19929_ | ~new_n19805_;
  assign new_n19931_ = ~new_n5702_ | ~pi424;
  assign new_n19932_ = ~new_n20000_ | ~new_n19930_ | ~new_n19931_ | ~new_n20001_;
  assign new_n19933_ = ~new_n5702_ | ~pi424;
  assign new_n19934_ = ~new_n19928_ | ~new_n19933_;
  assign new_n19935_ = new_n5702_ | pi424;
  assign new_n19936_ = ~new_n19934_ | ~new_n19935_ | ~new_n20004_;
  assign new_n19937_ = pi422 | new_n5696_;
  assign new_n19938_ = ~new_n19937_ | ~new_n19806_;
  assign new_n19939_ = ~new_n20012_ | ~new_n19938_ | ~new_n19787_ | ~new_n20013_;
  assign new_n19940_ = ~new_n19920_ | ~new_n19787_;
  assign new_n19941_ = ~pi423 | ~new_n5699_;
  assign new_n19942_ = ~new_n19940_ | ~new_n19941_ | ~new_n19749_;
  assign new_n19943_ = new_n5696_ | pi422;
  assign new_n19944_ = ~new_n19908_ | ~new_n19828_;
  assign new_n19945_ = ~new_n19807_;
  assign new_n19946_ = pi418 | new_n5684_;
  assign new_n19947_ = ~new_n19946_ | ~new_n19807_;
  assign new_n19948_ = ~new_n20033_ | ~new_n19947_ | ~new_n19831_ | ~new_n20034_;
  assign new_n19949_ = ~new_n19945_ | ~new_n19831_;
  assign new_n19950_ = ~new_n5687_ | ~pi419;
  assign new_n19951_ = ~new_n19949_ | ~new_n19950_ | ~new_n19748_;
  assign new_n19952_ = new_n5684_ | pi418;
  assign new_n19953_ = pi415 | new_n5675_;
  assign new_n19954_ = ~new_n19953_ | ~new_n19778_;
  assign new_n19955_ = ~new_n20045_ | ~new_n19954_ | ~new_n19830_ | ~new_n20046_;
  assign new_n19956_ = ~new_n19862_ | ~new_n19830_;
  assign new_n19957_ = ~new_n5678_ | ~pi416;
  assign new_n19958_ = ~new_n19956_ | ~new_n19957_ | ~new_n19747_;
  assign new_n19959_ = ~new_n19863_ | ~new_n19830_;
  assign new_n19960_ = ~new_n19860_ | ~new_n19789_;
  assign new_n19961_ = ~new_n19870_ | ~new_n19760_;
  assign new_n19962_ = ~new_n19884_ | ~new_n19772_;
  assign new_n19963_ = ~new_n19887_ | ~new_n19836_;
  assign new_n19964_ = ~new_n19943_ | ~new_n19787_;
  assign new_n19965_ = ~new_n19952_ | ~new_n19831_;
  assign new_n19966_ = ~new_n19908_ | ~new_n19796_;
  assign new_n19967_ = ~new_n5675_ | ~new_n19777_;
  assign new_n19968_ = ~pi415 | ~new_n19776_;
  assign new_n19969_ = ~new_n19968_ | ~new_n19967_;
  assign new_n19970_ = ~new_n19959_ | ~new_n19778_;
  assign new_n19971_ = ~new_n19969_ | ~new_n19862_;
  assign new_n19972_ = ~new_n5672_ | ~new_n19774_;
  assign new_n19973_ = ~pi414 | ~new_n19775_;
  assign new_n19974_ = ~new_n19973_ | ~new_n19972_;
  assign new_n19975_ = ~new_n19960_ | ~new_n19821_;
  assign new_n19976_ = ~new_n19859_ | ~new_n19974_;
  assign new_n19977_ = ~new_n5669_ | ~new_n19761_;
  assign new_n19978_ = ~pi413 | ~new_n19759_;
  assign new_n19979_ = ~new_n5666_ | ~new_n19757_;
  assign new_n19980_ = ~pi412 | ~new_n19758_;
  assign new_n19981_ = ~new_n19980_ | ~new_n19979_;
  assign new_n19982_ = ~new_n19961_ | ~new_n19779_;
  assign new_n19983_ = ~new_n19981_ | ~new_n19851_;
  assign new_n19984_ = ~new_n5663_ | ~new_n19773_;
  assign new_n19985_ = ~pi411 | ~new_n19764_;
  assign new_n19986_ = ~new_n5660_ | ~new_n19762_;
  assign new_n19987_ = ~pi410 | ~new_n19763_;
  assign new_n19988_ = ~new_n19987_ | ~new_n19986_;
  assign new_n19989_ = ~new_n19962_ | ~new_n19782_;
  assign new_n19990_ = ~new_n19988_ | ~new_n19877_;
  assign new_n19991_ = ~new_n5657_ | ~new_n19770_;
  assign new_n19992_ = ~pi409 | ~new_n19771_;
  assign new_n19993_ = ~new_n19992_ | ~new_n19991_;
  assign new_n19994_ = ~new_n19963_ | ~new_n19822_;
  assign new_n19995_ = ~new_n19886_ | ~new_n19993_;
  assign new_n19996_ = ~new_n5654_ | ~new_n19765_;
  assign new_n19997_ = ~pi408 | ~new_n19766_;
  assign new_n19998_ = ~new_n19838_ | ~new_n19823_;
  assign new_n19999_ = ~new_n19893_ | ~new_n19769_;
  assign new_n20000_ = ~new_n5644_ | ~new_n19825_;
  assign new_n20001_ = ~pi425 | ~new_n19824_;
  assign new_n20002_ = ~new_n5644_ | ~new_n19825_;
  assign new_n20003_ = ~pi425 | ~new_n19824_;
  assign new_n20004_ = ~new_n20003_ | ~new_n20002_;
  assign new_n20005_ = ~new_n5702_ | ~new_n19803_;
  assign new_n20006_ = ~pi424 | ~new_n19804_;
  assign new_n20007_ = ~new_n5702_ | ~new_n19803_;
  assign new_n20008_ = ~pi424 | ~new_n19804_;
  assign new_n20009_ = ~new_n20008_ | ~new_n20007_;
  assign new_n20010_ = ~new_n19805_ | ~new_n20006_ | ~new_n20005_;
  assign new_n20011_ = ~new_n20009_ | ~new_n19928_;
  assign new_n20012_ = ~new_n5699_ | ~new_n19788_;
  assign new_n20013_ = ~pi423 | ~new_n19786_;
  assign new_n20014_ = ~new_n5696_ | ~new_n19784_;
  assign new_n20015_ = ~pi422 | ~new_n19785_;
  assign new_n20016_ = ~new_n20015_ | ~new_n20014_;
  assign new_n20017_ = ~new_n19964_ | ~new_n19806_;
  assign new_n20018_ = ~new_n20016_ | ~new_n19920_;
  assign new_n20019_ = ~new_n5693_ | ~new_n19801_;
  assign new_n20020_ = ~pi421 | ~new_n19802_;
  assign new_n20021_ = ~new_n5693_ | ~new_n19801_;
  assign new_n20022_ = ~pi421 | ~new_n19802_;
  assign new_n20023_ = ~new_n20022_ | ~new_n20021_;
  assign new_n20024_ = ~new_n19826_ | ~new_n20020_ | ~new_n20019_;
  assign new_n20025_ = ~new_n19916_ | ~new_n20023_;
  assign new_n20026_ = ~new_n5690_ | ~new_n19799_;
  assign new_n20027_ = ~pi420 | ~new_n19800_;
  assign new_n20028_ = ~new_n5690_ | ~new_n19799_;
  assign new_n20029_ = ~pi420 | ~new_n19800_;
  assign new_n20030_ = ~new_n20029_ | ~new_n20028_;
  assign new_n20031_ = ~new_n19827_ | ~new_n20027_ | ~new_n20026_;
  assign new_n20032_ = ~new_n19912_ | ~new_n20030_;
  assign new_n20033_ = ~new_n5687_ | ~new_n19797_;
  assign new_n20034_ = ~pi419 | ~new_n19798_;
  assign new_n20035_ = ~new_n5684_ | ~new_n19792_;
  assign new_n20036_ = ~pi418 | ~new_n19793_;
  assign new_n20037_ = ~new_n20036_ | ~new_n20035_;
  assign new_n20038_ = ~new_n19965_ | ~new_n19807_;
  assign new_n20039_ = ~new_n20037_ | ~new_n19945_;
  assign new_n20040_ = ~new_n5681_ | ~new_n19794_;
  assign new_n20041_ = ~pi417 | ~new_n19795_;
  assign new_n20042_ = ~new_n20041_ | ~new_n20040_;
  assign new_n20043_ = ~new_n19966_ | ~new_n19828_;
  assign new_n20044_ = ~new_n19902_ | ~new_n20042_;
  assign new_n20045_ = ~new_n5678_ | ~new_n19790_;
  assign new_n20046_ = ~pi416 | ~new_n19791_;
  assign new_n20047_ = ~new_n5645_ | ~new_n19767_;
  assign new_n20048_ = ~pi406 | ~new_n19768_;
  assign new_n20049_ = new_n20178_ & new_n20078_;
  assign new_n20050_ = new_n20176_ & new_n20079_;
  assign new_n20051_ = new_n20175_ & new_n20080_;
  assign new_n20052_ = new_n20174_ & new_n20081_;
  assign new_n20053_ = new_n20172_ & new_n20082_;
  assign new_n20054_ = new_n20171_ & new_n20083_;
  assign new_n20055_ = new_n20170_ & new_n20084_;
  assign new_n20056_ = new_n20168_ & new_n20085_;
  assign new_n20057_ = new_n20166_ & new_n20086_;
  assign new_n20058_ = new_n20164_ & new_n20087_;
  assign new_n20059_ = new_n20162_ & new_n20088_;
  assign new_n20060_ = new_n20160_ & new_n20089_;
  assign new_n20061_ = new_n20158_ & new_n20068_;
  assign new_n20062_ = new_n20156_ & new_n20110_;
  assign new_n20063_ = new_n20141_ & new_n20069_;
  assign new_n20064_ = new_n20140_ & new_n20070_;
  assign new_n20065_ = new_n20139_ & new_n20071_;
  assign new_n20066_ = new_n20137_ & new_n20072_;
  assign new_n20067_ = new_n20136_ & new_n20073_;
  assign new_n20068_ = new_n5655_ | new_n5652_ | new_n5647_;
  assign new_n20069_ = ~new_n20130_ | ~new_n20077_;
  assign new_n20070_ = ~new_n20131_ | ~new_n20076_;
  assign new_n20071_ = ~new_n20099_ | ~new_n20132_;
  assign new_n20072_ = ~new_n20133_ | ~new_n20075_;
  assign new_n20073_ = ~new_n20134_ | ~new_n20074_;
  assign new_n20074_ = ~new_n5673_;
  assign new_n20075_ = ~new_n5670_;
  assign new_n20076_ = ~new_n5661_;
  assign new_n20077_ = ~new_n5658_;
  assign new_n20078_ = ~new_n20100_ | ~new_n20135_;
  assign new_n20079_ = ~new_n20142_ | ~new_n20097_;
  assign new_n20080_ = ~new_n20143_ | ~new_n20096_;
  assign new_n20081_ = ~new_n20101_ | ~new_n20144_;
  assign new_n20082_ = ~new_n20145_ | ~new_n20095_;
  assign new_n20083_ = ~new_n20146_ | ~new_n20094_;
  assign new_n20084_ = ~new_n20102_ | ~new_n20147_;
  assign new_n20085_ = ~new_n20103_ | ~new_n20148_;
  assign new_n20086_ = ~new_n20104_ | ~new_n20149_;
  assign new_n20087_ = ~new_n20093_ | ~new_n20150_ | ~new_n20118_;
  assign new_n20088_ = ~new_n20092_ | ~new_n20151_ | ~new_n20116_;
  assign new_n20089_ = ~new_n20091_ | ~new_n20152_ | ~new_n20114_;
  assign new_n20090_ = ~new_n6179_;
  assign new_n20091_ = ~new_n6169_;
  assign new_n20092_ = ~new_n6171_;
  assign new_n20093_ = ~new_n6173_;
  assign new_n20094_ = ~new_n5697_;
  assign new_n20095_ = ~new_n5694_;
  assign new_n20096_ = ~new_n5685_;
  assign new_n20097_ = ~new_n5682_;
  assign new_n20098_ = ~new_n20196_ | ~new_n20195_;
  assign new_n20099_ = ~new_n5664_ & ~new_n5667_;
  assign new_n20100_ = ~new_n5679_ & ~new_n5676_;
  assign new_n20101_ = ~new_n5688_ & ~new_n5691_;
  assign new_n20102_ = ~new_n5700_ & ~new_n5703_;
  assign new_n20103_ = ~new_n5705_ & ~new_n6177_;
  assign new_n20104_ = ~new_n6176_ & ~new_n6175_;
  assign new_n20105_ = ~new_n5676_;
  assign new_n20106_ = new_n20180_ & new_n20179_;
  assign new_n20107_ = ~new_n5664_;
  assign new_n20108_ = new_n20182_ & new_n20181_;
  assign new_n20109_ = ~new_n6178_;
  assign new_n20110_ = ~new_n20090_ | ~new_n20153_ | ~new_n20112_;
  assign new_n20111_ = new_n20184_ & new_n20183_;
  assign new_n20112_ = ~new_n6180_;
  assign new_n20113_ = new_n20186_ & new_n20185_;
  assign new_n20114_ = ~new_n6170_;
  assign new_n20115_ = new_n20188_ & new_n20187_;
  assign new_n20116_ = ~new_n6172_;
  assign new_n20117_ = new_n20190_ & new_n20189_;
  assign new_n20118_ = ~new_n6174_;
  assign new_n20119_ = new_n20192_ & new_n20191_;
  assign new_n20120_ = ~new_n6176_;
  assign new_n20121_ = new_n20194_ & new_n20193_;
  assign new_n20122_ = ~new_n5652_;
  assign new_n20123_ = ~new_n5647_;
  assign new_n20124_ = ~new_n5705_;
  assign new_n20125_ = new_n20198_ & new_n20197_;
  assign new_n20126_ = ~new_n5700_;
  assign new_n20127_ = new_n20200_ & new_n20199_;
  assign new_n20128_ = ~new_n5688_;
  assign new_n20129_ = new_n20202_ & new_n20201_;
  assign new_n20130_ = ~new_n20068_;
  assign new_n20131_ = ~new_n20069_;
  assign new_n20132_ = ~new_n20070_;
  assign new_n20133_ = ~new_n20071_;
  assign new_n20134_ = ~new_n20072_;
  assign new_n20135_ = ~new_n20073_;
  assign new_n20136_ = ~new_n5673_ | ~new_n20072_;
  assign new_n20137_ = ~new_n5670_ | ~new_n20071_;
  assign new_n20138_ = ~new_n20132_ | ~new_n20107_;
  assign new_n20139_ = ~new_n5667_ | ~new_n20138_;
  assign new_n20140_ = ~new_n5661_ | ~new_n20069_;
  assign new_n20141_ = ~new_n5658_ | ~new_n20068_;
  assign new_n20142_ = ~new_n20078_;
  assign new_n20143_ = ~new_n20079_;
  assign new_n20144_ = ~new_n20080_;
  assign new_n20145_ = ~new_n20081_;
  assign new_n20146_ = ~new_n20082_;
  assign new_n20147_ = ~new_n20083_;
  assign new_n20148_ = ~new_n20084_;
  assign new_n20149_ = ~new_n20085_;
  assign new_n20150_ = ~new_n20086_;
  assign new_n20151_ = ~new_n20087_;
  assign new_n20152_ = ~new_n20088_;
  assign new_n20153_ = ~new_n20089_;
  assign new_n20154_ = ~new_n20110_;
  assign new_n20155_ = ~new_n20153_ | ~new_n20112_;
  assign new_n20156_ = ~new_n6179_ | ~new_n20155_;
  assign new_n20157_ = new_n5652_ | new_n5647_;
  assign new_n20158_ = ~new_n5655_ | ~new_n20157_;
  assign new_n20159_ = ~new_n20152_ | ~new_n20114_;
  assign new_n20160_ = ~new_n6169_ | ~new_n20159_;
  assign new_n20161_ = ~new_n20151_ | ~new_n20116_;
  assign new_n20162_ = ~new_n6171_ | ~new_n20161_;
  assign new_n20163_ = ~new_n20150_ | ~new_n20118_;
  assign new_n20164_ = ~new_n6173_ | ~new_n20163_;
  assign new_n20165_ = ~new_n20149_ | ~new_n20120_;
  assign new_n20166_ = ~new_n6175_ | ~new_n20165_;
  assign new_n20167_ = ~new_n20148_ | ~new_n20124_;
  assign new_n20168_ = ~new_n6177_ | ~new_n20167_;
  assign new_n20169_ = ~new_n20147_ | ~new_n20126_;
  assign new_n20170_ = ~new_n5703_ | ~new_n20169_;
  assign new_n20171_ = ~new_n5697_ | ~new_n20082_;
  assign new_n20172_ = ~new_n5694_ | ~new_n20081_;
  assign new_n20173_ = ~new_n20144_ | ~new_n20128_;
  assign new_n20174_ = ~new_n5691_ | ~new_n20173_;
  assign new_n20175_ = ~new_n5685_ | ~new_n20079_;
  assign new_n20176_ = ~new_n5682_ | ~new_n20078_;
  assign new_n20177_ = ~new_n20135_ | ~new_n20105_;
  assign new_n20178_ = ~new_n5679_ | ~new_n20177_;
  assign new_n20179_ = ~new_n5676_ | ~new_n20073_;
  assign new_n20180_ = ~new_n20135_ | ~new_n20105_;
  assign new_n20181_ = ~new_n5664_ | ~new_n20070_;
  assign new_n20182_ = ~new_n20132_ | ~new_n20107_;
  assign new_n20183_ = ~new_n6178_ | ~new_n20110_;
  assign new_n20184_ = ~new_n20154_ | ~new_n20109_;
  assign new_n20185_ = ~new_n6180_ | ~new_n20089_;
  assign new_n20186_ = ~new_n20153_ | ~new_n20112_;
  assign new_n20187_ = ~new_n6170_ | ~new_n20088_;
  assign new_n20188_ = ~new_n20152_ | ~new_n20114_;
  assign new_n20189_ = ~new_n6172_ | ~new_n20087_;
  assign new_n20190_ = ~new_n20151_ | ~new_n20116_;
  assign new_n20191_ = ~new_n6174_ | ~new_n20086_;
  assign new_n20192_ = ~new_n20150_ | ~new_n20118_;
  assign new_n20193_ = ~new_n6176_ | ~new_n20085_;
  assign new_n20194_ = ~new_n20149_ | ~new_n20120_;
  assign new_n20195_ = ~new_n5652_ | ~new_n20123_;
  assign new_n20196_ = ~new_n5647_ | ~new_n20122_;
  assign new_n20197_ = ~new_n5705_ | ~new_n20084_;
  assign new_n20198_ = ~new_n20148_ | ~new_n20124_;
  assign new_n20199_ = ~new_n5700_ | ~new_n20083_;
  assign new_n20200_ = ~new_n20147_ | ~new_n20126_;
  assign new_n20201_ = ~new_n5688_ | ~new_n20080_;
  assign new_n20202_ = ~new_n20144_ | ~new_n20128_;
  assign new_n20203_ = new_n20399_ & new_n20398_;
  assign new_n20204_ = new_n20438_ & new_n20437_;
  assign new_n20205_ = new_n20378_ & new_n20453_;
  assign new_n20206_ = new_n20455_ & new_n20454_;
  assign new_n20207_ = new_n20379_ & new_n20479_;
  assign new_n20208_ = new_n20481_ & new_n20480_;
  assign new_n20209_ = ~new_n20541_ | ~new_n20544_;
  assign new_n20210_ = ~new_n20530_ | ~new_n20533_;
  assign new_n20211_ = ~new_n20519_ | ~new_n20522_;
  assign new_n20212_ = ~new_n20511_ | ~new_n20513_;
  assign new_n20213_ = ~new_n20549_ | ~new_n20509_;
  assign new_n20214_ = ~new_n20432_ | ~new_n20434_;
  assign new_n20215_ = ~new_n20424_ | ~new_n20427_;
  assign new_n20216_ = ~new_n20416_ | ~new_n20418_;
  assign new_n20217_ = ~new_n20363_ | ~new_n20547_;
  assign new_n20218_ = ~new_n5670_;
  assign new_n20219_ = ~new_n5664_;
  assign new_n20220_ = ~new_n5655_;
  assign new_n20221_ = ~new_n5647_;
  assign new_n20222_ = ~new_n5300_;
  assign new_n20223_ = ~new_n5658_;
  assign new_n20224_ = ~new_n5290_;
  assign new_n20225_ = ~new_n5290_ | ~new_n20220_;
  assign new_n20226_ = ~new_n5286_;
  assign new_n20227_ = ~new_n5667_;
  assign new_n20228_ = ~new_n5661_;
  assign new_n20229_ = ~new_n5293_;
  assign new_n20230_ = ~new_n5289_;
  assign new_n20231_ = ~new_n5282_;
  assign new_n20232_ = ~new_n5282_ | ~new_n20228_;
  assign new_n20233_ = ~new_n5673_;
  assign new_n20234_ = ~new_n5292_;
  assign new_n20235_ = ~new_n5292_ | ~new_n20218_;
  assign new_n20236_ = ~new_n5306_;
  assign new_n20237_ = ~new_n5676_;
  assign new_n20238_ = ~new_n5305_;
  assign new_n20239_ = ~new_n20405_ | ~new_n20404_;
  assign new_n20240_ = ~new_n20232_ | ~new_n20420_;
  assign new_n20241_ = ~new_n20548_ | ~new_n20389_ | ~new_n20373_;
  assign new_n20242_ = ~new_n6171_;
  assign new_n20243_ = ~new_n5679_;
  assign new_n20244_ = ~new_n5682_;
  assign new_n20245_ = ~new_n5285_;
  assign new_n20246_ = ~new_n5284_;
  assign new_n20247_ = ~new_n5305_ | ~new_n20237_;
  assign new_n20248_ = ~new_n5685_;
  assign new_n20249_ = ~new_n5294_;
  assign new_n20250_ = ~new_n5688_;
  assign new_n20251_ = ~new_n5302_;
  assign new_n20252_ = ~new_n5697_;
  assign new_n20253_ = ~new_n5694_;
  assign new_n20254_ = ~new_n5691_;
  assign new_n20255_ = ~new_n5295_;
  assign new_n20256_ = ~new_n5296_;
  assign new_n20257_ = ~new_n5301_;
  assign new_n20258_ = ~new_n5301_ | ~new_n20254_;
  assign new_n20259_ = ~new_n5700_;
  assign new_n20260_ = ~new_n5291_;
  assign new_n20261_ = ~new_n20465_ | ~new_n20464_;
  assign new_n20262_ = ~new_n5304_;
  assign new_n20263_ = ~new_n5705_;
  assign new_n20264_ = ~new_n5303_;
  assign new_n20265_ = ~new_n6177_;
  assign new_n20266_ = ~new_n5298_;
  assign new_n20267_ = ~new_n6174_;
  assign new_n20268_ = ~new_n6175_;
  assign new_n20269_ = ~new_n6176_;
  assign new_n20270_ = ~new_n5288_;
  assign new_n20271_ = ~new_n5283_;
  assign new_n20272_ = ~new_n5297_;
  assign new_n20273_ = ~new_n5297_ | ~new_n20269_;
  assign new_n20274_ = ~new_n6173_;
  assign new_n20275_ = ~new_n5287_;
  assign new_n20276_ = ~new_n6172_;
  assign new_n20277_ = ~new_n5280_;
  assign new_n20278_ = ~new_n6170_;
  assign new_n20279_ = ~new_n5279_;
  assign new_n20280_ = ~new_n5279_ | ~new_n20242_;
  assign new_n20281_ = ~new_n5275_;
  assign new_n20282_ = ~new_n6169_;
  assign new_n20283_ = ~new_n5276_;
  assign new_n20284_ = ~new_n20325_ | ~new_n20498_;
  assign new_n20285_ = ~new_n20495_ | ~new_n20494_;
  assign new_n20286_ = ~new_n20273_ | ~new_n20515_;
  assign new_n20287_ = ~new_n20258_ | ~new_n20526_;
  assign new_n20288_ = ~new_n20247_ | ~new_n20537_;
  assign new_n20289_ = ~new_n5299_;
  assign new_n20290_ = ~new_n20592_ | ~new_n20591_;
  assign new_n20291_ = ~new_n20606_ | ~new_n20605_;
  assign new_n20292_ = ~new_n20611_ | ~new_n20610_;
  assign new_n20293_ = ~new_n20627_ | ~new_n20626_;
  assign new_n20294_ = ~new_n20632_ | ~new_n20631_;
  assign new_n20295_ = ~new_n20637_ | ~new_n20636_;
  assign new_n20296_ = ~new_n20642_ | ~new_n20641_;
  assign new_n20297_ = ~new_n20647_ | ~new_n20646_;
  assign new_n20298_ = ~new_n20663_ | ~new_n20662_;
  assign new_n20299_ = ~new_n20668_ | ~new_n20667_;
  assign new_n20300_ = ~new_n20553_ | ~new_n20552_;
  assign new_n20301_ = ~new_n20562_ | ~new_n20561_;
  assign new_n20302_ = ~new_n20569_ | ~new_n20568_;
  assign new_n20303_ = ~new_n20573_ | ~new_n20572_;
  assign new_n20304_ = ~new_n20582_ | ~new_n20581_;
  assign new_n20305_ = ~new_n20601_ | ~new_n20600_;
  assign new_n20306_ = ~new_n20618_ | ~new_n20617_;
  assign new_n20307_ = ~new_n20622_ | ~new_n20621_;
  assign new_n20308_ = ~new_n20654_ | ~new_n20653_;
  assign new_n20309_ = ~new_n20658_ | ~new_n20657_;
  assign new_n20310_ = ~new_n20675_ | ~new_n20674_;
  assign new_n20311_ = new_n20391_ & new_n20381_;
  assign new_n20312_ = new_n20394_ & new_n20395_;
  assign new_n20313_ = new_n20382_ & new_n20402_ & new_n20397_;
  assign new_n20314_ = new_n20407_ & new_n20383_;
  assign new_n20315_ = new_n20410_ & new_n20411_;
  assign new_n20316_ = new_n20235_ & new_n20555_ & new_n20554_;
  assign new_n20317_ = new_n20558_ & new_n20383_;
  assign new_n20318_ = new_n20426_ & new_n20203_;
  assign new_n20319_ = new_n20565_ & new_n20382_;
  assign new_n20320_ = new_n20225_ & new_n20575_ & new_n20574_;
  assign new_n20321_ = new_n20578_ & new_n20381_;
  assign new_n20322_ = new_n20377_ & new_n20436_ & new_n20413_;
  assign new_n20323_ = new_n20458_ & new_n20205_;
  assign new_n20324_ = new_n20484_ & new_n20207_;
  assign new_n20325_ = new_n20500_ & new_n20501_;
  assign new_n20326_ = new_n20508_ & new_n20584_ & new_n20583_;
  assign new_n20327_ = new_n20505_ & new_n20587_;
  assign new_n20328_ = ~new_n20589_ | ~new_n20588_;
  assign new_n20329_ = new_n20280_ & new_n20594_ & new_n20593_;
  assign new_n20330_ = new_n20597_ & new_n20380_;
  assign new_n20331_ = ~new_n20603_ | ~new_n20602_;
  assign new_n20332_ = ~new_n20608_ | ~new_n20607_;
  assign new_n20333_ = new_n20521_ & new_n20208_;
  assign new_n20334_ = new_n20614_ & new_n20379_;
  assign new_n20335_ = ~new_n20624_ | ~new_n20623_;
  assign new_n20336_ = ~new_n20629_ | ~new_n20628_;
  assign new_n20337_ = ~new_n20634_ | ~new_n20633_;
  assign new_n20338_ = ~new_n20639_ | ~new_n20638_;
  assign new_n20339_ = ~new_n20644_ | ~new_n20643_;
  assign new_n20340_ = new_n20532_ & new_n20206_;
  assign new_n20341_ = new_n20650_ & new_n20378_;
  assign new_n20342_ = ~new_n20660_ | ~new_n20659_;
  assign new_n20343_ = ~new_n20665_ | ~new_n20664_;
  assign new_n20344_ = new_n20543_ & new_n20204_;
  assign new_n20345_ = new_n20671_ & new_n20377_;
  assign new_n20346_ = new_n20551_ & new_n20550_;
  assign new_n20347_ = ~new_n20315_ | ~new_n20408_;
  assign new_n20348_ = new_n20560_ & new_n20559_;
  assign new_n20349_ = new_n20567_ & new_n20566_;
  assign new_n20350_ = new_n20571_ & new_n20570_;
  assign new_n20351_ = ~new_n20312_ | ~new_n20392_;
  assign new_n20352_ = new_n20580_ & new_n20579_;
  assign new_n20353_ = ~new_n6180_;
  assign new_n20354_ = ~new_n5277_;
  assign new_n20355_ = new_n20599_ & new_n20598_;
  assign new_n20356_ = ~new_n20491_ | ~new_n20490_;
  assign new_n20357_ = ~new_n20487_ | ~new_n20486_;
  assign new_n20358_ = new_n20616_ & new_n20615_;
  assign new_n20359_ = new_n20620_ & new_n20619_;
  assign new_n20360_ = ~new_n20477_ | ~new_n20476_;
  assign new_n20361_ = ~new_n20473_ | ~new_n20472_;
  assign new_n20362_ = ~new_n5652_;
  assign new_n20363_ = ~new_n5647_ | ~new_n20289_;
  assign new_n20364_ = ~new_n20469_ | ~new_n20468_;
  assign new_n20365_ = ~new_n5703_;
  assign new_n20366_ = ~new_n20461_ | ~new_n20460_;
  assign new_n20367_ = new_n20652_ & new_n20651_;
  assign new_n20368_ = new_n20656_ & new_n20655_;
  assign new_n20369_ = ~new_n20451_ | ~new_n20450_;
  assign new_n20370_ = ~new_n20447_ | ~new_n20446_;
  assign new_n20371_ = ~new_n20443_ | ~new_n20442_;
  assign new_n20372_ = new_n20673_ & new_n20672_;
  assign new_n20373_ = ~new_n20363_ | ~new_n20362_;
  assign new_n20374_ = ~new_n20280_;
  assign new_n20375_ = ~new_n20225_;
  assign new_n20376_ = ~new_n20235_;
  assign new_n20377_ = ~new_n5679_ | ~new_n20246_;
  assign new_n20378_ = ~new_n5694_ | ~new_n20256_;
  assign new_n20379_ = ~new_n6175_ | ~new_n20271_;
  assign new_n20380_ = ~new_n6171_ | ~new_n20279_;
  assign new_n20381_ = ~new_n5655_ | ~new_n20224_;
  assign new_n20382_ = ~new_n5664_ | ~new_n20230_;
  assign new_n20383_ = ~new_n5670_ | ~new_n20234_;
  assign new_n20384_ = ~new_n20258_;
  assign new_n20385_ = ~new_n20273_;
  assign new_n20386_ = ~new_n20232_;
  assign new_n20387_ = ~new_n20247_;
  assign new_n20388_ = ~new_n20363_;
  assign new_n20389_ = ~new_n5300_ | ~new_n20363_;
  assign new_n20390_ = ~new_n20241_;
  assign new_n20391_ = ~new_n5658_ | ~new_n20226_;
  assign new_n20392_ = ~new_n20311_ | ~new_n20241_;
  assign new_n20393_ = ~new_n20226_ | ~new_n20225_;
  assign new_n20394_ = ~new_n20393_ | ~new_n20223_;
  assign new_n20395_ = ~new_n5286_ | ~new_n20375_;
  assign new_n20396_ = ~new_n20351_;
  assign new_n20397_ = ~new_n5667_ | ~new_n20229_;
  assign new_n20398_ = ~new_n5293_ | ~new_n20227_;
  assign new_n20399_ = ~new_n5289_ | ~new_n20219_;
  assign new_n20400_ = ~new_n20386_ | ~new_n20382_;
  assign new_n20401_ = ~new_n20203_ | ~new_n20400_;
  assign new_n20402_ = ~new_n5661_ | ~new_n20231_;
  assign new_n20403_ = ~new_n5667_ | ~new_n20229_;
  assign new_n20404_ = ~new_n20351_ | ~new_n20313_;
  assign new_n20405_ = ~new_n20403_ | ~new_n20401_;
  assign new_n20406_ = ~new_n20239_;
  assign new_n20407_ = ~new_n5673_ | ~new_n20236_;
  assign new_n20408_ = ~new_n20314_ | ~new_n20239_;
  assign new_n20409_ = ~new_n20236_ | ~new_n20235_;
  assign new_n20410_ = ~new_n20409_ | ~new_n20233_;
  assign new_n20411_ = ~new_n5306_ | ~new_n20376_;
  assign new_n20412_ = ~new_n20347_;
  assign new_n20413_ = ~new_n5676_ | ~new_n20238_;
  assign new_n20414_ = ~new_n20413_ | ~new_n20247_;
  assign new_n20415_ = ~new_n20406_ | ~new_n20235_;
  assign new_n20416_ = ~new_n20317_ | ~new_n20415_;
  assign new_n20417_ = ~new_n20239_ | ~new_n20383_;
  assign new_n20418_ = ~new_n20316_ | ~new_n20417_;
  assign new_n20419_ = ~new_n20235_ | ~new_n20383_;
  assign new_n20420_ = ~new_n20402_ | ~new_n20351_;
  assign new_n20421_ = ~new_n20240_;
  assign new_n20422_ = ~new_n5289_ | ~new_n20219_;
  assign new_n20423_ = ~new_n20421_ | ~new_n20422_;
  assign new_n20424_ = ~new_n20319_ | ~new_n20423_;
  assign new_n20425_ = ~new_n20240_ | ~new_n20382_;
  assign new_n20426_ = ~new_n5667_ | ~new_n20229_;
  assign new_n20427_ = ~new_n20318_ | ~new_n20425_;
  assign new_n20428_ = ~new_n5289_ | ~new_n20219_;
  assign new_n20429_ = ~new_n20382_ | ~new_n20428_;
  assign new_n20430_ = ~new_n20402_ | ~new_n20232_;
  assign new_n20431_ = ~new_n20390_ | ~new_n20225_;
  assign new_n20432_ = ~new_n20321_ | ~new_n20431_;
  assign new_n20433_ = ~new_n20241_ | ~new_n20381_;
  assign new_n20434_ = ~new_n20320_ | ~new_n20433_;
  assign new_n20435_ = ~new_n20225_ | ~new_n20381_;
  assign new_n20436_ = ~new_n5682_ | ~new_n20245_;
  assign new_n20437_ = ~new_n5285_ | ~new_n20244_;
  assign new_n20438_ = ~new_n5284_ | ~new_n20243_;
  assign new_n20439_ = ~new_n20387_ | ~new_n20377_;
  assign new_n20440_ = ~new_n20204_ | ~new_n20439_;
  assign new_n20441_ = ~new_n5682_ | ~new_n20245_;
  assign new_n20442_ = ~new_n20347_ | ~new_n20322_;
  assign new_n20443_ = ~new_n20441_ | ~new_n20440_;
  assign new_n20444_ = ~new_n20371_;
  assign new_n20445_ = ~new_n5685_ | ~new_n20249_;
  assign new_n20446_ = ~new_n20445_ | ~new_n20371_;
  assign new_n20447_ = ~new_n5294_ | ~new_n20248_;
  assign new_n20448_ = ~new_n20370_;
  assign new_n20449_ = ~new_n5688_ | ~new_n20251_;
  assign new_n20450_ = ~new_n20449_ | ~new_n20370_;
  assign new_n20451_ = ~new_n5302_ | ~new_n20250_;
  assign new_n20452_ = ~new_n20369_;
  assign new_n20453_ = ~new_n5697_ | ~new_n20255_;
  assign new_n20454_ = ~new_n5295_ | ~new_n20252_;
  assign new_n20455_ = ~new_n5296_ | ~new_n20253_;
  assign new_n20456_ = ~new_n20384_ | ~new_n20205_;
  assign new_n20457_ = ~new_n20206_ | ~new_n20456_;
  assign new_n20458_ = ~new_n5691_ | ~new_n20257_;
  assign new_n20459_ = ~new_n5697_ | ~new_n20255_;
  assign new_n20460_ = ~new_n20323_ | ~new_n20369_;
  assign new_n20461_ = ~new_n20459_ | ~new_n20457_;
  assign new_n20462_ = ~new_n20366_;
  assign new_n20463_ = ~new_n5700_ | ~new_n20260_;
  assign new_n20464_ = ~new_n20463_ | ~new_n20366_;
  assign new_n20465_ = ~new_n5291_ | ~new_n20259_;
  assign new_n20466_ = ~new_n20261_;
  assign new_n20467_ = ~new_n20466_ | ~new_n20262_;
  assign new_n20468_ = ~new_n20467_ | ~new_n20365_;
  assign new_n20469_ = ~new_n5304_ | ~new_n20261_;
  assign new_n20470_ = ~new_n20364_;
  assign new_n20471_ = ~new_n5705_ | ~new_n20264_;
  assign new_n20472_ = ~new_n20471_ | ~new_n20364_;
  assign new_n20473_ = ~new_n5303_ | ~new_n20263_;
  assign new_n20474_ = ~new_n20361_;
  assign new_n20475_ = ~new_n6177_ | ~new_n20266_;
  assign new_n20476_ = ~new_n20475_ | ~new_n20361_;
  assign new_n20477_ = ~new_n5298_ | ~new_n20265_;
  assign new_n20478_ = ~new_n20360_;
  assign new_n20479_ = ~new_n6174_ | ~new_n20270_;
  assign new_n20480_ = ~new_n5288_ | ~new_n20267_;
  assign new_n20481_ = ~new_n5283_ | ~new_n20268_;
  assign new_n20482_ = ~new_n20385_ | ~new_n20207_;
  assign new_n20483_ = ~new_n20208_ | ~new_n20482_;
  assign new_n20484_ = ~new_n6176_ | ~new_n20272_;
  assign new_n20485_ = ~new_n6174_ | ~new_n20270_;
  assign new_n20486_ = ~new_n20324_ | ~new_n20360_;
  assign new_n20487_ = ~new_n20485_ | ~new_n20483_;
  assign new_n20488_ = ~new_n20357_;
  assign new_n20489_ = ~new_n6173_ | ~new_n20275_;
  assign new_n20490_ = ~new_n20489_ | ~new_n20357_;
  assign new_n20491_ = ~new_n5287_ | ~new_n20274_;
  assign new_n20492_ = ~new_n20356_;
  assign new_n20493_ = ~new_n6172_ | ~new_n20277_;
  assign new_n20494_ = ~new_n20493_ | ~new_n20356_;
  assign new_n20495_ = ~new_n5280_ | ~new_n20276_;
  assign new_n20496_ = ~new_n20285_;
  assign new_n20497_ = ~new_n6170_ | ~new_n20281_;
  assign new_n20498_ = ~new_n20497_ | ~new_n20285_ | ~new_n20380_;
  assign new_n20499_ = ~new_n20281_ | ~new_n20280_;
  assign new_n20500_ = ~new_n20499_ | ~new_n20278_;
  assign new_n20501_ = ~new_n5275_ | ~new_n20374_;
  assign new_n20502_ = ~new_n20284_;
  assign new_n20503_ = ~new_n5276_ | ~new_n20282_;
  assign new_n20504_ = ~new_n20502_ | ~new_n20503_;
  assign new_n20505_ = ~new_n6169_ | ~new_n20283_;
  assign new_n20506_ = ~new_n6169_ | ~new_n20283_;
  assign new_n20507_ = ~new_n20506_ | ~new_n20284_;
  assign new_n20508_ = ~new_n5276_ | ~new_n20282_;
  assign new_n20509_ = ~new_n20326_ | ~new_n20507_;
  assign new_n20510_ = ~new_n20496_ | ~new_n20280_;
  assign new_n20511_ = ~new_n20330_ | ~new_n20510_;
  assign new_n20512_ = ~new_n20285_ | ~new_n20380_;
  assign new_n20513_ = ~new_n20329_ | ~new_n20512_;
  assign new_n20514_ = ~new_n20280_ | ~new_n20380_;
  assign new_n20515_ = ~new_n20484_ | ~new_n20360_;
  assign new_n20516_ = ~new_n20286_;
  assign new_n20517_ = ~new_n5283_ | ~new_n20268_;
  assign new_n20518_ = ~new_n20516_ | ~new_n20517_;
  assign new_n20519_ = ~new_n20334_ | ~new_n20518_;
  assign new_n20520_ = ~new_n20286_ | ~new_n20379_;
  assign new_n20521_ = ~new_n6174_ | ~new_n20270_;
  assign new_n20522_ = ~new_n20333_ | ~new_n20520_;
  assign new_n20523_ = ~new_n5283_ | ~new_n20268_;
  assign new_n20524_ = ~new_n20379_ | ~new_n20523_;
  assign new_n20525_ = ~new_n20484_ | ~new_n20273_;
  assign new_n20526_ = ~new_n20458_ | ~new_n20369_;
  assign new_n20527_ = ~new_n20287_;
  assign new_n20528_ = ~new_n5296_ | ~new_n20253_;
  assign new_n20529_ = ~new_n20527_ | ~new_n20528_;
  assign new_n20530_ = ~new_n20341_ | ~new_n20529_;
  assign new_n20531_ = ~new_n20287_ | ~new_n20378_;
  assign new_n20532_ = ~new_n5697_ | ~new_n20255_;
  assign new_n20533_ = ~new_n20340_ | ~new_n20531_;
  assign new_n20534_ = ~new_n5296_ | ~new_n20253_;
  assign new_n20535_ = ~new_n20378_ | ~new_n20534_;
  assign new_n20536_ = ~new_n20458_ | ~new_n20258_;
  assign new_n20537_ = ~new_n20413_ | ~new_n20347_;
  assign new_n20538_ = ~new_n20288_;
  assign new_n20539_ = ~new_n5284_ | ~new_n20243_;
  assign new_n20540_ = ~new_n20538_ | ~new_n20539_;
  assign new_n20541_ = ~new_n20345_ | ~new_n20540_;
  assign new_n20542_ = ~new_n20288_ | ~new_n20377_;
  assign new_n20543_ = ~new_n5682_ | ~new_n20245_;
  assign new_n20544_ = ~new_n20344_ | ~new_n20542_;
  assign new_n20545_ = ~new_n5284_ | ~new_n20243_;
  assign new_n20546_ = ~new_n20377_ | ~new_n20545_;
  assign new_n20547_ = ~new_n5299_ | ~new_n20221_;
  assign new_n20548_ = ~new_n5300_ | ~new_n20362_;
  assign new_n20549_ = ~new_n20327_ | ~new_n20504_;
  assign new_n20550_ = ~new_n5676_ | ~new_n20238_;
  assign new_n20551_ = ~new_n5305_ | ~new_n20237_;
  assign new_n20552_ = ~new_n20414_ | ~new_n20347_;
  assign new_n20553_ = ~new_n20412_ | ~new_n20346_;
  assign new_n20554_ = ~new_n5673_ | ~new_n20236_;
  assign new_n20555_ = ~new_n5306_ | ~new_n20233_;
  assign new_n20556_ = ~new_n5673_ | ~new_n20236_;
  assign new_n20557_ = ~new_n5306_ | ~new_n20233_;
  assign new_n20558_ = ~new_n20557_ | ~new_n20556_;
  assign new_n20559_ = ~new_n5670_ | ~new_n20234_;
  assign new_n20560_ = ~new_n5292_ | ~new_n20218_;
  assign new_n20561_ = ~new_n20419_ | ~new_n20239_;
  assign new_n20562_ = ~new_n20348_ | ~new_n20406_;
  assign new_n20563_ = ~new_n5667_ | ~new_n20229_;
  assign new_n20564_ = ~new_n5293_ | ~new_n20227_;
  assign new_n20565_ = ~new_n20564_ | ~new_n20563_;
  assign new_n20566_ = ~new_n5664_ | ~new_n20230_;
  assign new_n20567_ = ~new_n5289_ | ~new_n20219_;
  assign new_n20568_ = ~new_n20429_ | ~new_n20240_;
  assign new_n20569_ = ~new_n20349_ | ~new_n20421_;
  assign new_n20570_ = ~new_n5661_ | ~new_n20231_;
  assign new_n20571_ = ~new_n5282_ | ~new_n20228_;
  assign new_n20572_ = ~new_n20430_ | ~new_n20351_;
  assign new_n20573_ = ~new_n20396_ | ~new_n20350_;
  assign new_n20574_ = ~new_n5658_ | ~new_n20226_;
  assign new_n20575_ = ~new_n5286_ | ~new_n20223_;
  assign new_n20576_ = ~new_n5658_ | ~new_n20226_;
  assign new_n20577_ = ~new_n5286_ | ~new_n20223_;
  assign new_n20578_ = ~new_n20577_ | ~new_n20576_;
  assign new_n20579_ = ~new_n5655_ | ~new_n20224_;
  assign new_n20580_ = ~new_n5290_ | ~new_n20220_;
  assign new_n20581_ = ~new_n20435_ | ~new_n20241_;
  assign new_n20582_ = ~new_n20352_ | ~new_n20390_;
  assign new_n20583_ = ~new_n6180_ | ~new_n20354_;
  assign new_n20584_ = ~new_n5277_ | ~new_n20353_;
  assign new_n20585_ = ~new_n6180_ | ~new_n20354_;
  assign new_n20586_ = ~new_n5277_ | ~new_n20353_;
  assign new_n20587_ = ~new_n20586_ | ~new_n20585_;
  assign new_n20588_ = ~new_n6169_ | ~new_n20283_;
  assign new_n20589_ = ~new_n5276_ | ~new_n20282_;
  assign new_n20590_ = ~new_n20328_;
  assign new_n20591_ = ~new_n20590_ | ~new_n20502_;
  assign new_n20592_ = ~new_n20328_ | ~new_n20284_;
  assign new_n20593_ = ~new_n6170_ | ~new_n20281_;
  assign new_n20594_ = ~new_n5275_ | ~new_n20278_;
  assign new_n20595_ = ~new_n6170_ | ~new_n20281_;
  assign new_n20596_ = ~new_n5275_ | ~new_n20278_;
  assign new_n20597_ = ~new_n20596_ | ~new_n20595_;
  assign new_n20598_ = ~new_n6171_ | ~new_n20279_;
  assign new_n20599_ = ~new_n5279_ | ~new_n20242_;
  assign new_n20600_ = ~new_n20514_ | ~new_n20285_;
  assign new_n20601_ = ~new_n20355_ | ~new_n20496_;
  assign new_n20602_ = ~new_n6172_ | ~new_n20277_;
  assign new_n20603_ = ~new_n5280_ | ~new_n20276_;
  assign new_n20604_ = ~new_n20331_;
  assign new_n20605_ = ~new_n20492_ | ~new_n20604_;
  assign new_n20606_ = ~new_n20331_ | ~new_n20356_;
  assign new_n20607_ = ~new_n6173_ | ~new_n20275_;
  assign new_n20608_ = ~new_n5287_ | ~new_n20274_;
  assign new_n20609_ = ~new_n20332_;
  assign new_n20610_ = ~new_n20488_ | ~new_n20609_;
  assign new_n20611_ = ~new_n20332_ | ~new_n20357_;
  assign new_n20612_ = ~new_n6174_ | ~new_n20270_;
  assign new_n20613_ = ~new_n5288_ | ~new_n20267_;
  assign new_n20614_ = ~new_n20613_ | ~new_n20612_;
  assign new_n20615_ = ~new_n6175_ | ~new_n20271_;
  assign new_n20616_ = ~new_n5283_ | ~new_n20268_;
  assign new_n20617_ = ~new_n20524_ | ~new_n20286_;
  assign new_n20618_ = ~new_n20358_ | ~new_n20516_;
  assign new_n20619_ = ~new_n6176_ | ~new_n20272_;
  assign new_n20620_ = ~new_n5297_ | ~new_n20269_;
  assign new_n20621_ = ~new_n20525_ | ~new_n20360_;
  assign new_n20622_ = ~new_n20478_ | ~new_n20359_;
  assign new_n20623_ = ~new_n6177_ | ~new_n20266_;
  assign new_n20624_ = ~new_n5298_ | ~new_n20265_;
  assign new_n20625_ = ~new_n20335_;
  assign new_n20626_ = ~new_n20474_ | ~new_n20625_;
  assign new_n20627_ = ~new_n20335_ | ~new_n20361_;
  assign new_n20628_ = ~new_n5652_ | ~new_n20222_;
  assign new_n20629_ = ~new_n5300_ | ~new_n20362_;
  assign new_n20630_ = ~new_n20336_;
  assign new_n20631_ = ~new_n20388_ | ~new_n20630_;
  assign new_n20632_ = ~new_n20336_ | ~new_n20363_;
  assign new_n20633_ = ~new_n5705_ | ~new_n20264_;
  assign new_n20634_ = ~new_n5303_ | ~new_n20263_;
  assign new_n20635_ = ~new_n20337_;
  assign new_n20636_ = ~new_n20470_ | ~new_n20635_;
  assign new_n20637_ = ~new_n20337_ | ~new_n20364_;
  assign new_n20638_ = ~new_n5703_ | ~new_n20262_;
  assign new_n20639_ = ~new_n5304_ | ~new_n20365_;
  assign new_n20640_ = ~new_n20338_;
  assign new_n20641_ = ~new_n20640_ | ~new_n20466_;
  assign new_n20642_ = ~new_n20338_ | ~new_n20261_;
  assign new_n20643_ = ~new_n5700_ | ~new_n20260_;
  assign new_n20644_ = ~new_n5291_ | ~new_n20259_;
  assign new_n20645_ = ~new_n20339_;
  assign new_n20646_ = ~new_n20462_ | ~new_n20645_;
  assign new_n20647_ = ~new_n20339_ | ~new_n20366_;
  assign new_n20648_ = ~new_n5697_ | ~new_n20255_;
  assign new_n20649_ = ~new_n5295_ | ~new_n20252_;
  assign new_n20650_ = ~new_n20649_ | ~new_n20648_;
  assign new_n20651_ = ~new_n5694_ | ~new_n20256_;
  assign new_n20652_ = ~new_n5296_ | ~new_n20253_;
  assign new_n20653_ = ~new_n20535_ | ~new_n20287_;
  assign new_n20654_ = ~new_n20367_ | ~new_n20527_;
  assign new_n20655_ = ~new_n5691_ | ~new_n20257_;
  assign new_n20656_ = ~new_n5301_ | ~new_n20254_;
  assign new_n20657_ = ~new_n20536_ | ~new_n20369_;
  assign new_n20658_ = ~new_n20452_ | ~new_n20368_;
  assign new_n20659_ = ~new_n5688_ | ~new_n20251_;
  assign new_n20660_ = ~new_n5302_ | ~new_n20250_;
  assign new_n20661_ = ~new_n20342_;
  assign new_n20662_ = ~new_n20448_ | ~new_n20661_;
  assign new_n20663_ = ~new_n20342_ | ~new_n20370_;
  assign new_n20664_ = ~new_n5685_ | ~new_n20249_;
  assign new_n20665_ = ~new_n5294_ | ~new_n20248_;
  assign new_n20666_ = ~new_n20343_;
  assign new_n20667_ = ~new_n20444_ | ~new_n20666_;
  assign new_n20668_ = ~new_n20343_ | ~new_n20371_;
  assign new_n20669_ = ~new_n5682_ | ~new_n20245_;
  assign new_n20670_ = ~new_n5285_ | ~new_n20244_;
  assign new_n20671_ = ~new_n20670_ | ~new_n20669_;
  assign new_n20672_ = ~new_n5679_ | ~new_n20246_;
  assign new_n20673_ = ~new_n5284_ | ~new_n20243_;
  assign new_n20674_ = ~new_n20546_ | ~new_n20288_;
  assign new_n20675_ = ~new_n20372_ | ~new_n20538_;
  assign new_n20676_ = new_n20851_ & new_n20850_;
  assign new_n20677_ = new_n20852_ & new_n20853_;
  assign new_n20678_ = new_n20869_ & new_n20868_;
  assign new_n20679_ = new_n20909_ & new_n20908_;
  assign new_n20680_ = new_n20918_ & new_n20917_;
  assign new_n20681_ = new_n20936_ & new_n20935_;
  assign new_n20682_ = new_n20944_ & new_n20943_;
  assign new_n20683_ = new_n21023_ & new_n21020_;
  assign new_n20684_ = new_n21016_ & new_n21013_;
  assign new_n20685_ = new_n21007_ & new_n21004_;
  assign new_n20686_ = new_n20998_ & new_n20995_;
  assign new_n20687_ = new_n20992_ & new_n20990_;
  assign new_n20688_ = new_n20985_ & new_n20982_;
  assign new_n20689_ = new_n20907_ & new_n20904_;
  assign new_n20690_ = new_n20899_ & new_n20896_;
  assign new_n20691_ = new_n20885_ & new_n20882_;
  assign new_n20692_ = ~new_n5667_;
  assign new_n20693_ = ~new_n5293_;
  assign new_n20694_ = ~new_n5292_;
  assign new_n20695_ = ~new_n5293_ | ~new_n5667_;
  assign new_n20696_ = ~new_n5670_;
  assign new_n20697_ = ~new_n5661_;
  assign new_n20698_ = ~new_n5282_;
  assign new_n20699_ = ~new_n5289_;
  assign new_n20700_ = ~new_n5655_;
  assign new_n20701_ = ~new_n5290_;
  assign new_n20702_ = ~new_n5647_;
  assign new_n20703_ = ~new_n5299_;
  assign new_n20704_ = ~new_n5299_ | ~new_n5647_;
  assign new_n20705_ = ~new_n5658_;
  assign new_n20706_ = ~new_n5286_;
  assign new_n20707_ = ~new_n5282_ | ~new_n5661_;
  assign new_n20708_ = ~new_n5664_;
  assign new_n20709_ = ~new_n5673_;
  assign new_n20710_ = ~new_n5306_;
  assign new_n20711_ = ~new_n5305_;
  assign new_n20712_ = ~new_n5676_;
  assign new_n20713_ = ~new_n20734_ | ~new_n20877_;
  assign new_n20714_ = ~new_n20790_ | ~new_n20865_;
  assign new_n20715_ = ~new_n20854_ | ~new_n20855_;
  assign new_n20716_ = ~new_n5652_ | ~new_n5300_;
  assign new_n20717_ = ~new_n20794_ | ~new_n20891_;
  assign new_n20718_ = ~new_n20888_ | ~new_n20887_;
  assign new_n20719_ = ~new_n6170_;
  assign new_n20720_ = ~new_n5275_;
  assign new_n20721_ = ~new_n5279_;
  assign new_n20722_ = ~new_n6171_;
  assign new_n20723_ = ~new_n6172_;
  assign new_n20724_ = ~new_n5280_;
  assign new_n20725_ = ~new_n6173_;
  assign new_n20726_ = ~new_n5287_;
  assign new_n20727_ = ~new_n6176_;
  assign new_n20728_ = ~new_n5297_;
  assign new_n20729_ = ~new_n5697_;
  assign new_n20730_ = ~new_n5295_;
  assign new_n20731_ = ~new_n5291_;
  assign new_n20732_ = ~new_n5295_ | ~new_n5697_;
  assign new_n20733_ = ~new_n5700_;
  assign new_n20734_ = ~new_n5306_ | ~new_n5673_;
  assign new_n20735_ = ~new_n5679_;
  assign new_n20736_ = ~new_n5284_;
  assign new_n20737_ = ~new_n5685_;
  assign new_n20738_ = ~new_n5294_;
  assign new_n20739_ = ~new_n5682_;
  assign new_n20740_ = ~new_n5285_;
  assign new_n20741_ = ~new_n5285_ | ~new_n5682_;
  assign new_n20742_ = ~new_n5688_;
  assign new_n20743_ = ~new_n5302_;
  assign new_n20744_ = ~new_n5691_;
  assign new_n20745_ = ~new_n5301_;
  assign new_n20746_ = ~new_n5694_;
  assign new_n20747_ = ~new_n5296_;
  assign new_n20748_ = ~new_n5703_;
  assign new_n20749_ = ~new_n5304_;
  assign new_n20750_ = ~new_n5304_ | ~new_n5703_;
  assign new_n20751_ = ~new_n5705_;
  assign new_n20752_ = ~new_n5303_;
  assign new_n20753_ = ~new_n5303_ | ~new_n5705_;
  assign new_n20754_ = ~new_n6177_;
  assign new_n20755_ = ~new_n6175_;
  assign new_n20756_ = ~new_n5283_;
  assign new_n20757_ = ~new_n6174_;
  assign new_n20758_ = ~new_n5288_;
  assign new_n20759_ = ~new_n6171_ | ~new_n5279_;
  assign new_n20760_ = ~new_n5276_;
  assign new_n20761_ = ~new_n6169_;
  assign new_n20762_ = ~new_n20978_ | ~new_n20848_;
  assign new_n20763_ = ~new_n5298_;
  assign new_n20764_ = ~new_n20750_ | ~new_n20987_;
  assign new_n20765_ = ~new_n20933_ | ~new_n20932_;
  assign new_n20766_ = ~new_n20741_ | ~new_n21009_;
  assign new_n20767_ = ~new_n21129_ | ~new_n21128_;
  assign new_n20768_ = ~new_n21176_ | ~new_n21175_;
  assign new_n20769_ = ~new_n21047_ | ~new_n21046_;
  assign new_n20770_ = ~new_n21052_ | ~new_n21051_;
  assign new_n20771_ = ~new_n21059_ | ~new_n21058_;
  assign new_n20772_ = ~new_n21066_ | ~new_n21065_;
  assign new_n20773_ = ~new_n21071_ | ~new_n21070_;
  assign new_n20774_ = ~new_n21080_ | ~new_n21079_;
  assign new_n20775_ = ~new_n21087_ | ~new_n21086_;
  assign new_n20776_ = ~new_n21094_ | ~new_n21093_;
  assign new_n20777_ = ~new_n21101_ | ~new_n21100_;
  assign new_n20778_ = ~new_n21106_ | ~new_n21105_;
  assign new_n20779_ = ~new_n21113_ | ~new_n21112_;
  assign new_n20780_ = ~new_n21120_ | ~new_n21119_;
  assign new_n20781_ = ~new_n21134_ | ~new_n21133_;
  assign new_n20782_ = ~new_n21139_ | ~new_n21138_;
  assign new_n20783_ = ~new_n21146_ | ~new_n21145_;
  assign new_n20784_ = ~new_n21153_ | ~new_n21152_;
  assign new_n20785_ = ~new_n21160_ | ~new_n21159_;
  assign new_n20786_ = ~new_n21167_ | ~new_n21166_;
  assign new_n20787_ = ~new_n21172_ | ~new_n21171_;
  assign new_n20788_ = new_n5655_ & new_n5290_;
  assign new_n20789_ = new_n20861_ & new_n20859_;
  assign new_n20790_ = new_n20866_ & new_n20864_;
  assign new_n20791_ = new_n20873_ & new_n20872_;
  assign new_n20792_ = new_n20695_ & new_n21054_ & new_n21053_;
  assign new_n20793_ = new_n20884_ & new_n20678_;
  assign new_n20794_ = new_n20892_ & new_n20890_;
  assign new_n20795_ = new_n20707_ & new_n21061_ & new_n21060_;
  assign new_n20796_ = new_n20898_ & new_n20676_;
  assign new_n20797_ = new_n20906_ & new_n20853_;
  assign new_n20798_ = new_n20876_ & new_n20679_;
  assign new_n20799_ = new_n20911_ & new_n20843_;
  assign new_n20800_ = new_n20922_ & new_n20680_;
  assign new_n20801_ = new_n20920_ & new_n20844_;
  assign new_n20802_ = new_n20940_ & new_n20939_;
  assign new_n20803_ = new_n20682_ & new_n20954_;
  assign new_n20804_ = new_n20957_ & new_n20952_;
  assign new_n20805_ = new_n20973_ & new_n20970_;
  assign new_n20806_ = new_n21040_ & new_n20974_;
  assign new_n20807_ = new_n20832_ & new_n20950_;
  assign new_n20808_ = new_n20753_ & new_n21127_ & new_n21126_;
  assign new_n20809_ = new_n20997_ & new_n20682_;
  assign new_n20810_ = new_n20732_ & new_n21141_ & new_n21140_;
  assign new_n20811_ = new_n21006_ & new_n20681_;
  assign new_n20812_ = new_n20844_ & new_n21162_ & new_n21161_;
  assign new_n20813_ = new_n21015_ & new_n20680_;
  assign new_n20814_ = new_n20843_ & new_n21174_ & new_n21173_;
  assign new_n20815_ = new_n21022_ & new_n20679_;
  assign new_n20816_ = ~new_n20791_ | ~new_n20874_;
  assign new_n20817_ = ~new_n20889_ | ~new_n20901_;
  assign new_n20818_ = ~new_n5277_;
  assign new_n20819_ = ~new_n6180_;
  assign new_n20820_ = new_n21075_ & new_n21074_;
  assign new_n20821_ = ~new_n21036_ | ~new_n20976_ | ~new_n20841_;
  assign new_n20822_ = new_n21082_ & new_n21081_;
  assign new_n20823_ = ~new_n20806_ | ~new_n21042_ | ~new_n21041_;
  assign new_n20824_ = new_n21089_ & new_n21088_;
  assign new_n20825_ = ~new_n20759_ | ~new_n21037_ | ~new_n20971_;
  assign new_n20826_ = new_n21096_ & new_n21095_;
  assign new_n20827_ = ~new_n20965_ | ~new_n20964_;
  assign new_n20828_ = new_n21108_ & new_n21107_;
  assign new_n20829_ = ~new_n20961_ | ~new_n20960_;
  assign new_n20830_ = new_n21115_ & new_n21114_;
  assign new_n20831_ = ~new_n20804_ | ~new_n20956_;
  assign new_n20832_ = new_n21122_ & new_n21121_;
  assign new_n20833_ = ~new_n20716_ | ~new_n20999_;
  assign new_n20834_ = ~new_n20802_ | ~new_n20941_;
  assign new_n20835_ = new_n21148_ & new_n21147_;
  assign new_n20836_ = ~new_n20929_ | ~new_n20928_;
  assign new_n20837_ = new_n21155_ & new_n21154_;
  assign new_n20838_ = ~new_n20925_ | ~new_n20924_;
  assign new_n20839_ = ~new_n20915_ | ~new_n20914_;
  assign new_n20840_ = ~new_n21039_ | ~new_n21038_;
  assign new_n20841_ = ~new_n5276_ | ~new_n20823_;
  assign new_n20842_ = ~new_n20707_;
  assign new_n20843_ = ~new_n5676_ | ~new_n5305_;
  assign new_n20844_ = ~new_n5294_ | ~new_n5685_;
  assign new_n20845_ = ~new_n5280_ | ~new_n6172_;
  assign new_n20846_ = ~new_n20741_;
  assign new_n20847_ = ~new_n20750_;
  assign new_n20848_ = ~new_n5287_ | ~new_n6173_;
  assign new_n20849_ = ~new_n20734_;
  assign new_n20850_ = new_n5289_ | new_n5664_;
  assign new_n20851_ = new_n5282_ | new_n5661_;
  assign new_n20852_ = new_n5658_ | new_n5286_;
  assign new_n20853_ = new_n5655_ | new_n5290_;
  assign new_n20854_ = ~new_n20704_;
  assign new_n20855_ = new_n5652_ | new_n5300_;
  assign new_n20856_ = ~new_n20715_;
  assign new_n20857_ = ~new_n20716_;
  assign new_n20858_ = ~new_n20715_ | ~new_n20716_;
  assign new_n20859_ = ~new_n20788_ | ~new_n20852_;
  assign new_n20860_ = ~new_n20677_ | ~new_n20858_;
  assign new_n20861_ = ~new_n5286_ | ~new_n5658_;
  assign new_n20862_ = ~new_n20789_ | ~new_n20860_;
  assign new_n20863_ = ~new_n20708_ | ~new_n20707_;
  assign new_n20864_ = ~new_n5289_ | ~new_n20863_;
  assign new_n20865_ = ~new_n20676_ | ~new_n20862_;
  assign new_n20866_ = ~new_n5664_ | ~new_n20842_;
  assign new_n20867_ = ~new_n20714_;
  assign new_n20868_ = new_n5292_ | new_n5670_;
  assign new_n20869_ = new_n5293_ | new_n5667_;
  assign new_n20870_ = ~new_n20695_;
  assign new_n20871_ = ~new_n20696_ | ~new_n20695_;
  assign new_n20872_ = ~new_n5292_ | ~new_n20871_;
  assign new_n20873_ = ~new_n5670_ | ~new_n20870_;
  assign new_n20874_ = ~new_n20678_ | ~new_n20714_;
  assign new_n20875_ = ~new_n20816_;
  assign new_n20876_ = new_n5673_ | new_n5306_;
  assign new_n20877_ = ~new_n20876_ | ~new_n20816_;
  assign new_n20878_ = ~new_n20713_;
  assign new_n20879_ = new_n5305_ | new_n5676_;
  assign new_n20880_ = new_n5667_ | new_n5293_;
  assign new_n20881_ = ~new_n20880_ | ~new_n20714_;
  assign new_n20882_ = ~new_n20792_ | ~new_n20881_;
  assign new_n20883_ = ~new_n20867_ | ~new_n20695_;
  assign new_n20884_ = ~new_n5670_ | ~new_n5292_;
  assign new_n20885_ = ~new_n20793_ | ~new_n20883_;
  assign new_n20886_ = new_n5293_ | new_n5667_;
  assign new_n20887_ = ~new_n20857_ | ~new_n20853_;
  assign new_n20888_ = ~new_n5290_ | ~new_n5655_;
  assign new_n20889_ = ~new_n20718_;
  assign new_n20890_ = ~new_n20856_ | ~new_n20677_;
  assign new_n20891_ = ~new_n20718_ | ~new_n20852_;
  assign new_n20892_ = ~new_n5286_ | ~new_n5658_;
  assign new_n20893_ = ~new_n20717_;
  assign new_n20894_ = new_n5661_ | new_n5282_;
  assign new_n20895_ = ~new_n20894_ | ~new_n20717_;
  assign new_n20896_ = ~new_n20795_ | ~new_n20895_;
  assign new_n20897_ = ~new_n20893_ | ~new_n20707_;
  assign new_n20898_ = ~new_n5664_ | ~new_n5289_;
  assign new_n20899_ = ~new_n20796_ | ~new_n20897_;
  assign new_n20900_ = new_n5282_ | new_n5661_;
  assign new_n20901_ = ~new_n20856_ | ~new_n20853_;
  assign new_n20902_ = ~new_n20817_;
  assign new_n20903_ = ~new_n5286_ | ~new_n5658_;
  assign new_n20904_ = ~new_n21072_ | ~new_n20715_ | ~new_n20716_ | ~new_n21073_;
  assign new_n20905_ = ~new_n20716_ | ~new_n20715_;
  assign new_n20906_ = ~new_n5290_ | ~new_n5655_;
  assign new_n20907_ = ~new_n20797_ | ~new_n20905_;
  assign new_n20908_ = new_n5305_ | new_n5676_;
  assign new_n20909_ = new_n5284_ | new_n5679_;
  assign new_n20910_ = ~new_n20849_ | ~new_n20679_;
  assign new_n20911_ = ~new_n5284_ | ~new_n5679_;
  assign new_n20912_ = ~new_n20799_ | ~new_n20910_;
  assign new_n20913_ = new_n5679_ | new_n5284_;
  assign new_n20914_ = ~new_n20798_ | ~new_n20816_;
  assign new_n20915_ = ~new_n20913_ | ~new_n20912_;
  assign new_n20916_ = ~new_n20839_;
  assign new_n20917_ = new_n5302_ | new_n5688_;
  assign new_n20918_ = new_n5294_ | new_n5685_;
  assign new_n20919_ = ~new_n20846_ | ~new_n20680_;
  assign new_n20920_ = ~new_n5302_ | ~new_n5688_;
  assign new_n20921_ = ~new_n20801_ | ~new_n20919_;
  assign new_n20922_ = new_n5682_ | new_n5285_;
  assign new_n20923_ = new_n5688_ | new_n5302_;
  assign new_n20924_ = ~new_n20800_ | ~new_n20839_;
  assign new_n20925_ = ~new_n20923_ | ~new_n20921_;
  assign new_n20926_ = ~new_n20838_;
  assign new_n20927_ = new_n5691_ | new_n5301_;
  assign new_n20928_ = ~new_n20927_ | ~new_n20838_;
  assign new_n20929_ = ~new_n5301_ | ~new_n5691_;
  assign new_n20930_ = ~new_n20836_;
  assign new_n20931_ = new_n5694_ | new_n5296_;
  assign new_n20932_ = ~new_n20931_ | ~new_n20836_;
  assign new_n20933_ = ~new_n5296_ | ~new_n5694_;
  assign new_n20934_ = ~new_n20765_;
  assign new_n20935_ = new_n5291_ | new_n5700_;
  assign new_n20936_ = new_n5295_ | new_n5697_;
  assign new_n20937_ = ~new_n20732_;
  assign new_n20938_ = ~new_n20733_ | ~new_n20732_;
  assign new_n20939_ = ~new_n5291_ | ~new_n20938_;
  assign new_n20940_ = ~new_n5700_ | ~new_n20937_;
  assign new_n20941_ = ~new_n20681_ | ~new_n20765_;
  assign new_n20942_ = ~new_n20834_;
  assign new_n20943_ = new_n5298_ | new_n6177_;
  assign new_n20944_ = new_n5303_ | new_n5705_;
  assign new_n20945_ = new_n5297_ | new_n6176_;
  assign new_n20946_ = ~new_n20753_;
  assign new_n20947_ = ~new_n6177_ | ~new_n20946_;
  assign new_n20948_ = ~new_n20947_ | ~new_n20763_;
  assign new_n20949_ = ~new_n20753_ | ~new_n20754_;
  assign new_n20950_ = ~new_n20949_ | ~new_n20948_;
  assign new_n20951_ = ~new_n20847_ | ~new_n20682_;
  assign new_n20952_ = ~new_n5297_ | ~new_n6176_;
  assign new_n20953_ = ~new_n20950_ | ~new_n20951_;
  assign new_n20954_ = new_n5703_ | new_n5304_;
  assign new_n20955_ = new_n6176_ | new_n5297_;
  assign new_n20956_ = ~new_n20803_ | ~new_n20945_ | ~new_n20834_;
  assign new_n20957_ = ~new_n20955_ | ~new_n20953_;
  assign new_n20958_ = ~new_n20831_;
  assign new_n20959_ = new_n6175_ | new_n5283_;
  assign new_n20960_ = ~new_n20959_ | ~new_n20831_;
  assign new_n20961_ = ~new_n5283_ | ~new_n6175_;
  assign new_n20962_ = ~new_n20829_;
  assign new_n20963_ = new_n6174_ | new_n5288_;
  assign new_n20964_ = ~new_n20963_ | ~new_n20829_;
  assign new_n20965_ = ~new_n5288_ | ~new_n6174_;
  assign new_n20966_ = ~new_n20827_;
  assign new_n20967_ = new_n5280_ | new_n6172_;
  assign new_n20968_ = ~new_n20848_ | ~new_n20845_;
  assign new_n20969_ = ~new_n20759_;
  assign new_n20970_ = new_n6173_ | new_n5287_;
  assign new_n20971_ = ~new_n20840_ | ~new_n20827_ | ~new_n20970_;
  assign new_n20972_ = ~new_n20825_;
  assign new_n20973_ = new_n6170_ | new_n5275_;
  assign new_n20974_ = ~new_n5275_ | ~new_n6170_;
  assign new_n20975_ = ~new_n20823_;
  assign new_n20976_ = ~new_n6169_ | ~new_n20823_;
  assign new_n20977_ = ~new_n20821_;
  assign new_n20978_ = ~new_n20970_ | ~new_n20827_;
  assign new_n20979_ = ~new_n20762_;
  assign new_n20980_ = new_n6172_ | new_n5280_;
  assign new_n20981_ = ~new_n20980_ | ~new_n20762_;
  assign new_n20982_ = ~new_n20826_ | ~new_n20981_ | ~new_n20845_;
  assign new_n20983_ = ~new_n20979_ | ~new_n20845_;
  assign new_n20984_ = ~new_n6171_ | ~new_n5279_;
  assign new_n20985_ = ~new_n20840_ | ~new_n20983_ | ~new_n20984_;
  assign new_n20986_ = new_n5280_ | new_n6172_;
  assign new_n20987_ = ~new_n20954_ | ~new_n20834_;
  assign new_n20988_ = ~new_n20764_;
  assign new_n20989_ = ~new_n20682_ | ~new_n20764_;
  assign new_n20990_ = ~new_n20807_ | ~new_n20989_;
  assign new_n20991_ = ~new_n20989_ | ~new_n20950_;
  assign new_n20992_ = ~new_n21125_ | ~new_n20991_;
  assign new_n20993_ = new_n5705_ | new_n5303_;
  assign new_n20994_ = ~new_n20993_ | ~new_n20764_;
  assign new_n20995_ = ~new_n20808_ | ~new_n20994_;
  assign new_n20996_ = ~new_n20988_ | ~new_n20753_;
  assign new_n20997_ = ~new_n5298_ | ~new_n6177_;
  assign new_n20998_ = ~new_n20809_ | ~new_n20996_;
  assign new_n20999_ = new_n5652_ | new_n5300_;
  assign new_n21000_ = ~new_n20833_;
  assign new_n21001_ = new_n5303_ | new_n5705_;
  assign new_n21002_ = new_n5697_ | new_n5295_;
  assign new_n21003_ = ~new_n21002_ | ~new_n20765_;
  assign new_n21004_ = ~new_n20810_ | ~new_n21003_;
  assign new_n21005_ = ~new_n20934_ | ~new_n20732_;
  assign new_n21006_ = ~new_n5700_ | ~new_n5291_;
  assign new_n21007_ = ~new_n20811_ | ~new_n21005_;
  assign new_n21008_ = new_n5295_ | new_n5697_;
  assign new_n21009_ = ~new_n20922_ | ~new_n20839_;
  assign new_n21010_ = ~new_n20766_;
  assign new_n21011_ = new_n5685_ | new_n5294_;
  assign new_n21012_ = ~new_n21011_ | ~new_n20766_;
  assign new_n21013_ = ~new_n20812_ | ~new_n21012_;
  assign new_n21014_ = ~new_n21010_ | ~new_n20844_;
  assign new_n21015_ = ~new_n5302_ | ~new_n5688_;
  assign new_n21016_ = ~new_n20813_ | ~new_n21014_;
  assign new_n21017_ = new_n5294_ | new_n5685_;
  assign new_n21018_ = new_n5676_ | new_n5305_;
  assign new_n21019_ = ~new_n21018_ | ~new_n20713_;
  assign new_n21020_ = ~new_n20814_ | ~new_n21019_;
  assign new_n21021_ = ~new_n20878_ | ~new_n20843_;
  assign new_n21022_ = ~new_n5284_ | ~new_n5679_;
  assign new_n21023_ = ~new_n20815_ | ~new_n21021_;
  assign new_n21024_ = ~new_n20879_ | ~new_n20843_;
  assign new_n21025_ = ~new_n20876_ | ~new_n20734_;
  assign new_n21026_ = ~new_n20886_ | ~new_n20695_;
  assign new_n21027_ = ~new_n20900_ | ~new_n20707_;
  assign new_n21028_ = ~new_n20903_ | ~new_n20852_;
  assign new_n21029_ = ~new_n20986_ | ~new_n20845_;
  assign new_n21030_ = ~new_n20970_ | ~new_n20848_;
  assign new_n21031_ = ~new_n21001_ | ~new_n20753_;
  assign new_n21032_ = ~new_n20954_ | ~new_n20750_;
  assign new_n21033_ = ~new_n21008_ | ~new_n20732_;
  assign new_n21034_ = ~new_n21017_ | ~new_n20844_;
  assign new_n21035_ = ~new_n20922_ | ~new_n20741_;
  assign new_n21036_ = ~new_n6169_ | ~new_n5276_;
  assign new_n21037_ = ~new_n20968_ | ~new_n20840_;
  assign new_n21038_ = ~new_n5279_ | ~new_n20967_;
  assign new_n21039_ = ~new_n6171_ | ~new_n20967_;
  assign new_n21040_ = ~new_n20973_ | ~new_n20968_ | ~new_n20840_;
  assign new_n21041_ = ~new_n20805_ | ~new_n20827_ | ~new_n20840_;
  assign new_n21042_ = ~new_n20969_ | ~new_n20973_;
  assign new_n21043_ = ~new_n5305_ | ~new_n20712_;
  assign new_n21044_ = ~new_n5676_ | ~new_n20711_;
  assign new_n21045_ = ~new_n21044_ | ~new_n21043_;
  assign new_n21046_ = ~new_n21024_ | ~new_n20713_;
  assign new_n21047_ = ~new_n21045_ | ~new_n20878_;
  assign new_n21048_ = ~new_n5306_ | ~new_n20709_;
  assign new_n21049_ = ~new_n5673_ | ~new_n20710_;
  assign new_n21050_ = ~new_n21049_ | ~new_n21048_;
  assign new_n21051_ = ~new_n21025_ | ~new_n20816_;
  assign new_n21052_ = ~new_n20875_ | ~new_n21050_;
  assign new_n21053_ = ~new_n5292_ | ~new_n20696_;
  assign new_n21054_ = ~new_n5670_ | ~new_n20694_;
  assign new_n21055_ = ~new_n5293_ | ~new_n20692_;
  assign new_n21056_ = ~new_n5667_ | ~new_n20693_;
  assign new_n21057_ = ~new_n21056_ | ~new_n21055_;
  assign new_n21058_ = ~new_n21026_ | ~new_n20714_;
  assign new_n21059_ = ~new_n21057_ | ~new_n20867_;
  assign new_n21060_ = ~new_n5289_ | ~new_n20708_;
  assign new_n21061_ = ~new_n5664_ | ~new_n20699_;
  assign new_n21062_ = ~new_n5282_ | ~new_n20697_;
  assign new_n21063_ = ~new_n5661_ | ~new_n20698_;
  assign new_n21064_ = ~new_n21063_ | ~new_n21062_;
  assign new_n21065_ = ~new_n21027_ | ~new_n20717_;
  assign new_n21066_ = ~new_n21064_ | ~new_n20893_;
  assign new_n21067_ = ~new_n5286_ | ~new_n20705_;
  assign new_n21068_ = ~new_n5658_ | ~new_n20706_;
  assign new_n21069_ = ~new_n21068_ | ~new_n21067_;
  assign new_n21070_ = ~new_n21028_ | ~new_n20817_;
  assign new_n21071_ = ~new_n20902_ | ~new_n21069_;
  assign new_n21072_ = ~new_n5290_ | ~new_n20700_;
  assign new_n21073_ = ~new_n5655_ | ~new_n20701_;
  assign new_n21074_ = ~new_n5277_ | ~new_n20819_;
  assign new_n21075_ = ~new_n6180_ | ~new_n20818_;
  assign new_n21076_ = ~new_n5277_ | ~new_n20819_;
  assign new_n21077_ = ~new_n6180_ | ~new_n20818_;
  assign new_n21078_ = ~new_n21077_ | ~new_n21076_;
  assign new_n21079_ = ~new_n20820_ | ~new_n20821_;
  assign new_n21080_ = ~new_n20977_ | ~new_n21078_;
  assign new_n21081_ = ~new_n5276_ | ~new_n20761_;
  assign new_n21082_ = ~new_n6169_ | ~new_n20760_;
  assign new_n21083_ = ~new_n5276_ | ~new_n20761_;
  assign new_n21084_ = ~new_n6169_ | ~new_n20760_;
  assign new_n21085_ = ~new_n21084_ | ~new_n21083_;
  assign new_n21086_ = ~new_n20822_ | ~new_n20823_;
  assign new_n21087_ = ~new_n20975_ | ~new_n21085_;
  assign new_n21088_ = ~new_n5275_ | ~new_n20719_;
  assign new_n21089_ = ~new_n6170_ | ~new_n20720_;
  assign new_n21090_ = ~new_n5275_ | ~new_n20719_;
  assign new_n21091_ = ~new_n6170_ | ~new_n20720_;
  assign new_n21092_ = ~new_n21091_ | ~new_n21090_;
  assign new_n21093_ = ~new_n20824_ | ~new_n20825_;
  assign new_n21094_ = ~new_n20972_ | ~new_n21092_;
  assign new_n21095_ = ~new_n5279_ | ~new_n20722_;
  assign new_n21096_ = ~new_n6171_ | ~new_n20721_;
  assign new_n21097_ = ~new_n5280_ | ~new_n20723_;
  assign new_n21098_ = ~new_n6172_ | ~new_n20724_;
  assign new_n21099_ = ~new_n21098_ | ~new_n21097_;
  assign new_n21100_ = ~new_n21029_ | ~new_n20762_;
  assign new_n21101_ = ~new_n21099_ | ~new_n20979_;
  assign new_n21102_ = ~new_n5287_ | ~new_n20725_;
  assign new_n21103_ = ~new_n6173_ | ~new_n20726_;
  assign new_n21104_ = ~new_n21103_ | ~new_n21102_;
  assign new_n21105_ = ~new_n21030_ | ~new_n20827_;
  assign new_n21106_ = ~new_n20966_ | ~new_n21104_;
  assign new_n21107_ = ~new_n5288_ | ~new_n20757_;
  assign new_n21108_ = ~new_n6174_ | ~new_n20758_;
  assign new_n21109_ = ~new_n5288_ | ~new_n20757_;
  assign new_n21110_ = ~new_n6174_ | ~new_n20758_;
  assign new_n21111_ = ~new_n21110_ | ~new_n21109_;
  assign new_n21112_ = ~new_n20828_ | ~new_n20829_;
  assign new_n21113_ = ~new_n20962_ | ~new_n21111_;
  assign new_n21114_ = ~new_n5283_ | ~new_n20755_;
  assign new_n21115_ = ~new_n6175_ | ~new_n20756_;
  assign new_n21116_ = ~new_n5283_ | ~new_n20755_;
  assign new_n21117_ = ~new_n6175_ | ~new_n20756_;
  assign new_n21118_ = ~new_n21117_ | ~new_n21116_;
  assign new_n21119_ = ~new_n20830_ | ~new_n20831_;
  assign new_n21120_ = ~new_n20958_ | ~new_n21118_;
  assign new_n21121_ = ~new_n5297_ | ~new_n20727_;
  assign new_n21122_ = ~new_n6176_ | ~new_n20728_;
  assign new_n21123_ = ~new_n5297_ | ~new_n20727_;
  assign new_n21124_ = ~new_n6176_ | ~new_n20728_;
  assign new_n21125_ = ~new_n21124_ | ~new_n21123_;
  assign new_n21126_ = ~new_n5298_ | ~new_n20754_;
  assign new_n21127_ = ~new_n6177_ | ~new_n20763_;
  assign new_n21128_ = ~new_n20854_ | ~new_n20833_;
  assign new_n21129_ = ~new_n21000_ | ~new_n20704_;
  assign new_n21130_ = ~new_n5303_ | ~new_n20751_;
  assign new_n21131_ = ~new_n5705_ | ~new_n20752_;
  assign new_n21132_ = ~new_n21131_ | ~new_n21130_;
  assign new_n21133_ = ~new_n21031_ | ~new_n20764_;
  assign new_n21134_ = ~new_n21132_ | ~new_n20988_;
  assign new_n21135_ = ~new_n5304_ | ~new_n20748_;
  assign new_n21136_ = ~new_n5703_ | ~new_n20749_;
  assign new_n21137_ = ~new_n21136_ | ~new_n21135_;
  assign new_n21138_ = ~new_n21032_ | ~new_n20834_;
  assign new_n21139_ = ~new_n20942_ | ~new_n21137_;
  assign new_n21140_ = ~new_n5291_ | ~new_n20733_;
  assign new_n21141_ = ~new_n5700_ | ~new_n20731_;
  assign new_n21142_ = ~new_n5295_ | ~new_n20729_;
  assign new_n21143_ = ~new_n5697_ | ~new_n20730_;
  assign new_n21144_ = ~new_n21143_ | ~new_n21142_;
  assign new_n21145_ = ~new_n21033_ | ~new_n20765_;
  assign new_n21146_ = ~new_n21144_ | ~new_n20934_;
  assign new_n21147_ = ~new_n5296_ | ~new_n20746_;
  assign new_n21148_ = ~new_n5694_ | ~new_n20747_;
  assign new_n21149_ = ~new_n5296_ | ~new_n20746_;
  assign new_n21150_ = ~new_n5694_ | ~new_n20747_;
  assign new_n21151_ = ~new_n21150_ | ~new_n21149_;
  assign new_n21152_ = ~new_n20835_ | ~new_n20836_;
  assign new_n21153_ = ~new_n20930_ | ~new_n21151_;
  assign new_n21154_ = ~new_n5301_ | ~new_n20744_;
  assign new_n21155_ = ~new_n5691_ | ~new_n20745_;
  assign new_n21156_ = ~new_n5301_ | ~new_n20744_;
  assign new_n21157_ = ~new_n5691_ | ~new_n20745_;
  assign new_n21158_ = ~new_n21157_ | ~new_n21156_;
  assign new_n21159_ = ~new_n20837_ | ~new_n20838_;
  assign new_n21160_ = ~new_n20926_ | ~new_n21158_;
  assign new_n21161_ = ~new_n5302_ | ~new_n20742_;
  assign new_n21162_ = ~new_n5688_ | ~new_n20743_;
  assign new_n21163_ = ~new_n5294_ | ~new_n20737_;
  assign new_n21164_ = ~new_n5685_ | ~new_n20738_;
  assign new_n21165_ = ~new_n21164_ | ~new_n21163_;
  assign new_n21166_ = ~new_n21034_ | ~new_n20766_;
  assign new_n21167_ = ~new_n21165_ | ~new_n21010_;
  assign new_n21168_ = ~new_n5285_ | ~new_n20739_;
  assign new_n21169_ = ~new_n5682_ | ~new_n20740_;
  assign new_n21170_ = ~new_n21169_ | ~new_n21168_;
  assign new_n21171_ = ~new_n21035_ | ~new_n20839_;
  assign new_n21172_ = ~new_n20916_ | ~new_n21170_;
  assign new_n21173_ = ~new_n5284_ | ~new_n20735_;
  assign new_n21174_ = ~new_n5679_ | ~new_n20736_;
  assign new_n21175_ = ~new_n5299_ | ~new_n20702_;
  assign new_n21176_ = ~new_n5647_ | ~new_n20703_;
  assign new_n21177_ = new_n21352_ & new_n21351_;
  assign new_n21178_ = new_n21370_ & new_n21369_;
  assign new_n21179_ = new_n21410_ & new_n21409_;
  assign new_n21180_ = new_n21419_ & new_n21418_;
  assign new_n21181_ = new_n21437_ & new_n21436_;
  assign new_n21182_ = new_n21445_ & new_n21444_;
  assign new_n21183_ = new_n21524_ & new_n21521_;
  assign new_n21184_ = new_n21517_ & new_n21514_;
  assign new_n21185_ = new_n21508_ & new_n21505_;
  assign new_n21186_ = new_n21499_ & new_n21496_;
  assign new_n21187_ = new_n21493_ & new_n21491_;
  assign new_n21188_ = new_n21486_ & new_n21483_;
  assign new_n21189_ = new_n21408_ & new_n21405_;
  assign new_n21190_ = new_n21400_ & new_n21397_;
  assign new_n21191_ = new_n21386_ & new_n21383_;
  assign new_n21192_ = ~new_n5667_;
  assign new_n21193_ = ~new_n5293_;
  assign new_n21194_ = ~new_n5292_;
  assign new_n21195_ = ~new_n5293_ | ~new_n5667_;
  assign new_n21196_ = ~new_n5670_;
  assign new_n21197_ = ~new_n5661_;
  assign new_n21198_ = ~new_n5282_;
  assign new_n21199_ = ~new_n5289_;
  assign new_n21200_ = ~new_n5655_;
  assign new_n21201_ = ~new_n5290_;
  assign new_n21202_ = ~new_n5647_;
  assign new_n21203_ = ~new_n5299_;
  assign new_n21204_ = ~new_n5299_ | ~new_n5647_;
  assign new_n21205_ = ~new_n5658_;
  assign new_n21206_ = ~new_n5286_;
  assign new_n21207_ = ~new_n5282_ | ~new_n5661_;
  assign new_n21208_ = ~new_n5664_;
  assign new_n21209_ = ~new_n5673_;
  assign new_n21210_ = ~new_n5306_;
  assign new_n21211_ = ~new_n5305_;
  assign new_n21212_ = ~new_n5676_;
  assign new_n21213_ = ~new_n21234_ | ~new_n21378_;
  assign new_n21214_ = ~new_n21290_ | ~new_n21366_;
  assign new_n21215_ = ~new_n21355_ | ~new_n21356_;
  assign new_n21216_ = ~new_n5652_ | ~new_n5300_;
  assign new_n21217_ = ~new_n21295_ | ~new_n21392_;
  assign new_n21218_ = ~new_n21389_ | ~new_n21388_;
  assign new_n21219_ = ~new_n6170_;
  assign new_n21220_ = ~new_n5275_;
  assign new_n21221_ = ~new_n5279_;
  assign new_n21222_ = ~new_n6171_;
  assign new_n21223_ = ~new_n6172_;
  assign new_n21224_ = ~new_n5280_;
  assign new_n21225_ = ~new_n6173_;
  assign new_n21226_ = ~new_n5287_;
  assign new_n21227_ = ~new_n6176_;
  assign new_n21228_ = ~new_n5297_;
  assign new_n21229_ = ~new_n5697_;
  assign new_n21230_ = ~new_n5295_;
  assign new_n21231_ = ~new_n5291_;
  assign new_n21232_ = ~new_n5295_ | ~new_n5697_;
  assign new_n21233_ = ~new_n5700_;
  assign new_n21234_ = ~new_n5306_ | ~new_n5673_;
  assign new_n21235_ = ~new_n5679_;
  assign new_n21236_ = ~new_n5284_;
  assign new_n21237_ = ~new_n5685_;
  assign new_n21238_ = ~new_n5294_;
  assign new_n21239_ = ~new_n5682_;
  assign new_n21240_ = ~new_n5285_;
  assign new_n21241_ = ~new_n5285_ | ~new_n5682_;
  assign new_n21242_ = ~new_n5688_;
  assign new_n21243_ = ~new_n5302_;
  assign new_n21244_ = ~new_n5691_;
  assign new_n21245_ = ~new_n5301_;
  assign new_n21246_ = ~new_n5694_;
  assign new_n21247_ = ~new_n5296_;
  assign new_n21248_ = ~new_n5703_;
  assign new_n21249_ = ~new_n5304_;
  assign new_n21250_ = ~new_n5304_ | ~new_n5703_;
  assign new_n21251_ = ~new_n5705_;
  assign new_n21252_ = ~new_n5303_;
  assign new_n21253_ = ~new_n5303_ | ~new_n5705_;
  assign new_n21254_ = ~new_n6177_;
  assign new_n21255_ = ~new_n6175_;
  assign new_n21256_ = ~new_n5283_;
  assign new_n21257_ = ~new_n6174_;
  assign new_n21258_ = ~new_n5288_;
  assign new_n21259_ = ~new_n6171_ | ~new_n5279_;
  assign new_n21260_ = ~new_n5276_;
  assign new_n21261_ = ~new_n6169_;
  assign new_n21262_ = ~new_n21479_ | ~new_n21349_;
  assign new_n21263_ = ~new_n5298_;
  assign new_n21264_ = ~new_n21250_ | ~new_n21488_;
  assign new_n21265_ = ~new_n21434_ | ~new_n21433_;
  assign new_n21266_ = ~new_n21241_ | ~new_n21510_;
  assign new_n21267_ = ~new_n21630_ | ~new_n21629_;
  assign new_n21268_ = ~new_n21677_ | ~new_n21676_;
  assign new_n21269_ = ~new_n21548_ | ~new_n21547_;
  assign new_n21270_ = ~new_n21553_ | ~new_n21552_;
  assign new_n21271_ = ~new_n21560_ | ~new_n21559_;
  assign new_n21272_ = ~new_n21567_ | ~new_n21566_;
  assign new_n21273_ = ~new_n21572_ | ~new_n21571_;
  assign new_n21274_ = ~new_n21581_ | ~new_n21580_;
  assign new_n21275_ = ~new_n21588_ | ~new_n21587_;
  assign new_n21276_ = ~new_n21595_ | ~new_n21594_;
  assign new_n21277_ = ~new_n21602_ | ~new_n21601_;
  assign new_n21278_ = ~new_n21607_ | ~new_n21606_;
  assign new_n21279_ = ~new_n21614_ | ~new_n21613_;
  assign new_n21280_ = ~new_n21621_ | ~new_n21620_;
  assign new_n21281_ = ~new_n21635_ | ~new_n21634_;
  assign new_n21282_ = ~new_n21640_ | ~new_n21639_;
  assign new_n21283_ = ~new_n21647_ | ~new_n21646_;
  assign new_n21284_ = ~new_n21654_ | ~new_n21653_;
  assign new_n21285_ = ~new_n21661_ | ~new_n21660_;
  assign new_n21286_ = ~new_n21668_ | ~new_n21667_;
  assign new_n21287_ = ~new_n21673_ | ~new_n21672_;
  assign new_n21288_ = new_n21362_ & new_n21360_;
  assign new_n21289_ = new_n21177_ & new_n21353_;
  assign new_n21290_ = new_n21367_ & new_n21365_;
  assign new_n21291_ = new_n21374_ & new_n21373_;
  assign new_n21292_ = new_n21195_ & new_n21555_ & new_n21554_;
  assign new_n21293_ = new_n21385_ & new_n21178_;
  assign new_n21294_ = new_n21354_ & new_n21353_;
  assign new_n21295_ = new_n21393_ & new_n21391_;
  assign new_n21296_ = new_n21207_ & new_n21562_ & new_n21561_;
  assign new_n21297_ = new_n21399_ & new_n21177_;
  assign new_n21298_ = new_n21407_ & new_n21354_;
  assign new_n21299_ = new_n21377_ & new_n21179_;
  assign new_n21300_ = new_n21412_ & new_n21344_;
  assign new_n21301_ = new_n21423_ & new_n21180_;
  assign new_n21302_ = new_n21421_ & new_n21345_;
  assign new_n21303_ = new_n21441_ & new_n21440_;
  assign new_n21304_ = new_n21182_ & new_n21455_;
  assign new_n21305_ = new_n21458_ & new_n21453_;
  assign new_n21306_ = new_n21474_ & new_n21471_;
  assign new_n21307_ = new_n21541_ & new_n21475_;
  assign new_n21308_ = new_n21333_ & new_n21451_;
  assign new_n21309_ = new_n21253_ & new_n21628_ & new_n21627_;
  assign new_n21310_ = new_n21498_ & new_n21182_;
  assign new_n21311_ = new_n21232_ & new_n21642_ & new_n21641_;
  assign new_n21312_ = new_n21507_ & new_n21181_;
  assign new_n21313_ = new_n21345_ & new_n21663_ & new_n21662_;
  assign new_n21314_ = new_n21516_ & new_n21180_;
  assign new_n21315_ = new_n21344_ & new_n21675_ & new_n21674_;
  assign new_n21316_ = new_n21523_ & new_n21179_;
  assign new_n21317_ = ~new_n21291_ | ~new_n21375_;
  assign new_n21318_ = ~new_n21390_ | ~new_n21402_;
  assign new_n21319_ = ~new_n5277_;
  assign new_n21320_ = ~new_n6180_;
  assign new_n21321_ = new_n21576_ & new_n21575_;
  assign new_n21322_ = ~new_n21537_ | ~new_n21477_ | ~new_n21342_;
  assign new_n21323_ = new_n21583_ & new_n21582_;
  assign new_n21324_ = ~new_n21307_ | ~new_n21543_ | ~new_n21542_;
  assign new_n21325_ = new_n21590_ & new_n21589_;
  assign new_n21326_ = ~new_n21259_ | ~new_n21538_ | ~new_n21472_;
  assign new_n21327_ = new_n21597_ & new_n21596_;
  assign new_n21328_ = ~new_n21466_ | ~new_n21465_;
  assign new_n21329_ = new_n21609_ & new_n21608_;
  assign new_n21330_ = ~new_n21462_ | ~new_n21461_;
  assign new_n21331_ = new_n21616_ & new_n21615_;
  assign new_n21332_ = ~new_n21305_ | ~new_n21457_;
  assign new_n21333_ = new_n21623_ & new_n21622_;
  assign new_n21334_ = ~new_n21216_ | ~new_n21500_;
  assign new_n21335_ = ~new_n21303_ | ~new_n21442_;
  assign new_n21336_ = new_n21649_ & new_n21648_;
  assign new_n21337_ = ~new_n21430_ | ~new_n21429_;
  assign new_n21338_ = new_n21656_ & new_n21655_;
  assign new_n21339_ = ~new_n21426_ | ~new_n21425_;
  assign new_n21340_ = ~new_n21416_ | ~new_n21415_;
  assign new_n21341_ = ~new_n21540_ | ~new_n21539_;
  assign new_n21342_ = ~new_n5276_ | ~new_n21324_;
  assign new_n21343_ = ~new_n21207_;
  assign new_n21344_ = ~new_n5676_ | ~new_n5305_;
  assign new_n21345_ = ~new_n5294_ | ~new_n5685_;
  assign new_n21346_ = ~new_n5280_ | ~new_n6172_;
  assign new_n21347_ = ~new_n21241_;
  assign new_n21348_ = ~new_n21250_;
  assign new_n21349_ = ~new_n5287_ | ~new_n6173_;
  assign new_n21350_ = ~new_n21234_;
  assign new_n21351_ = new_n5289_ | new_n5664_;
  assign new_n21352_ = new_n5282_ | new_n5661_;
  assign new_n21353_ = new_n5658_ | new_n5286_;
  assign new_n21354_ = new_n5655_ | new_n5290_;
  assign new_n21355_ = ~new_n21204_;
  assign new_n21356_ = new_n5652_ | new_n5300_;
  assign new_n21357_ = ~new_n21215_;
  assign new_n21358_ = ~new_n21216_;
  assign new_n21359_ = ~new_n21215_ | ~new_n21216_;
  assign new_n21360_ = ~new_n5290_ | ~new_n5655_;
  assign new_n21361_ = ~new_n21359_ | ~new_n21354_;
  assign new_n21362_ = ~new_n5286_ | ~new_n5658_;
  assign new_n21363_ = ~new_n21288_ | ~new_n21361_;
  assign new_n21364_ = ~new_n21208_ | ~new_n21207_;
  assign new_n21365_ = ~new_n5289_ | ~new_n21364_;
  assign new_n21366_ = ~new_n21289_ | ~new_n21363_;
  assign new_n21367_ = ~new_n5664_ | ~new_n21343_;
  assign new_n21368_ = ~new_n21214_;
  assign new_n21369_ = new_n5292_ | new_n5670_;
  assign new_n21370_ = new_n5293_ | new_n5667_;
  assign new_n21371_ = ~new_n21195_;
  assign new_n21372_ = ~new_n21196_ | ~new_n21195_;
  assign new_n21373_ = ~new_n5292_ | ~new_n21372_;
  assign new_n21374_ = ~new_n5670_ | ~new_n21371_;
  assign new_n21375_ = ~new_n21178_ | ~new_n21214_;
  assign new_n21376_ = ~new_n21317_;
  assign new_n21377_ = new_n5673_ | new_n5306_;
  assign new_n21378_ = ~new_n21377_ | ~new_n21317_;
  assign new_n21379_ = ~new_n21213_;
  assign new_n21380_ = new_n5305_ | new_n5676_;
  assign new_n21381_ = new_n5667_ | new_n5293_;
  assign new_n21382_ = ~new_n21381_ | ~new_n21214_;
  assign new_n21383_ = ~new_n21292_ | ~new_n21382_;
  assign new_n21384_ = ~new_n21368_ | ~new_n21195_;
  assign new_n21385_ = ~new_n5670_ | ~new_n5292_;
  assign new_n21386_ = ~new_n21293_ | ~new_n21384_;
  assign new_n21387_ = new_n5293_ | new_n5667_;
  assign new_n21388_ = ~new_n21358_ | ~new_n21354_;
  assign new_n21389_ = ~new_n5290_ | ~new_n5655_;
  assign new_n21390_ = ~new_n21218_;
  assign new_n21391_ = ~new_n21294_ | ~new_n21357_;
  assign new_n21392_ = ~new_n21218_ | ~new_n21353_;
  assign new_n21393_ = ~new_n5286_ | ~new_n5658_;
  assign new_n21394_ = ~new_n21217_;
  assign new_n21395_ = new_n5661_ | new_n5282_;
  assign new_n21396_ = ~new_n21395_ | ~new_n21217_;
  assign new_n21397_ = ~new_n21296_ | ~new_n21396_;
  assign new_n21398_ = ~new_n21394_ | ~new_n21207_;
  assign new_n21399_ = ~new_n5664_ | ~new_n5289_;
  assign new_n21400_ = ~new_n21297_ | ~new_n21398_;
  assign new_n21401_ = new_n5282_ | new_n5661_;
  assign new_n21402_ = ~new_n21357_ | ~new_n21354_;
  assign new_n21403_ = ~new_n21318_;
  assign new_n21404_ = ~new_n5286_ | ~new_n5658_;
  assign new_n21405_ = ~new_n21573_ | ~new_n21215_ | ~new_n21216_ | ~new_n21574_;
  assign new_n21406_ = ~new_n21216_ | ~new_n21215_;
  assign new_n21407_ = ~new_n5290_ | ~new_n5655_;
  assign new_n21408_ = ~new_n21298_ | ~new_n21406_;
  assign new_n21409_ = new_n5305_ | new_n5676_;
  assign new_n21410_ = new_n5284_ | new_n5679_;
  assign new_n21411_ = ~new_n21350_ | ~new_n21179_;
  assign new_n21412_ = ~new_n5284_ | ~new_n5679_;
  assign new_n21413_ = ~new_n21300_ | ~new_n21411_;
  assign new_n21414_ = new_n5679_ | new_n5284_;
  assign new_n21415_ = ~new_n21299_ | ~new_n21317_;
  assign new_n21416_ = ~new_n21414_ | ~new_n21413_;
  assign new_n21417_ = ~new_n21340_;
  assign new_n21418_ = new_n5302_ | new_n5688_;
  assign new_n21419_ = new_n5294_ | new_n5685_;
  assign new_n21420_ = ~new_n21347_ | ~new_n21180_;
  assign new_n21421_ = ~new_n5302_ | ~new_n5688_;
  assign new_n21422_ = ~new_n21302_ | ~new_n21420_;
  assign new_n21423_ = new_n5682_ | new_n5285_;
  assign new_n21424_ = new_n5688_ | new_n5302_;
  assign new_n21425_ = ~new_n21301_ | ~new_n21340_;
  assign new_n21426_ = ~new_n21424_ | ~new_n21422_;
  assign new_n21427_ = ~new_n21339_;
  assign new_n21428_ = new_n5691_ | new_n5301_;
  assign new_n21429_ = ~new_n21428_ | ~new_n21339_;
  assign new_n21430_ = ~new_n5301_ | ~new_n5691_;
  assign new_n21431_ = ~new_n21337_;
  assign new_n21432_ = new_n5694_ | new_n5296_;
  assign new_n21433_ = ~new_n21432_ | ~new_n21337_;
  assign new_n21434_ = ~new_n5296_ | ~new_n5694_;
  assign new_n21435_ = ~new_n21265_;
  assign new_n21436_ = new_n5291_ | new_n5700_;
  assign new_n21437_ = new_n5295_ | new_n5697_;
  assign new_n21438_ = ~new_n21232_;
  assign new_n21439_ = ~new_n21233_ | ~new_n21232_;
  assign new_n21440_ = ~new_n5291_ | ~new_n21439_;
  assign new_n21441_ = ~new_n5700_ | ~new_n21438_;
  assign new_n21442_ = ~new_n21181_ | ~new_n21265_;
  assign new_n21443_ = ~new_n21335_;
  assign new_n21444_ = new_n5298_ | new_n6177_;
  assign new_n21445_ = new_n5303_ | new_n5705_;
  assign new_n21446_ = new_n5297_ | new_n6176_;
  assign new_n21447_ = ~new_n21253_;
  assign new_n21448_ = ~new_n6177_ | ~new_n21447_;
  assign new_n21449_ = ~new_n21448_ | ~new_n21263_;
  assign new_n21450_ = ~new_n21253_ | ~new_n21254_;
  assign new_n21451_ = ~new_n21450_ | ~new_n21449_;
  assign new_n21452_ = ~new_n21348_ | ~new_n21182_;
  assign new_n21453_ = ~new_n5297_ | ~new_n6176_;
  assign new_n21454_ = ~new_n21451_ | ~new_n21452_;
  assign new_n21455_ = new_n5703_ | new_n5304_;
  assign new_n21456_ = new_n6176_ | new_n5297_;
  assign new_n21457_ = ~new_n21304_ | ~new_n21446_ | ~new_n21335_;
  assign new_n21458_ = ~new_n21456_ | ~new_n21454_;
  assign new_n21459_ = ~new_n21332_;
  assign new_n21460_ = new_n6175_ | new_n5283_;
  assign new_n21461_ = ~new_n21460_ | ~new_n21332_;
  assign new_n21462_ = ~new_n5283_ | ~new_n6175_;
  assign new_n21463_ = ~new_n21330_;
  assign new_n21464_ = new_n6174_ | new_n5288_;
  assign new_n21465_ = ~new_n21464_ | ~new_n21330_;
  assign new_n21466_ = ~new_n5288_ | ~new_n6174_;
  assign new_n21467_ = ~new_n21328_;
  assign new_n21468_ = new_n5280_ | new_n6172_;
  assign new_n21469_ = ~new_n21349_ | ~new_n21346_;
  assign new_n21470_ = ~new_n21259_;
  assign new_n21471_ = new_n6173_ | new_n5287_;
  assign new_n21472_ = ~new_n21341_ | ~new_n21328_ | ~new_n21471_;
  assign new_n21473_ = ~new_n21326_;
  assign new_n21474_ = new_n6170_ | new_n5275_;
  assign new_n21475_ = ~new_n5275_ | ~new_n6170_;
  assign new_n21476_ = ~new_n21324_;
  assign new_n21477_ = ~new_n6169_ | ~new_n21324_;
  assign new_n21478_ = ~new_n21322_;
  assign new_n21479_ = ~new_n21471_ | ~new_n21328_;
  assign new_n21480_ = ~new_n21262_;
  assign new_n21481_ = new_n6172_ | new_n5280_;
  assign new_n21482_ = ~new_n21481_ | ~new_n21262_;
  assign new_n21483_ = ~new_n21327_ | ~new_n21482_ | ~new_n21346_;
  assign new_n21484_ = ~new_n21480_ | ~new_n21346_;
  assign new_n21485_ = ~new_n6171_ | ~new_n5279_;
  assign new_n21486_ = ~new_n21341_ | ~new_n21484_ | ~new_n21485_;
  assign new_n21487_ = new_n5280_ | new_n6172_;
  assign new_n21488_ = ~new_n21455_ | ~new_n21335_;
  assign new_n21489_ = ~new_n21264_;
  assign new_n21490_ = ~new_n21182_ | ~new_n21264_;
  assign new_n21491_ = ~new_n21308_ | ~new_n21490_;
  assign new_n21492_ = ~new_n21490_ | ~new_n21451_;
  assign new_n21493_ = ~new_n21626_ | ~new_n21492_;
  assign new_n21494_ = new_n5705_ | new_n5303_;
  assign new_n21495_ = ~new_n21494_ | ~new_n21264_;
  assign new_n21496_ = ~new_n21309_ | ~new_n21495_;
  assign new_n21497_ = ~new_n21489_ | ~new_n21253_;
  assign new_n21498_ = ~new_n5298_ | ~new_n6177_;
  assign new_n21499_ = ~new_n21310_ | ~new_n21497_;
  assign new_n21500_ = new_n5652_ | new_n5300_;
  assign new_n21501_ = ~new_n21334_;
  assign new_n21502_ = new_n5303_ | new_n5705_;
  assign new_n21503_ = new_n5697_ | new_n5295_;
  assign new_n21504_ = ~new_n21503_ | ~new_n21265_;
  assign new_n21505_ = ~new_n21311_ | ~new_n21504_;
  assign new_n21506_ = ~new_n21435_ | ~new_n21232_;
  assign new_n21507_ = ~new_n5700_ | ~new_n5291_;
  assign new_n21508_ = ~new_n21312_ | ~new_n21506_;
  assign new_n21509_ = new_n5295_ | new_n5697_;
  assign new_n21510_ = ~new_n21423_ | ~new_n21340_;
  assign new_n21511_ = ~new_n21266_;
  assign new_n21512_ = new_n5685_ | new_n5294_;
  assign new_n21513_ = ~new_n21512_ | ~new_n21266_;
  assign new_n21514_ = ~new_n21313_ | ~new_n21513_;
  assign new_n21515_ = ~new_n21511_ | ~new_n21345_;
  assign new_n21516_ = ~new_n5302_ | ~new_n5688_;
  assign new_n21517_ = ~new_n21314_ | ~new_n21515_;
  assign new_n21518_ = new_n5294_ | new_n5685_;
  assign new_n21519_ = new_n5676_ | new_n5305_;
  assign new_n21520_ = ~new_n21519_ | ~new_n21213_;
  assign new_n21521_ = ~new_n21315_ | ~new_n21520_;
  assign new_n21522_ = ~new_n21379_ | ~new_n21344_;
  assign new_n21523_ = ~new_n5284_ | ~new_n5679_;
  assign new_n21524_ = ~new_n21316_ | ~new_n21522_;
  assign new_n21525_ = ~new_n21380_ | ~new_n21344_;
  assign new_n21526_ = ~new_n21377_ | ~new_n21234_;
  assign new_n21527_ = ~new_n21387_ | ~new_n21195_;
  assign new_n21528_ = ~new_n21401_ | ~new_n21207_;
  assign new_n21529_ = ~new_n21404_ | ~new_n21353_;
  assign new_n21530_ = ~new_n21487_ | ~new_n21346_;
  assign new_n21531_ = ~new_n21471_ | ~new_n21349_;
  assign new_n21532_ = ~new_n21502_ | ~new_n21253_;
  assign new_n21533_ = ~new_n21455_ | ~new_n21250_;
  assign new_n21534_ = ~new_n21509_ | ~new_n21232_;
  assign new_n21535_ = ~new_n21518_ | ~new_n21345_;
  assign new_n21536_ = ~new_n21423_ | ~new_n21241_;
  assign new_n21537_ = ~new_n6169_ | ~new_n5276_;
  assign new_n21538_ = ~new_n21469_ | ~new_n21341_;
  assign new_n21539_ = ~new_n5279_ | ~new_n21468_;
  assign new_n21540_ = ~new_n6171_ | ~new_n21468_;
  assign new_n21541_ = ~new_n21474_ | ~new_n21469_ | ~new_n21341_;
  assign new_n21542_ = ~new_n21306_ | ~new_n21328_ | ~new_n21341_;
  assign new_n21543_ = ~new_n21470_ | ~new_n21474_;
  assign new_n21544_ = ~new_n5305_ | ~new_n21212_;
  assign new_n21545_ = ~new_n5676_ | ~new_n21211_;
  assign new_n21546_ = ~new_n21545_ | ~new_n21544_;
  assign new_n21547_ = ~new_n21525_ | ~new_n21213_;
  assign new_n21548_ = ~new_n21546_ | ~new_n21379_;
  assign new_n21549_ = ~new_n5306_ | ~new_n21209_;
  assign new_n21550_ = ~new_n5673_ | ~new_n21210_;
  assign new_n21551_ = ~new_n21550_ | ~new_n21549_;
  assign new_n21552_ = ~new_n21526_ | ~new_n21317_;
  assign new_n21553_ = ~new_n21376_ | ~new_n21551_;
  assign new_n21554_ = ~new_n5292_ | ~new_n21196_;
  assign new_n21555_ = ~new_n5670_ | ~new_n21194_;
  assign new_n21556_ = ~new_n5293_ | ~new_n21192_;
  assign new_n21557_ = ~new_n5667_ | ~new_n21193_;
  assign new_n21558_ = ~new_n21557_ | ~new_n21556_;
  assign new_n21559_ = ~new_n21527_ | ~new_n21214_;
  assign new_n21560_ = ~new_n21558_ | ~new_n21368_;
  assign new_n21561_ = ~new_n5289_ | ~new_n21208_;
  assign new_n21562_ = ~new_n5664_ | ~new_n21199_;
  assign new_n21563_ = ~new_n5282_ | ~new_n21197_;
  assign new_n21564_ = ~new_n5661_ | ~new_n21198_;
  assign new_n21565_ = ~new_n21564_ | ~new_n21563_;
  assign new_n21566_ = ~new_n21528_ | ~new_n21217_;
  assign new_n21567_ = ~new_n21565_ | ~new_n21394_;
  assign new_n21568_ = ~new_n5286_ | ~new_n21205_;
  assign new_n21569_ = ~new_n5658_ | ~new_n21206_;
  assign new_n21570_ = ~new_n21569_ | ~new_n21568_;
  assign new_n21571_ = ~new_n21529_ | ~new_n21318_;
  assign new_n21572_ = ~new_n21403_ | ~new_n21570_;
  assign new_n21573_ = ~new_n5290_ | ~new_n21200_;
  assign new_n21574_ = ~new_n5655_ | ~new_n21201_;
  assign new_n21575_ = ~new_n5277_ | ~new_n21320_;
  assign new_n21576_ = ~new_n6180_ | ~new_n21319_;
  assign new_n21577_ = ~new_n5277_ | ~new_n21320_;
  assign new_n21578_ = ~new_n6180_ | ~new_n21319_;
  assign new_n21579_ = ~new_n21578_ | ~new_n21577_;
  assign new_n21580_ = ~new_n21321_ | ~new_n21322_;
  assign new_n21581_ = ~new_n21478_ | ~new_n21579_;
  assign new_n21582_ = ~new_n5276_ | ~new_n21261_;
  assign new_n21583_ = ~new_n6169_ | ~new_n21260_;
  assign new_n21584_ = ~new_n5276_ | ~new_n21261_;
  assign new_n21585_ = ~new_n6169_ | ~new_n21260_;
  assign new_n21586_ = ~new_n21585_ | ~new_n21584_;
  assign new_n21587_ = ~new_n21323_ | ~new_n21324_;
  assign new_n21588_ = ~new_n21476_ | ~new_n21586_;
  assign new_n21589_ = ~new_n5275_ | ~new_n21219_;
  assign new_n21590_ = ~new_n6170_ | ~new_n21220_;
  assign new_n21591_ = ~new_n5275_ | ~new_n21219_;
  assign new_n21592_ = ~new_n6170_ | ~new_n21220_;
  assign new_n21593_ = ~new_n21592_ | ~new_n21591_;
  assign new_n21594_ = ~new_n21325_ | ~new_n21326_;
  assign new_n21595_ = ~new_n21473_ | ~new_n21593_;
  assign new_n21596_ = ~new_n5279_ | ~new_n21222_;
  assign new_n21597_ = ~new_n6171_ | ~new_n21221_;
  assign new_n21598_ = ~new_n5280_ | ~new_n21223_;
  assign new_n21599_ = ~new_n6172_ | ~new_n21224_;
  assign new_n21600_ = ~new_n21599_ | ~new_n21598_;
  assign new_n21601_ = ~new_n21530_ | ~new_n21262_;
  assign new_n21602_ = ~new_n21600_ | ~new_n21480_;
  assign new_n21603_ = ~new_n5287_ | ~new_n21225_;
  assign new_n21604_ = ~new_n6173_ | ~new_n21226_;
  assign new_n21605_ = ~new_n21604_ | ~new_n21603_;
  assign new_n21606_ = ~new_n21531_ | ~new_n21328_;
  assign new_n21607_ = ~new_n21467_ | ~new_n21605_;
  assign new_n21608_ = ~new_n5288_ | ~new_n21257_;
  assign new_n21609_ = ~new_n6174_ | ~new_n21258_;
  assign new_n21610_ = ~new_n5288_ | ~new_n21257_;
  assign new_n21611_ = ~new_n6174_ | ~new_n21258_;
  assign new_n21612_ = ~new_n21611_ | ~new_n21610_;
  assign new_n21613_ = ~new_n21329_ | ~new_n21330_;
  assign new_n21614_ = ~new_n21463_ | ~new_n21612_;
  assign new_n21615_ = ~new_n5283_ | ~new_n21255_;
  assign new_n21616_ = ~new_n6175_ | ~new_n21256_;
  assign new_n21617_ = ~new_n5283_ | ~new_n21255_;
  assign new_n21618_ = ~new_n6175_ | ~new_n21256_;
  assign new_n21619_ = ~new_n21618_ | ~new_n21617_;
  assign new_n21620_ = ~new_n21331_ | ~new_n21332_;
  assign new_n21621_ = ~new_n21459_ | ~new_n21619_;
  assign new_n21622_ = ~new_n5297_ | ~new_n21227_;
  assign new_n21623_ = ~new_n6176_ | ~new_n21228_;
  assign new_n21624_ = ~new_n5297_ | ~new_n21227_;
  assign new_n21625_ = ~new_n6176_ | ~new_n21228_;
  assign new_n21626_ = ~new_n21625_ | ~new_n21624_;
  assign new_n21627_ = ~new_n5298_ | ~new_n21254_;
  assign new_n21628_ = ~new_n6177_ | ~new_n21263_;
  assign new_n21629_ = ~new_n21355_ | ~new_n21334_;
  assign new_n21630_ = ~new_n21501_ | ~new_n21204_;
  assign new_n21631_ = ~new_n5303_ | ~new_n21251_;
  assign new_n21632_ = ~new_n5705_ | ~new_n21252_;
  assign new_n21633_ = ~new_n21632_ | ~new_n21631_;
  assign new_n21634_ = ~new_n21532_ | ~new_n21264_;
  assign new_n21635_ = ~new_n21633_ | ~new_n21489_;
  assign new_n21636_ = ~new_n5304_ | ~new_n21248_;
  assign new_n21637_ = ~new_n5703_ | ~new_n21249_;
  assign new_n21638_ = ~new_n21637_ | ~new_n21636_;
  assign new_n21639_ = ~new_n21533_ | ~new_n21335_;
  assign new_n21640_ = ~new_n21443_ | ~new_n21638_;
  assign new_n21641_ = ~new_n5291_ | ~new_n21233_;
  assign new_n21642_ = ~new_n5700_ | ~new_n21231_;
  assign new_n21643_ = ~new_n5295_ | ~new_n21229_;
  assign new_n21644_ = ~new_n5697_ | ~new_n21230_;
  assign new_n21645_ = ~new_n21644_ | ~new_n21643_;
  assign new_n21646_ = ~new_n21534_ | ~new_n21265_;
  assign new_n21647_ = ~new_n21645_ | ~new_n21435_;
  assign new_n21648_ = ~new_n5296_ | ~new_n21246_;
  assign new_n21649_ = ~new_n5694_ | ~new_n21247_;
  assign new_n21650_ = ~new_n5296_ | ~new_n21246_;
  assign new_n21651_ = ~new_n5694_ | ~new_n21247_;
  assign new_n21652_ = ~new_n21651_ | ~new_n21650_;
  assign new_n21653_ = ~new_n21336_ | ~new_n21337_;
  assign new_n21654_ = ~new_n21431_ | ~new_n21652_;
  assign new_n21655_ = ~new_n5301_ | ~new_n21244_;
  assign new_n21656_ = ~new_n5691_ | ~new_n21245_;
  assign new_n21657_ = ~new_n5301_ | ~new_n21244_;
  assign new_n21658_ = ~new_n5691_ | ~new_n21245_;
  assign new_n21659_ = ~new_n21658_ | ~new_n21657_;
  assign new_n21660_ = ~new_n21338_ | ~new_n21339_;
  assign new_n21661_ = ~new_n21427_ | ~new_n21659_;
  assign new_n21662_ = ~new_n5302_ | ~new_n21242_;
  assign new_n21663_ = ~new_n5688_ | ~new_n21243_;
  assign new_n21664_ = ~new_n5294_ | ~new_n21237_;
  assign new_n21665_ = ~new_n5685_ | ~new_n21238_;
  assign new_n21666_ = ~new_n21665_ | ~new_n21664_;
  assign new_n21667_ = ~new_n21535_ | ~new_n21266_;
  assign new_n21668_ = ~new_n21666_ | ~new_n21511_;
  assign new_n21669_ = ~new_n5285_ | ~new_n21239_;
  assign new_n21670_ = ~new_n5682_ | ~new_n21240_;
  assign new_n21671_ = ~new_n21670_ | ~new_n21669_;
  assign new_n21672_ = ~new_n21536_ | ~new_n21340_;
  assign new_n21673_ = ~new_n21417_ | ~new_n21671_;
  assign new_n21674_ = ~new_n5284_ | ~new_n21235_;
  assign new_n21675_ = ~new_n5679_ | ~new_n21236_;
  assign new_n21676_ = ~new_n5299_ | ~new_n21202_;
  assign new_n21677_ = ~new_n5647_ | ~new_n21203_;
  assign new_n21678_ = new_n21853_ & new_n21852_;
  assign new_n21679_ = new_n21871_ & new_n21870_;
  assign new_n21680_ = new_n21911_ & new_n21910_;
  assign new_n21681_ = new_n21920_ & new_n21919_;
  assign new_n21682_ = new_n21938_ & new_n21937_;
  assign new_n21683_ = new_n21946_ & new_n21945_;
  assign new_n21684_ = new_n22025_ & new_n22022_;
  assign new_n21685_ = new_n22018_ & new_n22015_;
  assign new_n21686_ = new_n22009_ & new_n22006_;
  assign new_n21687_ = new_n22000_ & new_n21997_;
  assign new_n21688_ = new_n21994_ & new_n21992_;
  assign new_n21689_ = new_n21987_ & new_n21984_;
  assign new_n21690_ = new_n21909_ & new_n21906_;
  assign new_n21691_ = new_n21901_ & new_n21898_;
  assign new_n21692_ = new_n21887_ & new_n21884_;
  assign new_n21693_ = ~new_n5667_;
  assign new_n21694_ = ~new_n5293_;
  assign new_n21695_ = ~new_n5292_;
  assign new_n21696_ = ~new_n5293_ | ~new_n5667_;
  assign new_n21697_ = ~new_n5670_;
  assign new_n21698_ = ~new_n5661_;
  assign new_n21699_ = ~new_n5282_;
  assign new_n21700_ = ~new_n5289_;
  assign new_n21701_ = ~new_n5655_;
  assign new_n21702_ = ~new_n5290_;
  assign new_n21703_ = ~new_n5647_;
  assign new_n21704_ = ~new_n5299_;
  assign new_n21705_ = ~new_n5299_ | ~new_n5647_;
  assign new_n21706_ = ~new_n5658_;
  assign new_n21707_ = ~new_n5286_;
  assign new_n21708_ = ~new_n5282_ | ~new_n5661_;
  assign new_n21709_ = ~new_n5664_;
  assign new_n21710_ = ~new_n5673_;
  assign new_n21711_ = ~new_n5306_;
  assign new_n21712_ = ~new_n5305_;
  assign new_n21713_ = ~new_n5676_;
  assign new_n21714_ = ~new_n21735_ | ~new_n21879_;
  assign new_n21715_ = ~new_n21791_ | ~new_n21867_;
  assign new_n21716_ = ~new_n21856_ | ~new_n21857_;
  assign new_n21717_ = ~new_n5652_ | ~new_n5300_;
  assign new_n21718_ = ~new_n21796_ | ~new_n21893_;
  assign new_n21719_ = ~new_n21890_ | ~new_n21889_;
  assign new_n21720_ = ~new_n6170_;
  assign new_n21721_ = ~new_n5275_;
  assign new_n21722_ = ~new_n5279_;
  assign new_n21723_ = ~new_n6171_;
  assign new_n21724_ = ~new_n6172_;
  assign new_n21725_ = ~new_n5280_;
  assign new_n21726_ = ~new_n6173_;
  assign new_n21727_ = ~new_n5287_;
  assign new_n21728_ = ~new_n6176_;
  assign new_n21729_ = ~new_n5297_;
  assign new_n21730_ = ~new_n5697_;
  assign new_n21731_ = ~new_n5295_;
  assign new_n21732_ = ~new_n5291_;
  assign new_n21733_ = ~new_n5295_ | ~new_n5697_;
  assign new_n21734_ = ~new_n5700_;
  assign new_n21735_ = ~new_n5306_ | ~new_n5673_;
  assign new_n21736_ = ~new_n5679_;
  assign new_n21737_ = ~new_n5284_;
  assign new_n21738_ = ~new_n5685_;
  assign new_n21739_ = ~new_n5294_;
  assign new_n21740_ = ~new_n5682_;
  assign new_n21741_ = ~new_n5285_;
  assign new_n21742_ = ~new_n5285_ | ~new_n5682_;
  assign new_n21743_ = ~new_n5688_;
  assign new_n21744_ = ~new_n5302_;
  assign new_n21745_ = ~new_n5691_;
  assign new_n21746_ = ~new_n5301_;
  assign new_n21747_ = ~new_n5694_;
  assign new_n21748_ = ~new_n5296_;
  assign new_n21749_ = ~new_n5703_;
  assign new_n21750_ = ~new_n5304_;
  assign new_n21751_ = ~new_n5304_ | ~new_n5703_;
  assign new_n21752_ = ~new_n5705_;
  assign new_n21753_ = ~new_n5303_;
  assign new_n21754_ = ~new_n5303_ | ~new_n5705_;
  assign new_n21755_ = ~new_n6177_;
  assign new_n21756_ = ~new_n6175_;
  assign new_n21757_ = ~new_n5283_;
  assign new_n21758_ = ~new_n6174_;
  assign new_n21759_ = ~new_n5288_;
  assign new_n21760_ = ~new_n6171_ | ~new_n5279_;
  assign new_n21761_ = ~new_n5276_;
  assign new_n21762_ = ~new_n6169_;
  assign new_n21763_ = ~new_n21980_ | ~new_n21850_;
  assign new_n21764_ = ~new_n5298_;
  assign new_n21765_ = ~new_n21751_ | ~new_n21989_;
  assign new_n21766_ = ~new_n21935_ | ~new_n21934_;
  assign new_n21767_ = ~new_n21742_ | ~new_n22011_;
  assign new_n21768_ = ~new_n22131_ | ~new_n22130_;
  assign new_n21769_ = ~new_n22178_ | ~new_n22177_;
  assign new_n21770_ = ~new_n22049_ | ~new_n22048_;
  assign new_n21771_ = ~new_n22054_ | ~new_n22053_;
  assign new_n21772_ = ~new_n22061_ | ~new_n22060_;
  assign new_n21773_ = ~new_n22068_ | ~new_n22067_;
  assign new_n21774_ = ~new_n22073_ | ~new_n22072_;
  assign new_n21775_ = ~new_n22082_ | ~new_n22081_;
  assign new_n21776_ = ~new_n22089_ | ~new_n22088_;
  assign new_n21777_ = ~new_n22096_ | ~new_n22095_;
  assign new_n21778_ = ~new_n22103_ | ~new_n22102_;
  assign new_n21779_ = ~new_n22108_ | ~new_n22107_;
  assign new_n21780_ = ~new_n22115_ | ~new_n22114_;
  assign new_n21781_ = ~new_n22122_ | ~new_n22121_;
  assign new_n21782_ = ~new_n22136_ | ~new_n22135_;
  assign new_n21783_ = ~new_n22141_ | ~new_n22140_;
  assign new_n21784_ = ~new_n22148_ | ~new_n22147_;
  assign new_n21785_ = ~new_n22155_ | ~new_n22154_;
  assign new_n21786_ = ~new_n22162_ | ~new_n22161_;
  assign new_n21787_ = ~new_n22169_ | ~new_n22168_;
  assign new_n21788_ = ~new_n22174_ | ~new_n22173_;
  assign new_n21789_ = new_n21863_ & new_n21861_;
  assign new_n21790_ = new_n21678_ & new_n21854_;
  assign new_n21791_ = new_n21868_ & new_n21866_;
  assign new_n21792_ = new_n21875_ & new_n21874_;
  assign new_n21793_ = new_n21696_ & new_n22056_ & new_n22055_;
  assign new_n21794_ = new_n21886_ & new_n21679_;
  assign new_n21795_ = new_n21855_ & new_n21854_;
  assign new_n21796_ = new_n21894_ & new_n21892_;
  assign new_n21797_ = new_n21708_ & new_n22063_ & new_n22062_;
  assign new_n21798_ = new_n21900_ & new_n21678_;
  assign new_n21799_ = new_n21908_ & new_n21855_;
  assign new_n21800_ = new_n21878_ & new_n21680_;
  assign new_n21801_ = new_n21913_ & new_n21845_;
  assign new_n21802_ = new_n21924_ & new_n21681_;
  assign new_n21803_ = new_n21922_ & new_n21846_;
  assign new_n21804_ = new_n21942_ & new_n21941_;
  assign new_n21805_ = new_n21683_ & new_n21956_;
  assign new_n21806_ = new_n21959_ & new_n21954_;
  assign new_n21807_ = new_n21975_ & new_n21972_;
  assign new_n21808_ = new_n22042_ & new_n21976_;
  assign new_n21809_ = new_n21834_ & new_n21952_;
  assign new_n21810_ = new_n21754_ & new_n22129_ & new_n22128_;
  assign new_n21811_ = new_n21999_ & new_n21683_;
  assign new_n21812_ = new_n21733_ & new_n22143_ & new_n22142_;
  assign new_n21813_ = new_n22008_ & new_n21682_;
  assign new_n21814_ = new_n21846_ & new_n22164_ & new_n22163_;
  assign new_n21815_ = new_n22017_ & new_n21681_;
  assign new_n21816_ = new_n21845_ & new_n22176_ & new_n22175_;
  assign new_n21817_ = new_n22024_ & new_n21680_;
  assign new_n21818_ = ~new_n21792_ | ~new_n21876_;
  assign new_n21819_ = ~new_n21891_ | ~new_n21903_;
  assign new_n21820_ = ~new_n5277_;
  assign new_n21821_ = ~new_n6180_;
  assign new_n21822_ = new_n22077_ & new_n22076_;
  assign new_n21823_ = ~new_n22038_ | ~new_n21978_ | ~new_n21843_;
  assign new_n21824_ = new_n22084_ & new_n22083_;
  assign new_n21825_ = ~new_n21808_ | ~new_n22044_ | ~new_n22043_;
  assign new_n21826_ = new_n22091_ & new_n22090_;
  assign new_n21827_ = ~new_n21760_ | ~new_n22039_ | ~new_n21973_;
  assign new_n21828_ = new_n22098_ & new_n22097_;
  assign new_n21829_ = ~new_n21967_ | ~new_n21966_;
  assign new_n21830_ = new_n22110_ & new_n22109_;
  assign new_n21831_ = ~new_n21963_ | ~new_n21962_;
  assign new_n21832_ = new_n22117_ & new_n22116_;
  assign new_n21833_ = ~new_n21806_ | ~new_n21958_;
  assign new_n21834_ = new_n22124_ & new_n22123_;
  assign new_n21835_ = ~new_n21717_ | ~new_n22001_;
  assign new_n21836_ = ~new_n21804_ | ~new_n21943_;
  assign new_n21837_ = new_n22150_ & new_n22149_;
  assign new_n21838_ = ~new_n21931_ | ~new_n21930_;
  assign new_n21839_ = new_n22157_ & new_n22156_;
  assign new_n21840_ = ~new_n21927_ | ~new_n21926_;
  assign new_n21841_ = ~new_n21917_ | ~new_n21916_;
  assign new_n21842_ = ~new_n22041_ | ~new_n22040_;
  assign new_n21843_ = ~new_n5276_ | ~new_n21825_;
  assign new_n21844_ = ~new_n21708_;
  assign new_n21845_ = ~new_n5676_ | ~new_n5305_;
  assign new_n21846_ = ~new_n5294_ | ~new_n5685_;
  assign new_n21847_ = ~new_n5280_ | ~new_n6172_;
  assign new_n21848_ = ~new_n21742_;
  assign new_n21849_ = ~new_n21751_;
  assign new_n21850_ = ~new_n5287_ | ~new_n6173_;
  assign new_n21851_ = ~new_n21735_;
  assign new_n21852_ = new_n5289_ | new_n5664_;
  assign new_n21853_ = new_n5282_ | new_n5661_;
  assign new_n21854_ = new_n5658_ | new_n5286_;
  assign new_n21855_ = new_n5655_ | new_n5290_;
  assign new_n21856_ = ~new_n21705_;
  assign new_n21857_ = new_n5652_ | new_n5300_;
  assign new_n21858_ = ~new_n21716_;
  assign new_n21859_ = ~new_n21717_;
  assign new_n21860_ = ~new_n21716_ | ~new_n21717_;
  assign new_n21861_ = ~new_n5290_ | ~new_n5655_;
  assign new_n21862_ = ~new_n21860_ | ~new_n21855_;
  assign new_n21863_ = ~new_n5286_ | ~new_n5658_;
  assign new_n21864_ = ~new_n21789_ | ~new_n21862_;
  assign new_n21865_ = ~new_n21709_ | ~new_n21708_;
  assign new_n21866_ = ~new_n5289_ | ~new_n21865_;
  assign new_n21867_ = ~new_n21790_ | ~new_n21864_;
  assign new_n21868_ = ~new_n5664_ | ~new_n21844_;
  assign new_n21869_ = ~new_n21715_;
  assign new_n21870_ = new_n5292_ | new_n5670_;
  assign new_n21871_ = new_n5293_ | new_n5667_;
  assign new_n21872_ = ~new_n21696_;
  assign new_n21873_ = ~new_n21697_ | ~new_n21696_;
  assign new_n21874_ = ~new_n5292_ | ~new_n21873_;
  assign new_n21875_ = ~new_n5670_ | ~new_n21872_;
  assign new_n21876_ = ~new_n21679_ | ~new_n21715_;
  assign new_n21877_ = ~new_n21818_;
  assign new_n21878_ = new_n5673_ | new_n5306_;
  assign new_n21879_ = ~new_n21878_ | ~new_n21818_;
  assign new_n21880_ = ~new_n21714_;
  assign new_n21881_ = new_n5305_ | new_n5676_;
  assign new_n21882_ = new_n5667_ | new_n5293_;
  assign new_n21883_ = ~new_n21882_ | ~new_n21715_;
  assign new_n21884_ = ~new_n21793_ | ~new_n21883_;
  assign new_n21885_ = ~new_n21869_ | ~new_n21696_;
  assign new_n21886_ = ~new_n5670_ | ~new_n5292_;
  assign new_n21887_ = ~new_n21794_ | ~new_n21885_;
  assign new_n21888_ = new_n5293_ | new_n5667_;
  assign new_n21889_ = ~new_n21859_ | ~new_n21855_;
  assign new_n21890_ = ~new_n5290_ | ~new_n5655_;
  assign new_n21891_ = ~new_n21719_;
  assign new_n21892_ = ~new_n21795_ | ~new_n21858_;
  assign new_n21893_ = ~new_n21719_ | ~new_n21854_;
  assign new_n21894_ = ~new_n5286_ | ~new_n5658_;
  assign new_n21895_ = ~new_n21718_;
  assign new_n21896_ = new_n5661_ | new_n5282_;
  assign new_n21897_ = ~new_n21896_ | ~new_n21718_;
  assign new_n21898_ = ~new_n21797_ | ~new_n21897_;
  assign new_n21899_ = ~new_n21895_ | ~new_n21708_;
  assign new_n21900_ = ~new_n5664_ | ~new_n5289_;
  assign new_n21901_ = ~new_n21798_ | ~new_n21899_;
  assign new_n21902_ = new_n5282_ | new_n5661_;
  assign new_n21903_ = ~new_n21858_ | ~new_n21855_;
  assign new_n21904_ = ~new_n21819_;
  assign new_n21905_ = ~new_n5286_ | ~new_n5658_;
  assign new_n21906_ = ~new_n22074_ | ~new_n21716_ | ~new_n21717_ | ~new_n22075_;
  assign new_n21907_ = ~new_n21717_ | ~new_n21716_;
  assign new_n21908_ = ~new_n5290_ | ~new_n5655_;
  assign new_n21909_ = ~new_n21799_ | ~new_n21907_;
  assign new_n21910_ = new_n5305_ | new_n5676_;
  assign new_n21911_ = new_n5284_ | new_n5679_;
  assign new_n21912_ = ~new_n21851_ | ~new_n21680_;
  assign new_n21913_ = ~new_n5284_ | ~new_n5679_;
  assign new_n21914_ = ~new_n21801_ | ~new_n21912_;
  assign new_n21915_ = new_n5679_ | new_n5284_;
  assign new_n21916_ = ~new_n21800_ | ~new_n21818_;
  assign new_n21917_ = ~new_n21915_ | ~new_n21914_;
  assign new_n21918_ = ~new_n21841_;
  assign new_n21919_ = new_n5302_ | new_n5688_;
  assign new_n21920_ = new_n5294_ | new_n5685_;
  assign new_n21921_ = ~new_n21848_ | ~new_n21681_;
  assign new_n21922_ = ~new_n5302_ | ~new_n5688_;
  assign new_n21923_ = ~new_n21803_ | ~new_n21921_;
  assign new_n21924_ = new_n5682_ | new_n5285_;
  assign new_n21925_ = new_n5688_ | new_n5302_;
  assign new_n21926_ = ~new_n21802_ | ~new_n21841_;
  assign new_n21927_ = ~new_n21925_ | ~new_n21923_;
  assign new_n21928_ = ~new_n21840_;
  assign new_n21929_ = new_n5691_ | new_n5301_;
  assign new_n21930_ = ~new_n21929_ | ~new_n21840_;
  assign new_n21931_ = ~new_n5301_ | ~new_n5691_;
  assign new_n21932_ = ~new_n21838_;
  assign new_n21933_ = new_n5694_ | new_n5296_;
  assign new_n21934_ = ~new_n21933_ | ~new_n21838_;
  assign new_n21935_ = ~new_n5296_ | ~new_n5694_;
  assign new_n21936_ = ~new_n21766_;
  assign new_n21937_ = new_n5291_ | new_n5700_;
  assign new_n21938_ = new_n5295_ | new_n5697_;
  assign new_n21939_ = ~new_n21733_;
  assign new_n21940_ = ~new_n21734_ | ~new_n21733_;
  assign new_n21941_ = ~new_n5291_ | ~new_n21940_;
  assign new_n21942_ = ~new_n5700_ | ~new_n21939_;
  assign new_n21943_ = ~new_n21682_ | ~new_n21766_;
  assign new_n21944_ = ~new_n21836_;
  assign new_n21945_ = new_n5298_ | new_n6177_;
  assign new_n21946_ = new_n5303_ | new_n5705_;
  assign new_n21947_ = new_n5297_ | new_n6176_;
  assign new_n21948_ = ~new_n21754_;
  assign new_n21949_ = ~new_n6177_ | ~new_n21948_;
  assign new_n21950_ = ~new_n21949_ | ~new_n21764_;
  assign new_n21951_ = ~new_n21754_ | ~new_n21755_;
  assign new_n21952_ = ~new_n21951_ | ~new_n21950_;
  assign new_n21953_ = ~new_n21849_ | ~new_n21683_;
  assign new_n21954_ = ~new_n5297_ | ~new_n6176_;
  assign new_n21955_ = ~new_n21952_ | ~new_n21953_;
  assign new_n21956_ = new_n5703_ | new_n5304_;
  assign new_n21957_ = new_n6176_ | new_n5297_;
  assign new_n21958_ = ~new_n21805_ | ~new_n21947_ | ~new_n21836_;
  assign new_n21959_ = ~new_n21957_ | ~new_n21955_;
  assign new_n21960_ = ~new_n21833_;
  assign new_n21961_ = new_n6175_ | new_n5283_;
  assign new_n21962_ = ~new_n21961_ | ~new_n21833_;
  assign new_n21963_ = ~new_n5283_ | ~new_n6175_;
  assign new_n21964_ = ~new_n21831_;
  assign new_n21965_ = new_n6174_ | new_n5288_;
  assign new_n21966_ = ~new_n21965_ | ~new_n21831_;
  assign new_n21967_ = ~new_n5288_ | ~new_n6174_;
  assign new_n21968_ = ~new_n21829_;
  assign new_n21969_ = new_n5280_ | new_n6172_;
  assign new_n21970_ = ~new_n21850_ | ~new_n21847_;
  assign new_n21971_ = ~new_n21760_;
  assign new_n21972_ = new_n6173_ | new_n5287_;
  assign new_n21973_ = ~new_n21842_ | ~new_n21829_ | ~new_n21972_;
  assign new_n21974_ = ~new_n21827_;
  assign new_n21975_ = new_n6170_ | new_n5275_;
  assign new_n21976_ = ~new_n5275_ | ~new_n6170_;
  assign new_n21977_ = ~new_n21825_;
  assign new_n21978_ = ~new_n6169_ | ~new_n21825_;
  assign new_n21979_ = ~new_n21823_;
  assign new_n21980_ = ~new_n21972_ | ~new_n21829_;
  assign new_n21981_ = ~new_n21763_;
  assign new_n21982_ = new_n6172_ | new_n5280_;
  assign new_n21983_ = ~new_n21982_ | ~new_n21763_;
  assign new_n21984_ = ~new_n21828_ | ~new_n21983_ | ~new_n21847_;
  assign new_n21985_ = ~new_n21981_ | ~new_n21847_;
  assign new_n21986_ = ~new_n6171_ | ~new_n5279_;
  assign new_n21987_ = ~new_n21842_ | ~new_n21985_ | ~new_n21986_;
  assign new_n21988_ = new_n5280_ | new_n6172_;
  assign new_n21989_ = ~new_n21956_ | ~new_n21836_;
  assign new_n21990_ = ~new_n21765_;
  assign new_n21991_ = ~new_n21683_ | ~new_n21765_;
  assign new_n21992_ = ~new_n21809_ | ~new_n21991_;
  assign new_n21993_ = ~new_n21991_ | ~new_n21952_;
  assign new_n21994_ = ~new_n22127_ | ~new_n21993_;
  assign new_n21995_ = new_n5705_ | new_n5303_;
  assign new_n21996_ = ~new_n21995_ | ~new_n21765_;
  assign new_n21997_ = ~new_n21810_ | ~new_n21996_;
  assign new_n21998_ = ~new_n21990_ | ~new_n21754_;
  assign new_n21999_ = ~new_n5298_ | ~new_n6177_;
  assign new_n22000_ = ~new_n21811_ | ~new_n21998_;
  assign new_n22001_ = new_n5652_ | new_n5300_;
  assign new_n22002_ = ~new_n21835_;
  assign new_n22003_ = new_n5303_ | new_n5705_;
  assign new_n22004_ = new_n5697_ | new_n5295_;
  assign new_n22005_ = ~new_n22004_ | ~new_n21766_;
  assign new_n22006_ = ~new_n21812_ | ~new_n22005_;
  assign new_n22007_ = ~new_n21936_ | ~new_n21733_;
  assign new_n22008_ = ~new_n5700_ | ~new_n5291_;
  assign new_n22009_ = ~new_n21813_ | ~new_n22007_;
  assign new_n22010_ = new_n5295_ | new_n5697_;
  assign new_n22011_ = ~new_n21924_ | ~new_n21841_;
  assign new_n22012_ = ~new_n21767_;
  assign new_n22013_ = new_n5685_ | new_n5294_;
  assign new_n22014_ = ~new_n22013_ | ~new_n21767_;
  assign new_n22015_ = ~new_n21814_ | ~new_n22014_;
  assign new_n22016_ = ~new_n22012_ | ~new_n21846_;
  assign new_n22017_ = ~new_n5302_ | ~new_n5688_;
  assign new_n22018_ = ~new_n21815_ | ~new_n22016_;
  assign new_n22019_ = new_n5294_ | new_n5685_;
  assign new_n22020_ = new_n5676_ | new_n5305_;
  assign new_n22021_ = ~new_n22020_ | ~new_n21714_;
  assign new_n22022_ = ~new_n21816_ | ~new_n22021_;
  assign new_n22023_ = ~new_n21880_ | ~new_n21845_;
  assign new_n22024_ = ~new_n5284_ | ~new_n5679_;
  assign new_n22025_ = ~new_n21817_ | ~new_n22023_;
  assign new_n22026_ = ~new_n21881_ | ~new_n21845_;
  assign new_n22027_ = ~new_n21878_ | ~new_n21735_;
  assign new_n22028_ = ~new_n21888_ | ~new_n21696_;
  assign new_n22029_ = ~new_n21902_ | ~new_n21708_;
  assign new_n22030_ = ~new_n21905_ | ~new_n21854_;
  assign new_n22031_ = ~new_n21988_ | ~new_n21847_;
  assign new_n22032_ = ~new_n21972_ | ~new_n21850_;
  assign new_n22033_ = ~new_n22003_ | ~new_n21754_;
  assign new_n22034_ = ~new_n21956_ | ~new_n21751_;
  assign new_n22035_ = ~new_n22010_ | ~new_n21733_;
  assign new_n22036_ = ~new_n22019_ | ~new_n21846_;
  assign new_n22037_ = ~new_n21924_ | ~new_n21742_;
  assign new_n22038_ = ~new_n6169_ | ~new_n5276_;
  assign new_n22039_ = ~new_n21970_ | ~new_n21842_;
  assign new_n22040_ = ~new_n5279_ | ~new_n21969_;
  assign new_n22041_ = ~new_n6171_ | ~new_n21969_;
  assign new_n22042_ = ~new_n21975_ | ~new_n21970_ | ~new_n21842_;
  assign new_n22043_ = ~new_n21807_ | ~new_n21829_ | ~new_n21842_;
  assign new_n22044_ = ~new_n21971_ | ~new_n21975_;
  assign new_n22045_ = ~new_n5305_ | ~new_n21713_;
  assign new_n22046_ = ~new_n5676_ | ~new_n21712_;
  assign new_n22047_ = ~new_n22046_ | ~new_n22045_;
  assign new_n22048_ = ~new_n22026_ | ~new_n21714_;
  assign new_n22049_ = ~new_n22047_ | ~new_n21880_;
  assign new_n22050_ = ~new_n5306_ | ~new_n21710_;
  assign new_n22051_ = ~new_n5673_ | ~new_n21711_;
  assign new_n22052_ = ~new_n22051_ | ~new_n22050_;
  assign new_n22053_ = ~new_n22027_ | ~new_n21818_;
  assign new_n22054_ = ~new_n21877_ | ~new_n22052_;
  assign new_n22055_ = ~new_n5292_ | ~new_n21697_;
  assign new_n22056_ = ~new_n5670_ | ~new_n21695_;
  assign new_n22057_ = ~new_n5293_ | ~new_n21693_;
  assign new_n22058_ = ~new_n5667_ | ~new_n21694_;
  assign new_n22059_ = ~new_n22058_ | ~new_n22057_;
  assign new_n22060_ = ~new_n22028_ | ~new_n21715_;
  assign new_n22061_ = ~new_n22059_ | ~new_n21869_;
  assign new_n22062_ = ~new_n5289_ | ~new_n21709_;
  assign new_n22063_ = ~new_n5664_ | ~new_n21700_;
  assign new_n22064_ = ~new_n5282_ | ~new_n21698_;
  assign new_n22065_ = ~new_n5661_ | ~new_n21699_;
  assign new_n22066_ = ~new_n22065_ | ~new_n22064_;
  assign new_n22067_ = ~new_n22029_ | ~new_n21718_;
  assign new_n22068_ = ~new_n22066_ | ~new_n21895_;
  assign new_n22069_ = ~new_n5286_ | ~new_n21706_;
  assign new_n22070_ = ~new_n5658_ | ~new_n21707_;
  assign new_n22071_ = ~new_n22070_ | ~new_n22069_;
  assign new_n22072_ = ~new_n22030_ | ~new_n21819_;
  assign new_n22073_ = ~new_n21904_ | ~new_n22071_;
  assign new_n22074_ = ~new_n5290_ | ~new_n21701_;
  assign new_n22075_ = ~new_n5655_ | ~new_n21702_;
  assign new_n22076_ = ~new_n5277_ | ~new_n21821_;
  assign new_n22077_ = ~new_n6180_ | ~new_n21820_;
  assign new_n22078_ = ~new_n5277_ | ~new_n21821_;
  assign new_n22079_ = ~new_n6180_ | ~new_n21820_;
  assign new_n22080_ = ~new_n22079_ | ~new_n22078_;
  assign new_n22081_ = ~new_n21822_ | ~new_n21823_;
  assign new_n22082_ = ~new_n21979_ | ~new_n22080_;
  assign new_n22083_ = ~new_n5276_ | ~new_n21762_;
  assign new_n22084_ = ~new_n6169_ | ~new_n21761_;
  assign new_n22085_ = ~new_n5276_ | ~new_n21762_;
  assign new_n22086_ = ~new_n6169_ | ~new_n21761_;
  assign new_n22087_ = ~new_n22086_ | ~new_n22085_;
  assign new_n22088_ = ~new_n21824_ | ~new_n21825_;
  assign new_n22089_ = ~new_n21977_ | ~new_n22087_;
  assign new_n22090_ = ~new_n5275_ | ~new_n21720_;
  assign new_n22091_ = ~new_n6170_ | ~new_n21721_;
  assign new_n22092_ = ~new_n5275_ | ~new_n21720_;
  assign new_n22093_ = ~new_n6170_ | ~new_n21721_;
  assign new_n22094_ = ~new_n22093_ | ~new_n22092_;
  assign new_n22095_ = ~new_n21826_ | ~new_n21827_;
  assign new_n22096_ = ~new_n21974_ | ~new_n22094_;
  assign new_n22097_ = ~new_n5279_ | ~new_n21723_;
  assign new_n22098_ = ~new_n6171_ | ~new_n21722_;
  assign new_n22099_ = ~new_n5280_ | ~new_n21724_;
  assign new_n22100_ = ~new_n6172_ | ~new_n21725_;
  assign new_n22101_ = ~new_n22100_ | ~new_n22099_;
  assign new_n22102_ = ~new_n22031_ | ~new_n21763_;
  assign new_n22103_ = ~new_n22101_ | ~new_n21981_;
  assign new_n22104_ = ~new_n5287_ | ~new_n21726_;
  assign new_n22105_ = ~new_n6173_ | ~new_n21727_;
  assign new_n22106_ = ~new_n22105_ | ~new_n22104_;
  assign new_n22107_ = ~new_n22032_ | ~new_n21829_;
  assign new_n22108_ = ~new_n21968_ | ~new_n22106_;
  assign new_n22109_ = ~new_n5288_ | ~new_n21758_;
  assign new_n22110_ = ~new_n6174_ | ~new_n21759_;
  assign new_n22111_ = ~new_n5288_ | ~new_n21758_;
  assign new_n22112_ = ~new_n6174_ | ~new_n21759_;
  assign new_n22113_ = ~new_n22112_ | ~new_n22111_;
  assign new_n22114_ = ~new_n21830_ | ~new_n21831_;
  assign new_n22115_ = ~new_n21964_ | ~new_n22113_;
  assign new_n22116_ = ~new_n5283_ | ~new_n21756_;
  assign new_n22117_ = ~new_n6175_ | ~new_n21757_;
  assign new_n22118_ = ~new_n5283_ | ~new_n21756_;
  assign new_n22119_ = ~new_n6175_ | ~new_n21757_;
  assign new_n22120_ = ~new_n22119_ | ~new_n22118_;
  assign new_n22121_ = ~new_n21832_ | ~new_n21833_;
  assign new_n22122_ = ~new_n21960_ | ~new_n22120_;
  assign new_n22123_ = ~new_n5297_ | ~new_n21728_;
  assign new_n22124_ = ~new_n6176_ | ~new_n21729_;
  assign new_n22125_ = ~new_n5297_ | ~new_n21728_;
  assign new_n22126_ = ~new_n6176_ | ~new_n21729_;
  assign new_n22127_ = ~new_n22126_ | ~new_n22125_;
  assign new_n22128_ = ~new_n5298_ | ~new_n21755_;
  assign new_n22129_ = ~new_n6177_ | ~new_n21764_;
  assign new_n22130_ = ~new_n21856_ | ~new_n21835_;
  assign new_n22131_ = ~new_n22002_ | ~new_n21705_;
  assign new_n22132_ = ~new_n5303_ | ~new_n21752_;
  assign new_n22133_ = ~new_n5705_ | ~new_n21753_;
  assign new_n22134_ = ~new_n22133_ | ~new_n22132_;
  assign new_n22135_ = ~new_n22033_ | ~new_n21765_;
  assign new_n22136_ = ~new_n22134_ | ~new_n21990_;
  assign new_n22137_ = ~new_n5304_ | ~new_n21749_;
  assign new_n22138_ = ~new_n5703_ | ~new_n21750_;
  assign new_n22139_ = ~new_n22138_ | ~new_n22137_;
  assign new_n22140_ = ~new_n22034_ | ~new_n21836_;
  assign new_n22141_ = ~new_n21944_ | ~new_n22139_;
  assign new_n22142_ = ~new_n5291_ | ~new_n21734_;
  assign new_n22143_ = ~new_n5700_ | ~new_n21732_;
  assign new_n22144_ = ~new_n5295_ | ~new_n21730_;
  assign new_n22145_ = ~new_n5697_ | ~new_n21731_;
  assign new_n22146_ = ~new_n22145_ | ~new_n22144_;
  assign new_n22147_ = ~new_n22035_ | ~new_n21766_;
  assign new_n22148_ = ~new_n22146_ | ~new_n21936_;
  assign new_n22149_ = ~new_n5296_ | ~new_n21747_;
  assign new_n22150_ = ~new_n5694_ | ~new_n21748_;
  assign new_n22151_ = ~new_n5296_ | ~new_n21747_;
  assign new_n22152_ = ~new_n5694_ | ~new_n21748_;
  assign new_n22153_ = ~new_n22152_ | ~new_n22151_;
  assign new_n22154_ = ~new_n21837_ | ~new_n21838_;
  assign new_n22155_ = ~new_n21932_ | ~new_n22153_;
  assign new_n22156_ = ~new_n5301_ | ~new_n21745_;
  assign new_n22157_ = ~new_n5691_ | ~new_n21746_;
  assign new_n22158_ = ~new_n5301_ | ~new_n21745_;
  assign new_n22159_ = ~new_n5691_ | ~new_n21746_;
  assign new_n22160_ = ~new_n22159_ | ~new_n22158_;
  assign new_n22161_ = ~new_n21839_ | ~new_n21840_;
  assign new_n22162_ = ~new_n21928_ | ~new_n22160_;
  assign new_n22163_ = ~new_n5302_ | ~new_n21743_;
  assign new_n22164_ = ~new_n5688_ | ~new_n21744_;
  assign new_n22165_ = ~new_n5294_ | ~new_n21738_;
  assign new_n22166_ = ~new_n5685_ | ~new_n21739_;
  assign new_n22167_ = ~new_n22166_ | ~new_n22165_;
  assign new_n22168_ = ~new_n22036_ | ~new_n21767_;
  assign new_n22169_ = ~new_n22167_ | ~new_n22012_;
  assign new_n22170_ = ~new_n5285_ | ~new_n21740_;
  assign new_n22171_ = ~new_n5682_ | ~new_n21741_;
  assign new_n22172_ = ~new_n22171_ | ~new_n22170_;
  assign new_n22173_ = ~new_n22037_ | ~new_n21841_;
  assign new_n22174_ = ~new_n21918_ | ~new_n22172_;
  assign new_n22175_ = ~new_n5284_ | ~new_n21736_;
  assign new_n22176_ = ~new_n5679_ | ~new_n21737_;
  assign new_n22177_ = ~new_n5299_ | ~new_n21703_;
  assign new_n22178_ = ~new_n5647_ | ~new_n21704_;
  assign new_n22179_ = new_n22396_ & new_n22395_;
  assign new_n22180_ = new_n22409_ & new_n22408_;
  assign new_n22181_ = new_n22439_ & new_n22438_;
  assign new_n22182_ = new_n22455_ & new_n22454_;
  assign new_n22183_ = new_n22467_ & new_n22466_;
  assign new_n22184_ = new_n22181_ & new_n22443_;
  assign new_n22185_ = new_n22180_ & new_n22404_;
  assign new_n22186_ = new_n22184_ & new_n22434_;
  assign new_n22187_ = new_n22703_ & new_n22702_;
  assign new_n22188_ = new_n22526_ & new_n22523_;
  assign new_n22189_ = new_n22517_ & new_n22514_;
  assign new_n22190_ = new_n22510_ & new_n22507_;
  assign new_n22191_ = new_n22560_ & new_n22501_ & new_n22498_;
  assign new_n22192_ = new_n22430_ & new_n22427_;
  assign new_n22193_ = new_n22423_ & new_n22420_;
  assign new_n22194_ = ~new_n5404_;
  assign new_n22195_ = ~new_n5395_;
  assign new_n22196_ = ~new_n5401_;
  assign new_n22197_ = ~new_n5401_ | ~new_n22241_;
  assign new_n22198_ = ~new_n5400_;
  assign new_n22199_ = ~new_n5402_;
  assign new_n22200_ = ~new_n5403_;
  assign new_n22201_ = ~new_n5404_ | ~new_n22244_;
  assign new_n22202_ = ~new_n5399_;
  assign new_n22203_ = ~new_n5397_;
  assign new_n22204_ = ~new_n5397_ | ~new_n22248_;
  assign new_n22205_ = ~new_n5396_;
  assign new_n22206_ = ~new_n5398_;
  assign new_n22207_ = ~new_n5398_ | ~new_n22246_;
  assign new_n22208_ = ~new_n5394_;
  assign new_n22209_ = ~new_n22544_ | ~new_n22413_ | ~new_n22412_;
  assign new_n22210_ = ~new_n22207_ | ~new_n22405_;
  assign new_n22211_ = ~new_n22540_ | ~new_n22541_ | ~new_n22393_;
  assign new_n22212_ = ~new_n5376_;
  assign new_n22213_ = ~new_n5378_;
  assign new_n22214_ = ~new_n5379_;
  assign new_n22215_ = ~new_n5377_;
  assign new_n22216_ = ~new_n5387_;
  assign new_n22217_ = ~new_n5387_ | ~new_n22253_;
  assign new_n22218_ = ~new_n5386_;
  assign new_n22219_ = ~new_n5389_;
  assign new_n22220_ = ~new_n5391_;
  assign new_n22221_ = ~new_n5392_;
  assign new_n22222_ = ~new_n5392_ | ~new_n22257_;
  assign new_n22223_ = ~new_n5390_;
  assign new_n22224_ = ~new_n5393_;
  assign new_n22225_ = ~new_n5393_ | ~new_n22256_;
  assign new_n22226_ = ~new_n5388_;
  assign new_n22227_ = ~new_n5385_;
  assign new_n22228_ = ~new_n5383_;
  assign new_n22229_ = ~new_n5384_;
  assign new_n22230_ = ~new_n5384_ | ~new_n22262_;
  assign new_n22231_ = ~new_n5382_;
  assign new_n22232_ = ~new_n5381_;
  assign new_n22233_ = ~new_n5380_;
  assign new_n22234_ = ~new_n22387_ | ~new_n22496_;
  assign new_n22235_ = ~new_n22230_ | ~new_n22503_;
  assign new_n22236_ = ~new_n22452_ | ~new_n22451_;
  assign new_n22237_ = ~new_n22549_ | ~new_n22445_;
  assign new_n22238_ = ~new_n22222_ | ~new_n22519_;
  assign new_n22239_ = ~new_n22562_ | ~new_n22561_;
  assign new_n22240_ = ~new_n22594_ | ~new_n22593_;
  assign new_n22241_ = ~new_n22582_ | ~new_n22581_;
  assign new_n22242_ = ~new_n22579_ | ~new_n22578_;
  assign new_n22243_ = ~new_n22573_ | ~new_n22572_;
  assign new_n22244_ = ~new_n22576_ | ~new_n22575_;
  assign new_n22245_ = ~new_n22570_ | ~new_n22569_;
  assign new_n22246_ = ~new_n22585_ | ~new_n22584_;
  assign new_n22247_ = ~new_n22588_ | ~new_n22587_;
  assign new_n22248_ = ~new_n22591_ | ~new_n22590_;
  assign new_n22249_ = ~new_n22634_ | ~new_n22633_;
  assign new_n22250_ = ~new_n22682_ | ~new_n22681_;
  assign new_n22251_ = ~new_n22685_ | ~new_n22684_;
  assign new_n22252_ = ~new_n22637_ | ~new_n22636_;
  assign new_n22253_ = ~new_n22661_ | ~new_n22660_;
  assign new_n22254_ = ~new_n22658_ | ~new_n22657_;
  assign new_n22255_ = ~new_n22652_ | ~new_n22651_;
  assign new_n22256_ = ~new_n22640_ | ~new_n22639_;
  assign new_n22257_ = ~new_n22643_ | ~new_n22642_;
  assign new_n22258_ = ~new_n22646_ | ~new_n22645_;
  assign new_n22259_ = ~new_n22649_ | ~new_n22648_;
  assign new_n22260_ = ~new_n22655_ | ~new_n22654_;
  assign new_n22261_ = ~new_n22664_ | ~new_n22663_;
  assign new_n22262_ = ~new_n22673_ | ~new_n22672_;
  assign new_n22263_ = ~new_n22667_ | ~new_n22666_;
  assign new_n22264_ = ~new_n22670_ | ~new_n22669_;
  assign new_n22265_ = ~new_n22676_ | ~new_n22675_;
  assign new_n22266_ = ~new_n22679_ | ~new_n22678_;
  assign new_n22267_ = ~new_n22691_ | ~new_n22690_;
  assign new_n22268_ = ~new_n22798_ | ~new_n22797_;
  assign new_n22269_ = ~new_n22597_ | ~new_n22596_;
  assign new_n22270_ = ~new_n22604_ | ~new_n22603_;
  assign new_n22271_ = ~new_n22611_ | ~new_n22610_;
  assign new_n22272_ = ~new_n22618_ | ~new_n22617_;
  assign new_n22273_ = ~new_n22625_ | ~new_n22624_;
  assign new_n22274_ = ~new_n22632_ | ~new_n22631_;
  assign new_n22275_ = ~new_n22694_ | ~new_n22693_;
  assign new_n22276_ = ~new_n22701_ | ~new_n22700_;
  assign new_n22277_ = ~new_n22708_ | ~new_n22707_;
  assign new_n22278_ = ~new_n22713_ | ~new_n22712_;
  assign new_n22279_ = ~new_n22720_ | ~new_n22719_;
  assign new_n22280_ = ~new_n22727_ | ~new_n22726_;
  assign new_n22281_ = ~new_n22734_ | ~new_n22733_;
  assign new_n22282_ = ~new_n22741_ | ~new_n22740_;
  assign new_n22283_ = ~new_n22746_ | ~new_n22745_;
  assign new_n22284_ = ~new_n22753_ | ~new_n22752_;
  assign new_n22285_ = ~new_n22760_ | ~new_n22759_;
  assign new_n22286_ = ~new_n22767_ | ~new_n22766_;
  assign new_n22287_ = ~new_n22774_ | ~new_n22773_;
  assign new_n22288_ = ~new_n22781_ | ~new_n22780_;
  assign new_n22289_ = ~new_n22786_ | ~new_n22785_;
  assign new_n22290_ = ~new_n22793_ | ~new_n22792_;
  assign new_n22291_ = new_n22399_ & new_n22398_;
  assign new_n22292_ = new_n22415_ & new_n22185_;
  assign new_n22293_ = new_n22547_ & new_n22416_;
  assign new_n22294_ = new_n22204_ & new_n22606_ & new_n22605_;
  assign new_n22295_ = new_n22422_ & new_n22180_;
  assign new_n22296_ = new_n22197_ & new_n22627_ & new_n22626_;
  assign new_n22297_ = new_n22429_ & new_n22179_;
  assign new_n22298_ = new_n22447_ & new_n22186_;
  assign new_n22299_ = new_n22441_ & new_n22382_;
  assign new_n22300_ = new_n22555_ & new_n22448_;
  assign new_n22301_ = new_n22459_ & new_n22458_;
  assign new_n22302_ = new_n22471_ & new_n22183_;
  assign new_n22303_ = new_n22469_ & new_n22383_;
  assign new_n22304_ = new_n22487_ & new_n22378_;
  assign new_n22305_ = new_n22558_ & new_n22493_;
  assign new_n22306_ = new_n22495_ & new_n22485_;
  assign new_n22307_ = new_n22495_ & new_n22487_;
  assign new_n22308_ = new_n22556_ & new_n22494_;
  assign new_n22309_ = ~new_n22688_ | ~new_n22687_;
  assign new_n22310_ = new_n22683_ & new_n22213_;
  assign new_n22311_ = new_n22387_ & new_n22384_;
  assign new_n22312_ = new_n22500_ & new_n22378_;
  assign new_n22313_ = new_n22187_ & new_n22384_;
  assign new_n22314_ = new_n22383_ & new_n22729_ & new_n22728_;
  assign new_n22315_ = new_n22509_ & new_n22183_;
  assign new_n22316_ = new_n22217_ & new_n22755_ & new_n22754_;
  assign new_n22317_ = new_n22516_ & new_n22182_;
  assign new_n22318_ = new_n22382_ & new_n22776_ & new_n22775_;
  assign new_n22319_ = new_n22525_ & new_n22181_;
  assign new_n22320_ = ~new_n22795_ | ~new_n22794_;
  assign new_n22321_ = ~new_n5676_;
  assign new_n22322_ = new_n22565_ & new_n22564_;
  assign new_n22323_ = ~new_n5661_;
  assign new_n22324_ = ~new_n5652_;
  assign new_n22325_ = ~new_n5647_;
  assign new_n22326_ = ~new_n5658_;
  assign new_n22327_ = ~new_n5655_;
  assign new_n22328_ = ~new_n5664_;
  assign new_n22329_ = ~new_n5670_;
  assign new_n22330_ = ~new_n5667_;
  assign new_n22331_ = ~new_n5673_;
  assign new_n22332_ = ~new_n22293_ | ~new_n22546_;
  assign new_n22333_ = new_n22599_ & new_n22598_;
  assign new_n22334_ = ~new_n22545_ | ~new_n22543_;
  assign new_n22335_ = new_n22613_ & new_n22612_;
  assign new_n22336_ = ~new_n22537_ | ~new_n22402_ | ~new_n22380_;
  assign new_n22337_ = new_n22620_ & new_n22619_;
  assign new_n22338_ = ~new_n22291_ | ~new_n22400_;
  assign new_n22339_ = ~new_n6170_;
  assign new_n22340_ = ~new_n6171_;
  assign new_n22341_ = ~new_n5679_;
  assign new_n22342_ = ~new_n5682_;
  assign new_n22343_ = ~new_n5688_;
  assign new_n22344_ = ~new_n5685_;
  assign new_n22345_ = ~new_n5691_;
  assign new_n22346_ = ~new_n5694_;
  assign new_n22347_ = ~new_n5700_;
  assign new_n22348_ = ~new_n5697_;
  assign new_n22349_ = ~new_n5703_;
  assign new_n22350_ = ~new_n6176_;
  assign new_n22351_ = ~new_n6177_;
  assign new_n22352_ = ~new_n5705_;
  assign new_n22353_ = ~new_n6175_;
  assign new_n22354_ = ~new_n6174_;
  assign new_n22355_ = ~new_n6172_;
  assign new_n22356_ = ~new_n6173_;
  assign new_n22357_ = ~new_n6169_;
  assign new_n22358_ = ~new_n5375_;
  assign new_n22359_ = new_n22696_ & new_n22695_;
  assign new_n22360_ = ~new_n22490_ | ~new_n22489_;
  assign new_n22361_ = ~new_n22482_ | ~new_n22481_;
  assign new_n22362_ = new_n22715_ & new_n22714_;
  assign new_n22363_ = ~new_n22478_ | ~new_n22477_;
  assign new_n22364_ = new_n22722_ & new_n22721_;
  assign new_n22365_ = ~new_n22474_ | ~new_n22473_;
  assign new_n22366_ = new_n22736_ & new_n22735_;
  assign new_n22367_ = ~new_n22201_ | ~new_n22389_;
  assign new_n22368_ = ~new_n22464_ | ~new_n22463_;
  assign new_n22369_ = new_n22748_ & new_n22747_;
  assign new_n22370_ = ~new_n22301_ | ~new_n22460_;
  assign new_n22371_ = new_n22762_ & new_n22761_;
  assign new_n22372_ = ~new_n22300_ | ~new_n22554_;
  assign new_n22373_ = new_n22769_ & new_n22768_;
  assign new_n22374_ = ~new_n22553_ | ~new_n22548_;
  assign new_n22375_ = ~new_n22225_ | ~new_n22435_;
  assign new_n22376_ = new_n22788_ & new_n22787_;
  assign new_n22377_ = ~new_n22538_ | ~new_n22432_ | ~new_n22379_;
  assign new_n22378_ = ~new_n22552_ | ~new_n22551_;
  assign new_n22379_ = ~new_n22239_ | ~new_n22332_;
  assign new_n22380_ = ~new_n22245_ | ~new_n22338_;
  assign new_n22381_ = ~new_n22197_;
  assign new_n22382_ = ~new_n5391_ | ~new_n22259_;
  assign new_n22383_ = ~new_n5383_ | ~new_n22264_;
  assign new_n22384_ = ~new_n5378_ | ~new_n22250_;
  assign new_n22385_ = ~new_n22222_;
  assign new_n22386_ = ~new_n22230_;
  assign new_n22387_ = ~new_n5379_ | ~new_n22251_;
  assign new_n22388_ = ~new_n22577_ | ~new_n22194_;
  assign new_n22389_ = ~new_n5403_ | ~new_n22388_;
  assign new_n22390_ = ~new_n22201_;
  assign new_n22391_ = ~new_n22367_;
  assign new_n22392_ = ~new_n22574_ | ~new_n22199_;
  assign new_n22393_ = ~new_n5402_ | ~new_n22243_;
  assign new_n22394_ = ~new_n22211_;
  assign new_n22395_ = ~new_n22580_ | ~new_n22198_;
  assign new_n22396_ = ~new_n22583_ | ~new_n22196_;
  assign new_n22397_ = ~new_n22198_ | ~new_n22197_;
  assign new_n22398_ = ~new_n22242_ | ~new_n22397_;
  assign new_n22399_ = ~new_n5400_ | ~new_n22381_;
  assign new_n22400_ = ~new_n22179_ | ~new_n22211_;
  assign new_n22401_ = ~new_n22338_;
  assign new_n22402_ = ~new_n5399_ | ~new_n22338_;
  assign new_n22403_ = ~new_n22336_;
  assign new_n22404_ = ~new_n22586_ | ~new_n22206_;
  assign new_n22405_ = ~new_n22404_ | ~new_n22336_;
  assign new_n22406_ = ~new_n22207_;
  assign new_n22407_ = ~new_n22210_;
  assign new_n22408_ = ~new_n22589_ | ~new_n22205_;
  assign new_n22409_ = ~new_n22592_ | ~new_n22203_;
  assign new_n22410_ = ~new_n22204_;
  assign new_n22411_ = ~new_n22205_ | ~new_n22204_;
  assign new_n22412_ = ~new_n22247_ | ~new_n22411_;
  assign new_n22413_ = ~new_n5396_ | ~new_n22410_;
  assign new_n22414_ = ~new_n22334_;
  assign new_n22415_ = ~new_n22595_ | ~new_n22195_;
  assign new_n22416_ = ~new_n5395_ | ~new_n22240_;
  assign new_n22417_ = ~new_n22332_;
  assign new_n22418_ = ~new_n22592_ | ~new_n22203_;
  assign new_n22419_ = ~new_n22418_ | ~new_n22210_;
  assign new_n22420_ = ~new_n22294_ | ~new_n22419_;
  assign new_n22421_ = ~new_n22407_ | ~new_n22204_;
  assign new_n22422_ = ~new_n5396_ | ~new_n22247_;
  assign new_n22423_ = ~new_n22295_ | ~new_n22421_;
  assign new_n22424_ = ~new_n22592_ | ~new_n22203_;
  assign new_n22425_ = ~new_n22583_ | ~new_n22196_;
  assign new_n22426_ = ~new_n22425_ | ~new_n22211_;
  assign new_n22427_ = ~new_n22296_ | ~new_n22426_;
  assign new_n22428_ = ~new_n22394_ | ~new_n22197_;
  assign new_n22429_ = ~new_n5400_ | ~new_n22242_;
  assign new_n22430_ = ~new_n22297_ | ~new_n22428_;
  assign new_n22431_ = ~new_n22583_ | ~new_n22196_;
  assign new_n22432_ = ~new_n5394_ | ~new_n22332_;
  assign new_n22433_ = ~new_n22377_;
  assign new_n22434_ = ~new_n22641_ | ~new_n22224_;
  assign new_n22435_ = ~new_n22434_ | ~new_n22377_;
  assign new_n22436_ = ~new_n22225_;
  assign new_n22437_ = ~new_n22375_;
  assign new_n22438_ = ~new_n22647_ | ~new_n22223_;
  assign new_n22439_ = ~new_n22650_ | ~new_n22220_;
  assign new_n22440_ = ~new_n22385_ | ~new_n22181_;
  assign new_n22441_ = ~new_n5390_ | ~new_n22258_;
  assign new_n22442_ = ~new_n22299_ | ~new_n22440_;
  assign new_n22443_ = ~new_n22644_ | ~new_n22221_;
  assign new_n22444_ = ~new_n22647_ | ~new_n22223_;
  assign new_n22445_ = ~new_n22444_ | ~new_n22442_;
  assign new_n22446_ = ~new_n22374_;
  assign new_n22447_ = ~new_n22653_ | ~new_n22219_;
  assign new_n22448_ = ~new_n5389_ | ~new_n22255_;
  assign new_n22449_ = ~new_n22372_;
  assign new_n22450_ = ~new_n22656_ | ~new_n22226_;
  assign new_n22451_ = ~new_n22450_ | ~new_n22372_;
  assign new_n22452_ = ~new_n5388_ | ~new_n22260_;
  assign new_n22453_ = ~new_n22236_;
  assign new_n22454_ = ~new_n22659_ | ~new_n22218_;
  assign new_n22455_ = ~new_n22662_ | ~new_n22216_;
  assign new_n22456_ = ~new_n22217_;
  assign new_n22457_ = ~new_n22218_ | ~new_n22217_;
  assign new_n22458_ = ~new_n22254_ | ~new_n22457_;
  assign new_n22459_ = ~new_n5386_ | ~new_n22456_;
  assign new_n22460_ = ~new_n22182_ | ~new_n22236_;
  assign new_n22461_ = ~new_n22370_;
  assign new_n22462_ = ~new_n22665_ | ~new_n22227_;
  assign new_n22463_ = ~new_n22462_ | ~new_n22370_;
  assign new_n22464_ = ~new_n5385_ | ~new_n22261_;
  assign new_n22465_ = ~new_n22368_;
  assign new_n22466_ = ~new_n22668_ | ~new_n22231_;
  assign new_n22467_ = ~new_n22671_ | ~new_n22228_;
  assign new_n22468_ = ~new_n22386_ | ~new_n22183_;
  assign new_n22469_ = ~new_n5382_ | ~new_n22263_;
  assign new_n22470_ = ~new_n22303_ | ~new_n22468_;
  assign new_n22471_ = ~new_n22674_ | ~new_n22229_;
  assign new_n22472_ = ~new_n22668_ | ~new_n22231_;
  assign new_n22473_ = ~new_n22302_ | ~new_n22368_;
  assign new_n22474_ = ~new_n22472_ | ~new_n22470_;
  assign new_n22475_ = ~new_n22365_;
  assign new_n22476_ = ~new_n22677_ | ~new_n22232_;
  assign new_n22477_ = ~new_n22476_ | ~new_n22365_;
  assign new_n22478_ = ~new_n5381_ | ~new_n22265_;
  assign new_n22479_ = ~new_n22363_;
  assign new_n22480_ = ~new_n22680_ | ~new_n22233_;
  assign new_n22481_ = ~new_n22480_ | ~new_n22363_;
  assign new_n22482_ = ~new_n5380_ | ~new_n22266_;
  assign new_n22483_ = ~new_n22361_;
  assign new_n22484_ = ~new_n22683_ | ~new_n22213_;
  assign new_n22485_ = ~new_n22486_ | ~new_n22387_ | ~new_n22384_;
  assign new_n22486_ = ~new_n5377_ | ~new_n22252_;
  assign new_n22487_ = ~new_n22686_ | ~new_n22214_;
  assign new_n22488_ = ~new_n22638_ | ~new_n22215_;
  assign new_n22489_ = ~new_n22304_ | ~new_n22361_;
  assign new_n22490_ = ~new_n22550_ | ~new_n22485_;
  assign new_n22491_ = ~new_n22360_;
  assign new_n22492_ = ~new_n22635_ | ~new_n22212_;
  assign new_n22493_ = ~new_n5376_ | ~new_n22249_;
  assign new_n22494_ = ~new_n5376_ | ~new_n22249_;
  assign new_n22495_ = ~new_n22635_ | ~new_n22212_;
  assign new_n22496_ = ~new_n22487_ | ~new_n22361_;
  assign new_n22497_ = ~new_n22234_;
  assign new_n22498_ = ~new_n22310_ | ~new_n22187_;
  assign new_n22499_ = ~new_n22311_ | ~new_n22496_;
  assign new_n22500_ = ~new_n5377_ | ~new_n22252_;
  assign new_n22501_ = ~new_n22312_ | ~new_n22499_;
  assign new_n22502_ = ~new_n22683_ | ~new_n22213_;
  assign new_n22503_ = ~new_n22471_ | ~new_n22368_;
  assign new_n22504_ = ~new_n22235_;
  assign new_n22505_ = ~new_n22671_ | ~new_n22228_;
  assign new_n22506_ = ~new_n22505_ | ~new_n22235_;
  assign new_n22507_ = ~new_n22314_ | ~new_n22506_;
  assign new_n22508_ = ~new_n22504_ | ~new_n22383_;
  assign new_n22509_ = ~new_n5382_ | ~new_n22263_;
  assign new_n22510_ = ~new_n22315_ | ~new_n22508_;
  assign new_n22511_ = ~new_n22671_ | ~new_n22228_;
  assign new_n22512_ = ~new_n22662_ | ~new_n22216_;
  assign new_n22513_ = ~new_n22512_ | ~new_n22236_;
  assign new_n22514_ = ~new_n22316_ | ~new_n22513_;
  assign new_n22515_ = ~new_n22453_ | ~new_n22217_;
  assign new_n22516_ = ~new_n5386_ | ~new_n22254_;
  assign new_n22517_ = ~new_n22317_ | ~new_n22515_;
  assign new_n22518_ = ~new_n22662_ | ~new_n22216_;
  assign new_n22519_ = ~new_n22443_ | ~new_n22375_;
  assign new_n22520_ = ~new_n22238_;
  assign new_n22521_ = ~new_n22650_ | ~new_n22220_;
  assign new_n22522_ = ~new_n22521_ | ~new_n22238_;
  assign new_n22523_ = ~new_n22318_ | ~new_n22522_;
  assign new_n22524_ = ~new_n22520_ | ~new_n22382_;
  assign new_n22525_ = ~new_n5390_ | ~new_n22258_;
  assign new_n22526_ = ~new_n22319_ | ~new_n22524_;
  assign new_n22527_ = ~new_n22650_ | ~new_n22220_;
  assign new_n22528_ = ~new_n22424_ | ~new_n22204_;
  assign new_n22529_ = ~new_n22431_ | ~new_n22197_;
  assign new_n22530_ = ~new_n22502_ | ~new_n22384_;
  assign new_n22531_ = ~new_n22487_ | ~new_n22387_;
  assign new_n22532_ = ~new_n22511_ | ~new_n22383_;
  assign new_n22533_ = ~new_n22471_ | ~new_n22230_;
  assign new_n22534_ = ~new_n22518_ | ~new_n22217_;
  assign new_n22535_ = ~new_n22527_ | ~new_n22382_;
  assign new_n22536_ = ~new_n22443_ | ~new_n22222_;
  assign new_n22537_ = ~new_n5399_ | ~new_n22245_;
  assign new_n22538_ = ~new_n5394_ | ~new_n22239_;
  assign new_n22539_ = ~new_n22305_ | ~new_n22489_ | ~new_n22486_;
  assign new_n22540_ = ~new_n22542_ | ~new_n5403_ | ~new_n22388_;
  assign new_n22541_ = ~new_n22390_ | ~new_n22392_;
  assign new_n22542_ = ~new_n22574_ | ~new_n22199_;
  assign new_n22543_ = ~new_n22185_ | ~new_n22336_;
  assign new_n22544_ = ~new_n22406_ | ~new_n22180_;
  assign new_n22545_ = ~new_n22209_;
  assign new_n22546_ = ~new_n22292_ | ~new_n22336_;
  assign new_n22547_ = ~new_n22209_ | ~new_n22415_;
  assign new_n22548_ = ~new_n22186_ | ~new_n22377_;
  assign new_n22549_ = ~new_n22436_ | ~new_n22184_;
  assign new_n22550_ = ~new_n22552_ | ~new_n22551_ | ~new_n22486_;
  assign new_n22551_ = ~new_n22252_ | ~new_n22484_;
  assign new_n22552_ = ~new_n5377_ | ~new_n22484_;
  assign new_n22553_ = ~new_n22237_;
  assign new_n22554_ = ~new_n22298_ | ~new_n22377_;
  assign new_n22555_ = ~new_n22237_ | ~new_n22447_;
  assign new_n22556_ = ~new_n22306_ | ~new_n22550_;
  assign new_n22557_ = ~new_n22307_ | ~new_n22361_ | ~new_n22378_;
  assign new_n22558_ = ~new_n22488_ | ~new_n22559_ | ~new_n22484_;
  assign new_n22559_ = ~new_n22387_ | ~new_n22384_;
  assign new_n22560_ = ~new_n22313_ | ~new_n22497_;
  assign new_n22561_ = ~new_n5404_ | ~new_n22321_;
  assign new_n22562_ = ~new_n5676_ | ~new_n22194_;
  assign new_n22563_ = ~new_n22239_;
  assign new_n22564_ = ~new_n22563_ | ~new_n5394_;
  assign new_n22565_ = ~new_n22239_ | ~new_n22208_;
  assign new_n22566_ = ~new_n22563_ | ~new_n5394_;
  assign new_n22567_ = ~new_n22239_ | ~new_n22208_;
  assign new_n22568_ = ~new_n22567_ | ~new_n22566_;
  assign new_n22569_ = ~new_n5404_ | ~new_n22323_;
  assign new_n22570_ = ~new_n5661_ | ~new_n22194_;
  assign new_n22571_ = ~new_n22245_;
  assign new_n22572_ = ~new_n5404_ | ~new_n22324_;
  assign new_n22573_ = ~new_n5652_ | ~new_n22194_;
  assign new_n22574_ = ~new_n22243_;
  assign new_n22575_ = ~new_n5404_ | ~new_n22325_;
  assign new_n22576_ = ~new_n5647_ | ~new_n22194_;
  assign new_n22577_ = ~new_n22244_;
  assign new_n22578_ = ~new_n5404_ | ~new_n22326_;
  assign new_n22579_ = ~new_n5658_ | ~new_n22194_;
  assign new_n22580_ = ~new_n22242_;
  assign new_n22581_ = ~new_n5404_ | ~new_n22327_;
  assign new_n22582_ = ~new_n5655_ | ~new_n22194_;
  assign new_n22583_ = ~new_n22241_;
  assign new_n22584_ = ~new_n5404_ | ~new_n22328_;
  assign new_n22585_ = ~new_n5664_ | ~new_n22194_;
  assign new_n22586_ = ~new_n22246_;
  assign new_n22587_ = ~new_n5404_ | ~new_n22329_;
  assign new_n22588_ = ~new_n5670_ | ~new_n22194_;
  assign new_n22589_ = ~new_n22247_;
  assign new_n22590_ = ~new_n5404_ | ~new_n22330_;
  assign new_n22591_ = ~new_n5667_ | ~new_n22194_;
  assign new_n22592_ = ~new_n22248_;
  assign new_n22593_ = ~new_n5404_ | ~new_n22331_;
  assign new_n22594_ = ~new_n5673_ | ~new_n22194_;
  assign new_n22595_ = ~new_n22240_;
  assign new_n22596_ = ~new_n22322_ | ~new_n22332_;
  assign new_n22597_ = ~new_n22417_ | ~new_n22568_;
  assign new_n22598_ = ~new_n22595_ | ~new_n5395_;
  assign new_n22599_ = ~new_n22240_ | ~new_n22195_;
  assign new_n22600_ = ~new_n22595_ | ~new_n5395_;
  assign new_n22601_ = ~new_n22240_ | ~new_n22195_;
  assign new_n22602_ = ~new_n22601_ | ~new_n22600_;
  assign new_n22603_ = ~new_n22333_ | ~new_n22334_;
  assign new_n22604_ = ~new_n22414_ | ~new_n22602_;
  assign new_n22605_ = ~new_n22589_ | ~new_n5396_;
  assign new_n22606_ = ~new_n22247_ | ~new_n22205_;
  assign new_n22607_ = ~new_n22592_ | ~new_n5397_;
  assign new_n22608_ = ~new_n22248_ | ~new_n22203_;
  assign new_n22609_ = ~new_n22608_ | ~new_n22607_;
  assign new_n22610_ = ~new_n22528_ | ~new_n22210_;
  assign new_n22611_ = ~new_n22609_ | ~new_n22407_;
  assign new_n22612_ = ~new_n22586_ | ~new_n5398_;
  assign new_n22613_ = ~new_n22246_ | ~new_n22206_;
  assign new_n22614_ = ~new_n22586_ | ~new_n5398_;
  assign new_n22615_ = ~new_n22246_ | ~new_n22206_;
  assign new_n22616_ = ~new_n22615_ | ~new_n22614_;
  assign new_n22617_ = ~new_n22335_ | ~new_n22336_;
  assign new_n22618_ = ~new_n22403_ | ~new_n22616_;
  assign new_n22619_ = ~new_n22571_ | ~new_n5399_;
  assign new_n22620_ = ~new_n22245_ | ~new_n22202_;
  assign new_n22621_ = ~new_n22571_ | ~new_n5399_;
  assign new_n22622_ = ~new_n22245_ | ~new_n22202_;
  assign new_n22623_ = ~new_n22622_ | ~new_n22621_;
  assign new_n22624_ = ~new_n22337_ | ~new_n22338_;
  assign new_n22625_ = ~new_n22401_ | ~new_n22623_;
  assign new_n22626_ = ~new_n22580_ | ~new_n5400_;
  assign new_n22627_ = ~new_n22242_ | ~new_n22198_;
  assign new_n22628_ = ~new_n22583_ | ~new_n5401_;
  assign new_n22629_ = ~new_n22241_ | ~new_n22196_;
  assign new_n22630_ = ~new_n22629_ | ~new_n22628_;
  assign new_n22631_ = ~new_n22529_ | ~new_n22211_;
  assign new_n22632_ = ~new_n22630_ | ~new_n22394_;
  assign new_n22633_ = ~new_n5404_ | ~new_n22339_;
  assign new_n22634_ = ~new_n6170_ | ~new_n22194_;
  assign new_n22635_ = ~new_n22249_;
  assign new_n22636_ = ~new_n5404_ | ~new_n22340_;
  assign new_n22637_ = ~new_n6171_ | ~new_n22194_;
  assign new_n22638_ = ~new_n22252_;
  assign new_n22639_ = ~new_n5404_ | ~new_n22341_;
  assign new_n22640_ = ~new_n5679_ | ~new_n22194_;
  assign new_n22641_ = ~new_n22256_;
  assign new_n22642_ = ~new_n5404_ | ~new_n22342_;
  assign new_n22643_ = ~new_n5682_ | ~new_n22194_;
  assign new_n22644_ = ~new_n22257_;
  assign new_n22645_ = ~new_n5404_ | ~new_n22343_;
  assign new_n22646_ = ~new_n5688_ | ~new_n22194_;
  assign new_n22647_ = ~new_n22258_;
  assign new_n22648_ = ~new_n5404_ | ~new_n22344_;
  assign new_n22649_ = ~new_n5685_ | ~new_n22194_;
  assign new_n22650_ = ~new_n22259_;
  assign new_n22651_ = ~new_n5404_ | ~new_n22345_;
  assign new_n22652_ = ~new_n5691_ | ~new_n22194_;
  assign new_n22653_ = ~new_n22255_;
  assign new_n22654_ = ~new_n5404_ | ~new_n22346_;
  assign new_n22655_ = ~new_n5694_ | ~new_n22194_;
  assign new_n22656_ = ~new_n22260_;
  assign new_n22657_ = ~new_n5404_ | ~new_n22347_;
  assign new_n22658_ = ~new_n5700_ | ~new_n22194_;
  assign new_n22659_ = ~new_n22254_;
  assign new_n22660_ = ~new_n5404_ | ~new_n22348_;
  assign new_n22661_ = ~new_n5697_ | ~new_n22194_;
  assign new_n22662_ = ~new_n22253_;
  assign new_n22663_ = ~new_n5404_ | ~new_n22349_;
  assign new_n22664_ = ~new_n5703_ | ~new_n22194_;
  assign new_n22665_ = ~new_n22261_;
  assign new_n22666_ = ~new_n5404_ | ~new_n22350_;
  assign new_n22667_ = ~new_n6176_ | ~new_n22194_;
  assign new_n22668_ = ~new_n22263_;
  assign new_n22669_ = ~new_n5404_ | ~new_n22351_;
  assign new_n22670_ = ~new_n6177_ | ~new_n22194_;
  assign new_n22671_ = ~new_n22264_;
  assign new_n22672_ = ~new_n5404_ | ~new_n22352_;
  assign new_n22673_ = ~new_n5705_ | ~new_n22194_;
  assign new_n22674_ = ~new_n22262_;
  assign new_n22675_ = ~new_n5404_ | ~new_n22353_;
  assign new_n22676_ = ~new_n6175_ | ~new_n22194_;
  assign new_n22677_ = ~new_n22265_;
  assign new_n22678_ = ~new_n5404_ | ~new_n22354_;
  assign new_n22679_ = ~new_n6174_ | ~new_n22194_;
  assign new_n22680_ = ~new_n22266_;
  assign new_n22681_ = ~new_n5404_ | ~new_n22355_;
  assign new_n22682_ = ~new_n6172_ | ~new_n22194_;
  assign new_n22683_ = ~new_n22250_;
  assign new_n22684_ = ~new_n5404_ | ~new_n22356_;
  assign new_n22685_ = ~new_n6173_ | ~new_n22194_;
  assign new_n22686_ = ~new_n22251_;
  assign new_n22687_ = ~new_n5404_ | ~new_n22357_;
  assign new_n22688_ = ~new_n6169_ | ~new_n22194_;
  assign new_n22689_ = ~new_n22309_;
  assign new_n22690_ = ~new_n5375_ | ~new_n22689_;
  assign new_n22691_ = ~new_n22309_ | ~new_n22358_;
  assign new_n22692_ = ~new_n22267_;
  assign new_n22693_ = ~new_n22692_ | ~new_n22539_ | ~new_n22492_;
  assign new_n22694_ = ~new_n22267_ | ~new_n22308_ | ~new_n22557_;
  assign new_n22695_ = ~new_n22635_ | ~new_n5376_;
  assign new_n22696_ = ~new_n22249_ | ~new_n22212_;
  assign new_n22697_ = ~new_n22635_ | ~new_n5376_;
  assign new_n22698_ = ~new_n22249_ | ~new_n22212_;
  assign new_n22699_ = ~new_n22698_ | ~new_n22697_;
  assign new_n22700_ = ~new_n22359_ | ~new_n22360_;
  assign new_n22701_ = ~new_n22491_ | ~new_n22699_;
  assign new_n22702_ = ~new_n22638_ | ~new_n5377_;
  assign new_n22703_ = ~new_n22252_ | ~new_n22215_;
  assign new_n22704_ = ~new_n22683_ | ~new_n5378_;
  assign new_n22705_ = ~new_n22250_ | ~new_n22213_;
  assign new_n22706_ = ~new_n22705_ | ~new_n22704_;
  assign new_n22707_ = ~new_n22530_ | ~new_n22234_;
  assign new_n22708_ = ~new_n22706_ | ~new_n22497_;
  assign new_n22709_ = ~new_n22686_ | ~new_n5379_;
  assign new_n22710_ = ~new_n22251_ | ~new_n22214_;
  assign new_n22711_ = ~new_n22710_ | ~new_n22709_;
  assign new_n22712_ = ~new_n22531_ | ~new_n22361_;
  assign new_n22713_ = ~new_n22483_ | ~new_n22711_;
  assign new_n22714_ = ~new_n22680_ | ~new_n5380_;
  assign new_n22715_ = ~new_n22266_ | ~new_n22233_;
  assign new_n22716_ = ~new_n22680_ | ~new_n5380_;
  assign new_n22717_ = ~new_n22266_ | ~new_n22233_;
  assign new_n22718_ = ~new_n22717_ | ~new_n22716_;
  assign new_n22719_ = ~new_n22362_ | ~new_n22363_;
  assign new_n22720_ = ~new_n22479_ | ~new_n22718_;
  assign new_n22721_ = ~new_n22677_ | ~new_n5381_;
  assign new_n22722_ = ~new_n22265_ | ~new_n22232_;
  assign new_n22723_ = ~new_n22677_ | ~new_n5381_;
  assign new_n22724_ = ~new_n22265_ | ~new_n22232_;
  assign new_n22725_ = ~new_n22724_ | ~new_n22723_;
  assign new_n22726_ = ~new_n22364_ | ~new_n22365_;
  assign new_n22727_ = ~new_n22475_ | ~new_n22725_;
  assign new_n22728_ = ~new_n22668_ | ~new_n5382_;
  assign new_n22729_ = ~new_n22263_ | ~new_n22231_;
  assign new_n22730_ = ~new_n22671_ | ~new_n5383_;
  assign new_n22731_ = ~new_n22264_ | ~new_n22228_;
  assign new_n22732_ = ~new_n22731_ | ~new_n22730_;
  assign new_n22733_ = ~new_n22532_ | ~new_n22235_;
  assign new_n22734_ = ~new_n22732_ | ~new_n22504_;
  assign new_n22735_ = ~new_n22574_ | ~new_n5402_;
  assign new_n22736_ = ~new_n22243_ | ~new_n22199_;
  assign new_n22737_ = ~new_n22574_ | ~new_n5402_;
  assign new_n22738_ = ~new_n22243_ | ~new_n22199_;
  assign new_n22739_ = ~new_n22738_ | ~new_n22737_;
  assign new_n22740_ = ~new_n22366_ | ~new_n22367_;
  assign new_n22741_ = ~new_n22391_ | ~new_n22739_;
  assign new_n22742_ = ~new_n22674_ | ~new_n5384_;
  assign new_n22743_ = ~new_n22262_ | ~new_n22229_;
  assign new_n22744_ = ~new_n22743_ | ~new_n22742_;
  assign new_n22745_ = ~new_n22533_ | ~new_n22368_;
  assign new_n22746_ = ~new_n22465_ | ~new_n22744_;
  assign new_n22747_ = ~new_n22665_ | ~new_n5385_;
  assign new_n22748_ = ~new_n22261_ | ~new_n22227_;
  assign new_n22749_ = ~new_n22665_ | ~new_n5385_;
  assign new_n22750_ = ~new_n22261_ | ~new_n22227_;
  assign new_n22751_ = ~new_n22750_ | ~new_n22749_;
  assign new_n22752_ = ~new_n22369_ | ~new_n22370_;
  assign new_n22753_ = ~new_n22461_ | ~new_n22751_;
  assign new_n22754_ = ~new_n22659_ | ~new_n5386_;
  assign new_n22755_ = ~new_n22254_ | ~new_n22218_;
  assign new_n22756_ = ~new_n22662_ | ~new_n5387_;
  assign new_n22757_ = ~new_n22253_ | ~new_n22216_;
  assign new_n22758_ = ~new_n22757_ | ~new_n22756_;
  assign new_n22759_ = ~new_n22534_ | ~new_n22236_;
  assign new_n22760_ = ~new_n22758_ | ~new_n22453_;
  assign new_n22761_ = ~new_n22656_ | ~new_n5388_;
  assign new_n22762_ = ~new_n22260_ | ~new_n22226_;
  assign new_n22763_ = ~new_n22656_ | ~new_n5388_;
  assign new_n22764_ = ~new_n22260_ | ~new_n22226_;
  assign new_n22765_ = ~new_n22764_ | ~new_n22763_;
  assign new_n22766_ = ~new_n22371_ | ~new_n22372_;
  assign new_n22767_ = ~new_n22449_ | ~new_n22765_;
  assign new_n22768_ = ~new_n22653_ | ~new_n5389_;
  assign new_n22769_ = ~new_n22255_ | ~new_n22219_;
  assign new_n22770_ = ~new_n22653_ | ~new_n5389_;
  assign new_n22771_ = ~new_n22255_ | ~new_n22219_;
  assign new_n22772_ = ~new_n22771_ | ~new_n22770_;
  assign new_n22773_ = ~new_n22373_ | ~new_n22374_;
  assign new_n22774_ = ~new_n22446_ | ~new_n22772_;
  assign new_n22775_ = ~new_n22647_ | ~new_n5390_;
  assign new_n22776_ = ~new_n22258_ | ~new_n22223_;
  assign new_n22777_ = ~new_n22650_ | ~new_n5391_;
  assign new_n22778_ = ~new_n22259_ | ~new_n22220_;
  assign new_n22779_ = ~new_n22778_ | ~new_n22777_;
  assign new_n22780_ = ~new_n22535_ | ~new_n22238_;
  assign new_n22781_ = ~new_n22779_ | ~new_n22520_;
  assign new_n22782_ = ~new_n22644_ | ~new_n5392_;
  assign new_n22783_ = ~new_n22257_ | ~new_n22221_;
  assign new_n22784_ = ~new_n22783_ | ~new_n22782_;
  assign new_n22785_ = ~new_n22536_ | ~new_n22375_;
  assign new_n22786_ = ~new_n22437_ | ~new_n22784_;
  assign new_n22787_ = ~new_n22641_ | ~new_n5393_;
  assign new_n22788_ = ~new_n22256_ | ~new_n22224_;
  assign new_n22789_ = ~new_n22641_ | ~new_n5393_;
  assign new_n22790_ = ~new_n22256_ | ~new_n22224_;
  assign new_n22791_ = ~new_n22790_ | ~new_n22789_;
  assign new_n22792_ = ~new_n22376_ | ~new_n22377_;
  assign new_n22793_ = ~new_n22433_ | ~new_n22791_;
  assign new_n22794_ = ~new_n22244_ | ~new_n22194_;
  assign new_n22795_ = ~new_n22577_ | ~new_n5404_;
  assign new_n22796_ = ~new_n22320_;
  assign new_n22797_ = ~new_n22796_ | ~new_n5403_;
  assign new_n22798_ = ~new_n22320_ | ~new_n22200_;
  assign new_n22799_ = new_n22974_ & new_n22973_;
  assign new_n22800_ = new_n22992_ & new_n22991_;
  assign new_n22801_ = new_n23032_ & new_n23031_;
  assign new_n22802_ = new_n23041_ & new_n23040_;
  assign new_n22803_ = new_n23059_ & new_n23058_;
  assign new_n22804_ = new_n23067_ & new_n23066_;
  assign new_n22805_ = new_n23146_ & new_n23143_;
  assign new_n22806_ = new_n23139_ & new_n23136_;
  assign new_n22807_ = new_n23130_ & new_n23127_;
  assign new_n22808_ = new_n23121_ & new_n23118_;
  assign new_n22809_ = new_n23115_ & new_n23113_;
  assign new_n22810_ = new_n23108_ & new_n23105_;
  assign new_n22811_ = new_n23030_ & new_n23027_;
  assign new_n22812_ = new_n23022_ & new_n23019_;
  assign new_n22813_ = new_n23008_ & new_n23005_;
  assign new_n22814_ = ~new_n5667_;
  assign new_n22815_ = ~new_n5293_;
  assign new_n22816_ = ~new_n5292_;
  assign new_n22817_ = ~new_n5293_ | ~new_n5667_;
  assign new_n22818_ = ~new_n5670_;
  assign new_n22819_ = ~new_n5661_;
  assign new_n22820_ = ~new_n5282_;
  assign new_n22821_ = ~new_n5289_;
  assign new_n22822_ = ~new_n5655_;
  assign new_n22823_ = ~new_n5290_;
  assign new_n22824_ = ~new_n5647_;
  assign new_n22825_ = ~new_n5299_;
  assign new_n22826_ = ~new_n5299_ | ~new_n5647_;
  assign new_n22827_ = ~new_n5658_;
  assign new_n22828_ = ~new_n5286_;
  assign new_n22829_ = ~new_n5282_ | ~new_n5661_;
  assign new_n22830_ = ~new_n5664_;
  assign new_n22831_ = ~new_n5673_;
  assign new_n22832_ = ~new_n5306_;
  assign new_n22833_ = ~new_n5305_;
  assign new_n22834_ = ~new_n5676_;
  assign new_n22835_ = ~new_n22856_ | ~new_n23000_;
  assign new_n22836_ = ~new_n22912_ | ~new_n22988_;
  assign new_n22837_ = ~new_n22977_ | ~new_n22978_;
  assign new_n22838_ = ~new_n5652_ | ~new_n5300_;
  assign new_n22839_ = ~new_n22917_ | ~new_n23014_;
  assign new_n22840_ = ~new_n23011_ | ~new_n23010_;
  assign new_n22841_ = ~new_n6170_;
  assign new_n22842_ = ~new_n5275_;
  assign new_n22843_ = ~new_n5279_;
  assign new_n22844_ = ~new_n6171_;
  assign new_n22845_ = ~new_n6172_;
  assign new_n22846_ = ~new_n5280_;
  assign new_n22847_ = ~new_n6173_;
  assign new_n22848_ = ~new_n5287_;
  assign new_n22849_ = ~new_n6176_;
  assign new_n22850_ = ~new_n5297_;
  assign new_n22851_ = ~new_n5697_;
  assign new_n22852_ = ~new_n5295_;
  assign new_n22853_ = ~new_n5291_;
  assign new_n22854_ = ~new_n5295_ | ~new_n5697_;
  assign new_n22855_ = ~new_n5700_;
  assign new_n22856_ = ~new_n5306_ | ~new_n5673_;
  assign new_n22857_ = ~new_n5679_;
  assign new_n22858_ = ~new_n5284_;
  assign new_n22859_ = ~new_n5685_;
  assign new_n22860_ = ~new_n5294_;
  assign new_n22861_ = ~new_n5682_;
  assign new_n22862_ = ~new_n5285_;
  assign new_n22863_ = ~new_n5285_ | ~new_n5682_;
  assign new_n22864_ = ~new_n5688_;
  assign new_n22865_ = ~new_n5302_;
  assign new_n22866_ = ~new_n5691_;
  assign new_n22867_ = ~new_n5301_;
  assign new_n22868_ = ~new_n5694_;
  assign new_n22869_ = ~new_n5296_;
  assign new_n22870_ = ~new_n5703_;
  assign new_n22871_ = ~new_n5304_;
  assign new_n22872_ = ~new_n5304_ | ~new_n5703_;
  assign new_n22873_ = ~new_n5705_;
  assign new_n22874_ = ~new_n5303_;
  assign new_n22875_ = ~new_n5303_ | ~new_n5705_;
  assign new_n22876_ = ~new_n6177_;
  assign new_n22877_ = ~new_n6175_;
  assign new_n22878_ = ~new_n5283_;
  assign new_n22879_ = ~new_n6174_;
  assign new_n22880_ = ~new_n5288_;
  assign new_n22881_ = ~new_n6171_ | ~new_n5279_;
  assign new_n22882_ = ~new_n5276_;
  assign new_n22883_ = ~new_n6169_;
  assign new_n22884_ = ~new_n23101_ | ~new_n22971_;
  assign new_n22885_ = ~new_n5298_;
  assign new_n22886_ = ~new_n22872_ | ~new_n23110_;
  assign new_n22887_ = ~new_n23056_ | ~new_n23055_;
  assign new_n22888_ = ~new_n22863_ | ~new_n23132_;
  assign new_n22889_ = ~new_n23252_ | ~new_n23251_;
  assign new_n22890_ = ~new_n23299_ | ~new_n23298_;
  assign new_n22891_ = ~new_n23170_ | ~new_n23169_;
  assign new_n22892_ = ~new_n23175_ | ~new_n23174_;
  assign new_n22893_ = ~new_n23182_ | ~new_n23181_;
  assign new_n22894_ = ~new_n23189_ | ~new_n23188_;
  assign new_n22895_ = ~new_n23194_ | ~new_n23193_;
  assign new_n22896_ = ~new_n23203_ | ~new_n23202_;
  assign new_n22897_ = ~new_n23210_ | ~new_n23209_;
  assign new_n22898_ = ~new_n23217_ | ~new_n23216_;
  assign new_n22899_ = ~new_n23224_ | ~new_n23223_;
  assign new_n22900_ = ~new_n23229_ | ~new_n23228_;
  assign new_n22901_ = ~new_n23236_ | ~new_n23235_;
  assign new_n22902_ = ~new_n23243_ | ~new_n23242_;
  assign new_n22903_ = ~new_n23257_ | ~new_n23256_;
  assign new_n22904_ = ~new_n23262_ | ~new_n23261_;
  assign new_n22905_ = ~new_n23269_ | ~new_n23268_;
  assign new_n22906_ = ~new_n23276_ | ~new_n23275_;
  assign new_n22907_ = ~new_n23283_ | ~new_n23282_;
  assign new_n22908_ = ~new_n23290_ | ~new_n23289_;
  assign new_n22909_ = ~new_n23295_ | ~new_n23294_;
  assign new_n22910_ = new_n22984_ & new_n22982_;
  assign new_n22911_ = new_n22799_ & new_n22975_;
  assign new_n22912_ = new_n22989_ & new_n22987_;
  assign new_n22913_ = new_n22996_ & new_n22995_;
  assign new_n22914_ = new_n22817_ & new_n23177_ & new_n23176_;
  assign new_n22915_ = new_n23007_ & new_n22800_;
  assign new_n22916_ = new_n22976_ & new_n22975_;
  assign new_n22917_ = new_n23015_ & new_n23013_;
  assign new_n22918_ = new_n22829_ & new_n23184_ & new_n23183_;
  assign new_n22919_ = new_n23021_ & new_n22799_;
  assign new_n22920_ = new_n23029_ & new_n22976_;
  assign new_n22921_ = new_n22999_ & new_n22801_;
  assign new_n22922_ = new_n23034_ & new_n22966_;
  assign new_n22923_ = new_n23045_ & new_n22802_;
  assign new_n22924_ = new_n23043_ & new_n22967_;
  assign new_n22925_ = new_n23063_ & new_n23062_;
  assign new_n22926_ = new_n22804_ & new_n23077_;
  assign new_n22927_ = new_n23080_ & new_n23075_;
  assign new_n22928_ = new_n23096_ & new_n23093_;
  assign new_n22929_ = new_n23163_ & new_n23097_;
  assign new_n22930_ = new_n22955_ & new_n23073_;
  assign new_n22931_ = new_n22875_ & new_n23250_ & new_n23249_;
  assign new_n22932_ = new_n23120_ & new_n22804_;
  assign new_n22933_ = new_n22854_ & new_n23264_ & new_n23263_;
  assign new_n22934_ = new_n23129_ & new_n22803_;
  assign new_n22935_ = new_n22967_ & new_n23285_ & new_n23284_;
  assign new_n22936_ = new_n23138_ & new_n22802_;
  assign new_n22937_ = new_n22966_ & new_n23297_ & new_n23296_;
  assign new_n22938_ = new_n23145_ & new_n22801_;
  assign new_n22939_ = ~new_n22913_ | ~new_n22997_;
  assign new_n22940_ = ~new_n23012_ | ~new_n23024_;
  assign new_n22941_ = ~new_n5277_;
  assign new_n22942_ = ~new_n6180_;
  assign new_n22943_ = new_n23198_ & new_n23197_;
  assign new_n22944_ = ~new_n23159_ | ~new_n23099_ | ~new_n22964_;
  assign new_n22945_ = new_n23205_ & new_n23204_;
  assign new_n22946_ = ~new_n22929_ | ~new_n23165_ | ~new_n23164_;
  assign new_n22947_ = new_n23212_ & new_n23211_;
  assign new_n22948_ = ~new_n22881_ | ~new_n23160_ | ~new_n23094_;
  assign new_n22949_ = new_n23219_ & new_n23218_;
  assign new_n22950_ = ~new_n23088_ | ~new_n23087_;
  assign new_n22951_ = new_n23231_ & new_n23230_;
  assign new_n22952_ = ~new_n23084_ | ~new_n23083_;
  assign new_n22953_ = new_n23238_ & new_n23237_;
  assign new_n22954_ = ~new_n22927_ | ~new_n23079_;
  assign new_n22955_ = new_n23245_ & new_n23244_;
  assign new_n22956_ = ~new_n22838_ | ~new_n23122_;
  assign new_n22957_ = ~new_n22925_ | ~new_n23064_;
  assign new_n22958_ = new_n23271_ & new_n23270_;
  assign new_n22959_ = ~new_n23052_ | ~new_n23051_;
  assign new_n22960_ = new_n23278_ & new_n23277_;
  assign new_n22961_ = ~new_n23048_ | ~new_n23047_;
  assign new_n22962_ = ~new_n23038_ | ~new_n23037_;
  assign new_n22963_ = ~new_n23162_ | ~new_n23161_;
  assign new_n22964_ = ~new_n5276_ | ~new_n22946_;
  assign new_n22965_ = ~new_n22829_;
  assign new_n22966_ = ~new_n5676_ | ~new_n5305_;
  assign new_n22967_ = ~new_n5294_ | ~new_n5685_;
  assign new_n22968_ = ~new_n5280_ | ~new_n6172_;
  assign new_n22969_ = ~new_n22863_;
  assign new_n22970_ = ~new_n22872_;
  assign new_n22971_ = ~new_n5287_ | ~new_n6173_;
  assign new_n22972_ = ~new_n22856_;
  assign new_n22973_ = new_n5289_ | new_n5664_;
  assign new_n22974_ = new_n5282_ | new_n5661_;
  assign new_n22975_ = new_n5658_ | new_n5286_;
  assign new_n22976_ = new_n5655_ | new_n5290_;
  assign new_n22977_ = ~new_n22826_;
  assign new_n22978_ = new_n5652_ | new_n5300_;
  assign new_n22979_ = ~new_n22837_;
  assign new_n22980_ = ~new_n22838_;
  assign new_n22981_ = ~new_n22837_ | ~new_n22838_;
  assign new_n22982_ = ~new_n5290_ | ~new_n5655_;
  assign new_n22983_ = ~new_n22981_ | ~new_n22976_;
  assign new_n22984_ = ~new_n5286_ | ~new_n5658_;
  assign new_n22985_ = ~new_n22910_ | ~new_n22983_;
  assign new_n22986_ = ~new_n22830_ | ~new_n22829_;
  assign new_n22987_ = ~new_n5289_ | ~new_n22986_;
  assign new_n22988_ = ~new_n22911_ | ~new_n22985_;
  assign new_n22989_ = ~new_n5664_ | ~new_n22965_;
  assign new_n22990_ = ~new_n22836_;
  assign new_n22991_ = new_n5292_ | new_n5670_;
  assign new_n22992_ = new_n5293_ | new_n5667_;
  assign new_n22993_ = ~new_n22817_;
  assign new_n22994_ = ~new_n22818_ | ~new_n22817_;
  assign new_n22995_ = ~new_n5292_ | ~new_n22994_;
  assign new_n22996_ = ~new_n5670_ | ~new_n22993_;
  assign new_n22997_ = ~new_n22800_ | ~new_n22836_;
  assign new_n22998_ = ~new_n22939_;
  assign new_n22999_ = new_n5673_ | new_n5306_;
  assign new_n23000_ = ~new_n22999_ | ~new_n22939_;
  assign new_n23001_ = ~new_n22835_;
  assign new_n23002_ = new_n5305_ | new_n5676_;
  assign new_n23003_ = new_n5667_ | new_n5293_;
  assign new_n23004_ = ~new_n23003_ | ~new_n22836_;
  assign new_n23005_ = ~new_n22914_ | ~new_n23004_;
  assign new_n23006_ = ~new_n22990_ | ~new_n22817_;
  assign new_n23007_ = ~new_n5670_ | ~new_n5292_;
  assign new_n23008_ = ~new_n22915_ | ~new_n23006_;
  assign new_n23009_ = new_n5293_ | new_n5667_;
  assign new_n23010_ = ~new_n22980_ | ~new_n22976_;
  assign new_n23011_ = ~new_n5290_ | ~new_n5655_;
  assign new_n23012_ = ~new_n22840_;
  assign new_n23013_ = ~new_n22916_ | ~new_n22979_;
  assign new_n23014_ = ~new_n22840_ | ~new_n22975_;
  assign new_n23015_ = ~new_n5286_ | ~new_n5658_;
  assign new_n23016_ = ~new_n22839_;
  assign new_n23017_ = new_n5661_ | new_n5282_;
  assign new_n23018_ = ~new_n23017_ | ~new_n22839_;
  assign new_n23019_ = ~new_n22918_ | ~new_n23018_;
  assign new_n23020_ = ~new_n23016_ | ~new_n22829_;
  assign new_n23021_ = ~new_n5664_ | ~new_n5289_;
  assign new_n23022_ = ~new_n22919_ | ~new_n23020_;
  assign new_n23023_ = new_n5282_ | new_n5661_;
  assign new_n23024_ = ~new_n22979_ | ~new_n22976_;
  assign new_n23025_ = ~new_n22940_;
  assign new_n23026_ = ~new_n5286_ | ~new_n5658_;
  assign new_n23027_ = ~new_n23195_ | ~new_n22837_ | ~new_n22838_ | ~new_n23196_;
  assign new_n23028_ = ~new_n22838_ | ~new_n22837_;
  assign new_n23029_ = ~new_n5290_ | ~new_n5655_;
  assign new_n23030_ = ~new_n22920_ | ~new_n23028_;
  assign new_n23031_ = new_n5305_ | new_n5676_;
  assign new_n23032_ = new_n5284_ | new_n5679_;
  assign new_n23033_ = ~new_n22972_ | ~new_n22801_;
  assign new_n23034_ = ~new_n5284_ | ~new_n5679_;
  assign new_n23035_ = ~new_n22922_ | ~new_n23033_;
  assign new_n23036_ = new_n5679_ | new_n5284_;
  assign new_n23037_ = ~new_n22921_ | ~new_n22939_;
  assign new_n23038_ = ~new_n23036_ | ~new_n23035_;
  assign new_n23039_ = ~new_n22962_;
  assign new_n23040_ = new_n5302_ | new_n5688_;
  assign new_n23041_ = new_n5294_ | new_n5685_;
  assign new_n23042_ = ~new_n22969_ | ~new_n22802_;
  assign new_n23043_ = ~new_n5302_ | ~new_n5688_;
  assign new_n23044_ = ~new_n22924_ | ~new_n23042_;
  assign new_n23045_ = new_n5682_ | new_n5285_;
  assign new_n23046_ = new_n5688_ | new_n5302_;
  assign new_n23047_ = ~new_n22923_ | ~new_n22962_;
  assign new_n23048_ = ~new_n23046_ | ~new_n23044_;
  assign new_n23049_ = ~new_n22961_;
  assign new_n23050_ = new_n5691_ | new_n5301_;
  assign new_n23051_ = ~new_n23050_ | ~new_n22961_;
  assign new_n23052_ = ~new_n5301_ | ~new_n5691_;
  assign new_n23053_ = ~new_n22959_;
  assign new_n23054_ = new_n5694_ | new_n5296_;
  assign new_n23055_ = ~new_n23054_ | ~new_n22959_;
  assign new_n23056_ = ~new_n5296_ | ~new_n5694_;
  assign new_n23057_ = ~new_n22887_;
  assign new_n23058_ = new_n5291_ | new_n5700_;
  assign new_n23059_ = new_n5295_ | new_n5697_;
  assign new_n23060_ = ~new_n22854_;
  assign new_n23061_ = ~new_n22855_ | ~new_n22854_;
  assign new_n23062_ = ~new_n5291_ | ~new_n23061_;
  assign new_n23063_ = ~new_n5700_ | ~new_n23060_;
  assign new_n23064_ = ~new_n22803_ | ~new_n22887_;
  assign new_n23065_ = ~new_n22957_;
  assign new_n23066_ = new_n5298_ | new_n6177_;
  assign new_n23067_ = new_n5303_ | new_n5705_;
  assign new_n23068_ = new_n5297_ | new_n6176_;
  assign new_n23069_ = ~new_n22875_;
  assign new_n23070_ = ~new_n6177_ | ~new_n23069_;
  assign new_n23071_ = ~new_n23070_ | ~new_n22885_;
  assign new_n23072_ = ~new_n22875_ | ~new_n22876_;
  assign new_n23073_ = ~new_n23072_ | ~new_n23071_;
  assign new_n23074_ = ~new_n22970_ | ~new_n22804_;
  assign new_n23075_ = ~new_n5297_ | ~new_n6176_;
  assign new_n23076_ = ~new_n23073_ | ~new_n23074_;
  assign new_n23077_ = new_n5703_ | new_n5304_;
  assign new_n23078_ = new_n6176_ | new_n5297_;
  assign new_n23079_ = ~new_n22926_ | ~new_n23068_ | ~new_n22957_;
  assign new_n23080_ = ~new_n23078_ | ~new_n23076_;
  assign new_n23081_ = ~new_n22954_;
  assign new_n23082_ = new_n6175_ | new_n5283_;
  assign new_n23083_ = ~new_n23082_ | ~new_n22954_;
  assign new_n23084_ = ~new_n5283_ | ~new_n6175_;
  assign new_n23085_ = ~new_n22952_;
  assign new_n23086_ = new_n6174_ | new_n5288_;
  assign new_n23087_ = ~new_n23086_ | ~new_n22952_;
  assign new_n23088_ = ~new_n5288_ | ~new_n6174_;
  assign new_n23089_ = ~new_n22950_;
  assign new_n23090_ = new_n5280_ | new_n6172_;
  assign new_n23091_ = ~new_n22971_ | ~new_n22968_;
  assign new_n23092_ = ~new_n22881_;
  assign new_n23093_ = new_n6173_ | new_n5287_;
  assign new_n23094_ = ~new_n22963_ | ~new_n22950_ | ~new_n23093_;
  assign new_n23095_ = ~new_n22948_;
  assign new_n23096_ = new_n6170_ | new_n5275_;
  assign new_n23097_ = ~new_n5275_ | ~new_n6170_;
  assign new_n23098_ = ~new_n22946_;
  assign new_n23099_ = ~new_n6169_ | ~new_n22946_;
  assign new_n23100_ = ~new_n22944_;
  assign new_n23101_ = ~new_n23093_ | ~new_n22950_;
  assign new_n23102_ = ~new_n22884_;
  assign new_n23103_ = new_n6172_ | new_n5280_;
  assign new_n23104_ = ~new_n23103_ | ~new_n22884_;
  assign new_n23105_ = ~new_n22949_ | ~new_n23104_ | ~new_n22968_;
  assign new_n23106_ = ~new_n23102_ | ~new_n22968_;
  assign new_n23107_ = ~new_n6171_ | ~new_n5279_;
  assign new_n23108_ = ~new_n22963_ | ~new_n23106_ | ~new_n23107_;
  assign new_n23109_ = new_n5280_ | new_n6172_;
  assign new_n23110_ = ~new_n23077_ | ~new_n22957_;
  assign new_n23111_ = ~new_n22886_;
  assign new_n23112_ = ~new_n22804_ | ~new_n22886_;
  assign new_n23113_ = ~new_n22930_ | ~new_n23112_;
  assign new_n23114_ = ~new_n23112_ | ~new_n23073_;
  assign new_n23115_ = ~new_n23248_ | ~new_n23114_;
  assign new_n23116_ = new_n5705_ | new_n5303_;
  assign new_n23117_ = ~new_n23116_ | ~new_n22886_;
  assign new_n23118_ = ~new_n22931_ | ~new_n23117_;
  assign new_n23119_ = ~new_n23111_ | ~new_n22875_;
  assign new_n23120_ = ~new_n5298_ | ~new_n6177_;
  assign new_n23121_ = ~new_n22932_ | ~new_n23119_;
  assign new_n23122_ = new_n5652_ | new_n5300_;
  assign new_n23123_ = ~new_n22956_;
  assign new_n23124_ = new_n5303_ | new_n5705_;
  assign new_n23125_ = new_n5697_ | new_n5295_;
  assign new_n23126_ = ~new_n23125_ | ~new_n22887_;
  assign new_n23127_ = ~new_n22933_ | ~new_n23126_;
  assign new_n23128_ = ~new_n23057_ | ~new_n22854_;
  assign new_n23129_ = ~new_n5700_ | ~new_n5291_;
  assign new_n23130_ = ~new_n22934_ | ~new_n23128_;
  assign new_n23131_ = new_n5295_ | new_n5697_;
  assign new_n23132_ = ~new_n23045_ | ~new_n22962_;
  assign new_n23133_ = ~new_n22888_;
  assign new_n23134_ = new_n5685_ | new_n5294_;
  assign new_n23135_ = ~new_n23134_ | ~new_n22888_;
  assign new_n23136_ = ~new_n22935_ | ~new_n23135_;
  assign new_n23137_ = ~new_n23133_ | ~new_n22967_;
  assign new_n23138_ = ~new_n5302_ | ~new_n5688_;
  assign new_n23139_ = ~new_n22936_ | ~new_n23137_;
  assign new_n23140_ = new_n5294_ | new_n5685_;
  assign new_n23141_ = new_n5676_ | new_n5305_;
  assign new_n23142_ = ~new_n23141_ | ~new_n22835_;
  assign new_n23143_ = ~new_n22937_ | ~new_n23142_;
  assign new_n23144_ = ~new_n23001_ | ~new_n22966_;
  assign new_n23145_ = ~new_n5284_ | ~new_n5679_;
  assign new_n23146_ = ~new_n22938_ | ~new_n23144_;
  assign new_n23147_ = ~new_n23002_ | ~new_n22966_;
  assign new_n23148_ = ~new_n22999_ | ~new_n22856_;
  assign new_n23149_ = ~new_n23009_ | ~new_n22817_;
  assign new_n23150_ = ~new_n23023_ | ~new_n22829_;
  assign new_n23151_ = ~new_n23026_ | ~new_n22975_;
  assign new_n23152_ = ~new_n23109_ | ~new_n22968_;
  assign new_n23153_ = ~new_n23093_ | ~new_n22971_;
  assign new_n23154_ = ~new_n23124_ | ~new_n22875_;
  assign new_n23155_ = ~new_n23077_ | ~new_n22872_;
  assign new_n23156_ = ~new_n23131_ | ~new_n22854_;
  assign new_n23157_ = ~new_n23140_ | ~new_n22967_;
  assign new_n23158_ = ~new_n23045_ | ~new_n22863_;
  assign new_n23159_ = ~new_n6169_ | ~new_n5276_;
  assign new_n23160_ = ~new_n23091_ | ~new_n22963_;
  assign new_n23161_ = ~new_n5279_ | ~new_n23090_;
  assign new_n23162_ = ~new_n6171_ | ~new_n23090_;
  assign new_n23163_ = ~new_n23096_ | ~new_n23091_ | ~new_n22963_;
  assign new_n23164_ = ~new_n22928_ | ~new_n22950_ | ~new_n22963_;
  assign new_n23165_ = ~new_n23092_ | ~new_n23096_;
  assign new_n23166_ = ~new_n5305_ | ~new_n22834_;
  assign new_n23167_ = ~new_n5676_ | ~new_n22833_;
  assign new_n23168_ = ~new_n23167_ | ~new_n23166_;
  assign new_n23169_ = ~new_n23147_ | ~new_n22835_;
  assign new_n23170_ = ~new_n23168_ | ~new_n23001_;
  assign new_n23171_ = ~new_n5306_ | ~new_n22831_;
  assign new_n23172_ = ~new_n5673_ | ~new_n22832_;
  assign new_n23173_ = ~new_n23172_ | ~new_n23171_;
  assign new_n23174_ = ~new_n23148_ | ~new_n22939_;
  assign new_n23175_ = ~new_n22998_ | ~new_n23173_;
  assign new_n23176_ = ~new_n5292_ | ~new_n22818_;
  assign new_n23177_ = ~new_n5670_ | ~new_n22816_;
  assign new_n23178_ = ~new_n5293_ | ~new_n22814_;
  assign new_n23179_ = ~new_n5667_ | ~new_n22815_;
  assign new_n23180_ = ~new_n23179_ | ~new_n23178_;
  assign new_n23181_ = ~new_n23149_ | ~new_n22836_;
  assign new_n23182_ = ~new_n23180_ | ~new_n22990_;
  assign new_n23183_ = ~new_n5289_ | ~new_n22830_;
  assign new_n23184_ = ~new_n5664_ | ~new_n22821_;
  assign new_n23185_ = ~new_n5282_ | ~new_n22819_;
  assign new_n23186_ = ~new_n5661_ | ~new_n22820_;
  assign new_n23187_ = ~new_n23186_ | ~new_n23185_;
  assign new_n23188_ = ~new_n23150_ | ~new_n22839_;
  assign new_n23189_ = ~new_n23187_ | ~new_n23016_;
  assign new_n23190_ = ~new_n5286_ | ~new_n22827_;
  assign new_n23191_ = ~new_n5658_ | ~new_n22828_;
  assign new_n23192_ = ~new_n23191_ | ~new_n23190_;
  assign new_n23193_ = ~new_n23151_ | ~new_n22940_;
  assign new_n23194_ = ~new_n23025_ | ~new_n23192_;
  assign new_n23195_ = ~new_n5290_ | ~new_n22822_;
  assign new_n23196_ = ~new_n5655_ | ~new_n22823_;
  assign new_n23197_ = ~new_n5277_ | ~new_n22942_;
  assign new_n23198_ = ~new_n6180_ | ~new_n22941_;
  assign new_n23199_ = ~new_n5277_ | ~new_n22942_;
  assign new_n23200_ = ~new_n6180_ | ~new_n22941_;
  assign new_n23201_ = ~new_n23200_ | ~new_n23199_;
  assign new_n23202_ = ~new_n22943_ | ~new_n22944_;
  assign new_n23203_ = ~new_n23100_ | ~new_n23201_;
  assign new_n23204_ = ~new_n5276_ | ~new_n22883_;
  assign new_n23205_ = ~new_n6169_ | ~new_n22882_;
  assign new_n23206_ = ~new_n5276_ | ~new_n22883_;
  assign new_n23207_ = ~new_n6169_ | ~new_n22882_;
  assign new_n23208_ = ~new_n23207_ | ~new_n23206_;
  assign new_n23209_ = ~new_n22945_ | ~new_n22946_;
  assign new_n23210_ = ~new_n23098_ | ~new_n23208_;
  assign new_n23211_ = ~new_n5275_ | ~new_n22841_;
  assign new_n23212_ = ~new_n6170_ | ~new_n22842_;
  assign new_n23213_ = ~new_n5275_ | ~new_n22841_;
  assign new_n23214_ = ~new_n6170_ | ~new_n22842_;
  assign new_n23215_ = ~new_n23214_ | ~new_n23213_;
  assign new_n23216_ = ~new_n22947_ | ~new_n22948_;
  assign new_n23217_ = ~new_n23095_ | ~new_n23215_;
  assign new_n23218_ = ~new_n5279_ | ~new_n22844_;
  assign new_n23219_ = ~new_n6171_ | ~new_n22843_;
  assign new_n23220_ = ~new_n5280_ | ~new_n22845_;
  assign new_n23221_ = ~new_n6172_ | ~new_n22846_;
  assign new_n23222_ = ~new_n23221_ | ~new_n23220_;
  assign new_n23223_ = ~new_n23152_ | ~new_n22884_;
  assign new_n23224_ = ~new_n23222_ | ~new_n23102_;
  assign new_n23225_ = ~new_n5287_ | ~new_n22847_;
  assign new_n23226_ = ~new_n6173_ | ~new_n22848_;
  assign new_n23227_ = ~new_n23226_ | ~new_n23225_;
  assign new_n23228_ = ~new_n23153_ | ~new_n22950_;
  assign new_n23229_ = ~new_n23089_ | ~new_n23227_;
  assign new_n23230_ = ~new_n5288_ | ~new_n22879_;
  assign new_n23231_ = ~new_n6174_ | ~new_n22880_;
  assign new_n23232_ = ~new_n5288_ | ~new_n22879_;
  assign new_n23233_ = ~new_n6174_ | ~new_n22880_;
  assign new_n23234_ = ~new_n23233_ | ~new_n23232_;
  assign new_n23235_ = ~new_n22951_ | ~new_n22952_;
  assign new_n23236_ = ~new_n23085_ | ~new_n23234_;
  assign new_n23237_ = ~new_n5283_ | ~new_n22877_;
  assign new_n23238_ = ~new_n6175_ | ~new_n22878_;
  assign new_n23239_ = ~new_n5283_ | ~new_n22877_;
  assign new_n23240_ = ~new_n6175_ | ~new_n22878_;
  assign new_n23241_ = ~new_n23240_ | ~new_n23239_;
  assign new_n23242_ = ~new_n22953_ | ~new_n22954_;
  assign new_n23243_ = ~new_n23081_ | ~new_n23241_;
  assign new_n23244_ = ~new_n5297_ | ~new_n22849_;
  assign new_n23245_ = ~new_n6176_ | ~new_n22850_;
  assign new_n23246_ = ~new_n5297_ | ~new_n22849_;
  assign new_n23247_ = ~new_n6176_ | ~new_n22850_;
  assign new_n23248_ = ~new_n23247_ | ~new_n23246_;
  assign new_n23249_ = ~new_n5298_ | ~new_n22876_;
  assign new_n23250_ = ~new_n6177_ | ~new_n22885_;
  assign new_n23251_ = ~new_n22977_ | ~new_n22956_;
  assign new_n23252_ = ~new_n23123_ | ~new_n22826_;
  assign new_n23253_ = ~new_n5303_ | ~new_n22873_;
  assign new_n23254_ = ~new_n5705_ | ~new_n22874_;
  assign new_n23255_ = ~new_n23254_ | ~new_n23253_;
  assign new_n23256_ = ~new_n23154_ | ~new_n22886_;
  assign new_n23257_ = ~new_n23255_ | ~new_n23111_;
  assign new_n23258_ = ~new_n5304_ | ~new_n22870_;
  assign new_n23259_ = ~new_n5703_ | ~new_n22871_;
  assign new_n23260_ = ~new_n23259_ | ~new_n23258_;
  assign new_n23261_ = ~new_n23155_ | ~new_n22957_;
  assign new_n23262_ = ~new_n23065_ | ~new_n23260_;
  assign new_n23263_ = ~new_n5291_ | ~new_n22855_;
  assign new_n23264_ = ~new_n5700_ | ~new_n22853_;
  assign new_n23265_ = ~new_n5295_ | ~new_n22851_;
  assign new_n23266_ = ~new_n5697_ | ~new_n22852_;
  assign new_n23267_ = ~new_n23266_ | ~new_n23265_;
  assign new_n23268_ = ~new_n23156_ | ~new_n22887_;
  assign new_n23269_ = ~new_n23267_ | ~new_n23057_;
  assign new_n23270_ = ~new_n5296_ | ~new_n22868_;
  assign new_n23271_ = ~new_n5694_ | ~new_n22869_;
  assign new_n23272_ = ~new_n5296_ | ~new_n22868_;
  assign new_n23273_ = ~new_n5694_ | ~new_n22869_;
  assign new_n23274_ = ~new_n23273_ | ~new_n23272_;
  assign new_n23275_ = ~new_n22958_ | ~new_n22959_;
  assign new_n23276_ = ~new_n23053_ | ~new_n23274_;
  assign new_n23277_ = ~new_n5301_ | ~new_n22866_;
  assign new_n23278_ = ~new_n5691_ | ~new_n22867_;
  assign new_n23279_ = ~new_n5301_ | ~new_n22866_;
  assign new_n23280_ = ~new_n5691_ | ~new_n22867_;
  assign new_n23281_ = ~new_n23280_ | ~new_n23279_;
  assign new_n23282_ = ~new_n22960_ | ~new_n22961_;
  assign new_n23283_ = ~new_n23049_ | ~new_n23281_;
  assign new_n23284_ = ~new_n5302_ | ~new_n22864_;
  assign new_n23285_ = ~new_n5688_ | ~new_n22865_;
  assign new_n23286_ = ~new_n5294_ | ~new_n22859_;
  assign new_n23287_ = ~new_n5685_ | ~new_n22860_;
  assign new_n23288_ = ~new_n23287_ | ~new_n23286_;
  assign new_n23289_ = ~new_n23157_ | ~new_n22888_;
  assign new_n23290_ = ~new_n23288_ | ~new_n23133_;
  assign new_n23291_ = ~new_n5285_ | ~new_n22861_;
  assign new_n23292_ = ~new_n5682_ | ~new_n22862_;
  assign new_n23293_ = ~new_n23292_ | ~new_n23291_;
  assign new_n23294_ = ~new_n23158_ | ~new_n22962_;
  assign new_n23295_ = ~new_n23039_ | ~new_n23293_;
  assign new_n23296_ = ~new_n5284_ | ~new_n22857_;
  assign new_n23297_ = ~new_n5679_ | ~new_n22858_;
  assign new_n23298_ = ~new_n5299_ | ~new_n22824_;
  assign new_n23299_ = ~new_n5647_ | ~new_n22825_;
  assign new_n23300_ = new_n23496_ & new_n23495_;
  assign new_n23301_ = new_n23535_ & new_n23534_;
  assign new_n23302_ = new_n23475_ & new_n23550_;
  assign new_n23303_ = new_n23552_ & new_n23551_;
  assign new_n23304_ = new_n23476_ & new_n23576_;
  assign new_n23305_ = new_n23578_ & new_n23577_;
  assign new_n23306_ = ~new_n23638_ | ~new_n23641_;
  assign new_n23307_ = ~new_n23627_ | ~new_n23630_;
  assign new_n23308_ = ~new_n23616_ | ~new_n23619_;
  assign new_n23309_ = ~new_n23608_ | ~new_n23610_;
  assign new_n23310_ = ~new_n23646_ | ~new_n23606_;
  assign new_n23311_ = ~new_n23529_ | ~new_n23531_;
  assign new_n23312_ = ~new_n23521_ | ~new_n23524_;
  assign new_n23313_ = ~new_n23513_ | ~new_n23515_;
  assign new_n23314_ = ~new_n23460_ | ~new_n23644_;
  assign new_n23315_ = ~new_n5670_;
  assign new_n23316_ = ~new_n5664_;
  assign new_n23317_ = ~new_n5655_;
  assign new_n23318_ = ~new_n5647_;
  assign new_n23319_ = ~new_n5300_;
  assign new_n23320_ = ~new_n5658_;
  assign new_n23321_ = ~new_n5290_;
  assign new_n23322_ = ~new_n5290_ | ~new_n23317_;
  assign new_n23323_ = ~new_n5286_;
  assign new_n23324_ = ~new_n5667_;
  assign new_n23325_ = ~new_n5661_;
  assign new_n23326_ = ~new_n5293_;
  assign new_n23327_ = ~new_n5289_;
  assign new_n23328_ = ~new_n5282_;
  assign new_n23329_ = ~new_n5282_ | ~new_n23325_;
  assign new_n23330_ = ~new_n5673_;
  assign new_n23331_ = ~new_n5292_;
  assign new_n23332_ = ~new_n5292_ | ~new_n23315_;
  assign new_n23333_ = ~new_n5306_;
  assign new_n23334_ = ~new_n5676_;
  assign new_n23335_ = ~new_n5305_;
  assign new_n23336_ = ~new_n23502_ | ~new_n23501_;
  assign new_n23337_ = ~new_n23329_ | ~new_n23517_;
  assign new_n23338_ = ~new_n23645_ | ~new_n23486_ | ~new_n23470_;
  assign new_n23339_ = ~new_n6171_;
  assign new_n23340_ = ~new_n5679_;
  assign new_n23341_ = ~new_n5682_;
  assign new_n23342_ = ~new_n5285_;
  assign new_n23343_ = ~new_n5284_;
  assign new_n23344_ = ~new_n5305_ | ~new_n23334_;
  assign new_n23345_ = ~new_n5685_;
  assign new_n23346_ = ~new_n5294_;
  assign new_n23347_ = ~new_n5688_;
  assign new_n23348_ = ~new_n5302_;
  assign new_n23349_ = ~new_n5697_;
  assign new_n23350_ = ~new_n5694_;
  assign new_n23351_ = ~new_n5691_;
  assign new_n23352_ = ~new_n5295_;
  assign new_n23353_ = ~new_n5296_;
  assign new_n23354_ = ~new_n5301_;
  assign new_n23355_ = ~new_n5301_ | ~new_n23351_;
  assign new_n23356_ = ~new_n5700_;
  assign new_n23357_ = ~new_n5291_;
  assign new_n23358_ = ~new_n23562_ | ~new_n23561_;
  assign new_n23359_ = ~new_n5304_;
  assign new_n23360_ = ~new_n5705_;
  assign new_n23361_ = ~new_n5303_;
  assign new_n23362_ = ~new_n6177_;
  assign new_n23363_ = ~new_n5298_;
  assign new_n23364_ = ~new_n6174_;
  assign new_n23365_ = ~new_n6175_;
  assign new_n23366_ = ~new_n6176_;
  assign new_n23367_ = ~new_n5288_;
  assign new_n23368_ = ~new_n5283_;
  assign new_n23369_ = ~new_n5297_;
  assign new_n23370_ = ~new_n5297_ | ~new_n23366_;
  assign new_n23371_ = ~new_n6173_;
  assign new_n23372_ = ~new_n5287_;
  assign new_n23373_ = ~new_n6172_;
  assign new_n23374_ = ~new_n5280_;
  assign new_n23375_ = ~new_n6170_;
  assign new_n23376_ = ~new_n5279_;
  assign new_n23377_ = ~new_n5279_ | ~new_n23339_;
  assign new_n23378_ = ~new_n5275_;
  assign new_n23379_ = ~new_n6169_;
  assign new_n23380_ = ~new_n5276_;
  assign new_n23381_ = ~new_n23422_ | ~new_n23595_;
  assign new_n23382_ = ~new_n23592_ | ~new_n23591_;
  assign new_n23383_ = ~new_n23370_ | ~new_n23612_;
  assign new_n23384_ = ~new_n23355_ | ~new_n23623_;
  assign new_n23385_ = ~new_n23344_ | ~new_n23634_;
  assign new_n23386_ = ~new_n5299_;
  assign new_n23387_ = ~new_n23689_ | ~new_n23688_;
  assign new_n23388_ = ~new_n23703_ | ~new_n23702_;
  assign new_n23389_ = ~new_n23708_ | ~new_n23707_;
  assign new_n23390_ = ~new_n23724_ | ~new_n23723_;
  assign new_n23391_ = ~new_n23729_ | ~new_n23728_;
  assign new_n23392_ = ~new_n23734_ | ~new_n23733_;
  assign new_n23393_ = ~new_n23739_ | ~new_n23738_;
  assign new_n23394_ = ~new_n23744_ | ~new_n23743_;
  assign new_n23395_ = ~new_n23760_ | ~new_n23759_;
  assign new_n23396_ = ~new_n23765_ | ~new_n23764_;
  assign new_n23397_ = ~new_n23650_ | ~new_n23649_;
  assign new_n23398_ = ~new_n23659_ | ~new_n23658_;
  assign new_n23399_ = ~new_n23666_ | ~new_n23665_;
  assign new_n23400_ = ~new_n23670_ | ~new_n23669_;
  assign new_n23401_ = ~new_n23679_ | ~new_n23678_;
  assign new_n23402_ = ~new_n23698_ | ~new_n23697_;
  assign new_n23403_ = ~new_n23715_ | ~new_n23714_;
  assign new_n23404_ = ~new_n23719_ | ~new_n23718_;
  assign new_n23405_ = ~new_n23751_ | ~new_n23750_;
  assign new_n23406_ = ~new_n23755_ | ~new_n23754_;
  assign new_n23407_ = ~new_n23772_ | ~new_n23771_;
  assign new_n23408_ = new_n23488_ & new_n23478_;
  assign new_n23409_ = new_n23491_ & new_n23492_;
  assign new_n23410_ = new_n23479_ & new_n23499_ & new_n23494_;
  assign new_n23411_ = new_n23504_ & new_n23480_;
  assign new_n23412_ = new_n23507_ & new_n23508_;
  assign new_n23413_ = new_n23332_ & new_n23652_ & new_n23651_;
  assign new_n23414_ = new_n23655_ & new_n23480_;
  assign new_n23415_ = new_n23523_ & new_n23300_;
  assign new_n23416_ = new_n23662_ & new_n23479_;
  assign new_n23417_ = new_n23322_ & new_n23672_ & new_n23671_;
  assign new_n23418_ = new_n23675_ & new_n23478_;
  assign new_n23419_ = new_n23474_ & new_n23533_ & new_n23510_;
  assign new_n23420_ = new_n23555_ & new_n23302_;
  assign new_n23421_ = new_n23581_ & new_n23304_;
  assign new_n23422_ = new_n23597_ & new_n23598_;
  assign new_n23423_ = new_n23605_ & new_n23681_ & new_n23680_;
  assign new_n23424_ = new_n23602_ & new_n23684_;
  assign new_n23425_ = ~new_n23686_ | ~new_n23685_;
  assign new_n23426_ = new_n23377_ & new_n23691_ & new_n23690_;
  assign new_n23427_ = new_n23694_ & new_n23477_;
  assign new_n23428_ = ~new_n23700_ | ~new_n23699_;
  assign new_n23429_ = ~new_n23705_ | ~new_n23704_;
  assign new_n23430_ = new_n23618_ & new_n23305_;
  assign new_n23431_ = new_n23711_ & new_n23476_;
  assign new_n23432_ = ~new_n23721_ | ~new_n23720_;
  assign new_n23433_ = ~new_n23726_ | ~new_n23725_;
  assign new_n23434_ = ~new_n23731_ | ~new_n23730_;
  assign new_n23435_ = ~new_n23736_ | ~new_n23735_;
  assign new_n23436_ = ~new_n23741_ | ~new_n23740_;
  assign new_n23437_ = new_n23629_ & new_n23303_;
  assign new_n23438_ = new_n23747_ & new_n23475_;
  assign new_n23439_ = ~new_n23757_ | ~new_n23756_;
  assign new_n23440_ = ~new_n23762_ | ~new_n23761_;
  assign new_n23441_ = new_n23640_ & new_n23301_;
  assign new_n23442_ = new_n23768_ & new_n23474_;
  assign new_n23443_ = new_n23648_ & new_n23647_;
  assign new_n23444_ = ~new_n23412_ | ~new_n23505_;
  assign new_n23445_ = new_n23657_ & new_n23656_;
  assign new_n23446_ = new_n23664_ & new_n23663_;
  assign new_n23447_ = new_n23668_ & new_n23667_;
  assign new_n23448_ = ~new_n23409_ | ~new_n23489_;
  assign new_n23449_ = new_n23677_ & new_n23676_;
  assign new_n23450_ = ~new_n6180_;
  assign new_n23451_ = ~new_n5277_;
  assign new_n23452_ = new_n23696_ & new_n23695_;
  assign new_n23453_ = ~new_n23588_ | ~new_n23587_;
  assign new_n23454_ = ~new_n23584_ | ~new_n23583_;
  assign new_n23455_ = new_n23713_ & new_n23712_;
  assign new_n23456_ = new_n23717_ & new_n23716_;
  assign new_n23457_ = ~new_n23574_ | ~new_n23573_;
  assign new_n23458_ = ~new_n23570_ | ~new_n23569_;
  assign new_n23459_ = ~new_n5652_;
  assign new_n23460_ = ~new_n5647_ | ~new_n23386_;
  assign new_n23461_ = ~new_n23566_ | ~new_n23565_;
  assign new_n23462_ = ~new_n5703_;
  assign new_n23463_ = ~new_n23558_ | ~new_n23557_;
  assign new_n23464_ = new_n23749_ & new_n23748_;
  assign new_n23465_ = new_n23753_ & new_n23752_;
  assign new_n23466_ = ~new_n23548_ | ~new_n23547_;
  assign new_n23467_ = ~new_n23544_ | ~new_n23543_;
  assign new_n23468_ = ~new_n23540_ | ~new_n23539_;
  assign new_n23469_ = new_n23770_ & new_n23769_;
  assign new_n23470_ = ~new_n23460_ | ~new_n23459_;
  assign new_n23471_ = ~new_n23377_;
  assign new_n23472_ = ~new_n23322_;
  assign new_n23473_ = ~new_n23332_;
  assign new_n23474_ = ~new_n5679_ | ~new_n23343_;
  assign new_n23475_ = ~new_n5694_ | ~new_n23353_;
  assign new_n23476_ = ~new_n6175_ | ~new_n23368_;
  assign new_n23477_ = ~new_n6171_ | ~new_n23376_;
  assign new_n23478_ = ~new_n5655_ | ~new_n23321_;
  assign new_n23479_ = ~new_n5664_ | ~new_n23327_;
  assign new_n23480_ = ~new_n5670_ | ~new_n23331_;
  assign new_n23481_ = ~new_n23355_;
  assign new_n23482_ = ~new_n23370_;
  assign new_n23483_ = ~new_n23329_;
  assign new_n23484_ = ~new_n23344_;
  assign new_n23485_ = ~new_n23460_;
  assign new_n23486_ = ~new_n5300_ | ~new_n23460_;
  assign new_n23487_ = ~new_n23338_;
  assign new_n23488_ = ~new_n5658_ | ~new_n23323_;
  assign new_n23489_ = ~new_n23408_ | ~new_n23338_;
  assign new_n23490_ = ~new_n23323_ | ~new_n23322_;
  assign new_n23491_ = ~new_n23490_ | ~new_n23320_;
  assign new_n23492_ = ~new_n5286_ | ~new_n23472_;
  assign new_n23493_ = ~new_n23448_;
  assign new_n23494_ = ~new_n5667_ | ~new_n23326_;
  assign new_n23495_ = ~new_n5293_ | ~new_n23324_;
  assign new_n23496_ = ~new_n5289_ | ~new_n23316_;
  assign new_n23497_ = ~new_n23483_ | ~new_n23479_;
  assign new_n23498_ = ~new_n23300_ | ~new_n23497_;
  assign new_n23499_ = ~new_n5661_ | ~new_n23328_;
  assign new_n23500_ = ~new_n5667_ | ~new_n23326_;
  assign new_n23501_ = ~new_n23448_ | ~new_n23410_;
  assign new_n23502_ = ~new_n23500_ | ~new_n23498_;
  assign new_n23503_ = ~new_n23336_;
  assign new_n23504_ = ~new_n5673_ | ~new_n23333_;
  assign new_n23505_ = ~new_n23411_ | ~new_n23336_;
  assign new_n23506_ = ~new_n23333_ | ~new_n23332_;
  assign new_n23507_ = ~new_n23506_ | ~new_n23330_;
  assign new_n23508_ = ~new_n5306_ | ~new_n23473_;
  assign new_n23509_ = ~new_n23444_;
  assign new_n23510_ = ~new_n5676_ | ~new_n23335_;
  assign new_n23511_ = ~new_n23510_ | ~new_n23344_;
  assign new_n23512_ = ~new_n23503_ | ~new_n23332_;
  assign new_n23513_ = ~new_n23414_ | ~new_n23512_;
  assign new_n23514_ = ~new_n23336_ | ~new_n23480_;
  assign new_n23515_ = ~new_n23413_ | ~new_n23514_;
  assign new_n23516_ = ~new_n23332_ | ~new_n23480_;
  assign new_n23517_ = ~new_n23499_ | ~new_n23448_;
  assign new_n23518_ = ~new_n23337_;
  assign new_n23519_ = ~new_n5289_ | ~new_n23316_;
  assign new_n23520_ = ~new_n23518_ | ~new_n23519_;
  assign new_n23521_ = ~new_n23416_ | ~new_n23520_;
  assign new_n23522_ = ~new_n23337_ | ~new_n23479_;
  assign new_n23523_ = ~new_n5667_ | ~new_n23326_;
  assign new_n23524_ = ~new_n23415_ | ~new_n23522_;
  assign new_n23525_ = ~new_n5289_ | ~new_n23316_;
  assign new_n23526_ = ~new_n23479_ | ~new_n23525_;
  assign new_n23527_ = ~new_n23499_ | ~new_n23329_;
  assign new_n23528_ = ~new_n23487_ | ~new_n23322_;
  assign new_n23529_ = ~new_n23418_ | ~new_n23528_;
  assign new_n23530_ = ~new_n23338_ | ~new_n23478_;
  assign new_n23531_ = ~new_n23417_ | ~new_n23530_;
  assign new_n23532_ = ~new_n23322_ | ~new_n23478_;
  assign new_n23533_ = ~new_n5682_ | ~new_n23342_;
  assign new_n23534_ = ~new_n5285_ | ~new_n23341_;
  assign new_n23535_ = ~new_n5284_ | ~new_n23340_;
  assign new_n23536_ = ~new_n23484_ | ~new_n23474_;
  assign new_n23537_ = ~new_n23301_ | ~new_n23536_;
  assign new_n23538_ = ~new_n5682_ | ~new_n23342_;
  assign new_n23539_ = ~new_n23444_ | ~new_n23419_;
  assign new_n23540_ = ~new_n23538_ | ~new_n23537_;
  assign new_n23541_ = ~new_n23468_;
  assign new_n23542_ = ~new_n5685_ | ~new_n23346_;
  assign new_n23543_ = ~new_n23542_ | ~new_n23468_;
  assign new_n23544_ = ~new_n5294_ | ~new_n23345_;
  assign new_n23545_ = ~new_n23467_;
  assign new_n23546_ = ~new_n5688_ | ~new_n23348_;
  assign new_n23547_ = ~new_n23546_ | ~new_n23467_;
  assign new_n23548_ = ~new_n5302_ | ~new_n23347_;
  assign new_n23549_ = ~new_n23466_;
  assign new_n23550_ = ~new_n5697_ | ~new_n23352_;
  assign new_n23551_ = ~new_n5295_ | ~new_n23349_;
  assign new_n23552_ = ~new_n5296_ | ~new_n23350_;
  assign new_n23553_ = ~new_n23481_ | ~new_n23302_;
  assign new_n23554_ = ~new_n23303_ | ~new_n23553_;
  assign new_n23555_ = ~new_n5691_ | ~new_n23354_;
  assign new_n23556_ = ~new_n5697_ | ~new_n23352_;
  assign new_n23557_ = ~new_n23420_ | ~new_n23466_;
  assign new_n23558_ = ~new_n23556_ | ~new_n23554_;
  assign new_n23559_ = ~new_n23463_;
  assign new_n23560_ = ~new_n5700_ | ~new_n23357_;
  assign new_n23561_ = ~new_n23560_ | ~new_n23463_;
  assign new_n23562_ = ~new_n5291_ | ~new_n23356_;
  assign new_n23563_ = ~new_n23358_;
  assign new_n23564_ = ~new_n23563_ | ~new_n23359_;
  assign new_n23565_ = ~new_n23564_ | ~new_n23462_;
  assign new_n23566_ = ~new_n5304_ | ~new_n23358_;
  assign new_n23567_ = ~new_n23461_;
  assign new_n23568_ = ~new_n5705_ | ~new_n23361_;
  assign new_n23569_ = ~new_n23568_ | ~new_n23461_;
  assign new_n23570_ = ~new_n5303_ | ~new_n23360_;
  assign new_n23571_ = ~new_n23458_;
  assign new_n23572_ = ~new_n6177_ | ~new_n23363_;
  assign new_n23573_ = ~new_n23572_ | ~new_n23458_;
  assign new_n23574_ = ~new_n5298_ | ~new_n23362_;
  assign new_n23575_ = ~new_n23457_;
  assign new_n23576_ = ~new_n6174_ | ~new_n23367_;
  assign new_n23577_ = ~new_n5288_ | ~new_n23364_;
  assign new_n23578_ = ~new_n5283_ | ~new_n23365_;
  assign new_n23579_ = ~new_n23482_ | ~new_n23304_;
  assign new_n23580_ = ~new_n23305_ | ~new_n23579_;
  assign new_n23581_ = ~new_n6176_ | ~new_n23369_;
  assign new_n23582_ = ~new_n6174_ | ~new_n23367_;
  assign new_n23583_ = ~new_n23421_ | ~new_n23457_;
  assign new_n23584_ = ~new_n23582_ | ~new_n23580_;
  assign new_n23585_ = ~new_n23454_;
  assign new_n23586_ = ~new_n6173_ | ~new_n23372_;
  assign new_n23587_ = ~new_n23586_ | ~new_n23454_;
  assign new_n23588_ = ~new_n5287_ | ~new_n23371_;
  assign new_n23589_ = ~new_n23453_;
  assign new_n23590_ = ~new_n6172_ | ~new_n23374_;
  assign new_n23591_ = ~new_n23590_ | ~new_n23453_;
  assign new_n23592_ = ~new_n5280_ | ~new_n23373_;
  assign new_n23593_ = ~new_n23382_;
  assign new_n23594_ = ~new_n6170_ | ~new_n23378_;
  assign new_n23595_ = ~new_n23594_ | ~new_n23382_ | ~new_n23477_;
  assign new_n23596_ = ~new_n23378_ | ~new_n23377_;
  assign new_n23597_ = ~new_n23596_ | ~new_n23375_;
  assign new_n23598_ = ~new_n5275_ | ~new_n23471_;
  assign new_n23599_ = ~new_n23381_;
  assign new_n23600_ = ~new_n5276_ | ~new_n23379_;
  assign new_n23601_ = ~new_n23599_ | ~new_n23600_;
  assign new_n23602_ = ~new_n6169_ | ~new_n23380_;
  assign new_n23603_ = ~new_n6169_ | ~new_n23380_;
  assign new_n23604_ = ~new_n23603_ | ~new_n23381_;
  assign new_n23605_ = ~new_n5276_ | ~new_n23379_;
  assign new_n23606_ = ~new_n23423_ | ~new_n23604_;
  assign new_n23607_ = ~new_n23593_ | ~new_n23377_;
  assign new_n23608_ = ~new_n23427_ | ~new_n23607_;
  assign new_n23609_ = ~new_n23382_ | ~new_n23477_;
  assign new_n23610_ = ~new_n23426_ | ~new_n23609_;
  assign new_n23611_ = ~new_n23377_ | ~new_n23477_;
  assign new_n23612_ = ~new_n23581_ | ~new_n23457_;
  assign new_n23613_ = ~new_n23383_;
  assign new_n23614_ = ~new_n5283_ | ~new_n23365_;
  assign new_n23615_ = ~new_n23613_ | ~new_n23614_;
  assign new_n23616_ = ~new_n23431_ | ~new_n23615_;
  assign new_n23617_ = ~new_n23383_ | ~new_n23476_;
  assign new_n23618_ = ~new_n6174_ | ~new_n23367_;
  assign new_n23619_ = ~new_n23430_ | ~new_n23617_;
  assign new_n23620_ = ~new_n5283_ | ~new_n23365_;
  assign new_n23621_ = ~new_n23476_ | ~new_n23620_;
  assign new_n23622_ = ~new_n23581_ | ~new_n23370_;
  assign new_n23623_ = ~new_n23555_ | ~new_n23466_;
  assign new_n23624_ = ~new_n23384_;
  assign new_n23625_ = ~new_n5296_ | ~new_n23350_;
  assign new_n23626_ = ~new_n23624_ | ~new_n23625_;
  assign new_n23627_ = ~new_n23438_ | ~new_n23626_;
  assign new_n23628_ = ~new_n23384_ | ~new_n23475_;
  assign new_n23629_ = ~new_n5697_ | ~new_n23352_;
  assign new_n23630_ = ~new_n23437_ | ~new_n23628_;
  assign new_n23631_ = ~new_n5296_ | ~new_n23350_;
  assign new_n23632_ = ~new_n23475_ | ~new_n23631_;
  assign new_n23633_ = ~new_n23555_ | ~new_n23355_;
  assign new_n23634_ = ~new_n23510_ | ~new_n23444_;
  assign new_n23635_ = ~new_n23385_;
  assign new_n23636_ = ~new_n5284_ | ~new_n23340_;
  assign new_n23637_ = ~new_n23635_ | ~new_n23636_;
  assign new_n23638_ = ~new_n23442_ | ~new_n23637_;
  assign new_n23639_ = ~new_n23385_ | ~new_n23474_;
  assign new_n23640_ = ~new_n5682_ | ~new_n23342_;
  assign new_n23641_ = ~new_n23441_ | ~new_n23639_;
  assign new_n23642_ = ~new_n5284_ | ~new_n23340_;
  assign new_n23643_ = ~new_n23474_ | ~new_n23642_;
  assign new_n23644_ = ~new_n5299_ | ~new_n23318_;
  assign new_n23645_ = ~new_n5300_ | ~new_n23459_;
  assign new_n23646_ = ~new_n23424_ | ~new_n23601_;
  assign new_n23647_ = ~new_n5676_ | ~new_n23335_;
  assign new_n23648_ = ~new_n5305_ | ~new_n23334_;
  assign new_n23649_ = ~new_n23511_ | ~new_n23444_;
  assign new_n23650_ = ~new_n23509_ | ~new_n23443_;
  assign new_n23651_ = ~new_n5673_ | ~new_n23333_;
  assign new_n23652_ = ~new_n5306_ | ~new_n23330_;
  assign new_n23653_ = ~new_n5673_ | ~new_n23333_;
  assign new_n23654_ = ~new_n5306_ | ~new_n23330_;
  assign new_n23655_ = ~new_n23654_ | ~new_n23653_;
  assign new_n23656_ = ~new_n5670_ | ~new_n23331_;
  assign new_n23657_ = ~new_n5292_ | ~new_n23315_;
  assign new_n23658_ = ~new_n23516_ | ~new_n23336_;
  assign new_n23659_ = ~new_n23445_ | ~new_n23503_;
  assign new_n23660_ = ~new_n5667_ | ~new_n23326_;
  assign new_n23661_ = ~new_n5293_ | ~new_n23324_;
  assign new_n23662_ = ~new_n23661_ | ~new_n23660_;
  assign new_n23663_ = ~new_n5664_ | ~new_n23327_;
  assign new_n23664_ = ~new_n5289_ | ~new_n23316_;
  assign new_n23665_ = ~new_n23526_ | ~new_n23337_;
  assign new_n23666_ = ~new_n23446_ | ~new_n23518_;
  assign new_n23667_ = ~new_n5661_ | ~new_n23328_;
  assign new_n23668_ = ~new_n5282_ | ~new_n23325_;
  assign new_n23669_ = ~new_n23527_ | ~new_n23448_;
  assign new_n23670_ = ~new_n23493_ | ~new_n23447_;
  assign new_n23671_ = ~new_n5658_ | ~new_n23323_;
  assign new_n23672_ = ~new_n5286_ | ~new_n23320_;
  assign new_n23673_ = ~new_n5658_ | ~new_n23323_;
  assign new_n23674_ = ~new_n5286_ | ~new_n23320_;
  assign new_n23675_ = ~new_n23674_ | ~new_n23673_;
  assign new_n23676_ = ~new_n5655_ | ~new_n23321_;
  assign new_n23677_ = ~new_n5290_ | ~new_n23317_;
  assign new_n23678_ = ~new_n23532_ | ~new_n23338_;
  assign new_n23679_ = ~new_n23449_ | ~new_n23487_;
  assign new_n23680_ = ~new_n6180_ | ~new_n23451_;
  assign new_n23681_ = ~new_n5277_ | ~new_n23450_;
  assign new_n23682_ = ~new_n6180_ | ~new_n23451_;
  assign new_n23683_ = ~new_n5277_ | ~new_n23450_;
  assign new_n23684_ = ~new_n23683_ | ~new_n23682_;
  assign new_n23685_ = ~new_n6169_ | ~new_n23380_;
  assign new_n23686_ = ~new_n5276_ | ~new_n23379_;
  assign new_n23687_ = ~new_n23425_;
  assign new_n23688_ = ~new_n23687_ | ~new_n23599_;
  assign new_n23689_ = ~new_n23425_ | ~new_n23381_;
  assign new_n23690_ = ~new_n6170_ | ~new_n23378_;
  assign new_n23691_ = ~new_n5275_ | ~new_n23375_;
  assign new_n23692_ = ~new_n6170_ | ~new_n23378_;
  assign new_n23693_ = ~new_n5275_ | ~new_n23375_;
  assign new_n23694_ = ~new_n23693_ | ~new_n23692_;
  assign new_n23695_ = ~new_n6171_ | ~new_n23376_;
  assign new_n23696_ = ~new_n5279_ | ~new_n23339_;
  assign new_n23697_ = ~new_n23611_ | ~new_n23382_;
  assign new_n23698_ = ~new_n23452_ | ~new_n23593_;
  assign new_n23699_ = ~new_n6172_ | ~new_n23374_;
  assign new_n23700_ = ~new_n5280_ | ~new_n23373_;
  assign new_n23701_ = ~new_n23428_;
  assign new_n23702_ = ~new_n23589_ | ~new_n23701_;
  assign new_n23703_ = ~new_n23428_ | ~new_n23453_;
  assign new_n23704_ = ~new_n6173_ | ~new_n23372_;
  assign new_n23705_ = ~new_n5287_ | ~new_n23371_;
  assign new_n23706_ = ~new_n23429_;
  assign new_n23707_ = ~new_n23585_ | ~new_n23706_;
  assign new_n23708_ = ~new_n23429_ | ~new_n23454_;
  assign new_n23709_ = ~new_n6174_ | ~new_n23367_;
  assign new_n23710_ = ~new_n5288_ | ~new_n23364_;
  assign new_n23711_ = ~new_n23710_ | ~new_n23709_;
  assign new_n23712_ = ~new_n6175_ | ~new_n23368_;
  assign new_n23713_ = ~new_n5283_ | ~new_n23365_;
  assign new_n23714_ = ~new_n23621_ | ~new_n23383_;
  assign new_n23715_ = ~new_n23455_ | ~new_n23613_;
  assign new_n23716_ = ~new_n6176_ | ~new_n23369_;
  assign new_n23717_ = ~new_n5297_ | ~new_n23366_;
  assign new_n23718_ = ~new_n23622_ | ~new_n23457_;
  assign new_n23719_ = ~new_n23575_ | ~new_n23456_;
  assign new_n23720_ = ~new_n6177_ | ~new_n23363_;
  assign new_n23721_ = ~new_n5298_ | ~new_n23362_;
  assign new_n23722_ = ~new_n23432_;
  assign new_n23723_ = ~new_n23571_ | ~new_n23722_;
  assign new_n23724_ = ~new_n23432_ | ~new_n23458_;
  assign new_n23725_ = ~new_n5652_ | ~new_n23319_;
  assign new_n23726_ = ~new_n5300_ | ~new_n23459_;
  assign new_n23727_ = ~new_n23433_;
  assign new_n23728_ = ~new_n23485_ | ~new_n23727_;
  assign new_n23729_ = ~new_n23433_ | ~new_n23460_;
  assign new_n23730_ = ~new_n5705_ | ~new_n23361_;
  assign new_n23731_ = ~new_n5303_ | ~new_n23360_;
  assign new_n23732_ = ~new_n23434_;
  assign new_n23733_ = ~new_n23567_ | ~new_n23732_;
  assign new_n23734_ = ~new_n23434_ | ~new_n23461_;
  assign new_n23735_ = ~new_n5703_ | ~new_n23359_;
  assign new_n23736_ = ~new_n5304_ | ~new_n23462_;
  assign new_n23737_ = ~new_n23435_;
  assign new_n23738_ = ~new_n23737_ | ~new_n23563_;
  assign new_n23739_ = ~new_n23435_ | ~new_n23358_;
  assign new_n23740_ = ~new_n5700_ | ~new_n23357_;
  assign new_n23741_ = ~new_n5291_ | ~new_n23356_;
  assign new_n23742_ = ~new_n23436_;
  assign new_n23743_ = ~new_n23559_ | ~new_n23742_;
  assign new_n23744_ = ~new_n23436_ | ~new_n23463_;
  assign new_n23745_ = ~new_n5697_ | ~new_n23352_;
  assign new_n23746_ = ~new_n5295_ | ~new_n23349_;
  assign new_n23747_ = ~new_n23746_ | ~new_n23745_;
  assign new_n23748_ = ~new_n5694_ | ~new_n23353_;
  assign new_n23749_ = ~new_n5296_ | ~new_n23350_;
  assign new_n23750_ = ~new_n23632_ | ~new_n23384_;
  assign new_n23751_ = ~new_n23464_ | ~new_n23624_;
  assign new_n23752_ = ~new_n5691_ | ~new_n23354_;
  assign new_n23753_ = ~new_n5301_ | ~new_n23351_;
  assign new_n23754_ = ~new_n23633_ | ~new_n23466_;
  assign new_n23755_ = ~new_n23549_ | ~new_n23465_;
  assign new_n23756_ = ~new_n5688_ | ~new_n23348_;
  assign new_n23757_ = ~new_n5302_ | ~new_n23347_;
  assign new_n23758_ = ~new_n23439_;
  assign new_n23759_ = ~new_n23545_ | ~new_n23758_;
  assign new_n23760_ = ~new_n23439_ | ~new_n23467_;
  assign new_n23761_ = ~new_n5685_ | ~new_n23346_;
  assign new_n23762_ = ~new_n5294_ | ~new_n23345_;
  assign new_n23763_ = ~new_n23440_;
  assign new_n23764_ = ~new_n23541_ | ~new_n23763_;
  assign new_n23765_ = ~new_n23440_ | ~new_n23468_;
  assign new_n23766_ = ~new_n5682_ | ~new_n23342_;
  assign new_n23767_ = ~new_n5285_ | ~new_n23341_;
  assign new_n23768_ = ~new_n23767_ | ~new_n23766_;
  assign new_n23769_ = ~new_n5679_ | ~new_n23343_;
  assign new_n23770_ = ~new_n5284_ | ~new_n23340_;
  assign new_n23771_ = ~new_n23643_ | ~new_n23385_;
  assign new_n23772_ = ~new_n23469_ | ~new_n23635_;
  assign new_n23773_ = new_n23969_ & new_n23968_;
  assign new_n23774_ = new_n24008_ & new_n24007_;
  assign new_n23775_ = new_n23948_ & new_n24023_;
  assign new_n23776_ = new_n24025_ & new_n24024_;
  assign new_n23777_ = new_n23949_ & new_n24049_;
  assign new_n23778_ = new_n24051_ & new_n24050_;
  assign new_n23779_ = ~new_n24111_ | ~new_n24114_;
  assign new_n23780_ = ~new_n24100_ | ~new_n24103_;
  assign new_n23781_ = ~new_n24089_ | ~new_n24092_;
  assign new_n23782_ = ~new_n24081_ | ~new_n24083_;
  assign new_n23783_ = ~new_n24119_ | ~new_n24079_;
  assign new_n23784_ = ~new_n24002_ | ~new_n24004_;
  assign new_n23785_ = ~new_n23994_ | ~new_n23997_;
  assign new_n23786_ = ~new_n23986_ | ~new_n23988_;
  assign new_n23787_ = ~new_n23933_ | ~new_n24117_;
  assign new_n23788_ = ~new_n5670_;
  assign new_n23789_ = ~new_n5664_;
  assign new_n23790_ = ~new_n5655_;
  assign new_n23791_ = ~new_n5647_;
  assign new_n23792_ = ~new_n5300_;
  assign new_n23793_ = ~new_n5658_;
  assign new_n23794_ = ~new_n5290_;
  assign new_n23795_ = ~new_n5290_ | ~new_n23790_;
  assign new_n23796_ = ~new_n5286_;
  assign new_n23797_ = ~new_n5667_;
  assign new_n23798_ = ~new_n5661_;
  assign new_n23799_ = ~new_n5293_;
  assign new_n23800_ = ~new_n5289_;
  assign new_n23801_ = ~new_n5282_;
  assign new_n23802_ = ~new_n5282_ | ~new_n23798_;
  assign new_n23803_ = ~new_n5673_;
  assign new_n23804_ = ~new_n5292_;
  assign new_n23805_ = ~new_n5292_ | ~new_n23788_;
  assign new_n23806_ = ~new_n5306_;
  assign new_n23807_ = ~new_n5676_;
  assign new_n23808_ = ~new_n5305_;
  assign new_n23809_ = ~new_n23975_ | ~new_n23974_;
  assign new_n23810_ = ~new_n23802_ | ~new_n23990_;
  assign new_n23811_ = ~new_n24118_ | ~new_n23959_ | ~new_n23943_;
  assign new_n23812_ = ~new_n6171_;
  assign new_n23813_ = ~new_n5679_;
  assign new_n23814_ = ~new_n5682_;
  assign new_n23815_ = ~new_n5285_;
  assign new_n23816_ = ~new_n5284_;
  assign new_n23817_ = ~new_n5305_ | ~new_n23807_;
  assign new_n23818_ = ~new_n5685_;
  assign new_n23819_ = ~new_n5294_;
  assign new_n23820_ = ~new_n5688_;
  assign new_n23821_ = ~new_n5302_;
  assign new_n23822_ = ~new_n5697_;
  assign new_n23823_ = ~new_n5694_;
  assign new_n23824_ = ~new_n5691_;
  assign new_n23825_ = ~new_n5295_;
  assign new_n23826_ = ~new_n5296_;
  assign new_n23827_ = ~new_n5301_;
  assign new_n23828_ = ~new_n5301_ | ~new_n23824_;
  assign new_n23829_ = ~new_n5700_;
  assign new_n23830_ = ~new_n5291_;
  assign new_n23831_ = ~new_n24035_ | ~new_n24034_;
  assign new_n23832_ = ~new_n5304_;
  assign new_n23833_ = ~new_n5705_;
  assign new_n23834_ = ~new_n5303_;
  assign new_n23835_ = ~new_n6177_;
  assign new_n23836_ = ~new_n5298_;
  assign new_n23837_ = ~new_n6174_;
  assign new_n23838_ = ~new_n6175_;
  assign new_n23839_ = ~new_n6176_;
  assign new_n23840_ = ~new_n5288_;
  assign new_n23841_ = ~new_n5283_;
  assign new_n23842_ = ~new_n5297_;
  assign new_n23843_ = ~new_n5297_ | ~new_n23839_;
  assign new_n23844_ = ~new_n6173_;
  assign new_n23845_ = ~new_n5287_;
  assign new_n23846_ = ~new_n6172_;
  assign new_n23847_ = ~new_n5280_;
  assign new_n23848_ = ~new_n6170_;
  assign new_n23849_ = ~new_n5279_;
  assign new_n23850_ = ~new_n5279_ | ~new_n23812_;
  assign new_n23851_ = ~new_n5275_;
  assign new_n23852_ = ~new_n6169_;
  assign new_n23853_ = ~new_n5276_;
  assign new_n23854_ = ~new_n23895_ | ~new_n24068_;
  assign new_n23855_ = ~new_n24065_ | ~new_n24064_;
  assign new_n23856_ = ~new_n23843_ | ~new_n24085_;
  assign new_n23857_ = ~new_n23828_ | ~new_n24096_;
  assign new_n23858_ = ~new_n23817_ | ~new_n24107_;
  assign new_n23859_ = ~new_n5299_;
  assign new_n23860_ = ~new_n24162_ | ~new_n24161_;
  assign new_n23861_ = ~new_n24176_ | ~new_n24175_;
  assign new_n23862_ = ~new_n24181_ | ~new_n24180_;
  assign new_n23863_ = ~new_n24197_ | ~new_n24196_;
  assign new_n23864_ = ~new_n24202_ | ~new_n24201_;
  assign new_n23865_ = ~new_n24207_ | ~new_n24206_;
  assign new_n23866_ = ~new_n24212_ | ~new_n24211_;
  assign new_n23867_ = ~new_n24217_ | ~new_n24216_;
  assign new_n23868_ = ~new_n24233_ | ~new_n24232_;
  assign new_n23869_ = ~new_n24238_ | ~new_n24237_;
  assign new_n23870_ = ~new_n24123_ | ~new_n24122_;
  assign new_n23871_ = ~new_n24132_ | ~new_n24131_;
  assign new_n23872_ = ~new_n24139_ | ~new_n24138_;
  assign new_n23873_ = ~new_n24143_ | ~new_n24142_;
  assign new_n23874_ = ~new_n24152_ | ~new_n24151_;
  assign new_n23875_ = ~new_n24171_ | ~new_n24170_;
  assign new_n23876_ = ~new_n24188_ | ~new_n24187_;
  assign new_n23877_ = ~new_n24192_ | ~new_n24191_;
  assign new_n23878_ = ~new_n24224_ | ~new_n24223_;
  assign new_n23879_ = ~new_n24228_ | ~new_n24227_;
  assign new_n23880_ = ~new_n24245_ | ~new_n24244_;
  assign new_n23881_ = new_n23961_ & new_n23951_;
  assign new_n23882_ = new_n23964_ & new_n23965_;
  assign new_n23883_ = new_n23952_ & new_n23972_ & new_n23967_;
  assign new_n23884_ = new_n23977_ & new_n23953_;
  assign new_n23885_ = new_n23980_ & new_n23981_;
  assign new_n23886_ = new_n23805_ & new_n24125_ & new_n24124_;
  assign new_n23887_ = new_n24128_ & new_n23953_;
  assign new_n23888_ = new_n23996_ & new_n23773_;
  assign new_n23889_ = new_n24135_ & new_n23952_;
  assign new_n23890_ = new_n23795_ & new_n24145_ & new_n24144_;
  assign new_n23891_ = new_n24148_ & new_n23951_;
  assign new_n23892_ = new_n23947_ & new_n24006_ & new_n23983_;
  assign new_n23893_ = new_n24028_ & new_n23775_;
  assign new_n23894_ = new_n24054_ & new_n23777_;
  assign new_n23895_ = new_n24070_ & new_n24071_;
  assign new_n23896_ = new_n24078_ & new_n24154_ & new_n24153_;
  assign new_n23897_ = new_n24075_ & new_n24157_;
  assign new_n23898_ = ~new_n24159_ | ~new_n24158_;
  assign new_n23899_ = new_n23850_ & new_n24164_ & new_n24163_;
  assign new_n23900_ = new_n24167_ & new_n23950_;
  assign new_n23901_ = ~new_n24173_ | ~new_n24172_;
  assign new_n23902_ = ~new_n24178_ | ~new_n24177_;
  assign new_n23903_ = new_n24091_ & new_n23778_;
  assign new_n23904_ = new_n24184_ & new_n23949_;
  assign new_n23905_ = ~new_n24194_ | ~new_n24193_;
  assign new_n23906_ = ~new_n24199_ | ~new_n24198_;
  assign new_n23907_ = ~new_n24204_ | ~new_n24203_;
  assign new_n23908_ = ~new_n24209_ | ~new_n24208_;
  assign new_n23909_ = ~new_n24214_ | ~new_n24213_;
  assign new_n23910_ = new_n24102_ & new_n23776_;
  assign new_n23911_ = new_n24220_ & new_n23948_;
  assign new_n23912_ = ~new_n24230_ | ~new_n24229_;
  assign new_n23913_ = ~new_n24235_ | ~new_n24234_;
  assign new_n23914_ = new_n24113_ & new_n23774_;
  assign new_n23915_ = new_n24241_ & new_n23947_;
  assign new_n23916_ = new_n24121_ & new_n24120_;
  assign new_n23917_ = ~new_n23885_ | ~new_n23978_;
  assign new_n23918_ = new_n24130_ & new_n24129_;
  assign new_n23919_ = new_n24137_ & new_n24136_;
  assign new_n23920_ = new_n24141_ & new_n24140_;
  assign new_n23921_ = ~new_n23882_ | ~new_n23962_;
  assign new_n23922_ = new_n24150_ & new_n24149_;
  assign new_n23923_ = ~new_n6180_;
  assign new_n23924_ = ~new_n5277_;
  assign new_n23925_ = new_n24169_ & new_n24168_;
  assign new_n23926_ = ~new_n24061_ | ~new_n24060_;
  assign new_n23927_ = ~new_n24057_ | ~new_n24056_;
  assign new_n23928_ = new_n24186_ & new_n24185_;
  assign new_n23929_ = new_n24190_ & new_n24189_;
  assign new_n23930_ = ~new_n24047_ | ~new_n24046_;
  assign new_n23931_ = ~new_n24043_ | ~new_n24042_;
  assign new_n23932_ = ~new_n5652_;
  assign new_n23933_ = ~new_n5647_ | ~new_n23859_;
  assign new_n23934_ = ~new_n24039_ | ~new_n24038_;
  assign new_n23935_ = ~new_n5703_;
  assign new_n23936_ = ~new_n24031_ | ~new_n24030_;
  assign new_n23937_ = new_n24222_ & new_n24221_;
  assign new_n23938_ = new_n24226_ & new_n24225_;
  assign new_n23939_ = ~new_n24021_ | ~new_n24020_;
  assign new_n23940_ = ~new_n24017_ | ~new_n24016_;
  assign new_n23941_ = ~new_n24013_ | ~new_n24012_;
  assign new_n23942_ = new_n24243_ & new_n24242_;
  assign new_n23943_ = ~new_n23933_ | ~new_n23932_;
  assign new_n23944_ = ~new_n23850_;
  assign new_n23945_ = ~new_n23795_;
  assign new_n23946_ = ~new_n23805_;
  assign new_n23947_ = ~new_n5679_ | ~new_n23816_;
  assign new_n23948_ = ~new_n5694_ | ~new_n23826_;
  assign new_n23949_ = ~new_n6175_ | ~new_n23841_;
  assign new_n23950_ = ~new_n6171_ | ~new_n23849_;
  assign new_n23951_ = ~new_n5655_ | ~new_n23794_;
  assign new_n23952_ = ~new_n5664_ | ~new_n23800_;
  assign new_n23953_ = ~new_n5670_ | ~new_n23804_;
  assign new_n23954_ = ~new_n23828_;
  assign new_n23955_ = ~new_n23843_;
  assign new_n23956_ = ~new_n23802_;
  assign new_n23957_ = ~new_n23817_;
  assign new_n23958_ = ~new_n23933_;
  assign new_n23959_ = ~new_n5300_ | ~new_n23933_;
  assign new_n23960_ = ~new_n23811_;
  assign new_n23961_ = ~new_n5658_ | ~new_n23796_;
  assign new_n23962_ = ~new_n23881_ | ~new_n23811_;
  assign new_n23963_ = ~new_n23796_ | ~new_n23795_;
  assign new_n23964_ = ~new_n23963_ | ~new_n23793_;
  assign new_n23965_ = ~new_n5286_ | ~new_n23945_;
  assign new_n23966_ = ~new_n23921_;
  assign new_n23967_ = ~new_n5667_ | ~new_n23799_;
  assign new_n23968_ = ~new_n5293_ | ~new_n23797_;
  assign new_n23969_ = ~new_n5289_ | ~new_n23789_;
  assign new_n23970_ = ~new_n23956_ | ~new_n23952_;
  assign new_n23971_ = ~new_n23773_ | ~new_n23970_;
  assign new_n23972_ = ~new_n5661_ | ~new_n23801_;
  assign new_n23973_ = ~new_n5667_ | ~new_n23799_;
  assign new_n23974_ = ~new_n23921_ | ~new_n23883_;
  assign new_n23975_ = ~new_n23973_ | ~new_n23971_;
  assign new_n23976_ = ~new_n23809_;
  assign new_n23977_ = ~new_n5673_ | ~new_n23806_;
  assign new_n23978_ = ~new_n23884_ | ~new_n23809_;
  assign new_n23979_ = ~new_n23806_ | ~new_n23805_;
  assign new_n23980_ = ~new_n23979_ | ~new_n23803_;
  assign new_n23981_ = ~new_n5306_ | ~new_n23946_;
  assign new_n23982_ = ~new_n23917_;
  assign new_n23983_ = ~new_n5676_ | ~new_n23808_;
  assign new_n23984_ = ~new_n23983_ | ~new_n23817_;
  assign new_n23985_ = ~new_n23976_ | ~new_n23805_;
  assign new_n23986_ = ~new_n23887_ | ~new_n23985_;
  assign new_n23987_ = ~new_n23809_ | ~new_n23953_;
  assign new_n23988_ = ~new_n23886_ | ~new_n23987_;
  assign new_n23989_ = ~new_n23805_ | ~new_n23953_;
  assign new_n23990_ = ~new_n23972_ | ~new_n23921_;
  assign new_n23991_ = ~new_n23810_;
  assign new_n23992_ = ~new_n5289_ | ~new_n23789_;
  assign new_n23993_ = ~new_n23991_ | ~new_n23992_;
  assign new_n23994_ = ~new_n23889_ | ~new_n23993_;
  assign new_n23995_ = ~new_n23810_ | ~new_n23952_;
  assign new_n23996_ = ~new_n5667_ | ~new_n23799_;
  assign new_n23997_ = ~new_n23888_ | ~new_n23995_;
  assign new_n23998_ = ~new_n5289_ | ~new_n23789_;
  assign new_n23999_ = ~new_n23952_ | ~new_n23998_;
  assign new_n24000_ = ~new_n23972_ | ~new_n23802_;
  assign new_n24001_ = ~new_n23960_ | ~new_n23795_;
  assign new_n24002_ = ~new_n23891_ | ~new_n24001_;
  assign new_n24003_ = ~new_n23811_ | ~new_n23951_;
  assign new_n24004_ = ~new_n23890_ | ~new_n24003_;
  assign new_n24005_ = ~new_n23795_ | ~new_n23951_;
  assign new_n24006_ = ~new_n5682_ | ~new_n23815_;
  assign new_n24007_ = ~new_n5285_ | ~new_n23814_;
  assign new_n24008_ = ~new_n5284_ | ~new_n23813_;
  assign new_n24009_ = ~new_n23957_ | ~new_n23947_;
  assign new_n24010_ = ~new_n23774_ | ~new_n24009_;
  assign new_n24011_ = ~new_n5682_ | ~new_n23815_;
  assign new_n24012_ = ~new_n23917_ | ~new_n23892_;
  assign new_n24013_ = ~new_n24011_ | ~new_n24010_;
  assign new_n24014_ = ~new_n23941_;
  assign new_n24015_ = ~new_n5685_ | ~new_n23819_;
  assign new_n24016_ = ~new_n24015_ | ~new_n23941_;
  assign new_n24017_ = ~new_n5294_ | ~new_n23818_;
  assign new_n24018_ = ~new_n23940_;
  assign new_n24019_ = ~new_n5688_ | ~new_n23821_;
  assign new_n24020_ = ~new_n24019_ | ~new_n23940_;
  assign new_n24021_ = ~new_n5302_ | ~new_n23820_;
  assign new_n24022_ = ~new_n23939_;
  assign new_n24023_ = ~new_n5697_ | ~new_n23825_;
  assign new_n24024_ = ~new_n5295_ | ~new_n23822_;
  assign new_n24025_ = ~new_n5296_ | ~new_n23823_;
  assign new_n24026_ = ~new_n23954_ | ~new_n23775_;
  assign new_n24027_ = ~new_n23776_ | ~new_n24026_;
  assign new_n24028_ = ~new_n5691_ | ~new_n23827_;
  assign new_n24029_ = ~new_n5697_ | ~new_n23825_;
  assign new_n24030_ = ~new_n23893_ | ~new_n23939_;
  assign new_n24031_ = ~new_n24029_ | ~new_n24027_;
  assign new_n24032_ = ~new_n23936_;
  assign new_n24033_ = ~new_n5700_ | ~new_n23830_;
  assign new_n24034_ = ~new_n24033_ | ~new_n23936_;
  assign new_n24035_ = ~new_n5291_ | ~new_n23829_;
  assign new_n24036_ = ~new_n23831_;
  assign new_n24037_ = ~new_n24036_ | ~new_n23832_;
  assign new_n24038_ = ~new_n24037_ | ~new_n23935_;
  assign new_n24039_ = ~new_n5304_ | ~new_n23831_;
  assign new_n24040_ = ~new_n23934_;
  assign new_n24041_ = ~new_n5705_ | ~new_n23834_;
  assign new_n24042_ = ~new_n24041_ | ~new_n23934_;
  assign new_n24043_ = ~new_n5303_ | ~new_n23833_;
  assign new_n24044_ = ~new_n23931_;
  assign new_n24045_ = ~new_n6177_ | ~new_n23836_;
  assign new_n24046_ = ~new_n24045_ | ~new_n23931_;
  assign new_n24047_ = ~new_n5298_ | ~new_n23835_;
  assign new_n24048_ = ~new_n23930_;
  assign new_n24049_ = ~new_n6174_ | ~new_n23840_;
  assign new_n24050_ = ~new_n5288_ | ~new_n23837_;
  assign new_n24051_ = ~new_n5283_ | ~new_n23838_;
  assign new_n24052_ = ~new_n23955_ | ~new_n23777_;
  assign new_n24053_ = ~new_n23778_ | ~new_n24052_;
  assign new_n24054_ = ~new_n6176_ | ~new_n23842_;
  assign new_n24055_ = ~new_n6174_ | ~new_n23840_;
  assign new_n24056_ = ~new_n23894_ | ~new_n23930_;
  assign new_n24057_ = ~new_n24055_ | ~new_n24053_;
  assign new_n24058_ = ~new_n23927_;
  assign new_n24059_ = ~new_n6173_ | ~new_n23845_;
  assign new_n24060_ = ~new_n24059_ | ~new_n23927_;
  assign new_n24061_ = ~new_n5287_ | ~new_n23844_;
  assign new_n24062_ = ~new_n23926_;
  assign new_n24063_ = ~new_n6172_ | ~new_n23847_;
  assign new_n24064_ = ~new_n24063_ | ~new_n23926_;
  assign new_n24065_ = ~new_n5280_ | ~new_n23846_;
  assign new_n24066_ = ~new_n23855_;
  assign new_n24067_ = ~new_n6170_ | ~new_n23851_;
  assign new_n24068_ = ~new_n24067_ | ~new_n23855_ | ~new_n23950_;
  assign new_n24069_ = ~new_n23851_ | ~new_n23850_;
  assign new_n24070_ = ~new_n24069_ | ~new_n23848_;
  assign new_n24071_ = ~new_n5275_ | ~new_n23944_;
  assign new_n24072_ = ~new_n23854_;
  assign new_n24073_ = ~new_n5276_ | ~new_n23852_;
  assign new_n24074_ = ~new_n24072_ | ~new_n24073_;
  assign new_n24075_ = ~new_n6169_ | ~new_n23853_;
  assign new_n24076_ = ~new_n6169_ | ~new_n23853_;
  assign new_n24077_ = ~new_n24076_ | ~new_n23854_;
  assign new_n24078_ = ~new_n5276_ | ~new_n23852_;
  assign new_n24079_ = ~new_n23896_ | ~new_n24077_;
  assign new_n24080_ = ~new_n24066_ | ~new_n23850_;
  assign new_n24081_ = ~new_n23900_ | ~new_n24080_;
  assign new_n24082_ = ~new_n23855_ | ~new_n23950_;
  assign new_n24083_ = ~new_n23899_ | ~new_n24082_;
  assign new_n24084_ = ~new_n23850_ | ~new_n23950_;
  assign new_n24085_ = ~new_n24054_ | ~new_n23930_;
  assign new_n24086_ = ~new_n23856_;
  assign new_n24087_ = ~new_n5283_ | ~new_n23838_;
  assign new_n24088_ = ~new_n24086_ | ~new_n24087_;
  assign new_n24089_ = ~new_n23904_ | ~new_n24088_;
  assign new_n24090_ = ~new_n23856_ | ~new_n23949_;
  assign new_n24091_ = ~new_n6174_ | ~new_n23840_;
  assign new_n24092_ = ~new_n23903_ | ~new_n24090_;
  assign new_n24093_ = ~new_n5283_ | ~new_n23838_;
  assign new_n24094_ = ~new_n23949_ | ~new_n24093_;
  assign new_n24095_ = ~new_n24054_ | ~new_n23843_;
  assign new_n24096_ = ~new_n24028_ | ~new_n23939_;
  assign new_n24097_ = ~new_n23857_;
  assign new_n24098_ = ~new_n5296_ | ~new_n23823_;
  assign new_n24099_ = ~new_n24097_ | ~new_n24098_;
  assign new_n24100_ = ~new_n23911_ | ~new_n24099_;
  assign new_n24101_ = ~new_n23857_ | ~new_n23948_;
  assign new_n24102_ = ~new_n5697_ | ~new_n23825_;
  assign new_n24103_ = ~new_n23910_ | ~new_n24101_;
  assign new_n24104_ = ~new_n5296_ | ~new_n23823_;
  assign new_n24105_ = ~new_n23948_ | ~new_n24104_;
  assign new_n24106_ = ~new_n24028_ | ~new_n23828_;
  assign new_n24107_ = ~new_n23983_ | ~new_n23917_;
  assign new_n24108_ = ~new_n23858_;
  assign new_n24109_ = ~new_n5284_ | ~new_n23813_;
  assign new_n24110_ = ~new_n24108_ | ~new_n24109_;
  assign new_n24111_ = ~new_n23915_ | ~new_n24110_;
  assign new_n24112_ = ~new_n23858_ | ~new_n23947_;
  assign new_n24113_ = ~new_n5682_ | ~new_n23815_;
  assign new_n24114_ = ~new_n23914_ | ~new_n24112_;
  assign new_n24115_ = ~new_n5284_ | ~new_n23813_;
  assign new_n24116_ = ~new_n23947_ | ~new_n24115_;
  assign new_n24117_ = ~new_n5299_ | ~new_n23791_;
  assign new_n24118_ = ~new_n5300_ | ~new_n23932_;
  assign new_n24119_ = ~new_n23897_ | ~new_n24074_;
  assign new_n24120_ = ~new_n5676_ | ~new_n23808_;
  assign new_n24121_ = ~new_n5305_ | ~new_n23807_;
  assign new_n24122_ = ~new_n23984_ | ~new_n23917_;
  assign new_n24123_ = ~new_n23982_ | ~new_n23916_;
  assign new_n24124_ = ~new_n5673_ | ~new_n23806_;
  assign new_n24125_ = ~new_n5306_ | ~new_n23803_;
  assign new_n24126_ = ~new_n5673_ | ~new_n23806_;
  assign new_n24127_ = ~new_n5306_ | ~new_n23803_;
  assign new_n24128_ = ~new_n24127_ | ~new_n24126_;
  assign new_n24129_ = ~new_n5670_ | ~new_n23804_;
  assign new_n24130_ = ~new_n5292_ | ~new_n23788_;
  assign new_n24131_ = ~new_n23989_ | ~new_n23809_;
  assign new_n24132_ = ~new_n23918_ | ~new_n23976_;
  assign new_n24133_ = ~new_n5667_ | ~new_n23799_;
  assign new_n24134_ = ~new_n5293_ | ~new_n23797_;
  assign new_n24135_ = ~new_n24134_ | ~new_n24133_;
  assign new_n24136_ = ~new_n5664_ | ~new_n23800_;
  assign new_n24137_ = ~new_n5289_ | ~new_n23789_;
  assign new_n24138_ = ~new_n23999_ | ~new_n23810_;
  assign new_n24139_ = ~new_n23919_ | ~new_n23991_;
  assign new_n24140_ = ~new_n5661_ | ~new_n23801_;
  assign new_n24141_ = ~new_n5282_ | ~new_n23798_;
  assign new_n24142_ = ~new_n24000_ | ~new_n23921_;
  assign new_n24143_ = ~new_n23966_ | ~new_n23920_;
  assign new_n24144_ = ~new_n5658_ | ~new_n23796_;
  assign new_n24145_ = ~new_n5286_ | ~new_n23793_;
  assign new_n24146_ = ~new_n5658_ | ~new_n23796_;
  assign new_n24147_ = ~new_n5286_ | ~new_n23793_;
  assign new_n24148_ = ~new_n24147_ | ~new_n24146_;
  assign new_n24149_ = ~new_n5655_ | ~new_n23794_;
  assign new_n24150_ = ~new_n5290_ | ~new_n23790_;
  assign new_n24151_ = ~new_n24005_ | ~new_n23811_;
  assign new_n24152_ = ~new_n23922_ | ~new_n23960_;
  assign new_n24153_ = ~new_n6180_ | ~new_n23924_;
  assign new_n24154_ = ~new_n5277_ | ~new_n23923_;
  assign new_n24155_ = ~new_n6180_ | ~new_n23924_;
  assign new_n24156_ = ~new_n5277_ | ~new_n23923_;
  assign new_n24157_ = ~new_n24156_ | ~new_n24155_;
  assign new_n24158_ = ~new_n6169_ | ~new_n23853_;
  assign new_n24159_ = ~new_n5276_ | ~new_n23852_;
  assign new_n24160_ = ~new_n23898_;
  assign new_n24161_ = ~new_n24160_ | ~new_n24072_;
  assign new_n24162_ = ~new_n23898_ | ~new_n23854_;
  assign new_n24163_ = ~new_n6170_ | ~new_n23851_;
  assign new_n24164_ = ~new_n5275_ | ~new_n23848_;
  assign new_n24165_ = ~new_n6170_ | ~new_n23851_;
  assign new_n24166_ = ~new_n5275_ | ~new_n23848_;
  assign new_n24167_ = ~new_n24166_ | ~new_n24165_;
  assign new_n24168_ = ~new_n6171_ | ~new_n23849_;
  assign new_n24169_ = ~new_n5279_ | ~new_n23812_;
  assign new_n24170_ = ~new_n24084_ | ~new_n23855_;
  assign new_n24171_ = ~new_n23925_ | ~new_n24066_;
  assign new_n24172_ = ~new_n6172_ | ~new_n23847_;
  assign new_n24173_ = ~new_n5280_ | ~new_n23846_;
  assign new_n24174_ = ~new_n23901_;
  assign new_n24175_ = ~new_n24062_ | ~new_n24174_;
  assign new_n24176_ = ~new_n23901_ | ~new_n23926_;
  assign new_n24177_ = ~new_n6173_ | ~new_n23845_;
  assign new_n24178_ = ~new_n5287_ | ~new_n23844_;
  assign new_n24179_ = ~new_n23902_;
  assign new_n24180_ = ~new_n24058_ | ~new_n24179_;
  assign new_n24181_ = ~new_n23902_ | ~new_n23927_;
  assign new_n24182_ = ~new_n6174_ | ~new_n23840_;
  assign new_n24183_ = ~new_n5288_ | ~new_n23837_;
  assign new_n24184_ = ~new_n24183_ | ~new_n24182_;
  assign new_n24185_ = ~new_n6175_ | ~new_n23841_;
  assign new_n24186_ = ~new_n5283_ | ~new_n23838_;
  assign new_n24187_ = ~new_n24094_ | ~new_n23856_;
  assign new_n24188_ = ~new_n23928_ | ~new_n24086_;
  assign new_n24189_ = ~new_n6176_ | ~new_n23842_;
  assign new_n24190_ = ~new_n5297_ | ~new_n23839_;
  assign new_n24191_ = ~new_n24095_ | ~new_n23930_;
  assign new_n24192_ = ~new_n24048_ | ~new_n23929_;
  assign new_n24193_ = ~new_n6177_ | ~new_n23836_;
  assign new_n24194_ = ~new_n5298_ | ~new_n23835_;
  assign new_n24195_ = ~new_n23905_;
  assign new_n24196_ = ~new_n24044_ | ~new_n24195_;
  assign new_n24197_ = ~new_n23905_ | ~new_n23931_;
  assign new_n24198_ = ~new_n5652_ | ~new_n23792_;
  assign new_n24199_ = ~new_n5300_ | ~new_n23932_;
  assign new_n24200_ = ~new_n23906_;
  assign new_n24201_ = ~new_n23958_ | ~new_n24200_;
  assign new_n24202_ = ~new_n23906_ | ~new_n23933_;
  assign new_n24203_ = ~new_n5705_ | ~new_n23834_;
  assign new_n24204_ = ~new_n5303_ | ~new_n23833_;
  assign new_n24205_ = ~new_n23907_;
  assign new_n24206_ = ~new_n24040_ | ~new_n24205_;
  assign new_n24207_ = ~new_n23907_ | ~new_n23934_;
  assign new_n24208_ = ~new_n5703_ | ~new_n23832_;
  assign new_n24209_ = ~new_n5304_ | ~new_n23935_;
  assign new_n24210_ = ~new_n23908_;
  assign new_n24211_ = ~new_n24210_ | ~new_n24036_;
  assign new_n24212_ = ~new_n23908_ | ~new_n23831_;
  assign new_n24213_ = ~new_n5700_ | ~new_n23830_;
  assign new_n24214_ = ~new_n5291_ | ~new_n23829_;
  assign new_n24215_ = ~new_n23909_;
  assign new_n24216_ = ~new_n24032_ | ~new_n24215_;
  assign new_n24217_ = ~new_n23909_ | ~new_n23936_;
  assign new_n24218_ = ~new_n5697_ | ~new_n23825_;
  assign new_n24219_ = ~new_n5295_ | ~new_n23822_;
  assign new_n24220_ = ~new_n24219_ | ~new_n24218_;
  assign new_n24221_ = ~new_n5694_ | ~new_n23826_;
  assign new_n24222_ = ~new_n5296_ | ~new_n23823_;
  assign new_n24223_ = ~new_n24105_ | ~new_n23857_;
  assign new_n24224_ = ~new_n23937_ | ~new_n24097_;
  assign new_n24225_ = ~new_n5691_ | ~new_n23827_;
  assign new_n24226_ = ~new_n5301_ | ~new_n23824_;
  assign new_n24227_ = ~new_n24106_ | ~new_n23939_;
  assign new_n24228_ = ~new_n24022_ | ~new_n23938_;
  assign new_n24229_ = ~new_n5688_ | ~new_n23821_;
  assign new_n24230_ = ~new_n5302_ | ~new_n23820_;
  assign new_n24231_ = ~new_n23912_;
  assign new_n24232_ = ~new_n24018_ | ~new_n24231_;
  assign new_n24233_ = ~new_n23912_ | ~new_n23940_;
  assign new_n24234_ = ~new_n5685_ | ~new_n23819_;
  assign new_n24235_ = ~new_n5294_ | ~new_n23818_;
  assign new_n24236_ = ~new_n23913_;
  assign new_n24237_ = ~new_n24014_ | ~new_n24236_;
  assign new_n24238_ = ~new_n23913_ | ~new_n23941_;
  assign new_n24239_ = ~new_n5682_ | ~new_n23815_;
  assign new_n24240_ = ~new_n5285_ | ~new_n23814_;
  assign new_n24241_ = ~new_n24240_ | ~new_n24239_;
  assign new_n24242_ = ~new_n5679_ | ~new_n23816_;
  assign new_n24243_ = ~new_n5284_ | ~new_n23813_;
  assign new_n24244_ = ~new_n24116_ | ~new_n23858_;
  assign new_n24245_ = ~new_n23942_ | ~new_n24108_;
  assign new_n24246_ = new_n24442_ & new_n24441_;
  assign new_n24247_ = new_n24481_ & new_n24480_;
  assign new_n24248_ = new_n24421_ & new_n24496_;
  assign new_n24249_ = new_n24498_ & new_n24497_;
  assign new_n24250_ = new_n24422_ & new_n24522_;
  assign new_n24251_ = new_n24524_ & new_n24523_;
  assign new_n24252_ = ~new_n24584_ | ~new_n24587_;
  assign new_n24253_ = ~new_n24573_ | ~new_n24576_;
  assign new_n24254_ = ~new_n24562_ | ~new_n24565_;
  assign new_n24255_ = ~new_n24554_ | ~new_n24556_;
  assign new_n24256_ = ~new_n24592_ | ~new_n24552_;
  assign new_n24257_ = ~new_n24475_ | ~new_n24477_;
  assign new_n24258_ = ~new_n24467_ | ~new_n24470_;
  assign new_n24259_ = ~new_n24459_ | ~new_n24461_;
  assign new_n24260_ = ~new_n24406_ | ~new_n24590_;
  assign new_n24261_ = ~new_n5670_;
  assign new_n24262_ = ~new_n5664_;
  assign new_n24263_ = ~new_n5655_;
  assign new_n24264_ = ~new_n5647_;
  assign new_n24265_ = ~new_n5300_;
  assign new_n24266_ = ~new_n5658_;
  assign new_n24267_ = ~new_n5290_;
  assign new_n24268_ = ~new_n5290_ | ~new_n24263_;
  assign new_n24269_ = ~new_n5286_;
  assign new_n24270_ = ~new_n5667_;
  assign new_n24271_ = ~new_n5661_;
  assign new_n24272_ = ~new_n5293_;
  assign new_n24273_ = ~new_n5289_;
  assign new_n24274_ = ~new_n5282_;
  assign new_n24275_ = ~new_n5282_ | ~new_n24271_;
  assign new_n24276_ = ~new_n5673_;
  assign new_n24277_ = ~new_n5292_;
  assign new_n24278_ = ~new_n5292_ | ~new_n24261_;
  assign new_n24279_ = ~new_n5306_;
  assign new_n24280_ = ~new_n5676_;
  assign new_n24281_ = ~new_n5305_;
  assign new_n24282_ = ~new_n24448_ | ~new_n24447_;
  assign new_n24283_ = ~new_n24275_ | ~new_n24463_;
  assign new_n24284_ = ~new_n24591_ | ~new_n24432_ | ~new_n24416_;
  assign new_n24285_ = ~new_n6171_;
  assign new_n24286_ = ~new_n5679_;
  assign new_n24287_ = ~new_n5682_;
  assign new_n24288_ = ~new_n5285_;
  assign new_n24289_ = ~new_n5284_;
  assign new_n24290_ = ~new_n5305_ | ~new_n24280_;
  assign new_n24291_ = ~new_n5685_;
  assign new_n24292_ = ~new_n5294_;
  assign new_n24293_ = ~new_n5688_;
  assign new_n24294_ = ~new_n5302_;
  assign new_n24295_ = ~new_n5697_;
  assign new_n24296_ = ~new_n5694_;
  assign new_n24297_ = ~new_n5691_;
  assign new_n24298_ = ~new_n5295_;
  assign new_n24299_ = ~new_n5296_;
  assign new_n24300_ = ~new_n5301_;
  assign new_n24301_ = ~new_n5301_ | ~new_n24297_;
  assign new_n24302_ = ~new_n5700_;
  assign new_n24303_ = ~new_n5291_;
  assign new_n24304_ = ~new_n24508_ | ~new_n24507_;
  assign new_n24305_ = ~new_n5304_;
  assign new_n24306_ = ~new_n5705_;
  assign new_n24307_ = ~new_n5303_;
  assign new_n24308_ = ~new_n6177_;
  assign new_n24309_ = ~new_n5298_;
  assign new_n24310_ = ~new_n6174_;
  assign new_n24311_ = ~new_n6175_;
  assign new_n24312_ = ~new_n6176_;
  assign new_n24313_ = ~new_n5288_;
  assign new_n24314_ = ~new_n5283_;
  assign new_n24315_ = ~new_n5297_;
  assign new_n24316_ = ~new_n5297_ | ~new_n24312_;
  assign new_n24317_ = ~new_n6173_;
  assign new_n24318_ = ~new_n5287_;
  assign new_n24319_ = ~new_n6172_;
  assign new_n24320_ = ~new_n5280_;
  assign new_n24321_ = ~new_n6170_;
  assign new_n24322_ = ~new_n5279_;
  assign new_n24323_ = ~new_n5279_ | ~new_n24285_;
  assign new_n24324_ = ~new_n5275_;
  assign new_n24325_ = ~new_n6169_;
  assign new_n24326_ = ~new_n5276_;
  assign new_n24327_ = ~new_n24368_ | ~new_n24541_;
  assign new_n24328_ = ~new_n24538_ | ~new_n24537_;
  assign new_n24329_ = ~new_n24316_ | ~new_n24558_;
  assign new_n24330_ = ~new_n24301_ | ~new_n24569_;
  assign new_n24331_ = ~new_n24290_ | ~new_n24580_;
  assign new_n24332_ = ~new_n5299_;
  assign new_n24333_ = ~new_n24635_ | ~new_n24634_;
  assign new_n24334_ = ~new_n24649_ | ~new_n24648_;
  assign new_n24335_ = ~new_n24654_ | ~new_n24653_;
  assign new_n24336_ = ~new_n24670_ | ~new_n24669_;
  assign new_n24337_ = ~new_n24675_ | ~new_n24674_;
  assign new_n24338_ = ~new_n24680_ | ~new_n24679_;
  assign new_n24339_ = ~new_n24685_ | ~new_n24684_;
  assign new_n24340_ = ~new_n24690_ | ~new_n24689_;
  assign new_n24341_ = ~new_n24706_ | ~new_n24705_;
  assign new_n24342_ = ~new_n24711_ | ~new_n24710_;
  assign new_n24343_ = ~new_n24596_ | ~new_n24595_;
  assign new_n24344_ = ~new_n24605_ | ~new_n24604_;
  assign new_n24345_ = ~new_n24612_ | ~new_n24611_;
  assign new_n24346_ = ~new_n24616_ | ~new_n24615_;
  assign new_n24347_ = ~new_n24625_ | ~new_n24624_;
  assign new_n24348_ = ~new_n24644_ | ~new_n24643_;
  assign new_n24349_ = ~new_n24661_ | ~new_n24660_;
  assign new_n24350_ = ~new_n24665_ | ~new_n24664_;
  assign new_n24351_ = ~new_n24697_ | ~new_n24696_;
  assign new_n24352_ = ~new_n24701_ | ~new_n24700_;
  assign new_n24353_ = ~new_n24718_ | ~new_n24717_;
  assign new_n24354_ = new_n24434_ & new_n24424_;
  assign new_n24355_ = new_n24437_ & new_n24438_;
  assign new_n24356_ = new_n24425_ & new_n24445_ & new_n24440_;
  assign new_n24357_ = new_n24450_ & new_n24426_;
  assign new_n24358_ = new_n24453_ & new_n24454_;
  assign new_n24359_ = new_n24278_ & new_n24598_ & new_n24597_;
  assign new_n24360_ = new_n24601_ & new_n24426_;
  assign new_n24361_ = new_n24469_ & new_n24246_;
  assign new_n24362_ = new_n24608_ & new_n24425_;
  assign new_n24363_ = new_n24268_ & new_n24618_ & new_n24617_;
  assign new_n24364_ = new_n24621_ & new_n24424_;
  assign new_n24365_ = new_n24420_ & new_n24479_ & new_n24456_;
  assign new_n24366_ = new_n24501_ & new_n24248_;
  assign new_n24367_ = new_n24527_ & new_n24250_;
  assign new_n24368_ = new_n24543_ & new_n24544_;
  assign new_n24369_ = new_n24551_ & new_n24627_ & new_n24626_;
  assign new_n24370_ = new_n24548_ & new_n24630_;
  assign new_n24371_ = ~new_n24632_ | ~new_n24631_;
  assign new_n24372_ = new_n24323_ & new_n24637_ & new_n24636_;
  assign new_n24373_ = new_n24640_ & new_n24423_;
  assign new_n24374_ = ~new_n24646_ | ~new_n24645_;
  assign new_n24375_ = ~new_n24651_ | ~new_n24650_;
  assign new_n24376_ = new_n24564_ & new_n24251_;
  assign new_n24377_ = new_n24657_ & new_n24422_;
  assign new_n24378_ = ~new_n24667_ | ~new_n24666_;
  assign new_n24379_ = ~new_n24672_ | ~new_n24671_;
  assign new_n24380_ = ~new_n24677_ | ~new_n24676_;
  assign new_n24381_ = ~new_n24682_ | ~new_n24681_;
  assign new_n24382_ = ~new_n24687_ | ~new_n24686_;
  assign new_n24383_ = new_n24575_ & new_n24249_;
  assign new_n24384_ = new_n24693_ & new_n24421_;
  assign new_n24385_ = ~new_n24703_ | ~new_n24702_;
  assign new_n24386_ = ~new_n24708_ | ~new_n24707_;
  assign new_n24387_ = new_n24586_ & new_n24247_;
  assign new_n24388_ = new_n24714_ & new_n24420_;
  assign new_n24389_ = new_n24594_ & new_n24593_;
  assign new_n24390_ = ~new_n24358_ | ~new_n24451_;
  assign new_n24391_ = new_n24603_ & new_n24602_;
  assign new_n24392_ = new_n24610_ & new_n24609_;
  assign new_n24393_ = new_n24614_ & new_n24613_;
  assign new_n24394_ = ~new_n24355_ | ~new_n24435_;
  assign new_n24395_ = new_n24623_ & new_n24622_;
  assign new_n24396_ = ~new_n6180_;
  assign new_n24397_ = ~new_n5277_;
  assign new_n24398_ = new_n24642_ & new_n24641_;
  assign new_n24399_ = ~new_n24534_ | ~new_n24533_;
  assign new_n24400_ = ~new_n24530_ | ~new_n24529_;
  assign new_n24401_ = new_n24659_ & new_n24658_;
  assign new_n24402_ = new_n24663_ & new_n24662_;
  assign new_n24403_ = ~new_n24520_ | ~new_n24519_;
  assign new_n24404_ = ~new_n24516_ | ~new_n24515_;
  assign new_n24405_ = ~new_n5652_;
  assign new_n24406_ = ~new_n5647_ | ~new_n24332_;
  assign new_n24407_ = ~new_n24512_ | ~new_n24511_;
  assign new_n24408_ = ~new_n5703_;
  assign new_n24409_ = ~new_n24504_ | ~new_n24503_;
  assign new_n24410_ = new_n24695_ & new_n24694_;
  assign new_n24411_ = new_n24699_ & new_n24698_;
  assign new_n24412_ = ~new_n24494_ | ~new_n24493_;
  assign new_n24413_ = ~new_n24490_ | ~new_n24489_;
  assign new_n24414_ = ~new_n24486_ | ~new_n24485_;
  assign new_n24415_ = new_n24716_ & new_n24715_;
  assign new_n24416_ = ~new_n24406_ | ~new_n24405_;
  assign new_n24417_ = ~new_n24323_;
  assign new_n24418_ = ~new_n24268_;
  assign new_n24419_ = ~new_n24278_;
  assign new_n24420_ = ~new_n5679_ | ~new_n24289_;
  assign new_n24421_ = ~new_n5694_ | ~new_n24299_;
  assign new_n24422_ = ~new_n6175_ | ~new_n24314_;
  assign new_n24423_ = ~new_n6171_ | ~new_n24322_;
  assign new_n24424_ = ~new_n5655_ | ~new_n24267_;
  assign new_n24425_ = ~new_n5664_ | ~new_n24273_;
  assign new_n24426_ = ~new_n5670_ | ~new_n24277_;
  assign new_n24427_ = ~new_n24301_;
  assign new_n24428_ = ~new_n24316_;
  assign new_n24429_ = ~new_n24275_;
  assign new_n24430_ = ~new_n24290_;
  assign new_n24431_ = ~new_n24406_;
  assign new_n24432_ = ~new_n5300_ | ~new_n24406_;
  assign new_n24433_ = ~new_n24284_;
  assign new_n24434_ = ~new_n5658_ | ~new_n24269_;
  assign new_n24435_ = ~new_n24354_ | ~new_n24284_;
  assign new_n24436_ = ~new_n24269_ | ~new_n24268_;
  assign new_n24437_ = ~new_n24436_ | ~new_n24266_;
  assign new_n24438_ = ~new_n5286_ | ~new_n24418_;
  assign new_n24439_ = ~new_n24394_;
  assign new_n24440_ = ~new_n5667_ | ~new_n24272_;
  assign new_n24441_ = ~new_n5293_ | ~new_n24270_;
  assign new_n24442_ = ~new_n5289_ | ~new_n24262_;
  assign new_n24443_ = ~new_n24429_ | ~new_n24425_;
  assign new_n24444_ = ~new_n24246_ | ~new_n24443_;
  assign new_n24445_ = ~new_n5661_ | ~new_n24274_;
  assign new_n24446_ = ~new_n5667_ | ~new_n24272_;
  assign new_n24447_ = ~new_n24394_ | ~new_n24356_;
  assign new_n24448_ = ~new_n24446_ | ~new_n24444_;
  assign new_n24449_ = ~new_n24282_;
  assign new_n24450_ = ~new_n5673_ | ~new_n24279_;
  assign new_n24451_ = ~new_n24357_ | ~new_n24282_;
  assign new_n24452_ = ~new_n24279_ | ~new_n24278_;
  assign new_n24453_ = ~new_n24452_ | ~new_n24276_;
  assign new_n24454_ = ~new_n5306_ | ~new_n24419_;
  assign new_n24455_ = ~new_n24390_;
  assign new_n24456_ = ~new_n5676_ | ~new_n24281_;
  assign new_n24457_ = ~new_n24456_ | ~new_n24290_;
  assign new_n24458_ = ~new_n24449_ | ~new_n24278_;
  assign new_n24459_ = ~new_n24360_ | ~new_n24458_;
  assign new_n24460_ = ~new_n24282_ | ~new_n24426_;
  assign new_n24461_ = ~new_n24359_ | ~new_n24460_;
  assign new_n24462_ = ~new_n24278_ | ~new_n24426_;
  assign new_n24463_ = ~new_n24445_ | ~new_n24394_;
  assign new_n24464_ = ~new_n24283_;
  assign new_n24465_ = ~new_n5289_ | ~new_n24262_;
  assign new_n24466_ = ~new_n24464_ | ~new_n24465_;
  assign new_n24467_ = ~new_n24362_ | ~new_n24466_;
  assign new_n24468_ = ~new_n24283_ | ~new_n24425_;
  assign new_n24469_ = ~new_n5667_ | ~new_n24272_;
  assign new_n24470_ = ~new_n24361_ | ~new_n24468_;
  assign new_n24471_ = ~new_n5289_ | ~new_n24262_;
  assign new_n24472_ = ~new_n24425_ | ~new_n24471_;
  assign new_n24473_ = ~new_n24445_ | ~new_n24275_;
  assign new_n24474_ = ~new_n24433_ | ~new_n24268_;
  assign new_n24475_ = ~new_n24364_ | ~new_n24474_;
  assign new_n24476_ = ~new_n24284_ | ~new_n24424_;
  assign new_n24477_ = ~new_n24363_ | ~new_n24476_;
  assign new_n24478_ = ~new_n24268_ | ~new_n24424_;
  assign new_n24479_ = ~new_n5682_ | ~new_n24288_;
  assign new_n24480_ = ~new_n5285_ | ~new_n24287_;
  assign new_n24481_ = ~new_n5284_ | ~new_n24286_;
  assign new_n24482_ = ~new_n24430_ | ~new_n24420_;
  assign new_n24483_ = ~new_n24247_ | ~new_n24482_;
  assign new_n24484_ = ~new_n5682_ | ~new_n24288_;
  assign new_n24485_ = ~new_n24390_ | ~new_n24365_;
  assign new_n24486_ = ~new_n24484_ | ~new_n24483_;
  assign new_n24487_ = ~new_n24414_;
  assign new_n24488_ = ~new_n5685_ | ~new_n24292_;
  assign new_n24489_ = ~new_n24488_ | ~new_n24414_;
  assign new_n24490_ = ~new_n5294_ | ~new_n24291_;
  assign new_n24491_ = ~new_n24413_;
  assign new_n24492_ = ~new_n5688_ | ~new_n24294_;
  assign new_n24493_ = ~new_n24492_ | ~new_n24413_;
  assign new_n24494_ = ~new_n5302_ | ~new_n24293_;
  assign new_n24495_ = ~new_n24412_;
  assign new_n24496_ = ~new_n5697_ | ~new_n24298_;
  assign new_n24497_ = ~new_n5295_ | ~new_n24295_;
  assign new_n24498_ = ~new_n5296_ | ~new_n24296_;
  assign new_n24499_ = ~new_n24427_ | ~new_n24248_;
  assign new_n24500_ = ~new_n24249_ | ~new_n24499_;
  assign new_n24501_ = ~new_n5691_ | ~new_n24300_;
  assign new_n24502_ = ~new_n5697_ | ~new_n24298_;
  assign new_n24503_ = ~new_n24366_ | ~new_n24412_;
  assign new_n24504_ = ~new_n24502_ | ~new_n24500_;
  assign new_n24505_ = ~new_n24409_;
  assign new_n24506_ = ~new_n5700_ | ~new_n24303_;
  assign new_n24507_ = ~new_n24506_ | ~new_n24409_;
  assign new_n24508_ = ~new_n5291_ | ~new_n24302_;
  assign new_n24509_ = ~new_n24304_;
  assign new_n24510_ = ~new_n24509_ | ~new_n24305_;
  assign new_n24511_ = ~new_n24510_ | ~new_n24408_;
  assign new_n24512_ = ~new_n5304_ | ~new_n24304_;
  assign new_n24513_ = ~new_n24407_;
  assign new_n24514_ = ~new_n5705_ | ~new_n24307_;
  assign new_n24515_ = ~new_n24514_ | ~new_n24407_;
  assign new_n24516_ = ~new_n5303_ | ~new_n24306_;
  assign new_n24517_ = ~new_n24404_;
  assign new_n24518_ = ~new_n6177_ | ~new_n24309_;
  assign new_n24519_ = ~new_n24518_ | ~new_n24404_;
  assign new_n24520_ = ~new_n5298_ | ~new_n24308_;
  assign new_n24521_ = ~new_n24403_;
  assign new_n24522_ = ~new_n6174_ | ~new_n24313_;
  assign new_n24523_ = ~new_n5288_ | ~new_n24310_;
  assign new_n24524_ = ~new_n5283_ | ~new_n24311_;
  assign new_n24525_ = ~new_n24428_ | ~new_n24250_;
  assign new_n24526_ = ~new_n24251_ | ~new_n24525_;
  assign new_n24527_ = ~new_n6176_ | ~new_n24315_;
  assign new_n24528_ = ~new_n6174_ | ~new_n24313_;
  assign new_n24529_ = ~new_n24367_ | ~new_n24403_;
  assign new_n24530_ = ~new_n24528_ | ~new_n24526_;
  assign new_n24531_ = ~new_n24400_;
  assign new_n24532_ = ~new_n6173_ | ~new_n24318_;
  assign new_n24533_ = ~new_n24532_ | ~new_n24400_;
  assign new_n24534_ = ~new_n5287_ | ~new_n24317_;
  assign new_n24535_ = ~new_n24399_;
  assign new_n24536_ = ~new_n6172_ | ~new_n24320_;
  assign new_n24537_ = ~new_n24536_ | ~new_n24399_;
  assign new_n24538_ = ~new_n5280_ | ~new_n24319_;
  assign new_n24539_ = ~new_n24328_;
  assign new_n24540_ = ~new_n6170_ | ~new_n24324_;
  assign new_n24541_ = ~new_n24540_ | ~new_n24328_ | ~new_n24423_;
  assign new_n24542_ = ~new_n24324_ | ~new_n24323_;
  assign new_n24543_ = ~new_n24542_ | ~new_n24321_;
  assign new_n24544_ = ~new_n5275_ | ~new_n24417_;
  assign new_n24545_ = ~new_n24327_;
  assign new_n24546_ = ~new_n5276_ | ~new_n24325_;
  assign new_n24547_ = ~new_n24545_ | ~new_n24546_;
  assign new_n24548_ = ~new_n6169_ | ~new_n24326_;
  assign new_n24549_ = ~new_n6169_ | ~new_n24326_;
  assign new_n24550_ = ~new_n24549_ | ~new_n24327_;
  assign new_n24551_ = ~new_n5276_ | ~new_n24325_;
  assign new_n24552_ = ~new_n24369_ | ~new_n24550_;
  assign new_n24553_ = ~new_n24539_ | ~new_n24323_;
  assign new_n24554_ = ~new_n24373_ | ~new_n24553_;
  assign new_n24555_ = ~new_n24328_ | ~new_n24423_;
  assign new_n24556_ = ~new_n24372_ | ~new_n24555_;
  assign new_n24557_ = ~new_n24323_ | ~new_n24423_;
  assign new_n24558_ = ~new_n24527_ | ~new_n24403_;
  assign new_n24559_ = ~new_n24329_;
  assign new_n24560_ = ~new_n5283_ | ~new_n24311_;
  assign new_n24561_ = ~new_n24559_ | ~new_n24560_;
  assign new_n24562_ = ~new_n24377_ | ~new_n24561_;
  assign new_n24563_ = ~new_n24329_ | ~new_n24422_;
  assign new_n24564_ = ~new_n6174_ | ~new_n24313_;
  assign new_n24565_ = ~new_n24376_ | ~new_n24563_;
  assign new_n24566_ = ~new_n5283_ | ~new_n24311_;
  assign new_n24567_ = ~new_n24422_ | ~new_n24566_;
  assign new_n24568_ = ~new_n24527_ | ~new_n24316_;
  assign new_n24569_ = ~new_n24501_ | ~new_n24412_;
  assign new_n24570_ = ~new_n24330_;
  assign new_n24571_ = ~new_n5296_ | ~new_n24296_;
  assign new_n24572_ = ~new_n24570_ | ~new_n24571_;
  assign new_n24573_ = ~new_n24384_ | ~new_n24572_;
  assign new_n24574_ = ~new_n24330_ | ~new_n24421_;
  assign new_n24575_ = ~new_n5697_ | ~new_n24298_;
  assign new_n24576_ = ~new_n24383_ | ~new_n24574_;
  assign new_n24577_ = ~new_n5296_ | ~new_n24296_;
  assign new_n24578_ = ~new_n24421_ | ~new_n24577_;
  assign new_n24579_ = ~new_n24501_ | ~new_n24301_;
  assign new_n24580_ = ~new_n24456_ | ~new_n24390_;
  assign new_n24581_ = ~new_n24331_;
  assign new_n24582_ = ~new_n5284_ | ~new_n24286_;
  assign new_n24583_ = ~new_n24581_ | ~new_n24582_;
  assign new_n24584_ = ~new_n24388_ | ~new_n24583_;
  assign new_n24585_ = ~new_n24331_ | ~new_n24420_;
  assign new_n24586_ = ~new_n5682_ | ~new_n24288_;
  assign new_n24587_ = ~new_n24387_ | ~new_n24585_;
  assign new_n24588_ = ~new_n5284_ | ~new_n24286_;
  assign new_n24589_ = ~new_n24420_ | ~new_n24588_;
  assign new_n24590_ = ~new_n5299_ | ~new_n24264_;
  assign new_n24591_ = ~new_n5300_ | ~new_n24405_;
  assign new_n24592_ = ~new_n24370_ | ~new_n24547_;
  assign new_n24593_ = ~new_n5676_ | ~new_n24281_;
  assign new_n24594_ = ~new_n5305_ | ~new_n24280_;
  assign new_n24595_ = ~new_n24457_ | ~new_n24390_;
  assign new_n24596_ = ~new_n24455_ | ~new_n24389_;
  assign new_n24597_ = ~new_n5673_ | ~new_n24279_;
  assign new_n24598_ = ~new_n5306_ | ~new_n24276_;
  assign new_n24599_ = ~new_n5673_ | ~new_n24279_;
  assign new_n24600_ = ~new_n5306_ | ~new_n24276_;
  assign new_n24601_ = ~new_n24600_ | ~new_n24599_;
  assign new_n24602_ = ~new_n5670_ | ~new_n24277_;
  assign new_n24603_ = ~new_n5292_ | ~new_n24261_;
  assign new_n24604_ = ~new_n24462_ | ~new_n24282_;
  assign new_n24605_ = ~new_n24391_ | ~new_n24449_;
  assign new_n24606_ = ~new_n5667_ | ~new_n24272_;
  assign new_n24607_ = ~new_n5293_ | ~new_n24270_;
  assign new_n24608_ = ~new_n24607_ | ~new_n24606_;
  assign new_n24609_ = ~new_n5664_ | ~new_n24273_;
  assign new_n24610_ = ~new_n5289_ | ~new_n24262_;
  assign new_n24611_ = ~new_n24472_ | ~new_n24283_;
  assign new_n24612_ = ~new_n24392_ | ~new_n24464_;
  assign new_n24613_ = ~new_n5661_ | ~new_n24274_;
  assign new_n24614_ = ~new_n5282_ | ~new_n24271_;
  assign new_n24615_ = ~new_n24473_ | ~new_n24394_;
  assign new_n24616_ = ~new_n24439_ | ~new_n24393_;
  assign new_n24617_ = ~new_n5658_ | ~new_n24269_;
  assign new_n24618_ = ~new_n5286_ | ~new_n24266_;
  assign new_n24619_ = ~new_n5658_ | ~new_n24269_;
  assign new_n24620_ = ~new_n5286_ | ~new_n24266_;
  assign new_n24621_ = ~new_n24620_ | ~new_n24619_;
  assign new_n24622_ = ~new_n5655_ | ~new_n24267_;
  assign new_n24623_ = ~new_n5290_ | ~new_n24263_;
  assign new_n24624_ = ~new_n24478_ | ~new_n24284_;
  assign new_n24625_ = ~new_n24395_ | ~new_n24433_;
  assign new_n24626_ = ~new_n6180_ | ~new_n24397_;
  assign new_n24627_ = ~new_n5277_ | ~new_n24396_;
  assign new_n24628_ = ~new_n6180_ | ~new_n24397_;
  assign new_n24629_ = ~new_n5277_ | ~new_n24396_;
  assign new_n24630_ = ~new_n24629_ | ~new_n24628_;
  assign new_n24631_ = ~new_n6169_ | ~new_n24326_;
  assign new_n24632_ = ~new_n5276_ | ~new_n24325_;
  assign new_n24633_ = ~new_n24371_;
  assign new_n24634_ = ~new_n24633_ | ~new_n24545_;
  assign new_n24635_ = ~new_n24371_ | ~new_n24327_;
  assign new_n24636_ = ~new_n6170_ | ~new_n24324_;
  assign new_n24637_ = ~new_n5275_ | ~new_n24321_;
  assign new_n24638_ = ~new_n6170_ | ~new_n24324_;
  assign new_n24639_ = ~new_n5275_ | ~new_n24321_;
  assign new_n24640_ = ~new_n24639_ | ~new_n24638_;
  assign new_n24641_ = ~new_n6171_ | ~new_n24322_;
  assign new_n24642_ = ~new_n5279_ | ~new_n24285_;
  assign new_n24643_ = ~new_n24557_ | ~new_n24328_;
  assign new_n24644_ = ~new_n24398_ | ~new_n24539_;
  assign new_n24645_ = ~new_n6172_ | ~new_n24320_;
  assign new_n24646_ = ~new_n5280_ | ~new_n24319_;
  assign new_n24647_ = ~new_n24374_;
  assign new_n24648_ = ~new_n24535_ | ~new_n24647_;
  assign new_n24649_ = ~new_n24374_ | ~new_n24399_;
  assign new_n24650_ = ~new_n6173_ | ~new_n24318_;
  assign new_n24651_ = ~new_n5287_ | ~new_n24317_;
  assign new_n24652_ = ~new_n24375_;
  assign new_n24653_ = ~new_n24531_ | ~new_n24652_;
  assign new_n24654_ = ~new_n24375_ | ~new_n24400_;
  assign new_n24655_ = ~new_n6174_ | ~new_n24313_;
  assign new_n24656_ = ~new_n5288_ | ~new_n24310_;
  assign new_n24657_ = ~new_n24656_ | ~new_n24655_;
  assign new_n24658_ = ~new_n6175_ | ~new_n24314_;
  assign new_n24659_ = ~new_n5283_ | ~new_n24311_;
  assign new_n24660_ = ~new_n24567_ | ~new_n24329_;
  assign new_n24661_ = ~new_n24401_ | ~new_n24559_;
  assign new_n24662_ = ~new_n6176_ | ~new_n24315_;
  assign new_n24663_ = ~new_n5297_ | ~new_n24312_;
  assign new_n24664_ = ~new_n24568_ | ~new_n24403_;
  assign new_n24665_ = ~new_n24521_ | ~new_n24402_;
  assign new_n24666_ = ~new_n6177_ | ~new_n24309_;
  assign new_n24667_ = ~new_n5298_ | ~new_n24308_;
  assign new_n24668_ = ~new_n24378_;
  assign new_n24669_ = ~new_n24517_ | ~new_n24668_;
  assign new_n24670_ = ~new_n24378_ | ~new_n24404_;
  assign new_n24671_ = ~new_n5652_ | ~new_n24265_;
  assign new_n24672_ = ~new_n5300_ | ~new_n24405_;
  assign new_n24673_ = ~new_n24379_;
  assign new_n24674_ = ~new_n24431_ | ~new_n24673_;
  assign new_n24675_ = ~new_n24379_ | ~new_n24406_;
  assign new_n24676_ = ~new_n5705_ | ~new_n24307_;
  assign new_n24677_ = ~new_n5303_ | ~new_n24306_;
  assign new_n24678_ = ~new_n24380_;
  assign new_n24679_ = ~new_n24513_ | ~new_n24678_;
  assign new_n24680_ = ~new_n24380_ | ~new_n24407_;
  assign new_n24681_ = ~new_n5703_ | ~new_n24305_;
  assign new_n24682_ = ~new_n5304_ | ~new_n24408_;
  assign new_n24683_ = ~new_n24381_;
  assign new_n24684_ = ~new_n24683_ | ~new_n24509_;
  assign new_n24685_ = ~new_n24381_ | ~new_n24304_;
  assign new_n24686_ = ~new_n5700_ | ~new_n24303_;
  assign new_n24687_ = ~new_n5291_ | ~new_n24302_;
  assign new_n24688_ = ~new_n24382_;
  assign new_n24689_ = ~new_n24505_ | ~new_n24688_;
  assign new_n24690_ = ~new_n24382_ | ~new_n24409_;
  assign new_n24691_ = ~new_n5697_ | ~new_n24298_;
  assign new_n24692_ = ~new_n5295_ | ~new_n24295_;
  assign new_n24693_ = ~new_n24692_ | ~new_n24691_;
  assign new_n24694_ = ~new_n5694_ | ~new_n24299_;
  assign new_n24695_ = ~new_n5296_ | ~new_n24296_;
  assign new_n24696_ = ~new_n24578_ | ~new_n24330_;
  assign new_n24697_ = ~new_n24410_ | ~new_n24570_;
  assign new_n24698_ = ~new_n5691_ | ~new_n24300_;
  assign new_n24699_ = ~new_n5301_ | ~new_n24297_;
  assign new_n24700_ = ~new_n24579_ | ~new_n24412_;
  assign new_n24701_ = ~new_n24495_ | ~new_n24411_;
  assign new_n24702_ = ~new_n5688_ | ~new_n24294_;
  assign new_n24703_ = ~new_n5302_ | ~new_n24293_;
  assign new_n24704_ = ~new_n24385_;
  assign new_n24705_ = ~new_n24491_ | ~new_n24704_;
  assign new_n24706_ = ~new_n24385_ | ~new_n24413_;
  assign new_n24707_ = ~new_n5685_ | ~new_n24292_;
  assign new_n24708_ = ~new_n5294_ | ~new_n24291_;
  assign new_n24709_ = ~new_n24386_;
  assign new_n24710_ = ~new_n24487_ | ~new_n24709_;
  assign new_n24711_ = ~new_n24386_ | ~new_n24414_;
  assign new_n24712_ = ~new_n5682_ | ~new_n24288_;
  assign new_n24713_ = ~new_n5285_ | ~new_n24287_;
  assign new_n24714_ = ~new_n24713_ | ~new_n24712_;
  assign new_n24715_ = ~new_n5679_ | ~new_n24289_;
  assign new_n24716_ = ~new_n5284_ | ~new_n24286_;
  assign new_n24717_ = ~new_n24589_ | ~new_n24331_;
  assign new_n24718_ = ~new_n24415_ | ~new_n24581_;
  assign new_n24719_ = ~pi543 & ~pi541 & ~pi540 & ~pi542;
  assign new_n24720_ = new_n24849_ & new_n24762_;
  assign new_n24721_ = new_n24847_ & new_n24815_;
  assign new_n24722_ = new_n24846_ & new_n24759_;
  assign new_n24723_ = new_n24845_ & new_n24760_;
  assign new_n24724_ = new_n24843_ & new_n24818_;
  assign new_n24725_ = new_n24842_ & new_n24747_;
  assign new_n24726_ = new_n24841_ & new_n24757_;
  assign new_n24727_ = new_n24839_ & new_n24821_;
  assign new_n24728_ = new_n24838_ & new_n24753_;
  assign new_n24729_ = new_n24837_ & new_n24754_;
  assign new_n24730_ = new_n24835_ & new_n24824_;
  assign new_n24731_ = new_n24834_ & new_n24748_;
  assign new_n24732_ = new_n24833_ & new_n24791_;
  assign new_n24733_ = new_n24778_ & new_n24852_;
  assign new_n24734_ = new_n24831_ & new_n24750_;
  assign new_n24735_ = new_n24830_ & new_n24741_;
  assign new_n24736_ = new_n24813_ & new_n24803_;
  assign new_n24737_ = new_n24812_ & new_n24743_;
  assign new_n24738_ = new_n24811_ & new_n24744_;
  assign new_n24739_ = new_n24809_ & new_n24806_;
  assign new_n24740_ = new_n24808_ & new_n24742_;
  assign new_n24741_ = pi525 | pi524 | pi523;
  assign new_n24742_ = ~new_n24766_ | ~new_n24767_ | ~new_n24853_;
  assign new_n24743_ = ~new_n24768_ | ~new_n24853_;
  assign new_n24744_ = ~new_n24769_ | ~new_n24804_;
  assign new_n24745_ = ~pi530;
  assign new_n24746_ = ~pi526;
  assign new_n24747_ = ~new_n24772_ | ~new_n24770_ | ~new_n24771_ | ~new_n24773_;
  assign new_n24748_ = ~new_n24775_ | ~new_n24819_;
  assign new_n24749_ = ~new_n24776_ | ~new_n24825_;
  assign new_n24750_ = ~new_n24827_ | ~new_n24751_;
  assign new_n24751_ = ~pi552;
  assign new_n24752_ = ~pi550;
  assign new_n24753_ = ~new_n24819_ | ~new_n24719_;
  assign new_n24754_ = ~new_n24779_ | ~new_n24822_;
  assign new_n24755_ = ~pi547;
  assign new_n24756_ = ~pi546;
  assign new_n24757_ = ~new_n24780_ | ~new_n24819_;
  assign new_n24758_ = ~pi542;
  assign new_n24759_ = ~new_n24781_ | ~new_n24807_;
  assign new_n24760_ = ~new_n24782_ | ~new_n24816_;
  assign new_n24761_ = ~pi538;
  assign new_n24762_ = ~new_n24783_ | ~new_n24807_;
  assign new_n24763_ = ~pi534;
  assign new_n24764_ = ~new_n24869_ | ~new_n24868_;
  assign new_n24765_ = ~new_n24859_ | ~new_n24858_;
  assign new_n24766_ = ~pi527 & ~pi529 & ~pi528 & ~pi526;
  assign new_n24767_ = ~pi530 & ~pi531;
  assign new_n24768_ = ~pi526 & ~pi527;
  assign new_n24769_ = ~pi528 & ~pi529;
  assign new_n24770_ = ~pi537 & ~pi536 & ~pi534 & ~pi533 & ~pi535;
  assign new_n24771_ = ~pi539 & ~pi523 & ~pi524 & ~pi538;
  assign new_n24772_ = ~pi526 & ~pi528 & ~pi527 & ~pi525;
  assign new_n24773_ = ~pi530 & ~pi532 & ~pi531 & ~pi529;
  assign new_n24774_ = ~pi545 & ~pi546 & ~pi544;
  assign new_n24775_ = new_n24774_ & new_n24719_ & new_n24755_;
  assign new_n24776_ = ~pi549 & ~pi551 & ~pi550 & ~pi548;
  assign new_n24777_ = ~pi548 & ~pi549;
  assign new_n24778_ = new_n24851_ & new_n24749_;
  assign new_n24779_ = ~pi544 & ~pi545;
  assign new_n24780_ = ~pi540 & ~pi541;
  assign new_n24781_ = ~pi534 & ~pi532 & ~pi535 & ~pi533;
  assign new_n24782_ = ~pi536 & ~pi537;
  assign new_n24783_ = ~pi533 & ~pi532;
  assign new_n24784_ = ~pi532;
  assign new_n24785_ = new_n24855_ & new_n24854_;
  assign new_n24786_ = ~pi528;
  assign new_n24787_ = new_n24857_ & new_n24856_;
  assign new_n24788_ = ~pi554;
  assign new_n24789_ = ~pi553;
  assign new_n24790_ = new_n24861_ & new_n24860_;
  assign new_n24791_ = ~new_n24777_ | ~new_n24825_;
  assign new_n24792_ = new_n24863_ & new_n24862_;
  assign new_n24793_ = ~pi548;
  assign new_n24794_ = new_n24865_ & new_n24864_;
  assign new_n24795_ = ~pi544;
  assign new_n24796_ = new_n24867_ & new_n24866_;
  assign new_n24797_ = ~pi524;
  assign new_n24798_ = ~pi523;
  assign new_n24799_ = ~pi540;
  assign new_n24800_ = new_n24871_ & new_n24870_;
  assign new_n24801_ = ~pi536;
  assign new_n24802_ = new_n24873_ & new_n24872_;
  assign new_n24803_ = ~new_n24853_ | ~new_n24746_;
  assign new_n24804_ = ~new_n24743_;
  assign new_n24805_ = ~new_n24744_;
  assign new_n24806_ = ~new_n24805_ | ~new_n24745_;
  assign new_n24807_ = ~new_n24742_;
  assign new_n24808_ = ~pi531 | ~new_n24806_;
  assign new_n24809_ = ~pi530 | ~new_n24744_;
  assign new_n24810_ = ~new_n24804_ | ~new_n24786_;
  assign new_n24811_ = ~pi529 | ~new_n24810_;
  assign new_n24812_ = ~pi527 | ~new_n24803_;
  assign new_n24813_ = ~pi526 | ~new_n24741_;
  assign new_n24814_ = ~new_n24762_;
  assign new_n24815_ = ~new_n24814_ | ~new_n24763_;
  assign new_n24816_ = ~new_n24759_;
  assign new_n24817_ = ~new_n24760_;
  assign new_n24818_ = ~new_n24817_ | ~new_n24761_;
  assign new_n24819_ = ~new_n24747_;
  assign new_n24820_ = ~new_n24757_;
  assign new_n24821_ = ~new_n24820_ | ~new_n24758_;
  assign new_n24822_ = ~new_n24753_;
  assign new_n24823_ = ~new_n24754_;
  assign new_n24824_ = ~new_n24823_ | ~new_n24756_;
  assign new_n24825_ = ~new_n24748_;
  assign new_n24826_ = ~new_n24791_;
  assign new_n24827_ = ~new_n24749_;
  assign new_n24828_ = ~new_n24750_;
  assign new_n24829_ = pi524 | pi523;
  assign new_n24830_ = ~pi525 | ~new_n24829_;
  assign new_n24831_ = ~pi552 | ~new_n24749_;
  assign new_n24832_ = ~new_n24825_ | ~new_n24793_;
  assign new_n24833_ = ~pi549 | ~new_n24832_;
  assign new_n24834_ = ~pi547 | ~new_n24824_;
  assign new_n24835_ = ~pi546 | ~new_n24754_;
  assign new_n24836_ = ~new_n24822_ | ~new_n24795_;
  assign new_n24837_ = ~pi545 | ~new_n24836_;
  assign new_n24838_ = ~pi543 | ~new_n24821_;
  assign new_n24839_ = ~pi542 | ~new_n24757_;
  assign new_n24840_ = ~new_n24819_ | ~new_n24799_;
  assign new_n24841_ = ~pi541 | ~new_n24840_;
  assign new_n24842_ = ~pi539 | ~new_n24818_;
  assign new_n24843_ = ~pi538 | ~new_n24760_;
  assign new_n24844_ = ~new_n24816_ | ~new_n24801_;
  assign new_n24845_ = ~pi537 | ~new_n24844_;
  assign new_n24846_ = ~pi535 | ~new_n24815_;
  assign new_n24847_ = ~pi534 | ~new_n24762_;
  assign new_n24848_ = ~new_n24807_ | ~new_n24784_;
  assign new_n24849_ = ~pi533 | ~new_n24848_;
  assign new_n24850_ = ~new_n24828_ | ~new_n24789_;
  assign new_n24851_ = ~pi550 | ~pi551;
  assign new_n24852_ = ~pi551 | ~new_n24791_;
  assign new_n24853_ = ~new_n24741_;
  assign new_n24854_ = ~pi532 | ~new_n24742_;
  assign new_n24855_ = ~new_n24807_ | ~new_n24784_;
  assign new_n24856_ = ~pi528 | ~new_n24743_;
  assign new_n24857_ = ~new_n24804_ | ~new_n24786_;
  assign new_n24858_ = ~new_n24850_ | ~new_n24788_;
  assign new_n24859_ = ~pi554 | ~new_n24828_ | ~new_n24789_;
  assign new_n24860_ = ~pi553 | ~new_n24750_;
  assign new_n24861_ = ~new_n24828_ | ~new_n24789_;
  assign new_n24862_ = ~pi550 | ~new_n24791_;
  assign new_n24863_ = ~new_n24826_ | ~new_n24752_;
  assign new_n24864_ = ~pi548 | ~new_n24748_;
  assign new_n24865_ = ~new_n24825_ | ~new_n24793_;
  assign new_n24866_ = ~pi544 | ~new_n24753_;
  assign new_n24867_ = ~new_n24822_ | ~new_n24795_;
  assign new_n24868_ = ~pi524 | ~new_n24798_;
  assign new_n24869_ = ~pi523 | ~new_n24797_;
  assign new_n24870_ = ~pi540 | ~new_n24747_;
  assign new_n24871_ = ~new_n24819_ | ~new_n24799_;
  assign new_n24872_ = ~pi536 | ~new_n24759_;
  assign new_n24873_ = ~new_n24816_ | ~new_n24801_;
  assign new_n24874_ = new_n24981_ & new_n24982_;
  assign new_n24875_ = new_n24983_ & new_n24984_;
  assign new_n24876_ = new_n24986_ & new_n24875_ & new_n24988_ & new_n24948_;
  assign new_n24877_ = new_n24994_ & new_n24993_;
  assign new_n24878_ = new_n24998_ & new_n24999_;
  assign new_n24879_ = new_n24952_ & new_n24878_;
  assign new_n24880_ = new_n25010_ & new_n25009_;
  assign new_n24881_ = new_n25045_ & new_n25046_ & new_n25047_;
  assign new_n24882_ = new_n25056_ & new_n24977_ & new_n24976_ & new_n25057_;
  assign new_n24883_ = ~new_n8907_;
  assign new_n24884_ = ~new_n8915_;
  assign new_n24885_ = ~new_n8914_;
  assign new_n24886_ = ~new_n9283_;
  assign new_n24887_ = ~new_n8918_;
  assign new_n24888_ = ~new_n9284_;
  assign new_n24889_ = ~new_n8919_;
  assign new_n24890_ = ~new_n8921_;
  assign new_n24891_ = ~new_n8821_;
  assign new_n24892_ = ~new_n8922_;
  assign new_n24893_ = ~new_n8818_;
  assign new_n24894_ = ~new_n8823_;
  assign new_n24895_ = ~new_n9285_;
  assign new_n24896_ = ~new_n8923_;
  assign new_n24897_ = ~new_n8924_;
  assign new_n24898_ = ~new_n8815_;
  assign new_n24899_ = ~new_n8812_;
  assign new_n24900_ = ~new_n8904_;
  assign new_n24901_ = ~new_n8903_;
  assign new_n24902_ = ~new_n8782_;
  assign new_n24903_ = ~new_n8785_;
  assign new_n24904_ = ~new_n8794_;
  assign new_n24905_ = ~new_n8797_;
  assign new_n24906_ = ~new_n8788_;
  assign new_n24907_ = ~new_n8791_;
  assign new_n24908_ = ~new_n8776_;
  assign new_n24909_ = ~new_n8779_;
  assign new_n24910_ = ~new_n8931_;
  assign new_n24911_ = ~new_n8773_;
  assign new_n24912_ = ~new_n8770_;
  assign new_n24913_ = ~new_n8928_;
  assign new_n24914_ = ~new_n8927_;
  assign new_n24915_ = ~new_n8920_;
  assign new_n24916_ = ~new_n8909_;
  assign new_n24917_ = ~new_n8906_;
  assign new_n24918_ = ~new_n8905_;
  assign new_n24919_ = ~new_n8901_;
  assign new_n24920_ = ~new_n8902_;
  assign new_n24921_ = ~new_n8930_;
  assign new_n24922_ = ~new_n8929_;
  assign new_n24923_ = ~new_n8803_;
  assign new_n24924_ = ~new_n8800_;
  assign new_n24925_ = ~new_n8809_;
  assign new_n24926_ = ~new_n8806_;
  assign new_n24927_ = ~new_n8926_;
  assign new_n24928_ = ~new_n8925_;
  assign new_n24929_ = ~new_n8917_;
  assign new_n24930_ = ~new_n8916_;
  assign new_n24931_ = ~new_n9286_;
  assign new_n24932_ = ~new_n9278_;
  assign new_n24933_ = ~new_n9277_;
  assign new_n24934_ = ~new_n9282_;
  assign new_n24935_ = ~new_n9281_;
  assign new_n24936_ = ~new_n9280_;
  assign new_n24937_ = ~new_n9279_;
  assign new_n24938_ = ~new_n8911_;
  assign new_n24939_ = ~new_n8912_;
  assign new_n24940_ = ~new_n9250_;
  assign new_n24941_ = ~new_n8910_;
  assign new_n24942_ = ~new_n8913_;
  assign new_n24943_ = new_n8918_ & new_n24888_;
  assign new_n24944_ = new_n8919_ & new_n24895_;
  assign new_n24945_ = new_n25036_ & new_n25035_;
  assign new_n24946_ = new_n8821_ & new_n24892_;
  assign new_n24947_ = new_n8818_ & new_n24896_;
  assign new_n24948_ = new_n24987_ & new_n24985_;
  assign new_n24949_ = new_n8782_ & new_n24918_;
  assign new_n24950_ = new_n8785_ & new_n24900_;
  assign new_n24951_ = new_n8765_ & new_n24979_;
  assign new_n24952_ = new_n25001_ & new_n25000_;
  assign new_n24953_ = new_n24997_ & new_n24954_;
  assign new_n24954_ = new_n25003_ & new_n25002_;
  assign new_n24955_ = new_n25006_ & new_n25005_;
  assign new_n24956_ = new_n25003_ & new_n25002_;
  assign new_n24957_ = new_n24877_ & new_n25016_;
  assign new_n24958_ = new_n24879_ & new_n24997_ & new_n24995_;
  assign new_n24959_ = new_n8901_ & new_n24904_;
  assign new_n24960_ = new_n8902_ & new_n24907_;
  assign new_n24961_ = new_n24963_ & new_n25020_ & new_n25019_;
  assign new_n24962_ = new_n25022_ & new_n25021_;
  assign new_n24963_ = new_n24962_ & new_n24880_;
  assign new_n24964_ = new_n8803_ & new_n24913_;
  assign new_n24965_ = new_n8800_ & new_n24922_;
  assign new_n24966_ = new_n25025_ & new_n24968_;
  assign new_n24967_ = new_n24966_ & new_n25026_;
  assign new_n24968_ = new_n25028_ & new_n25027_;
  assign new_n24969_ = new_n25038_ & new_n24991_ & new_n24990_ & new_n25039_;
  assign new_n24970_ = new_n25043_ & new_n25042_;
  assign new_n24971_ = new_n25055_ & new_n25054_;
  assign new_n24972_ = new_n24971_ & new_n24881_;
  assign new_n24973_ = new_n24974_ & new_n25058_;
  assign new_n24974_ = new_n8911_ & new_n24933_;
  assign new_n24975_ = new_n8910_ & new_n24931_;
  assign new_n24976_ = new_n25060_ & new_n25059_;
  assign new_n24977_ = new_n25063_ & new_n25062_ & new_n25061_;
  assign new_n24978_ = ~new_n9251_;
  assign new_n24979_ = ~new_n8932_;
  assign new_n24980_ = ~new_n25049_ | ~new_n25064_;
  assign new_n24981_ = ~new_n8921_ | ~new_n24894_;
  assign new_n24982_ = ~new_n8922_ | ~new_n24891_;
  assign new_n24983_ = ~new_n9283_ | ~new_n24929_;
  assign new_n24984_ = ~new_n9284_ | ~new_n24887_;
  assign new_n24985_ = ~new_n24946_ | ~new_n24981_;
  assign new_n24986_ = ~new_n24947_ | ~new_n24874_;
  assign new_n24987_ = ~new_n8823_ | ~new_n24890_;
  assign new_n24988_ = ~new_n9285_ | ~new_n24889_;
  assign new_n24989_ = ~new_n8815_ | ~new_n24897_;
  assign new_n24990_ = ~new_n8915_ | ~new_n24935_;
  assign new_n24991_ = ~new_n8914_ | ~new_n24936_;
  assign new_n24992_ = ~new_n8812_ | ~new_n24928_;
  assign new_n24993_ = ~new_n8904_ | ~new_n24903_;
  assign new_n24994_ = ~new_n8903_ | ~new_n24906_;
  assign new_n24995_ = ~new_n24949_ | ~new_n24877_;
  assign new_n24996_ = ~new_n8903_ | ~new_n24906_;
  assign new_n24997_ = ~new_n24950_ | ~new_n24996_;
  assign new_n24998_ = ~new_n8797_ | ~new_n24921_;
  assign new_n24999_ = ~new_n8794_ | ~new_n24919_;
  assign new_n25000_ = ~new_n8788_ | ~new_n24901_;
  assign new_n25001_ = ~new_n8791_ | ~new_n24920_;
  assign new_n25002_ = ~new_n8776_ | ~new_n24916_;
  assign new_n25003_ = ~new_n8779_ | ~new_n24917_;
  assign new_n25004_ = ~new_n8931_ | ~new_n24912_;
  assign new_n25005_ = ~new_n24951_ | ~new_n25004_;
  assign new_n25006_ = ~new_n8773_ | ~new_n24915_;
  assign new_n25007_ = ~new_n8770_ | ~new_n24910_;
  assign new_n25008_ = ~new_n24879_ | ~new_n24953_ | ~new_n24995_ | ~new_n24955_ | ~new_n25007_;
  assign new_n25009_ = ~new_n8928_ | ~new_n24923_;
  assign new_n25010_ = ~new_n8927_ | ~new_n24926_;
  assign new_n25011_ = ~new_n8920_ | ~new_n24911_;
  assign new_n25012_ = ~new_n8909_ | ~new_n24908_;
  assign new_n25013_ = ~new_n25012_ | ~new_n25011_;
  assign new_n25014_ = ~new_n24956_ | ~new_n25013_;
  assign new_n25015_ = ~new_n8906_ | ~new_n24909_;
  assign new_n25016_ = ~new_n8905_ | ~new_n24902_;
  assign new_n25017_ = ~new_n24957_ | ~new_n25015_ | ~new_n25014_;
  assign new_n25018_ = ~new_n24958_ | ~new_n25017_;
  assign new_n25019_ = ~new_n24959_ | ~new_n24998_;
  assign new_n25020_ = ~new_n24960_ | ~new_n24878_;
  assign new_n25021_ = ~new_n8930_ | ~new_n24905_;
  assign new_n25022_ = ~new_n8929_ | ~new_n24924_;
  assign new_n25023_ = ~new_n24961_ | ~new_n25018_ | ~new_n25008_;
  assign new_n25024_ = ~new_n8927_ | ~new_n24926_;
  assign new_n25025_ = ~new_n24964_ | ~new_n25024_;
  assign new_n25026_ = ~new_n24965_ | ~new_n24880_;
  assign new_n25027_ = ~new_n8809_ | ~new_n24927_;
  assign new_n25028_ = ~new_n8806_ | ~new_n24914_;
  assign new_n25029_ = ~new_n25023_ | ~new_n24967_;
  assign new_n25030_ = ~new_n8926_ | ~new_n24925_;
  assign new_n25031_ = ~new_n25030_ | ~new_n25029_;
  assign new_n25032_ = ~new_n25031_ | ~new_n24992_;
  assign new_n25033_ = ~new_n8925_ | ~new_n24899_;
  assign new_n25034_ = ~new_n25033_ | ~new_n25032_;
  assign new_n25035_ = ~new_n8923_ | ~new_n24893_;
  assign new_n25036_ = ~new_n8924_ | ~new_n24898_;
  assign new_n25037_ = ~new_n24945_ | ~new_n24874_;
  assign new_n25038_ = ~new_n24943_ | ~new_n24983_;
  assign new_n25039_ = ~new_n24944_ | ~new_n24875_;
  assign new_n25040_ = ~new_n24876_ | ~new_n25037_;
  assign new_n25041_ = ~new_n24876_ | ~new_n25034_ | ~new_n24989_;
  assign new_n25042_ = ~new_n8917_ | ~new_n24886_;
  assign new_n25043_ = ~new_n8916_ | ~new_n24934_;
  assign new_n25044_ = ~new_n25040_ | ~new_n24969_ | ~new_n24970_ | ~new_n25041_;
  assign new_n25045_ = ~new_n9286_ | ~new_n24941_;
  assign new_n25046_ = ~new_n9278_ | ~new_n24939_;
  assign new_n25047_ = ~new_n9277_ | ~new_n24938_;
  assign new_n25048_ = ~new_n8907_ | ~new_n24940_;
  assign new_n25049_ = ~new_n25048_ | ~new_n24978_;
  assign new_n25050_ = ~new_n9282_ | ~new_n24930_;
  assign new_n25051_ = ~new_n9281_ | ~new_n24884_;
  assign new_n25052_ = ~new_n25051_ | ~new_n25050_;
  assign new_n25053_ = ~new_n24991_ | ~new_n25052_ | ~new_n24990_;
  assign new_n25054_ = ~new_n9280_ | ~new_n24885_;
  assign new_n25055_ = ~new_n9279_ | ~new_n24942_;
  assign new_n25056_ = ~new_n25053_ | ~new_n24972_ | ~new_n24980_ | ~new_n25044_;
  assign new_n25057_ = ~new_n24978_ | ~new_n25048_ | ~new_n8908_;
  assign new_n25058_ = ~new_n9286_ | ~new_n24941_;
  assign new_n25059_ = ~new_n24980_ | ~new_n24973_;
  assign new_n25060_ = ~new_n24881_ | ~new_n24932_ | ~new_n24980_ | ~new_n8912_;
  assign new_n25061_ = ~new_n9250_ | ~new_n24883_;
  assign new_n25062_ = ~new_n24975_ | ~new_n24980_;
  assign new_n25063_ = ~new_n24881_ | ~new_n24937_ | ~new_n24980_ | ~new_n8913_;
  assign new_n25064_ = ~new_n8908_ | ~new_n25048_;
  assign new_n25065_ = ~new_n25099_ | ~new_n25157_;
  assign new_n25066_ = ~new_n25138_ | ~new_n25164_;
  assign new_n25067_ = ~new_n25124_ | ~new_n25172_;
  assign new_n25068_ = ~new_n25093_ | ~new_n25169_;
  assign new_n25069_ = ~new_n25146_ | ~new_n25156_;
  assign new_n25070_ = ~new_n25140_ | ~new_n25162_;
  assign new_n25071_ = ~new_n25126_ | ~new_n25129_;
  assign new_n25072_ = ~new_n25132_ | ~new_n25170_;
  assign new_n25073_ = ~new_n25092_ | ~new_n25128_;
  assign new_n25074_ = ~new_n25097_ | ~new_n25161_;
  assign new_n25075_ = ~new_n25100_ | ~new_n25155_;
  assign new_n25076_ = ~new_n25144_ | ~new_n25158_;
  assign new_n25077_ = ~new_n25090_ | ~new_n25130_;
  assign new_n25078_ = ~new_n25096_ | ~new_n25163_;
  assign new_n25079_ = ~new_n25142_ | ~new_n25160_;
  assign new_n25080_ = ~new_n25095_ | ~new_n25165_;
  assign new_n25081_ = ~new_n25101_ | ~new_n25153_;
  assign new_n25082_ = ~new_n25134_ | ~new_n25168_;
  assign new_n25083_ = ~new_n25094_ | ~new_n25167_;
  assign new_n25084_ = ~pi759;
  assign new_n25085_ = ~new_n25148_ | ~new_n25154_;
  assign new_n25086_ = ~new_n25098_ | ~new_n25159_;
  assign new_n25087_ = ~new_n25150_ | ~new_n25152_;
  assign new_n25088_ = ~new_n25123_ | ~new_n25131_;
  assign new_n25089_ = ~new_n25136_ | ~new_n25166_;
  assign new_n25090_ = pi759 | pi747 | pi764 | pi738 | pi750;
  assign new_n25091_ = ~pi756;
  assign new_n25092_ = ~new_n25113_ | ~new_n25125_;
  assign new_n25093_ = ~new_n25114_ | ~new_n25127_;
  assign new_n25094_ = ~new_n25115_ | ~new_n25133_;
  assign new_n25095_ = ~new_n25116_ | ~new_n25135_;
  assign new_n25096_ = ~new_n25117_ | ~new_n25137_;
  assign new_n25097_ = ~new_n25118_ | ~new_n25139_;
  assign new_n25098_ = ~new_n25119_ | ~new_n25141_;
  assign new_n25099_ = ~new_n25120_ | ~new_n25143_;
  assign new_n25100_ = ~new_n25121_ | ~new_n25145_;
  assign new_n25101_ = ~new_n25122_ | ~new_n25147_;
  assign new_n25102_ = ~pi757;
  assign new_n25103_ = ~pi737;
  assign new_n25104_ = ~pi748;
  assign new_n25105_ = ~pi742;
  assign new_n25106_ = ~pi744;
  assign new_n25107_ = ~pi739;
  assign new_n25108_ = ~pi751;
  assign new_n25109_ = ~pi762;
  assign new_n25110_ = ~pi753;
  assign new_n25111_ = ~pi760;
  assign new_n25112_ = ~new_n25174_ | ~new_n25173_;
  assign new_n25113_ = ~pi756 & ~pi746;
  assign new_n25114_ = ~pi760 & ~pi741;
  assign new_n25115_ = ~pi753 & ~pi743;
  assign new_n25116_ = ~pi762 & ~pi736;
  assign new_n25117_ = ~pi751 & ~pi749;
  assign new_n25118_ = ~pi739 & ~pi758;
  assign new_n25119_ = ~pi744 & ~pi754;
  assign new_n25120_ = ~pi742 & ~pi761;
  assign new_n25121_ = ~pi748 & ~pi752;
  assign new_n25122_ = ~pi737 & ~pi763;
  assign new_n25123_ = pi759 | pi747;
  assign new_n25124_ = pi738 | pi759 | pi747 | pi750;
  assign new_n25125_ = ~new_n25090_;
  assign new_n25126_ = ~new_n25125_ | ~new_n25091_;
  assign new_n25127_ = ~new_n25092_;
  assign new_n25128_ = ~pi746 | ~new_n25126_;
  assign new_n25129_ = ~pi756 | ~new_n25090_;
  assign new_n25130_ = ~pi764 | ~new_n25124_;
  assign new_n25131_ = ~pi747 | ~pi759;
  assign new_n25132_ = ~new_n25127_ | ~new_n25111_;
  assign new_n25133_ = ~new_n25093_;
  assign new_n25134_ = ~new_n25133_ | ~new_n25110_;
  assign new_n25135_ = ~new_n25094_;
  assign new_n25136_ = ~new_n25135_ | ~new_n25109_;
  assign new_n25137_ = ~new_n25095_;
  assign new_n25138_ = ~new_n25137_ | ~new_n25108_;
  assign new_n25139_ = ~new_n25096_;
  assign new_n25140_ = ~new_n25139_ | ~new_n25107_;
  assign new_n25141_ = ~new_n25097_;
  assign new_n25142_ = ~new_n25141_ | ~new_n25106_;
  assign new_n25143_ = ~new_n25098_;
  assign new_n25144_ = ~new_n25143_ | ~new_n25105_;
  assign new_n25145_ = ~new_n25099_;
  assign new_n25146_ = ~new_n25145_ | ~new_n25104_;
  assign new_n25147_ = ~new_n25100_;
  assign new_n25148_ = ~new_n25147_ | ~new_n25103_;
  assign new_n25149_ = ~new_n25101_;
  assign new_n25150_ = ~new_n25149_ | ~new_n25102_;
  assign new_n25151_ = ~new_n25150_;
  assign new_n25152_ = ~pi757 | ~new_n25101_;
  assign new_n25153_ = ~pi763 | ~new_n25148_;
  assign new_n25154_ = ~pi737 | ~new_n25100_;
  assign new_n25155_ = ~pi752 | ~new_n25146_;
  assign new_n25156_ = ~pi748 | ~new_n25099_;
  assign new_n25157_ = ~pi761 | ~new_n25144_;
  assign new_n25158_ = ~pi742 | ~new_n25098_;
  assign new_n25159_ = ~pi754 | ~new_n25142_;
  assign new_n25160_ = ~pi744 | ~new_n25097_;
  assign new_n25161_ = ~pi758 | ~new_n25140_;
  assign new_n25162_ = ~pi739 | ~new_n25096_;
  assign new_n25163_ = ~pi749 | ~new_n25138_;
  assign new_n25164_ = ~pi751 | ~new_n25095_;
  assign new_n25165_ = ~pi736 | ~new_n25136_;
  assign new_n25166_ = ~pi762 | ~new_n25094_;
  assign new_n25167_ = ~pi743 | ~new_n25134_;
  assign new_n25168_ = ~pi753 | ~new_n25093_;
  assign new_n25169_ = ~pi741 | ~new_n25132_;
  assign new_n25170_ = ~pi760 | ~new_n25092_;
  assign new_n25171_ = pi750 | pi747 | pi759;
  assign new_n25172_ = ~pi738 | ~new_n25171_;
  assign new_n25173_ = ~pi750 | ~new_n25123_;
  assign new_n25174_ = pi750 | pi747 | pi759;
  assign new_n25175_ = new_n25379_ & new_n25378_;
  assign new_n25176_ = new_n25358_ & new_n25414_;
  assign new_n25177_ = new_n25416_ & new_n25415_;
  assign new_n25178_ = new_n25359_ & new_n25431_;
  assign new_n25179_ = new_n25433_ & new_n25432_;
  assign new_n25180_ = new_n25360_ & new_n25455_;
  assign new_n25181_ = new_n25457_ & new_n25456_;
  assign new_n25182_ = new_n25382_ & new_n25377_ & new_n25363_;
  assign new_n25183_ = new_n25387_ & new_n25364_;
  assign new_n25184_ = new_n25561_ & new_n25560_;
  assign new_n25185_ = ~new_n25511_ | ~new_n25514_;
  assign new_n25186_ = ~new_n25500_ | ~new_n25503_;
  assign new_n25187_ = ~new_n25489_ | ~new_n25492_;
  assign new_n25188_ = ~new_n25481_ | ~new_n25483_;
  assign new_n25189_ = ~new_n25520_ | ~new_n25331_ | ~new_n25352_;
  assign new_n25190_ = ~new_n25410_ | ~new_n25412_;
  assign new_n25191_ = ~new_n25402_ | ~new_n25405_;
  assign new_n25192_ = ~new_n25394_ | ~new_n25396_;
  assign new_n25193_ = ~new_n25341_ | ~new_n25517_;
  assign new_n25194_ = ~new_n8447_;
  assign new_n25195_ = ~new_n8447_ | ~new_n25208_;
  assign new_n25196_ = ~new_n8461_;
  assign new_n25197_ = ~new_n8791_;
  assign new_n25198_ = ~new_n8773_;
  assign new_n25199_ = ~new_n8765_;
  assign new_n25200_ = ~new_n8455_;
  assign new_n25201_ = ~new_n8776_;
  assign new_n25202_ = ~new_n8445_;
  assign new_n25203_ = ~new_n8445_ | ~new_n25198_;
  assign new_n25204_ = ~new_n8441_;
  assign new_n25205_ = ~new_n8782_;
  assign new_n25206_ = ~new_n8785_;
  assign new_n25207_ = ~new_n8779_;
  assign new_n25208_ = ~new_n8788_;
  assign new_n25209_ = ~new_n8448_;
  assign new_n25210_ = ~new_n8444_;
  assign new_n25211_ = ~new_n8437_;
  assign new_n25212_ = ~new_n8437_ | ~new_n25207_;
  assign new_n25213_ = ~new_n25383_ | ~new_n25381_;
  assign new_n25214_ = ~new_n8794_;
  assign new_n25215_ = ~new_n8460_;
  assign new_n25216_ = ~new_n25213_ | ~new_n25384_;
  assign new_n25217_ = ~new_n25212_ | ~new_n25398_;
  assign new_n25218_ = ~new_n25518_ | ~new_n25370_ | ~new_n25354_;
  assign new_n25219_ = ~new_n9279_;
  assign new_n25220_ = ~new_n8800_;
  assign new_n25221_ = ~new_n8797_;
  assign new_n25222_ = ~new_n8440_;
  assign new_n25223_ = ~new_n8439_;
  assign new_n25224_ = ~new_n8460_ | ~new_n25214_;
  assign new_n25225_ = ~new_n8803_;
  assign new_n25226_ = ~new_n8449_;
  assign new_n25227_ = ~new_n8806_;
  assign new_n25228_ = ~new_n8457_;
  assign new_n25229_ = ~new_n8815_;
  assign new_n25230_ = ~new_n8812_;
  assign new_n25231_ = ~new_n8809_;
  assign new_n25232_ = ~new_n8450_;
  assign new_n25233_ = ~new_n8451_;
  assign new_n25234_ = ~new_n8456_;
  assign new_n25235_ = ~new_n8456_ | ~new_n25231_;
  assign new_n25236_ = ~new_n8818_;
  assign new_n25237_ = ~new_n8446_;
  assign new_n25238_ = ~new_n8459_;
  assign new_n25239_ = ~new_n8823_;
  assign new_n25240_ = ~new_n8458_;
  assign new_n25241_ = ~new_n9285_;
  assign new_n25242_ = ~new_n8453_;
  assign new_n25243_ = ~new_n9282_;
  assign new_n25244_ = ~new_n9283_;
  assign new_n25245_ = ~new_n9284_;
  assign new_n25246_ = ~new_n8443_;
  assign new_n25247_ = ~new_n8438_;
  assign new_n25248_ = ~new_n8452_;
  assign new_n25249_ = ~new_n8452_ | ~new_n25245_;
  assign new_n25250_ = ~new_n9281_;
  assign new_n25251_ = ~new_n8442_;
  assign new_n25252_ = ~new_n9280_;
  assign new_n25253_ = ~new_n8435_;
  assign new_n25254_ = ~new_n9278_;
  assign new_n25255_ = ~new_n8434_;
  assign new_n25256_ = ~new_n8434_ | ~new_n25219_;
  assign new_n25257_ = ~new_n8430_;
  assign new_n25258_ = ~new_n9277_;
  assign new_n25259_ = ~new_n8431_;
  assign new_n25260_ = ~new_n25471_ | ~new_n25470_;
  assign new_n25261_ = ~new_n25249_ | ~new_n25485_;
  assign new_n25262_ = ~new_n25235_ | ~new_n25496_;
  assign new_n25263_ = ~new_n25224_ | ~new_n25507_;
  assign new_n25264_ = ~new_n8454_;
  assign new_n25265_ = ~new_n25571_ | ~new_n25570_;
  assign new_n25266_ = ~new_n25585_ | ~new_n25584_;
  assign new_n25267_ = ~new_n25590_ | ~new_n25589_;
  assign new_n25268_ = ~new_n25606_ | ~new_n25605_;
  assign new_n25269_ = ~new_n25611_ | ~new_n25610_;
  assign new_n25270_ = ~new_n25616_ | ~new_n25615_;
  assign new_n25271_ = ~new_n25621_ | ~new_n25620_;
  assign new_n25272_ = ~new_n25626_ | ~new_n25625_;
  assign new_n25273_ = ~new_n25642_ | ~new_n25641_;
  assign new_n25274_ = ~new_n25647_ | ~new_n25646_;
  assign new_n25275_ = ~new_n25530_ | ~new_n25529_;
  assign new_n25276_ = ~new_n25539_ | ~new_n25538_;
  assign new_n25277_ = ~new_n25546_ | ~new_n25545_;
  assign new_n25278_ = ~new_n25550_ | ~new_n25549_;
  assign new_n25279_ = ~new_n25559_ | ~new_n25558_;
  assign new_n25280_ = ~new_n25580_ | ~new_n25579_;
  assign new_n25281_ = ~new_n25597_ | ~new_n25596_;
  assign new_n25282_ = ~new_n25601_ | ~new_n25600_;
  assign new_n25283_ = ~new_n25633_ | ~new_n25632_;
  assign new_n25284_ = ~new_n25637_ | ~new_n25636_;
  assign new_n25285_ = ~new_n25654_ | ~new_n25653_;
  assign new_n25286_ = new_n25521_ & new_n25362_;
  assign new_n25287_ = new_n25374_ & new_n25375_;
  assign new_n25288_ = new_n25183_ & new_n25182_;
  assign new_n25289_ = new_n25526_ & new_n25523_;
  assign new_n25290_ = new_n25195_ & new_n25532_ & new_n25531_;
  assign new_n25291_ = new_n25535_ & new_n25364_;
  assign new_n25292_ = new_n25404_ & new_n25175_;
  assign new_n25293_ = new_n25542_ & new_n25363_;
  assign new_n25294_ = new_n25203_ & new_n25552_ & new_n25551_;
  assign new_n25295_ = new_n25555_ & new_n25362_;
  assign new_n25296_ = new_n25391_ & new_n25176_;
  assign new_n25297_ = new_n25436_ & new_n25178_;
  assign new_n25298_ = new_n25460_ & new_n25180_;
  assign new_n25299_ = new_n25524_ & new_n25361_;
  assign new_n25300_ = new_n25475_ & new_n25476_;
  assign new_n25301_ = new_n25478_ & new_n25564_;
  assign new_n25302_ = new_n25475_ & new_n25476_;
  assign new_n25303_ = new_n25184_ & new_n25479_;
  assign new_n25304_ = ~new_n25568_ | ~new_n25567_;
  assign new_n25305_ = new_n25256_ & new_n25573_ & new_n25572_;
  assign new_n25306_ = new_n25576_ & new_n25361_;
  assign new_n25307_ = ~new_n25582_ | ~new_n25581_;
  assign new_n25308_ = ~new_n25587_ | ~new_n25586_;
  assign new_n25309_ = new_n25491_ & new_n25181_;
  assign new_n25310_ = new_n25593_ & new_n25360_;
  assign new_n25311_ = ~new_n25603_ | ~new_n25602_;
  assign new_n25312_ = ~new_n25608_ | ~new_n25607_;
  assign new_n25313_ = ~new_n25613_ | ~new_n25612_;
  assign new_n25314_ = ~new_n25618_ | ~new_n25617_;
  assign new_n25315_ = ~new_n25623_ | ~new_n25622_;
  assign new_n25316_ = new_n25502_ & new_n25179_;
  assign new_n25317_ = new_n25629_ & new_n25359_;
  assign new_n25318_ = ~new_n25639_ | ~new_n25638_;
  assign new_n25319_ = ~new_n25644_ | ~new_n25643_;
  assign new_n25320_ = new_n25513_ & new_n25177_;
  assign new_n25321_ = new_n25650_ & new_n25358_;
  assign new_n25322_ = new_n25528_ & new_n25527_;
  assign new_n25323_ = ~new_n25289_ | ~new_n25525_;
  assign new_n25324_ = new_n25537_ & new_n25536_;
  assign new_n25325_ = new_n25544_ & new_n25543_;
  assign new_n25326_ = new_n25548_ & new_n25547_;
  assign new_n25327_ = ~new_n25287_ | ~new_n25372_;
  assign new_n25328_ = new_n25557_ & new_n25556_;
  assign new_n25329_ = ~new_n9286_;
  assign new_n25330_ = ~new_n8432_;
  assign new_n25331_ = new_n25566_ & new_n25565_;
  assign new_n25332_ = ~new_n25300_ | ~new_n25473_;
  assign new_n25333_ = new_n25578_ & new_n25577_;
  assign new_n25334_ = ~new_n25467_ | ~new_n25466_;
  assign new_n25335_ = ~new_n25463_ | ~new_n25462_;
  assign new_n25336_ = new_n25595_ & new_n25594_;
  assign new_n25337_ = new_n25599_ & new_n25598_;
  assign new_n25338_ = ~new_n25453_ | ~new_n25452_;
  assign new_n25339_ = ~new_n25449_ | ~new_n25448_;
  assign new_n25340_ = ~new_n8770_;
  assign new_n25341_ = ~new_n8765_ | ~new_n25264_;
  assign new_n25342_ = ~new_n25519_ | ~new_n25445_ | ~new_n25353_;
  assign new_n25343_ = ~new_n8821_;
  assign new_n25344_ = ~new_n25443_ | ~new_n25442_;
  assign new_n25345_ = ~new_n25439_ | ~new_n25438_;
  assign new_n25346_ = new_n25631_ & new_n25630_;
  assign new_n25347_ = new_n25635_ & new_n25634_;
  assign new_n25348_ = ~new_n25429_ | ~new_n25428_;
  assign new_n25349_ = ~new_n25425_ | ~new_n25424_;
  assign new_n25350_ = ~new_n25421_ | ~new_n25420_;
  assign new_n25351_ = new_n25652_ & new_n25651_;
  assign new_n25352_ = ~new_n25301_ | ~new_n25332_;
  assign new_n25353_ = ~new_n25344_ | ~new_n25343_;
  assign new_n25354_ = ~new_n25341_ | ~new_n25340_;
  assign new_n25355_ = ~new_n25256_;
  assign new_n25356_ = ~new_n25203_;
  assign new_n25357_ = ~new_n25195_;
  assign new_n25358_ = ~new_n8797_ | ~new_n25223_;
  assign new_n25359_ = ~new_n8812_ | ~new_n25233_;
  assign new_n25360_ = ~new_n9283_ | ~new_n25247_;
  assign new_n25361_ = ~new_n9279_ | ~new_n25255_;
  assign new_n25362_ = ~new_n8773_ | ~new_n25202_;
  assign new_n25363_ = ~new_n8782_ | ~new_n25210_;
  assign new_n25364_ = ~new_n8788_ | ~new_n25194_;
  assign new_n25365_ = ~new_n25235_;
  assign new_n25366_ = ~new_n25249_;
  assign new_n25367_ = ~new_n25212_;
  assign new_n25368_ = ~new_n25224_;
  assign new_n25369_ = ~new_n25341_;
  assign new_n25370_ = ~new_n8455_ | ~new_n25341_;
  assign new_n25371_ = ~new_n25218_;
  assign new_n25372_ = ~new_n25286_ | ~new_n25218_;
  assign new_n25373_ = ~new_n25204_ | ~new_n25203_;
  assign new_n25374_ = ~new_n25373_ | ~new_n25201_;
  assign new_n25375_ = ~new_n8441_ | ~new_n25356_;
  assign new_n25376_ = ~new_n25327_;
  assign new_n25377_ = ~new_n8785_ | ~new_n25209_;
  assign new_n25378_ = ~new_n8448_ | ~new_n25206_;
  assign new_n25379_ = ~new_n8444_ | ~new_n25205_;
  assign new_n25380_ = ~new_n25367_ | ~new_n25363_;
  assign new_n25381_ = ~new_n25175_ | ~new_n25380_;
  assign new_n25382_ = ~new_n8779_ | ~new_n25211_;
  assign new_n25383_ = ~new_n8785_ | ~new_n25209_;
  assign new_n25384_ = ~new_n25182_ | ~new_n25327_;
  assign new_n25385_ = ~new_n25213_;
  assign new_n25386_ = ~new_n25216_;
  assign new_n25387_ = ~new_n8791_ | ~new_n25196_;
  assign new_n25388_ = ~new_n25196_ | ~new_n25195_;
  assign new_n25389_ = ~new_n8461_ | ~new_n25357_;
  assign new_n25390_ = ~new_n25323_;
  assign new_n25391_ = ~new_n8794_ | ~new_n25215_;
  assign new_n25392_ = ~new_n25391_ | ~new_n25224_;
  assign new_n25393_ = ~new_n25386_ | ~new_n25195_;
  assign new_n25394_ = ~new_n25291_ | ~new_n25393_;
  assign new_n25395_ = ~new_n25216_ | ~new_n25364_;
  assign new_n25396_ = ~new_n25290_ | ~new_n25395_;
  assign new_n25397_ = ~new_n25195_ | ~new_n25364_;
  assign new_n25398_ = ~new_n25382_ | ~new_n25327_;
  assign new_n25399_ = ~new_n25217_;
  assign new_n25400_ = ~new_n8444_ | ~new_n25205_;
  assign new_n25401_ = ~new_n25399_ | ~new_n25400_;
  assign new_n25402_ = ~new_n25293_ | ~new_n25401_;
  assign new_n25403_ = ~new_n25217_ | ~new_n25363_;
  assign new_n25404_ = ~new_n8785_ | ~new_n25209_;
  assign new_n25405_ = ~new_n25292_ | ~new_n25403_;
  assign new_n25406_ = ~new_n8444_ | ~new_n25205_;
  assign new_n25407_ = ~new_n25363_ | ~new_n25406_;
  assign new_n25408_ = ~new_n25382_ | ~new_n25212_;
  assign new_n25409_ = ~new_n25371_ | ~new_n25203_;
  assign new_n25410_ = ~new_n25295_ | ~new_n25409_;
  assign new_n25411_ = ~new_n25218_ | ~new_n25362_;
  assign new_n25412_ = ~new_n25294_ | ~new_n25411_;
  assign new_n25413_ = ~new_n25362_ | ~new_n25203_;
  assign new_n25414_ = ~new_n8800_ | ~new_n25222_;
  assign new_n25415_ = ~new_n8440_ | ~new_n25220_;
  assign new_n25416_ = ~new_n8439_ | ~new_n25221_;
  assign new_n25417_ = ~new_n25368_ | ~new_n25176_;
  assign new_n25418_ = ~new_n25177_ | ~new_n25417_;
  assign new_n25419_ = ~new_n8800_ | ~new_n25222_;
  assign new_n25420_ = ~new_n25296_ | ~new_n25323_;
  assign new_n25421_ = ~new_n25419_ | ~new_n25418_;
  assign new_n25422_ = ~new_n25350_;
  assign new_n25423_ = ~new_n8803_ | ~new_n25226_;
  assign new_n25424_ = ~new_n25423_ | ~new_n25350_;
  assign new_n25425_ = ~new_n8449_ | ~new_n25225_;
  assign new_n25426_ = ~new_n25349_;
  assign new_n25427_ = ~new_n8806_ | ~new_n25228_;
  assign new_n25428_ = ~new_n25427_ | ~new_n25349_;
  assign new_n25429_ = ~new_n8457_ | ~new_n25227_;
  assign new_n25430_ = ~new_n25348_;
  assign new_n25431_ = ~new_n8815_ | ~new_n25232_;
  assign new_n25432_ = ~new_n8450_ | ~new_n25229_;
  assign new_n25433_ = ~new_n8451_ | ~new_n25230_;
  assign new_n25434_ = ~new_n25365_ | ~new_n25178_;
  assign new_n25435_ = ~new_n25179_ | ~new_n25434_;
  assign new_n25436_ = ~new_n8809_ | ~new_n25234_;
  assign new_n25437_ = ~new_n8815_ | ~new_n25232_;
  assign new_n25438_ = ~new_n25297_ | ~new_n25348_;
  assign new_n25439_ = ~new_n25437_ | ~new_n25435_;
  assign new_n25440_ = ~new_n25345_;
  assign new_n25441_ = ~new_n8818_ | ~new_n25237_;
  assign new_n25442_ = ~new_n25441_ | ~new_n25345_;
  assign new_n25443_ = ~new_n8446_ | ~new_n25236_;
  assign new_n25444_ = ~new_n25344_;
  assign new_n25445_ = ~new_n8459_ | ~new_n25344_;
  assign new_n25446_ = ~new_n25342_;
  assign new_n25447_ = ~new_n8823_ | ~new_n25240_;
  assign new_n25448_ = ~new_n25447_ | ~new_n25342_;
  assign new_n25449_ = ~new_n8458_ | ~new_n25239_;
  assign new_n25450_ = ~new_n25339_;
  assign new_n25451_ = ~new_n9285_ | ~new_n25242_;
  assign new_n25452_ = ~new_n25451_ | ~new_n25339_;
  assign new_n25453_ = ~new_n8453_ | ~new_n25241_;
  assign new_n25454_ = ~new_n25338_;
  assign new_n25455_ = ~new_n9282_ | ~new_n25246_;
  assign new_n25456_ = ~new_n8443_ | ~new_n25243_;
  assign new_n25457_ = ~new_n8438_ | ~new_n25244_;
  assign new_n25458_ = ~new_n25366_ | ~new_n25180_;
  assign new_n25459_ = ~new_n25181_ | ~new_n25458_;
  assign new_n25460_ = ~new_n9284_ | ~new_n25248_;
  assign new_n25461_ = ~new_n9282_ | ~new_n25246_;
  assign new_n25462_ = ~new_n25298_ | ~new_n25338_;
  assign new_n25463_ = ~new_n25461_ | ~new_n25459_;
  assign new_n25464_ = ~new_n25335_;
  assign new_n25465_ = ~new_n9281_ | ~new_n25251_;
  assign new_n25466_ = ~new_n25465_ | ~new_n25335_;
  assign new_n25467_ = ~new_n8442_ | ~new_n25250_;
  assign new_n25468_ = ~new_n25334_;
  assign new_n25469_ = ~new_n9280_ | ~new_n25253_;
  assign new_n25470_ = ~new_n25469_ | ~new_n25334_;
  assign new_n25471_ = ~new_n8435_ | ~new_n25252_;
  assign new_n25472_ = ~new_n25260_;
  assign new_n25473_ = ~new_n25299_ | ~new_n25260_;
  assign new_n25474_ = ~new_n25257_ | ~new_n25256_;
  assign new_n25475_ = ~new_n25474_ | ~new_n25254_;
  assign new_n25476_ = ~new_n8430_ | ~new_n25355_;
  assign new_n25477_ = ~new_n25332_;
  assign new_n25478_ = ~new_n9277_ | ~new_n25259_;
  assign new_n25479_ = ~new_n8431_ | ~new_n25258_;
  assign new_n25480_ = ~new_n25472_ | ~new_n25256_;
  assign new_n25481_ = ~new_n25306_ | ~new_n25480_;
  assign new_n25482_ = ~new_n25260_ | ~new_n25361_;
  assign new_n25483_ = ~new_n25305_ | ~new_n25482_;
  assign new_n25484_ = ~new_n25361_ | ~new_n25256_;
  assign new_n25485_ = ~new_n25460_ | ~new_n25338_;
  assign new_n25486_ = ~new_n25261_;
  assign new_n25487_ = ~new_n8438_ | ~new_n25244_;
  assign new_n25488_ = ~new_n25486_ | ~new_n25487_;
  assign new_n25489_ = ~new_n25310_ | ~new_n25488_;
  assign new_n25490_ = ~new_n25261_ | ~new_n25360_;
  assign new_n25491_ = ~new_n9282_ | ~new_n25246_;
  assign new_n25492_ = ~new_n25309_ | ~new_n25490_;
  assign new_n25493_ = ~new_n8438_ | ~new_n25244_;
  assign new_n25494_ = ~new_n25360_ | ~new_n25493_;
  assign new_n25495_ = ~new_n25460_ | ~new_n25249_;
  assign new_n25496_ = ~new_n25436_ | ~new_n25348_;
  assign new_n25497_ = ~new_n25262_;
  assign new_n25498_ = ~new_n8451_ | ~new_n25230_;
  assign new_n25499_ = ~new_n25497_ | ~new_n25498_;
  assign new_n25500_ = ~new_n25317_ | ~new_n25499_;
  assign new_n25501_ = ~new_n25262_ | ~new_n25359_;
  assign new_n25502_ = ~new_n8815_ | ~new_n25232_;
  assign new_n25503_ = ~new_n25316_ | ~new_n25501_;
  assign new_n25504_ = ~new_n8451_ | ~new_n25230_;
  assign new_n25505_ = ~new_n25359_ | ~new_n25504_;
  assign new_n25506_ = ~new_n25436_ | ~new_n25235_;
  assign new_n25507_ = ~new_n25391_ | ~new_n25323_;
  assign new_n25508_ = ~new_n25263_;
  assign new_n25509_ = ~new_n8439_ | ~new_n25221_;
  assign new_n25510_ = ~new_n25508_ | ~new_n25509_;
  assign new_n25511_ = ~new_n25321_ | ~new_n25510_;
  assign new_n25512_ = ~new_n25263_ | ~new_n25358_;
  assign new_n25513_ = ~new_n8800_ | ~new_n25222_;
  assign new_n25514_ = ~new_n25320_ | ~new_n25512_;
  assign new_n25515_ = ~new_n8439_ | ~new_n25221_;
  assign new_n25516_ = ~new_n25358_ | ~new_n25515_;
  assign new_n25517_ = ~new_n8454_ | ~new_n25199_;
  assign new_n25518_ = ~new_n8455_ | ~new_n25340_;
  assign new_n25519_ = ~new_n8459_ | ~new_n25343_;
  assign new_n25520_ = ~new_n25303_ | ~new_n25302_ | ~new_n25473_;
  assign new_n25521_ = ~new_n8776_ | ~new_n25204_;
  assign new_n25522_ = ~new_n8791_ | ~new_n25389_;
  assign new_n25523_ = ~new_n25522_ | ~new_n25388_;
  assign new_n25524_ = ~new_n9278_ | ~new_n25257_;
  assign new_n25525_ = ~new_n25288_ | ~new_n25327_;
  assign new_n25526_ = ~new_n25385_ | ~new_n25183_;
  assign new_n25527_ = ~new_n8794_ | ~new_n25215_;
  assign new_n25528_ = ~new_n8460_ | ~new_n25214_;
  assign new_n25529_ = ~new_n25392_ | ~new_n25323_;
  assign new_n25530_ = ~new_n25390_ | ~new_n25322_;
  assign new_n25531_ = ~new_n8791_ | ~new_n25196_;
  assign new_n25532_ = ~new_n8461_ | ~new_n25197_;
  assign new_n25533_ = ~new_n8791_ | ~new_n25196_;
  assign new_n25534_ = ~new_n8461_ | ~new_n25197_;
  assign new_n25535_ = ~new_n25534_ | ~new_n25533_;
  assign new_n25536_ = ~new_n8788_ | ~new_n25194_;
  assign new_n25537_ = ~new_n8447_ | ~new_n25208_;
  assign new_n25538_ = ~new_n25397_ | ~new_n25216_;
  assign new_n25539_ = ~new_n25324_ | ~new_n25386_;
  assign new_n25540_ = ~new_n8785_ | ~new_n25209_;
  assign new_n25541_ = ~new_n8448_ | ~new_n25206_;
  assign new_n25542_ = ~new_n25541_ | ~new_n25540_;
  assign new_n25543_ = ~new_n8782_ | ~new_n25210_;
  assign new_n25544_ = ~new_n8444_ | ~new_n25205_;
  assign new_n25545_ = ~new_n25407_ | ~new_n25217_;
  assign new_n25546_ = ~new_n25325_ | ~new_n25399_;
  assign new_n25547_ = ~new_n8779_ | ~new_n25211_;
  assign new_n25548_ = ~new_n8437_ | ~new_n25207_;
  assign new_n25549_ = ~new_n25408_ | ~new_n25327_;
  assign new_n25550_ = ~new_n25376_ | ~new_n25326_;
  assign new_n25551_ = ~new_n8776_ | ~new_n25204_;
  assign new_n25552_ = ~new_n8441_ | ~new_n25201_;
  assign new_n25553_ = ~new_n8776_ | ~new_n25204_;
  assign new_n25554_ = ~new_n8441_ | ~new_n25201_;
  assign new_n25555_ = ~new_n25554_ | ~new_n25553_;
  assign new_n25556_ = ~new_n8773_ | ~new_n25202_;
  assign new_n25557_ = ~new_n8445_ | ~new_n25198_;
  assign new_n25558_ = ~new_n25413_ | ~new_n25218_;
  assign new_n25559_ = ~new_n25328_ | ~new_n25371_;
  assign new_n25560_ = ~new_n9286_ | ~new_n25330_;
  assign new_n25561_ = ~new_n8432_ | ~new_n25329_;
  assign new_n25562_ = ~new_n9286_ | ~new_n25330_;
  assign new_n25563_ = ~new_n8432_ | ~new_n25329_;
  assign new_n25564_ = ~new_n25563_ | ~new_n25562_;
  assign new_n25565_ = ~new_n25258_ | ~new_n8431_ | ~new_n25564_;
  assign new_n25566_ = ~new_n9277_ | ~new_n25184_ | ~new_n25259_;
  assign new_n25567_ = ~new_n9277_ | ~new_n25259_;
  assign new_n25568_ = ~new_n8431_ | ~new_n25258_;
  assign new_n25569_ = ~new_n25304_;
  assign new_n25570_ = ~new_n25477_ | ~new_n25569_;
  assign new_n25571_ = ~new_n25304_ | ~new_n25332_;
  assign new_n25572_ = ~new_n9278_ | ~new_n25257_;
  assign new_n25573_ = ~new_n8430_ | ~new_n25254_;
  assign new_n25574_ = ~new_n9278_ | ~new_n25257_;
  assign new_n25575_ = ~new_n8430_ | ~new_n25254_;
  assign new_n25576_ = ~new_n25575_ | ~new_n25574_;
  assign new_n25577_ = ~new_n9279_ | ~new_n25255_;
  assign new_n25578_ = ~new_n8434_ | ~new_n25219_;
  assign new_n25579_ = ~new_n25484_ | ~new_n25260_;
  assign new_n25580_ = ~new_n25333_ | ~new_n25472_;
  assign new_n25581_ = ~new_n9280_ | ~new_n25253_;
  assign new_n25582_ = ~new_n8435_ | ~new_n25252_;
  assign new_n25583_ = ~new_n25307_;
  assign new_n25584_ = ~new_n25468_ | ~new_n25583_;
  assign new_n25585_ = ~new_n25307_ | ~new_n25334_;
  assign new_n25586_ = ~new_n9281_ | ~new_n25251_;
  assign new_n25587_ = ~new_n8442_ | ~new_n25250_;
  assign new_n25588_ = ~new_n25308_;
  assign new_n25589_ = ~new_n25464_ | ~new_n25588_;
  assign new_n25590_ = ~new_n25308_ | ~new_n25335_;
  assign new_n25591_ = ~new_n9282_ | ~new_n25246_;
  assign new_n25592_ = ~new_n8443_ | ~new_n25243_;
  assign new_n25593_ = ~new_n25592_ | ~new_n25591_;
  assign new_n25594_ = ~new_n9283_ | ~new_n25247_;
  assign new_n25595_ = ~new_n8438_ | ~new_n25244_;
  assign new_n25596_ = ~new_n25494_ | ~new_n25261_;
  assign new_n25597_ = ~new_n25336_ | ~new_n25486_;
  assign new_n25598_ = ~new_n9284_ | ~new_n25248_;
  assign new_n25599_ = ~new_n8452_ | ~new_n25245_;
  assign new_n25600_ = ~new_n25495_ | ~new_n25338_;
  assign new_n25601_ = ~new_n25454_ | ~new_n25337_;
  assign new_n25602_ = ~new_n9285_ | ~new_n25242_;
  assign new_n25603_ = ~new_n8453_ | ~new_n25241_;
  assign new_n25604_ = ~new_n25311_;
  assign new_n25605_ = ~new_n25450_ | ~new_n25604_;
  assign new_n25606_ = ~new_n25311_ | ~new_n25339_;
  assign new_n25607_ = ~new_n8770_ | ~new_n25200_;
  assign new_n25608_ = ~new_n8455_ | ~new_n25340_;
  assign new_n25609_ = ~new_n25312_;
  assign new_n25610_ = ~new_n25369_ | ~new_n25609_;
  assign new_n25611_ = ~new_n25312_ | ~new_n25341_;
  assign new_n25612_ = ~new_n8823_ | ~new_n25240_;
  assign new_n25613_ = ~new_n8458_ | ~new_n25239_;
  assign new_n25614_ = ~new_n25313_;
  assign new_n25615_ = ~new_n25446_ | ~new_n25614_;
  assign new_n25616_ = ~new_n25313_ | ~new_n25342_;
  assign new_n25617_ = ~new_n8821_ | ~new_n25238_;
  assign new_n25618_ = ~new_n8459_ | ~new_n25343_;
  assign new_n25619_ = ~new_n25314_;
  assign new_n25620_ = ~new_n25444_ | ~new_n25619_;
  assign new_n25621_ = ~new_n25314_ | ~new_n25344_;
  assign new_n25622_ = ~new_n8818_ | ~new_n25237_;
  assign new_n25623_ = ~new_n8446_ | ~new_n25236_;
  assign new_n25624_ = ~new_n25315_;
  assign new_n25625_ = ~new_n25440_ | ~new_n25624_;
  assign new_n25626_ = ~new_n25315_ | ~new_n25345_;
  assign new_n25627_ = ~new_n8815_ | ~new_n25232_;
  assign new_n25628_ = ~new_n8450_ | ~new_n25229_;
  assign new_n25629_ = ~new_n25628_ | ~new_n25627_;
  assign new_n25630_ = ~new_n8812_ | ~new_n25233_;
  assign new_n25631_ = ~new_n8451_ | ~new_n25230_;
  assign new_n25632_ = ~new_n25505_ | ~new_n25262_;
  assign new_n25633_ = ~new_n25346_ | ~new_n25497_;
  assign new_n25634_ = ~new_n8809_ | ~new_n25234_;
  assign new_n25635_ = ~new_n8456_ | ~new_n25231_;
  assign new_n25636_ = ~new_n25506_ | ~new_n25348_;
  assign new_n25637_ = ~new_n25430_ | ~new_n25347_;
  assign new_n25638_ = ~new_n8806_ | ~new_n25228_;
  assign new_n25639_ = ~new_n8457_ | ~new_n25227_;
  assign new_n25640_ = ~new_n25318_;
  assign new_n25641_ = ~new_n25426_ | ~new_n25640_;
  assign new_n25642_ = ~new_n25318_ | ~new_n25349_;
  assign new_n25643_ = ~new_n8803_ | ~new_n25226_;
  assign new_n25644_ = ~new_n8449_ | ~new_n25225_;
  assign new_n25645_ = ~new_n25319_;
  assign new_n25646_ = ~new_n25422_ | ~new_n25645_;
  assign new_n25647_ = ~new_n25319_ | ~new_n25350_;
  assign new_n25648_ = ~new_n8800_ | ~new_n25222_;
  assign new_n25649_ = ~new_n8440_ | ~new_n25220_;
  assign new_n25650_ = ~new_n25649_ | ~new_n25648_;
  assign new_n25651_ = ~new_n8797_ | ~new_n25223_;
  assign new_n25652_ = ~new_n8439_ | ~new_n25221_;
  assign new_n25653_ = ~new_n25516_ | ~new_n25263_;
  assign new_n25654_ = ~new_n25351_ | ~new_n25508_;
  assign new_n25655_ = ~new_n25825_ | ~new_n25829_;
  assign new_n25656_ = ~new_n25658_ | ~new_n25830_;
  assign new_n25657_ = ~pi651;
  assign new_n25658_ = ~pi651 | ~new_n25697_;
  assign new_n25659_ = ~pi652;
  assign new_n25660_ = ~new_n8769_;
  assign new_n25661_ = ~pi653;
  assign new_n25662_ = ~new_n8772_;
  assign new_n25663_ = ~pi654;
  assign new_n25664_ = ~new_n8775_;
  assign new_n25665_ = ~pi655;
  assign new_n25666_ = ~new_n8778_;
  assign new_n25667_ = ~pi656;
  assign new_n25668_ = ~new_n8781_;
  assign new_n25669_ = ~pi657;
  assign new_n25670_ = ~new_n8784_;
  assign new_n25671_ = ~pi658;
  assign new_n25672_ = ~new_n8787_;
  assign new_n25673_ = ~pi659;
  assign new_n25674_ = ~new_n8790_;
  assign new_n25675_ = ~pi660;
  assign new_n25676_ = ~new_n8793_;
  assign new_n25677_ = ~pi661;
  assign new_n25678_ = ~new_n8796_;
  assign new_n25679_ = ~pi662;
  assign new_n25680_ = ~new_n8799_;
  assign new_n25681_ = ~pi663;
  assign new_n25682_ = ~new_n8802_;
  assign new_n25683_ = ~pi664;
  assign new_n25684_ = ~new_n8805_;
  assign new_n25685_ = ~pi665;
  assign new_n25686_ = ~new_n8808_;
  assign new_n25687_ = ~new_n25808_ | ~new_n25807_;
  assign new_n25688_ = ~pi666;
  assign new_n25689_ = ~new_n8811_;
  assign new_n25690_ = ~pi667;
  assign new_n25691_ = ~new_n8814_;
  assign new_n25692_ = ~pi668;
  assign new_n25693_ = ~new_n8817_;
  assign new_n25694_ = ~pi669;
  assign new_n25695_ = ~new_n8820_;
  assign new_n25696_ = ~new_n25820_ | ~new_n25819_;
  assign new_n25697_ = ~new_n8764_;
  assign new_n25698_ = ~new_n25835_ | ~new_n25834_;
  assign new_n25699_ = ~new_n25840_ | ~new_n25839_;
  assign new_n25700_ = ~new_n25845_ | ~new_n25844_;
  assign new_n25701_ = ~new_n25850_ | ~new_n25849_;
  assign new_n25702_ = ~new_n25855_ | ~new_n25854_;
  assign new_n25703_ = ~new_n25860_ | ~new_n25859_;
  assign new_n25704_ = ~new_n25865_ | ~new_n25864_;
  assign new_n25705_ = ~new_n25870_ | ~new_n25869_;
  assign new_n25706_ = ~new_n25875_ | ~new_n25874_;
  assign new_n25707_ = ~new_n25885_ | ~new_n25884_;
  assign new_n25708_ = ~new_n25890_ | ~new_n25889_;
  assign new_n25709_ = ~new_n25895_ | ~new_n25894_;
  assign new_n25710_ = ~new_n25900_ | ~new_n25899_;
  assign new_n25711_ = ~new_n25905_ | ~new_n25904_;
  assign new_n25712_ = ~new_n25910_ | ~new_n25909_;
  assign new_n25713_ = ~new_n25915_ | ~new_n25914_;
  assign new_n25714_ = ~new_n25920_ | ~new_n25919_;
  assign new_n25715_ = ~new_n25925_ | ~new_n25924_;
  assign new_n25716_ = ~new_n25832_ | ~new_n25831_;
  assign new_n25717_ = ~new_n25837_ | ~new_n25836_;
  assign new_n25718_ = ~new_n25842_ | ~new_n25841_;
  assign new_n25719_ = ~new_n25847_ | ~new_n25846_;
  assign new_n25720_ = ~new_n25852_ | ~new_n25851_;
  assign new_n25721_ = ~new_n25857_ | ~new_n25856_;
  assign new_n25722_ = ~new_n25862_ | ~new_n25861_;
  assign new_n25723_ = ~new_n25867_ | ~new_n25866_;
  assign new_n25724_ = ~new_n25872_ | ~new_n25871_;
  assign new_n25725_ = new_n25828_ & new_n25877_ & new_n25876_;
  assign new_n25726_ = new_n25824_ & new_n25880_;
  assign new_n25727_ = ~new_n25882_ | ~new_n25881_;
  assign new_n25728_ = ~new_n25887_ | ~new_n25886_;
  assign new_n25729_ = ~new_n25892_ | ~new_n25891_;
  assign new_n25730_ = ~new_n25897_ | ~new_n25896_;
  assign new_n25731_ = ~new_n25902_ | ~new_n25901_;
  assign new_n25732_ = ~new_n25907_ | ~new_n25906_;
  assign new_n25733_ = ~new_n25912_ | ~new_n25911_;
  assign new_n25734_ = ~new_n25917_ | ~new_n25916_;
  assign new_n25735_ = ~new_n25922_ | ~new_n25921_;
  assign new_n25736_ = ~new_n25784_ | ~new_n25783_;
  assign new_n25737_ = ~new_n25780_ | ~new_n25779_;
  assign new_n25738_ = ~new_n25776_ | ~new_n25775_;
  assign new_n25739_ = ~new_n25772_ | ~new_n25771_;
  assign new_n25740_ = ~new_n25768_ | ~new_n25767_;
  assign new_n25741_ = ~new_n25764_ | ~new_n25763_;
  assign new_n25742_ = ~new_n25760_ | ~new_n25759_;
  assign new_n25743_ = ~new_n25756_ | ~new_n25755_;
  assign new_n25744_ = ~pi670;
  assign new_n25745_ = ~new_n8757_;
  assign new_n25746_ = ~new_n25816_ | ~new_n25815_;
  assign new_n25747_ = ~new_n25812_ | ~new_n25811_;
  assign new_n25748_ = ~new_n25804_ | ~new_n25803_;
  assign new_n25749_ = ~new_n25800_ | ~new_n25799_;
  assign new_n25750_ = ~new_n25796_ | ~new_n25795_;
  assign new_n25751_ = ~new_n25792_ | ~new_n25791_;
  assign new_n25752_ = ~new_n25788_ | ~new_n25787_;
  assign new_n25753_ = ~new_n25658_;
  assign new_n25754_ = ~pi652 | ~new_n25753_;
  assign new_n25755_ = ~new_n8769_ | ~new_n25754_;
  assign new_n25756_ = ~new_n25658_ | ~new_n25659_;
  assign new_n25757_ = ~new_n25743_;
  assign new_n25758_ = ~pi653 | ~new_n25662_;
  assign new_n25759_ = ~new_n25758_ | ~new_n25743_;
  assign new_n25760_ = ~new_n8772_ | ~new_n25661_;
  assign new_n25761_ = ~new_n25742_;
  assign new_n25762_ = ~pi654 | ~new_n25664_;
  assign new_n25763_ = ~new_n25762_ | ~new_n25742_;
  assign new_n25764_ = ~new_n8775_ | ~new_n25663_;
  assign new_n25765_ = ~new_n25741_;
  assign new_n25766_ = ~pi655 | ~new_n25666_;
  assign new_n25767_ = ~new_n25766_ | ~new_n25741_;
  assign new_n25768_ = ~new_n8778_ | ~new_n25665_;
  assign new_n25769_ = ~new_n25740_;
  assign new_n25770_ = ~pi656 | ~new_n25668_;
  assign new_n25771_ = ~new_n25770_ | ~new_n25740_;
  assign new_n25772_ = ~new_n8781_ | ~new_n25667_;
  assign new_n25773_ = ~new_n25739_;
  assign new_n25774_ = ~pi657 | ~new_n25670_;
  assign new_n25775_ = ~new_n25774_ | ~new_n25739_;
  assign new_n25776_ = ~new_n8784_ | ~new_n25669_;
  assign new_n25777_ = ~new_n25738_;
  assign new_n25778_ = ~pi658 | ~new_n25672_;
  assign new_n25779_ = ~new_n25778_ | ~new_n25738_;
  assign new_n25780_ = ~new_n8787_ | ~new_n25671_;
  assign new_n25781_ = ~new_n25737_;
  assign new_n25782_ = ~pi659 | ~new_n25674_;
  assign new_n25783_ = ~new_n25782_ | ~new_n25737_;
  assign new_n25784_ = ~new_n8790_ | ~new_n25673_;
  assign new_n25785_ = ~new_n25736_;
  assign new_n25786_ = ~pi660 | ~new_n25676_;
  assign new_n25787_ = ~new_n25786_ | ~new_n25736_;
  assign new_n25788_ = ~new_n8793_ | ~new_n25675_;
  assign new_n25789_ = ~new_n25752_;
  assign new_n25790_ = ~pi661 | ~new_n25678_;
  assign new_n25791_ = ~new_n25790_ | ~new_n25752_;
  assign new_n25792_ = ~new_n8796_ | ~new_n25677_;
  assign new_n25793_ = ~new_n25751_;
  assign new_n25794_ = ~pi662 | ~new_n25680_;
  assign new_n25795_ = ~new_n25794_ | ~new_n25751_;
  assign new_n25796_ = ~new_n8799_ | ~new_n25679_;
  assign new_n25797_ = ~new_n25750_;
  assign new_n25798_ = ~pi663 | ~new_n25682_;
  assign new_n25799_ = ~new_n25798_ | ~new_n25750_;
  assign new_n25800_ = ~new_n8802_ | ~new_n25681_;
  assign new_n25801_ = ~new_n25749_;
  assign new_n25802_ = ~pi664 | ~new_n25684_;
  assign new_n25803_ = ~new_n25802_ | ~new_n25749_;
  assign new_n25804_ = ~new_n8805_ | ~new_n25683_;
  assign new_n25805_ = ~new_n25748_;
  assign new_n25806_ = ~pi665 | ~new_n25686_;
  assign new_n25807_ = ~new_n25806_ | ~new_n25748_;
  assign new_n25808_ = ~new_n8808_ | ~new_n25685_;
  assign new_n25809_ = ~new_n25687_;
  assign new_n25810_ = ~pi666 | ~new_n25809_;
  assign new_n25811_ = ~new_n8811_ | ~new_n25810_;
  assign new_n25812_ = ~new_n25687_ | ~new_n25688_;
  assign new_n25813_ = ~new_n25747_;
  assign new_n25814_ = ~pi667 | ~new_n25691_;
  assign new_n25815_ = ~new_n25814_ | ~new_n25747_;
  assign new_n25816_ = ~new_n8814_ | ~new_n25690_;
  assign new_n25817_ = ~new_n25746_;
  assign new_n25818_ = ~pi668 | ~new_n25693_;
  assign new_n25819_ = ~new_n25818_ | ~new_n25746_;
  assign new_n25820_ = ~new_n8817_ | ~new_n25692_;
  assign new_n25821_ = ~new_n25696_;
  assign new_n25822_ = ~new_n8820_ | ~new_n25694_;
  assign new_n25823_ = ~new_n25821_ | ~new_n25822_;
  assign new_n25824_ = ~pi669 | ~new_n25695_;
  assign new_n25825_ = ~new_n25726_ | ~new_n25823_;
  assign new_n25826_ = ~pi669 | ~new_n25695_;
  assign new_n25827_ = ~new_n25826_ | ~new_n25696_;
  assign new_n25828_ = ~new_n8820_ | ~new_n25694_;
  assign new_n25829_ = ~new_n25725_ | ~new_n25827_;
  assign new_n25830_ = ~new_n8764_ | ~new_n25657_;
  assign new_n25831_ = ~pi660 | ~new_n25676_;
  assign new_n25832_ = ~new_n8793_ | ~new_n25675_;
  assign new_n25833_ = ~new_n25716_;
  assign new_n25834_ = ~new_n25785_ | ~new_n25833_;
  assign new_n25835_ = ~new_n25716_ | ~new_n25736_;
  assign new_n25836_ = ~pi659 | ~new_n25674_;
  assign new_n25837_ = ~new_n8790_ | ~new_n25673_;
  assign new_n25838_ = ~new_n25717_;
  assign new_n25839_ = ~new_n25781_ | ~new_n25838_;
  assign new_n25840_ = ~new_n25717_ | ~new_n25737_;
  assign new_n25841_ = ~pi658 | ~new_n25672_;
  assign new_n25842_ = ~new_n8787_ | ~new_n25671_;
  assign new_n25843_ = ~new_n25718_;
  assign new_n25844_ = ~new_n25777_ | ~new_n25843_;
  assign new_n25845_ = ~new_n25718_ | ~new_n25738_;
  assign new_n25846_ = ~pi657 | ~new_n25670_;
  assign new_n25847_ = ~new_n8784_ | ~new_n25669_;
  assign new_n25848_ = ~new_n25719_;
  assign new_n25849_ = ~new_n25773_ | ~new_n25848_;
  assign new_n25850_ = ~new_n25719_ | ~new_n25739_;
  assign new_n25851_ = ~pi656 | ~new_n25668_;
  assign new_n25852_ = ~new_n8781_ | ~new_n25667_;
  assign new_n25853_ = ~new_n25720_;
  assign new_n25854_ = ~new_n25769_ | ~new_n25853_;
  assign new_n25855_ = ~new_n25720_ | ~new_n25740_;
  assign new_n25856_ = ~pi655 | ~new_n25666_;
  assign new_n25857_ = ~new_n8778_ | ~new_n25665_;
  assign new_n25858_ = ~new_n25721_;
  assign new_n25859_ = ~new_n25765_ | ~new_n25858_;
  assign new_n25860_ = ~new_n25721_ | ~new_n25741_;
  assign new_n25861_ = ~pi654 | ~new_n25664_;
  assign new_n25862_ = ~new_n8775_ | ~new_n25663_;
  assign new_n25863_ = ~new_n25722_;
  assign new_n25864_ = ~new_n25761_ | ~new_n25863_;
  assign new_n25865_ = ~new_n25722_ | ~new_n25742_;
  assign new_n25866_ = ~pi653 | ~new_n25662_;
  assign new_n25867_ = ~new_n8772_ | ~new_n25661_;
  assign new_n25868_ = ~new_n25723_;
  assign new_n25869_ = ~new_n25757_ | ~new_n25868_;
  assign new_n25870_ = ~new_n25723_ | ~new_n25743_;
  assign new_n25871_ = ~new_n25753_ | ~new_n25659_;
  assign new_n25872_ = ~pi652 | ~new_n25658_;
  assign new_n25873_ = ~new_n25724_;
  assign new_n25874_ = ~new_n25873_ | ~new_n8769_;
  assign new_n25875_ = ~new_n25724_ | ~new_n25660_;
  assign new_n25876_ = ~pi670 | ~new_n25745_;
  assign new_n25877_ = ~new_n8757_ | ~new_n25744_;
  assign new_n25878_ = ~pi670 | ~new_n25745_;
  assign new_n25879_ = ~new_n8757_ | ~new_n25744_;
  assign new_n25880_ = ~new_n25879_ | ~new_n25878_;
  assign new_n25881_ = ~pi669 | ~new_n25695_;
  assign new_n25882_ = ~new_n8820_ | ~new_n25694_;
  assign new_n25883_ = ~new_n25727_;
  assign new_n25884_ = ~new_n25883_ | ~new_n25821_;
  assign new_n25885_ = ~new_n25727_ | ~new_n25696_;
  assign new_n25886_ = ~pi668 | ~new_n25693_;
  assign new_n25887_ = ~new_n8817_ | ~new_n25692_;
  assign new_n25888_ = ~new_n25728_;
  assign new_n25889_ = ~new_n25817_ | ~new_n25888_;
  assign new_n25890_ = ~new_n25728_ | ~new_n25746_;
  assign new_n25891_ = ~pi667 | ~new_n25691_;
  assign new_n25892_ = ~new_n8814_ | ~new_n25690_;
  assign new_n25893_ = ~new_n25729_;
  assign new_n25894_ = ~new_n25813_ | ~new_n25893_;
  assign new_n25895_ = ~new_n25729_ | ~new_n25747_;
  assign new_n25896_ = ~new_n8811_ | ~new_n25688_;
  assign new_n25897_ = ~pi666 | ~new_n25689_;
  assign new_n25898_ = ~new_n25730_;
  assign new_n25899_ = ~new_n25898_ | ~new_n25809_;
  assign new_n25900_ = ~new_n25730_ | ~new_n25687_;
  assign new_n25901_ = ~pi665 | ~new_n25686_;
  assign new_n25902_ = ~new_n8808_ | ~new_n25685_;
  assign new_n25903_ = ~new_n25731_;
  assign new_n25904_ = ~new_n25805_ | ~new_n25903_;
  assign new_n25905_ = ~new_n25731_ | ~new_n25748_;
  assign new_n25906_ = ~pi664 | ~new_n25684_;
  assign new_n25907_ = ~new_n8805_ | ~new_n25683_;
  assign new_n25908_ = ~new_n25732_;
  assign new_n25909_ = ~new_n25801_ | ~new_n25908_;
  assign new_n25910_ = ~new_n25732_ | ~new_n25749_;
  assign new_n25911_ = ~pi663 | ~new_n25682_;
  assign new_n25912_ = ~new_n8802_ | ~new_n25681_;
  assign new_n25913_ = ~new_n25733_;
  assign new_n25914_ = ~new_n25797_ | ~new_n25913_;
  assign new_n25915_ = ~new_n25733_ | ~new_n25750_;
  assign new_n25916_ = ~pi662 | ~new_n25680_;
  assign new_n25917_ = ~new_n8799_ | ~new_n25679_;
  assign new_n25918_ = ~new_n25734_;
  assign new_n25919_ = ~new_n25793_ | ~new_n25918_;
  assign new_n25920_ = ~new_n25734_ | ~new_n25751_;
  assign new_n25921_ = ~pi661 | ~new_n25678_;
  assign new_n25922_ = ~new_n8796_ | ~new_n25677_;
  assign new_n25923_ = ~new_n25735_;
  assign new_n25924_ = ~new_n25789_ | ~new_n25923_;
  assign new_n25925_ = ~new_n25735_ | ~new_n25752_;
  assign new_n25926_ = ~new_n26096_ | ~new_n26100_;
  assign new_n25927_ = ~new_n25929_ | ~new_n26101_;
  assign new_n25928_ = ~pi619;
  assign new_n25929_ = ~pi619 | ~new_n25968_;
  assign new_n25930_ = ~pi620;
  assign new_n25931_ = ~new_n8769_;
  assign new_n25932_ = ~pi621;
  assign new_n25933_ = ~new_n8772_;
  assign new_n25934_ = ~pi622;
  assign new_n25935_ = ~new_n8775_;
  assign new_n25936_ = ~pi623;
  assign new_n25937_ = ~new_n8778_;
  assign new_n25938_ = ~pi624;
  assign new_n25939_ = ~new_n8781_;
  assign new_n25940_ = ~pi625;
  assign new_n25941_ = ~new_n8784_;
  assign new_n25942_ = ~pi626;
  assign new_n25943_ = ~new_n8787_;
  assign new_n25944_ = ~pi627;
  assign new_n25945_ = ~new_n8790_;
  assign new_n25946_ = ~pi628;
  assign new_n25947_ = ~new_n8793_;
  assign new_n25948_ = ~pi629;
  assign new_n25949_ = ~new_n8796_;
  assign new_n25950_ = ~pi630;
  assign new_n25951_ = ~new_n8799_;
  assign new_n25952_ = ~pi631;
  assign new_n25953_ = ~new_n8802_;
  assign new_n25954_ = ~pi632;
  assign new_n25955_ = ~new_n8805_;
  assign new_n25956_ = ~pi633;
  assign new_n25957_ = ~new_n8808_;
  assign new_n25958_ = ~new_n26079_ | ~new_n26078_;
  assign new_n25959_ = ~pi634;
  assign new_n25960_ = ~new_n8811_;
  assign new_n25961_ = ~pi635;
  assign new_n25962_ = ~new_n8814_;
  assign new_n25963_ = ~pi636;
  assign new_n25964_ = ~new_n8817_;
  assign new_n25965_ = ~pi637;
  assign new_n25966_ = ~new_n8820_;
  assign new_n25967_ = ~new_n26091_ | ~new_n26090_;
  assign new_n25968_ = ~new_n8764_;
  assign new_n25969_ = ~new_n26106_ | ~new_n26105_;
  assign new_n25970_ = ~new_n26111_ | ~new_n26110_;
  assign new_n25971_ = ~new_n26116_ | ~new_n26115_;
  assign new_n25972_ = ~new_n26121_ | ~new_n26120_;
  assign new_n25973_ = ~new_n26126_ | ~new_n26125_;
  assign new_n25974_ = ~new_n26131_ | ~new_n26130_;
  assign new_n25975_ = ~new_n26136_ | ~new_n26135_;
  assign new_n25976_ = ~new_n26141_ | ~new_n26140_;
  assign new_n25977_ = ~new_n26146_ | ~new_n26145_;
  assign new_n25978_ = ~new_n26156_ | ~new_n26155_;
  assign new_n25979_ = ~new_n26161_ | ~new_n26160_;
  assign new_n25980_ = ~new_n26166_ | ~new_n26165_;
  assign new_n25981_ = ~new_n26171_ | ~new_n26170_;
  assign new_n25982_ = ~new_n26176_ | ~new_n26175_;
  assign new_n25983_ = ~new_n26181_ | ~new_n26180_;
  assign new_n25984_ = ~new_n26186_ | ~new_n26185_;
  assign new_n25985_ = ~new_n26191_ | ~new_n26190_;
  assign new_n25986_ = ~new_n26196_ | ~new_n26195_;
  assign new_n25987_ = ~new_n26103_ | ~new_n26102_;
  assign new_n25988_ = ~new_n26108_ | ~new_n26107_;
  assign new_n25989_ = ~new_n26113_ | ~new_n26112_;
  assign new_n25990_ = ~new_n26118_ | ~new_n26117_;
  assign new_n25991_ = ~new_n26123_ | ~new_n26122_;
  assign new_n25992_ = ~new_n26128_ | ~new_n26127_;
  assign new_n25993_ = ~new_n26133_ | ~new_n26132_;
  assign new_n25994_ = ~new_n26138_ | ~new_n26137_;
  assign new_n25995_ = ~new_n26143_ | ~new_n26142_;
  assign new_n25996_ = new_n26099_ & new_n26148_ & new_n26147_;
  assign new_n25997_ = new_n26095_ & new_n26151_;
  assign new_n25998_ = ~new_n26153_ | ~new_n26152_;
  assign new_n25999_ = ~new_n26158_ | ~new_n26157_;
  assign new_n26000_ = ~new_n26163_ | ~new_n26162_;
  assign new_n26001_ = ~new_n26168_ | ~new_n26167_;
  assign new_n26002_ = ~new_n26173_ | ~new_n26172_;
  assign new_n26003_ = ~new_n26178_ | ~new_n26177_;
  assign new_n26004_ = ~new_n26183_ | ~new_n26182_;
  assign new_n26005_ = ~new_n26188_ | ~new_n26187_;
  assign new_n26006_ = ~new_n26193_ | ~new_n26192_;
  assign new_n26007_ = ~new_n26055_ | ~new_n26054_;
  assign new_n26008_ = ~new_n26051_ | ~new_n26050_;
  assign new_n26009_ = ~new_n26047_ | ~new_n26046_;
  assign new_n26010_ = ~new_n26043_ | ~new_n26042_;
  assign new_n26011_ = ~new_n26039_ | ~new_n26038_;
  assign new_n26012_ = ~new_n26035_ | ~new_n26034_;
  assign new_n26013_ = ~new_n26031_ | ~new_n26030_;
  assign new_n26014_ = ~new_n26027_ | ~new_n26026_;
  assign new_n26015_ = ~pi638;
  assign new_n26016_ = ~new_n8757_;
  assign new_n26017_ = ~new_n26087_ | ~new_n26086_;
  assign new_n26018_ = ~new_n26083_ | ~new_n26082_;
  assign new_n26019_ = ~new_n26075_ | ~new_n26074_;
  assign new_n26020_ = ~new_n26071_ | ~new_n26070_;
  assign new_n26021_ = ~new_n26067_ | ~new_n26066_;
  assign new_n26022_ = ~new_n26063_ | ~new_n26062_;
  assign new_n26023_ = ~new_n26059_ | ~new_n26058_;
  assign new_n26024_ = ~new_n25929_;
  assign new_n26025_ = ~pi620 | ~new_n26024_;
  assign new_n26026_ = ~new_n8769_ | ~new_n26025_;
  assign new_n26027_ = ~new_n25929_ | ~new_n25930_;
  assign new_n26028_ = ~new_n26014_;
  assign new_n26029_ = ~pi621 | ~new_n25933_;
  assign new_n26030_ = ~new_n26029_ | ~new_n26014_;
  assign new_n26031_ = ~new_n8772_ | ~new_n25932_;
  assign new_n26032_ = ~new_n26013_;
  assign new_n26033_ = ~pi622 | ~new_n25935_;
  assign new_n26034_ = ~new_n26033_ | ~new_n26013_;
  assign new_n26035_ = ~new_n8775_ | ~new_n25934_;
  assign new_n26036_ = ~new_n26012_;
  assign new_n26037_ = ~pi623 | ~new_n25937_;
  assign new_n26038_ = ~new_n26037_ | ~new_n26012_;
  assign new_n26039_ = ~new_n8778_ | ~new_n25936_;
  assign new_n26040_ = ~new_n26011_;
  assign new_n26041_ = ~pi624 | ~new_n25939_;
  assign new_n26042_ = ~new_n26041_ | ~new_n26011_;
  assign new_n26043_ = ~new_n8781_ | ~new_n25938_;
  assign new_n26044_ = ~new_n26010_;
  assign new_n26045_ = ~pi625 | ~new_n25941_;
  assign new_n26046_ = ~new_n26045_ | ~new_n26010_;
  assign new_n26047_ = ~new_n8784_ | ~new_n25940_;
  assign new_n26048_ = ~new_n26009_;
  assign new_n26049_ = ~pi626 | ~new_n25943_;
  assign new_n26050_ = ~new_n26049_ | ~new_n26009_;
  assign new_n26051_ = ~new_n8787_ | ~new_n25942_;
  assign new_n26052_ = ~new_n26008_;
  assign new_n26053_ = ~pi627 | ~new_n25945_;
  assign new_n26054_ = ~new_n26053_ | ~new_n26008_;
  assign new_n26055_ = ~new_n8790_ | ~new_n25944_;
  assign new_n26056_ = ~new_n26007_;
  assign new_n26057_ = ~pi628 | ~new_n25947_;
  assign new_n26058_ = ~new_n26057_ | ~new_n26007_;
  assign new_n26059_ = ~new_n8793_ | ~new_n25946_;
  assign new_n26060_ = ~new_n26023_;
  assign new_n26061_ = ~pi629 | ~new_n25949_;
  assign new_n26062_ = ~new_n26061_ | ~new_n26023_;
  assign new_n26063_ = ~new_n8796_ | ~new_n25948_;
  assign new_n26064_ = ~new_n26022_;
  assign new_n26065_ = ~pi630 | ~new_n25951_;
  assign new_n26066_ = ~new_n26065_ | ~new_n26022_;
  assign new_n26067_ = ~new_n8799_ | ~new_n25950_;
  assign new_n26068_ = ~new_n26021_;
  assign new_n26069_ = ~pi631 | ~new_n25953_;
  assign new_n26070_ = ~new_n26069_ | ~new_n26021_;
  assign new_n26071_ = ~new_n8802_ | ~new_n25952_;
  assign new_n26072_ = ~new_n26020_;
  assign new_n26073_ = ~pi632 | ~new_n25955_;
  assign new_n26074_ = ~new_n26073_ | ~new_n26020_;
  assign new_n26075_ = ~new_n8805_ | ~new_n25954_;
  assign new_n26076_ = ~new_n26019_;
  assign new_n26077_ = ~pi633 | ~new_n25957_;
  assign new_n26078_ = ~new_n26077_ | ~new_n26019_;
  assign new_n26079_ = ~new_n8808_ | ~new_n25956_;
  assign new_n26080_ = ~new_n25958_;
  assign new_n26081_ = ~pi634 | ~new_n26080_;
  assign new_n26082_ = ~new_n8811_ | ~new_n26081_;
  assign new_n26083_ = ~new_n25958_ | ~new_n25959_;
  assign new_n26084_ = ~new_n26018_;
  assign new_n26085_ = ~pi635 | ~new_n25962_;
  assign new_n26086_ = ~new_n26085_ | ~new_n26018_;
  assign new_n26087_ = ~new_n8814_ | ~new_n25961_;
  assign new_n26088_ = ~new_n26017_;
  assign new_n26089_ = ~pi636 | ~new_n25964_;
  assign new_n26090_ = ~new_n26089_ | ~new_n26017_;
  assign new_n26091_ = ~new_n8817_ | ~new_n25963_;
  assign new_n26092_ = ~new_n25967_;
  assign new_n26093_ = ~new_n8820_ | ~new_n25965_;
  assign new_n26094_ = ~new_n26092_ | ~new_n26093_;
  assign new_n26095_ = ~pi637 | ~new_n25966_;
  assign new_n26096_ = ~new_n25997_ | ~new_n26094_;
  assign new_n26097_ = ~pi637 | ~new_n25966_;
  assign new_n26098_ = ~new_n26097_ | ~new_n25967_;
  assign new_n26099_ = ~new_n8820_ | ~new_n25965_;
  assign new_n26100_ = ~new_n25996_ | ~new_n26098_;
  assign new_n26101_ = ~new_n8764_ | ~new_n25928_;
  assign new_n26102_ = ~pi628 | ~new_n25947_;
  assign new_n26103_ = ~new_n8793_ | ~new_n25946_;
  assign new_n26104_ = ~new_n25987_;
  assign new_n26105_ = ~new_n26056_ | ~new_n26104_;
  assign new_n26106_ = ~new_n25987_ | ~new_n26007_;
  assign new_n26107_ = ~pi627 | ~new_n25945_;
  assign new_n26108_ = ~new_n8790_ | ~new_n25944_;
  assign new_n26109_ = ~new_n25988_;
  assign new_n26110_ = ~new_n26052_ | ~new_n26109_;
  assign new_n26111_ = ~new_n25988_ | ~new_n26008_;
  assign new_n26112_ = ~pi626 | ~new_n25943_;
  assign new_n26113_ = ~new_n8787_ | ~new_n25942_;
  assign new_n26114_ = ~new_n25989_;
  assign new_n26115_ = ~new_n26048_ | ~new_n26114_;
  assign new_n26116_ = ~new_n25989_ | ~new_n26009_;
  assign new_n26117_ = ~pi625 | ~new_n25941_;
  assign new_n26118_ = ~new_n8784_ | ~new_n25940_;
  assign new_n26119_ = ~new_n25990_;
  assign new_n26120_ = ~new_n26044_ | ~new_n26119_;
  assign new_n26121_ = ~new_n25990_ | ~new_n26010_;
  assign new_n26122_ = ~pi624 | ~new_n25939_;
  assign new_n26123_ = ~new_n8781_ | ~new_n25938_;
  assign new_n26124_ = ~new_n25991_;
  assign new_n26125_ = ~new_n26040_ | ~new_n26124_;
  assign new_n26126_ = ~new_n25991_ | ~new_n26011_;
  assign new_n26127_ = ~pi623 | ~new_n25937_;
  assign new_n26128_ = ~new_n8778_ | ~new_n25936_;
  assign new_n26129_ = ~new_n25992_;
  assign new_n26130_ = ~new_n26036_ | ~new_n26129_;
  assign new_n26131_ = ~new_n25992_ | ~new_n26012_;
  assign new_n26132_ = ~pi622 | ~new_n25935_;
  assign new_n26133_ = ~new_n8775_ | ~new_n25934_;
  assign new_n26134_ = ~new_n25993_;
  assign new_n26135_ = ~new_n26032_ | ~new_n26134_;
  assign new_n26136_ = ~new_n25993_ | ~new_n26013_;
  assign new_n26137_ = ~pi621 | ~new_n25933_;
  assign new_n26138_ = ~new_n8772_ | ~new_n25932_;
  assign new_n26139_ = ~new_n25994_;
  assign new_n26140_ = ~new_n26028_ | ~new_n26139_;
  assign new_n26141_ = ~new_n25994_ | ~new_n26014_;
  assign new_n26142_ = ~new_n26024_ | ~new_n25930_;
  assign new_n26143_ = ~pi620 | ~new_n25929_;
  assign new_n26144_ = ~new_n25995_;
  assign new_n26145_ = ~new_n26144_ | ~new_n8769_;
  assign new_n26146_ = ~new_n25995_ | ~new_n25931_;
  assign new_n26147_ = ~pi638 | ~new_n26016_;
  assign new_n26148_ = ~new_n8757_ | ~new_n26015_;
  assign new_n26149_ = ~pi638 | ~new_n26016_;
  assign new_n26150_ = ~new_n8757_ | ~new_n26015_;
  assign new_n26151_ = ~new_n26150_ | ~new_n26149_;
  assign new_n26152_ = ~pi637 | ~new_n25966_;
  assign new_n26153_ = ~new_n8820_ | ~new_n25965_;
  assign new_n26154_ = ~new_n25998_;
  assign new_n26155_ = ~new_n26154_ | ~new_n26092_;
  assign new_n26156_ = ~new_n25998_ | ~new_n25967_;
  assign new_n26157_ = ~pi636 | ~new_n25964_;
  assign new_n26158_ = ~new_n8817_ | ~new_n25963_;
  assign new_n26159_ = ~new_n25999_;
  assign new_n26160_ = ~new_n26088_ | ~new_n26159_;
  assign new_n26161_ = ~new_n25999_ | ~new_n26017_;
  assign new_n26162_ = ~pi635 | ~new_n25962_;
  assign new_n26163_ = ~new_n8814_ | ~new_n25961_;
  assign new_n26164_ = ~new_n26000_;
  assign new_n26165_ = ~new_n26084_ | ~new_n26164_;
  assign new_n26166_ = ~new_n26000_ | ~new_n26018_;
  assign new_n26167_ = ~new_n8811_ | ~new_n25959_;
  assign new_n26168_ = ~pi634 | ~new_n25960_;
  assign new_n26169_ = ~new_n26001_;
  assign new_n26170_ = ~new_n26169_ | ~new_n26080_;
  assign new_n26171_ = ~new_n26001_ | ~new_n25958_;
  assign new_n26172_ = ~pi633 | ~new_n25957_;
  assign new_n26173_ = ~new_n8808_ | ~new_n25956_;
  assign new_n26174_ = ~new_n26002_;
  assign new_n26175_ = ~new_n26076_ | ~new_n26174_;
  assign new_n26176_ = ~new_n26002_ | ~new_n26019_;
  assign new_n26177_ = ~pi632 | ~new_n25955_;
  assign new_n26178_ = ~new_n8805_ | ~new_n25954_;
  assign new_n26179_ = ~new_n26003_;
  assign new_n26180_ = ~new_n26072_ | ~new_n26179_;
  assign new_n26181_ = ~new_n26003_ | ~new_n26020_;
  assign new_n26182_ = ~pi631 | ~new_n25953_;
  assign new_n26183_ = ~new_n8802_ | ~new_n25952_;
  assign new_n26184_ = ~new_n26004_;
  assign new_n26185_ = ~new_n26068_ | ~new_n26184_;
  assign new_n26186_ = ~new_n26004_ | ~new_n26021_;
  assign new_n26187_ = ~pi630 | ~new_n25951_;
  assign new_n26188_ = ~new_n8799_ | ~new_n25950_;
  assign new_n26189_ = ~new_n26005_;
  assign new_n26190_ = ~new_n26064_ | ~new_n26189_;
  assign new_n26191_ = ~new_n26005_ | ~new_n26022_;
  assign new_n26192_ = ~pi629 | ~new_n25949_;
  assign new_n26193_ = ~new_n8796_ | ~new_n25948_;
  assign new_n26194_ = ~new_n26006_;
  assign new_n26195_ = ~new_n26060_ | ~new_n26194_;
  assign new_n26196_ = ~new_n26006_ | ~new_n26023_;
  assign new_n26197_ = ~new_n8436_;
  assign new_n26198_ = ~new_n8433_;
  assign new_n26199_ = new_n26201_ & new_n26200_;
  assign new_n26200_ = ~new_n8433_ | ~new_n26197_;
  assign new_n26201_ = ~new_n8436_ | ~new_n26198_;
  assign new_n26202_ = new_n26406_ & new_n26405_;
  assign new_n26203_ = new_n26385_ & new_n26441_;
  assign new_n26204_ = new_n26443_ & new_n26442_;
  assign new_n26205_ = new_n26386_ & new_n26458_;
  assign new_n26206_ = new_n26460_ & new_n26459_;
  assign new_n26207_ = new_n26387_ & new_n26482_;
  assign new_n26208_ = new_n26484_ & new_n26483_;
  assign new_n26209_ = new_n26409_ & new_n26404_ & new_n26390_;
  assign new_n26210_ = new_n26414_ & new_n26391_;
  assign new_n26211_ = new_n26588_ & new_n26587_;
  assign new_n26212_ = ~new_n26538_ | ~new_n26541_;
  assign new_n26213_ = ~new_n26527_ | ~new_n26530_;
  assign new_n26214_ = ~new_n26516_ | ~new_n26519_;
  assign new_n26215_ = ~new_n26508_ | ~new_n26510_;
  assign new_n26216_ = ~new_n26547_ | ~new_n26358_ | ~new_n26379_;
  assign new_n26217_ = ~new_n26437_ | ~new_n26439_;
  assign new_n26218_ = ~new_n26429_ | ~new_n26432_;
  assign new_n26219_ = ~new_n26421_ | ~new_n26423_;
  assign new_n26220_ = ~new_n26368_ | ~new_n26544_;
  assign new_n26221_ = ~new_n8447_;
  assign new_n26222_ = ~new_n8447_ | ~new_n26235_;
  assign new_n26223_ = ~new_n8461_;
  assign new_n26224_ = ~new_n8791_;
  assign new_n26225_ = ~new_n8773_;
  assign new_n26226_ = ~new_n8765_;
  assign new_n26227_ = ~new_n8455_;
  assign new_n26228_ = ~new_n8776_;
  assign new_n26229_ = ~new_n8445_;
  assign new_n26230_ = ~new_n8445_ | ~new_n26225_;
  assign new_n26231_ = ~new_n8441_;
  assign new_n26232_ = ~new_n8782_;
  assign new_n26233_ = ~new_n8785_;
  assign new_n26234_ = ~new_n8779_;
  assign new_n26235_ = ~new_n8788_;
  assign new_n26236_ = ~new_n8448_;
  assign new_n26237_ = ~new_n8444_;
  assign new_n26238_ = ~new_n8437_;
  assign new_n26239_ = ~new_n8437_ | ~new_n26234_;
  assign new_n26240_ = ~new_n26410_ | ~new_n26408_;
  assign new_n26241_ = ~new_n8794_;
  assign new_n26242_ = ~new_n8460_;
  assign new_n26243_ = ~new_n26240_ | ~new_n26411_;
  assign new_n26244_ = ~new_n26239_ | ~new_n26425_;
  assign new_n26245_ = ~new_n26545_ | ~new_n26397_ | ~new_n26381_;
  assign new_n26246_ = ~new_n9279_;
  assign new_n26247_ = ~new_n8800_;
  assign new_n26248_ = ~new_n8797_;
  assign new_n26249_ = ~new_n8440_;
  assign new_n26250_ = ~new_n8439_;
  assign new_n26251_ = ~new_n8460_ | ~new_n26241_;
  assign new_n26252_ = ~new_n8803_;
  assign new_n26253_ = ~new_n8449_;
  assign new_n26254_ = ~new_n8806_;
  assign new_n26255_ = ~new_n8457_;
  assign new_n26256_ = ~new_n8815_;
  assign new_n26257_ = ~new_n8812_;
  assign new_n26258_ = ~new_n8809_;
  assign new_n26259_ = ~new_n8450_;
  assign new_n26260_ = ~new_n8451_;
  assign new_n26261_ = ~new_n8456_;
  assign new_n26262_ = ~new_n8456_ | ~new_n26258_;
  assign new_n26263_ = ~new_n8818_;
  assign new_n26264_ = ~new_n8446_;
  assign new_n26265_ = ~new_n8459_;
  assign new_n26266_ = ~new_n8823_;
  assign new_n26267_ = ~new_n8458_;
  assign new_n26268_ = ~new_n9285_;
  assign new_n26269_ = ~new_n8453_;
  assign new_n26270_ = ~new_n9282_;
  assign new_n26271_ = ~new_n9283_;
  assign new_n26272_ = ~new_n9284_;
  assign new_n26273_ = ~new_n8443_;
  assign new_n26274_ = ~new_n8438_;
  assign new_n26275_ = ~new_n8452_;
  assign new_n26276_ = ~new_n8452_ | ~new_n26272_;
  assign new_n26277_ = ~new_n9281_;
  assign new_n26278_ = ~new_n8442_;
  assign new_n26279_ = ~new_n9280_;
  assign new_n26280_ = ~new_n8435_;
  assign new_n26281_ = ~new_n9278_;
  assign new_n26282_ = ~new_n8434_;
  assign new_n26283_ = ~new_n8434_ | ~new_n26246_;
  assign new_n26284_ = ~new_n8430_;
  assign new_n26285_ = ~new_n9277_;
  assign new_n26286_ = ~new_n8431_;
  assign new_n26287_ = ~new_n26498_ | ~new_n26497_;
  assign new_n26288_ = ~new_n26276_ | ~new_n26512_;
  assign new_n26289_ = ~new_n26262_ | ~new_n26523_;
  assign new_n26290_ = ~new_n26251_ | ~new_n26534_;
  assign new_n26291_ = ~new_n8454_;
  assign new_n26292_ = ~new_n26598_ | ~new_n26597_;
  assign new_n26293_ = ~new_n26612_ | ~new_n26611_;
  assign new_n26294_ = ~new_n26617_ | ~new_n26616_;
  assign new_n26295_ = ~new_n26633_ | ~new_n26632_;
  assign new_n26296_ = ~new_n26638_ | ~new_n26637_;
  assign new_n26297_ = ~new_n26643_ | ~new_n26642_;
  assign new_n26298_ = ~new_n26648_ | ~new_n26647_;
  assign new_n26299_ = ~new_n26653_ | ~new_n26652_;
  assign new_n26300_ = ~new_n26669_ | ~new_n26668_;
  assign new_n26301_ = ~new_n26674_ | ~new_n26673_;
  assign new_n26302_ = ~new_n26557_ | ~new_n26556_;
  assign new_n26303_ = ~new_n26566_ | ~new_n26565_;
  assign new_n26304_ = ~new_n26573_ | ~new_n26572_;
  assign new_n26305_ = ~new_n26577_ | ~new_n26576_;
  assign new_n26306_ = ~new_n26586_ | ~new_n26585_;
  assign new_n26307_ = ~new_n26607_ | ~new_n26606_;
  assign new_n26308_ = ~new_n26624_ | ~new_n26623_;
  assign new_n26309_ = ~new_n26628_ | ~new_n26627_;
  assign new_n26310_ = ~new_n26660_ | ~new_n26659_;
  assign new_n26311_ = ~new_n26664_ | ~new_n26663_;
  assign new_n26312_ = ~new_n26681_ | ~new_n26680_;
  assign new_n26313_ = new_n26548_ & new_n26389_;
  assign new_n26314_ = new_n26401_ & new_n26402_;
  assign new_n26315_ = new_n26210_ & new_n26209_;
  assign new_n26316_ = new_n26553_ & new_n26550_;
  assign new_n26317_ = new_n26222_ & new_n26559_ & new_n26558_;
  assign new_n26318_ = new_n26562_ & new_n26391_;
  assign new_n26319_ = new_n26431_ & new_n26202_;
  assign new_n26320_ = new_n26569_ & new_n26390_;
  assign new_n26321_ = new_n26230_ & new_n26579_ & new_n26578_;
  assign new_n26322_ = new_n26582_ & new_n26389_;
  assign new_n26323_ = new_n26418_ & new_n26203_;
  assign new_n26324_ = new_n26463_ & new_n26205_;
  assign new_n26325_ = new_n26487_ & new_n26207_;
  assign new_n26326_ = new_n26551_ & new_n26388_;
  assign new_n26327_ = new_n26502_ & new_n26503_;
  assign new_n26328_ = new_n26505_ & new_n26591_;
  assign new_n26329_ = new_n26502_ & new_n26503_;
  assign new_n26330_ = new_n26211_ & new_n26506_;
  assign new_n26331_ = ~new_n26595_ | ~new_n26594_;
  assign new_n26332_ = new_n26283_ & new_n26600_ & new_n26599_;
  assign new_n26333_ = new_n26603_ & new_n26388_;
  assign new_n26334_ = ~new_n26609_ | ~new_n26608_;
  assign new_n26335_ = ~new_n26614_ | ~new_n26613_;
  assign new_n26336_ = new_n26518_ & new_n26208_;
  assign new_n26337_ = new_n26620_ & new_n26387_;
  assign new_n26338_ = ~new_n26630_ | ~new_n26629_;
  assign new_n26339_ = ~new_n26635_ | ~new_n26634_;
  assign new_n26340_ = ~new_n26640_ | ~new_n26639_;
  assign new_n26341_ = ~new_n26645_ | ~new_n26644_;
  assign new_n26342_ = ~new_n26650_ | ~new_n26649_;
  assign new_n26343_ = new_n26529_ & new_n26206_;
  assign new_n26344_ = new_n26656_ & new_n26386_;
  assign new_n26345_ = ~new_n26666_ | ~new_n26665_;
  assign new_n26346_ = ~new_n26671_ | ~new_n26670_;
  assign new_n26347_ = new_n26540_ & new_n26204_;
  assign new_n26348_ = new_n26677_ & new_n26385_;
  assign new_n26349_ = new_n26555_ & new_n26554_;
  assign new_n26350_ = ~new_n26316_ | ~new_n26552_;
  assign new_n26351_ = new_n26564_ & new_n26563_;
  assign new_n26352_ = new_n26571_ & new_n26570_;
  assign new_n26353_ = new_n26575_ & new_n26574_;
  assign new_n26354_ = ~new_n26314_ | ~new_n26399_;
  assign new_n26355_ = new_n26584_ & new_n26583_;
  assign new_n26356_ = ~new_n9286_;
  assign new_n26357_ = ~new_n8432_;
  assign new_n26358_ = new_n26593_ & new_n26592_;
  assign new_n26359_ = ~new_n26327_ | ~new_n26500_;
  assign new_n26360_ = new_n26605_ & new_n26604_;
  assign new_n26361_ = ~new_n26494_ | ~new_n26493_;
  assign new_n26362_ = ~new_n26490_ | ~new_n26489_;
  assign new_n26363_ = new_n26622_ & new_n26621_;
  assign new_n26364_ = new_n26626_ & new_n26625_;
  assign new_n26365_ = ~new_n26480_ | ~new_n26479_;
  assign new_n26366_ = ~new_n26476_ | ~new_n26475_;
  assign new_n26367_ = ~new_n8770_;
  assign new_n26368_ = ~new_n8765_ | ~new_n26291_;
  assign new_n26369_ = ~new_n26546_ | ~new_n26472_ | ~new_n26380_;
  assign new_n26370_ = ~new_n8821_;
  assign new_n26371_ = ~new_n26470_ | ~new_n26469_;
  assign new_n26372_ = ~new_n26466_ | ~new_n26465_;
  assign new_n26373_ = new_n26658_ & new_n26657_;
  assign new_n26374_ = new_n26662_ & new_n26661_;
  assign new_n26375_ = ~new_n26456_ | ~new_n26455_;
  assign new_n26376_ = ~new_n26452_ | ~new_n26451_;
  assign new_n26377_ = ~new_n26448_ | ~new_n26447_;
  assign new_n26378_ = new_n26679_ & new_n26678_;
  assign new_n26379_ = ~new_n26328_ | ~new_n26359_;
  assign new_n26380_ = ~new_n26371_ | ~new_n26370_;
  assign new_n26381_ = ~new_n26368_ | ~new_n26367_;
  assign new_n26382_ = ~new_n26283_;
  assign new_n26383_ = ~new_n26230_;
  assign new_n26384_ = ~new_n26222_;
  assign new_n26385_ = ~new_n8797_ | ~new_n26250_;
  assign new_n26386_ = ~new_n8812_ | ~new_n26260_;
  assign new_n26387_ = ~new_n9283_ | ~new_n26274_;
  assign new_n26388_ = ~new_n9279_ | ~new_n26282_;
  assign new_n26389_ = ~new_n8773_ | ~new_n26229_;
  assign new_n26390_ = ~new_n8782_ | ~new_n26237_;
  assign new_n26391_ = ~new_n8788_ | ~new_n26221_;
  assign new_n26392_ = ~new_n26262_;
  assign new_n26393_ = ~new_n26276_;
  assign new_n26394_ = ~new_n26239_;
  assign new_n26395_ = ~new_n26251_;
  assign new_n26396_ = ~new_n26368_;
  assign new_n26397_ = ~new_n8455_ | ~new_n26368_;
  assign new_n26398_ = ~new_n26245_;
  assign new_n26399_ = ~new_n26313_ | ~new_n26245_;
  assign new_n26400_ = ~new_n26231_ | ~new_n26230_;
  assign new_n26401_ = ~new_n26400_ | ~new_n26228_;
  assign new_n26402_ = ~new_n8441_ | ~new_n26383_;
  assign new_n26403_ = ~new_n26354_;
  assign new_n26404_ = ~new_n8785_ | ~new_n26236_;
  assign new_n26405_ = ~new_n8448_ | ~new_n26233_;
  assign new_n26406_ = ~new_n8444_ | ~new_n26232_;
  assign new_n26407_ = ~new_n26394_ | ~new_n26390_;
  assign new_n26408_ = ~new_n26202_ | ~new_n26407_;
  assign new_n26409_ = ~new_n8779_ | ~new_n26238_;
  assign new_n26410_ = ~new_n8785_ | ~new_n26236_;
  assign new_n26411_ = ~new_n26209_ | ~new_n26354_;
  assign new_n26412_ = ~new_n26240_;
  assign new_n26413_ = ~new_n26243_;
  assign new_n26414_ = ~new_n8791_ | ~new_n26223_;
  assign new_n26415_ = ~new_n26223_ | ~new_n26222_;
  assign new_n26416_ = ~new_n8461_ | ~new_n26384_;
  assign new_n26417_ = ~new_n26350_;
  assign new_n26418_ = ~new_n8794_ | ~new_n26242_;
  assign new_n26419_ = ~new_n26418_ | ~new_n26251_;
  assign new_n26420_ = ~new_n26413_ | ~new_n26222_;
  assign new_n26421_ = ~new_n26318_ | ~new_n26420_;
  assign new_n26422_ = ~new_n26243_ | ~new_n26391_;
  assign new_n26423_ = ~new_n26317_ | ~new_n26422_;
  assign new_n26424_ = ~new_n26222_ | ~new_n26391_;
  assign new_n26425_ = ~new_n26409_ | ~new_n26354_;
  assign new_n26426_ = ~new_n26244_;
  assign new_n26427_ = ~new_n8444_ | ~new_n26232_;
  assign new_n26428_ = ~new_n26426_ | ~new_n26427_;
  assign new_n26429_ = ~new_n26320_ | ~new_n26428_;
  assign new_n26430_ = ~new_n26244_ | ~new_n26390_;
  assign new_n26431_ = ~new_n8785_ | ~new_n26236_;
  assign new_n26432_ = ~new_n26319_ | ~new_n26430_;
  assign new_n26433_ = ~new_n8444_ | ~new_n26232_;
  assign new_n26434_ = ~new_n26390_ | ~new_n26433_;
  assign new_n26435_ = ~new_n26409_ | ~new_n26239_;
  assign new_n26436_ = ~new_n26398_ | ~new_n26230_;
  assign new_n26437_ = ~new_n26322_ | ~new_n26436_;
  assign new_n26438_ = ~new_n26245_ | ~new_n26389_;
  assign new_n26439_ = ~new_n26321_ | ~new_n26438_;
  assign new_n26440_ = ~new_n26389_ | ~new_n26230_;
  assign new_n26441_ = ~new_n8800_ | ~new_n26249_;
  assign new_n26442_ = ~new_n8440_ | ~new_n26247_;
  assign new_n26443_ = ~new_n8439_ | ~new_n26248_;
  assign new_n26444_ = ~new_n26395_ | ~new_n26203_;
  assign new_n26445_ = ~new_n26204_ | ~new_n26444_;
  assign new_n26446_ = ~new_n8800_ | ~new_n26249_;
  assign new_n26447_ = ~new_n26323_ | ~new_n26350_;
  assign new_n26448_ = ~new_n26446_ | ~new_n26445_;
  assign new_n26449_ = ~new_n26377_;
  assign new_n26450_ = ~new_n8803_ | ~new_n26253_;
  assign new_n26451_ = ~new_n26450_ | ~new_n26377_;
  assign new_n26452_ = ~new_n8449_ | ~new_n26252_;
  assign new_n26453_ = ~new_n26376_;
  assign new_n26454_ = ~new_n8806_ | ~new_n26255_;
  assign new_n26455_ = ~new_n26454_ | ~new_n26376_;
  assign new_n26456_ = ~new_n8457_ | ~new_n26254_;
  assign new_n26457_ = ~new_n26375_;
  assign new_n26458_ = ~new_n8815_ | ~new_n26259_;
  assign new_n26459_ = ~new_n8450_ | ~new_n26256_;
  assign new_n26460_ = ~new_n8451_ | ~new_n26257_;
  assign new_n26461_ = ~new_n26392_ | ~new_n26205_;
  assign new_n26462_ = ~new_n26206_ | ~new_n26461_;
  assign new_n26463_ = ~new_n8809_ | ~new_n26261_;
  assign new_n26464_ = ~new_n8815_ | ~new_n26259_;
  assign new_n26465_ = ~new_n26324_ | ~new_n26375_;
  assign new_n26466_ = ~new_n26464_ | ~new_n26462_;
  assign new_n26467_ = ~new_n26372_;
  assign new_n26468_ = ~new_n8818_ | ~new_n26264_;
  assign new_n26469_ = ~new_n26468_ | ~new_n26372_;
  assign new_n26470_ = ~new_n8446_ | ~new_n26263_;
  assign new_n26471_ = ~new_n26371_;
  assign new_n26472_ = ~new_n8459_ | ~new_n26371_;
  assign new_n26473_ = ~new_n26369_;
  assign new_n26474_ = ~new_n8823_ | ~new_n26267_;
  assign new_n26475_ = ~new_n26474_ | ~new_n26369_;
  assign new_n26476_ = ~new_n8458_ | ~new_n26266_;
  assign new_n26477_ = ~new_n26366_;
  assign new_n26478_ = ~new_n9285_ | ~new_n26269_;
  assign new_n26479_ = ~new_n26478_ | ~new_n26366_;
  assign new_n26480_ = ~new_n8453_ | ~new_n26268_;
  assign new_n26481_ = ~new_n26365_;
  assign new_n26482_ = ~new_n9282_ | ~new_n26273_;
  assign new_n26483_ = ~new_n8443_ | ~new_n26270_;
  assign new_n26484_ = ~new_n8438_ | ~new_n26271_;
  assign new_n26485_ = ~new_n26393_ | ~new_n26207_;
  assign new_n26486_ = ~new_n26208_ | ~new_n26485_;
  assign new_n26487_ = ~new_n9284_ | ~new_n26275_;
  assign new_n26488_ = ~new_n9282_ | ~new_n26273_;
  assign new_n26489_ = ~new_n26325_ | ~new_n26365_;
  assign new_n26490_ = ~new_n26488_ | ~new_n26486_;
  assign new_n26491_ = ~new_n26362_;
  assign new_n26492_ = ~new_n9281_ | ~new_n26278_;
  assign new_n26493_ = ~new_n26492_ | ~new_n26362_;
  assign new_n26494_ = ~new_n8442_ | ~new_n26277_;
  assign new_n26495_ = ~new_n26361_;
  assign new_n26496_ = ~new_n9280_ | ~new_n26280_;
  assign new_n26497_ = ~new_n26496_ | ~new_n26361_;
  assign new_n26498_ = ~new_n8435_ | ~new_n26279_;
  assign new_n26499_ = ~new_n26287_;
  assign new_n26500_ = ~new_n26326_ | ~new_n26287_;
  assign new_n26501_ = ~new_n26284_ | ~new_n26283_;
  assign new_n26502_ = ~new_n26501_ | ~new_n26281_;
  assign new_n26503_ = ~new_n8430_ | ~new_n26382_;
  assign new_n26504_ = ~new_n26359_;
  assign new_n26505_ = ~new_n9277_ | ~new_n26286_;
  assign new_n26506_ = ~new_n8431_ | ~new_n26285_;
  assign new_n26507_ = ~new_n26499_ | ~new_n26283_;
  assign new_n26508_ = ~new_n26333_ | ~new_n26507_;
  assign new_n26509_ = ~new_n26287_ | ~new_n26388_;
  assign new_n26510_ = ~new_n26332_ | ~new_n26509_;
  assign new_n26511_ = ~new_n26388_ | ~new_n26283_;
  assign new_n26512_ = ~new_n26487_ | ~new_n26365_;
  assign new_n26513_ = ~new_n26288_;
  assign new_n26514_ = ~new_n8438_ | ~new_n26271_;
  assign new_n26515_ = ~new_n26513_ | ~new_n26514_;
  assign new_n26516_ = ~new_n26337_ | ~new_n26515_;
  assign new_n26517_ = ~new_n26288_ | ~new_n26387_;
  assign new_n26518_ = ~new_n9282_ | ~new_n26273_;
  assign new_n26519_ = ~new_n26336_ | ~new_n26517_;
  assign new_n26520_ = ~new_n8438_ | ~new_n26271_;
  assign new_n26521_ = ~new_n26387_ | ~new_n26520_;
  assign new_n26522_ = ~new_n26487_ | ~new_n26276_;
  assign new_n26523_ = ~new_n26463_ | ~new_n26375_;
  assign new_n26524_ = ~new_n26289_;
  assign new_n26525_ = ~new_n8451_ | ~new_n26257_;
  assign new_n26526_ = ~new_n26524_ | ~new_n26525_;
  assign new_n26527_ = ~new_n26344_ | ~new_n26526_;
  assign new_n26528_ = ~new_n26289_ | ~new_n26386_;
  assign new_n26529_ = ~new_n8815_ | ~new_n26259_;
  assign new_n26530_ = ~new_n26343_ | ~new_n26528_;
  assign new_n26531_ = ~new_n8451_ | ~new_n26257_;
  assign new_n26532_ = ~new_n26386_ | ~new_n26531_;
  assign new_n26533_ = ~new_n26463_ | ~new_n26262_;
  assign new_n26534_ = ~new_n26418_ | ~new_n26350_;
  assign new_n26535_ = ~new_n26290_;
  assign new_n26536_ = ~new_n8439_ | ~new_n26248_;
  assign new_n26537_ = ~new_n26535_ | ~new_n26536_;
  assign new_n26538_ = ~new_n26348_ | ~new_n26537_;
  assign new_n26539_ = ~new_n26290_ | ~new_n26385_;
  assign new_n26540_ = ~new_n8800_ | ~new_n26249_;
  assign new_n26541_ = ~new_n26347_ | ~new_n26539_;
  assign new_n26542_ = ~new_n8439_ | ~new_n26248_;
  assign new_n26543_ = ~new_n26385_ | ~new_n26542_;
  assign new_n26544_ = ~new_n8454_ | ~new_n26226_;
  assign new_n26545_ = ~new_n8455_ | ~new_n26367_;
  assign new_n26546_ = ~new_n8459_ | ~new_n26370_;
  assign new_n26547_ = ~new_n26330_ | ~new_n26329_ | ~new_n26500_;
  assign new_n26548_ = ~new_n8776_ | ~new_n26231_;
  assign new_n26549_ = ~new_n8791_ | ~new_n26416_;
  assign new_n26550_ = ~new_n26549_ | ~new_n26415_;
  assign new_n26551_ = ~new_n9278_ | ~new_n26284_;
  assign new_n26552_ = ~new_n26315_ | ~new_n26354_;
  assign new_n26553_ = ~new_n26412_ | ~new_n26210_;
  assign new_n26554_ = ~new_n8794_ | ~new_n26242_;
  assign new_n26555_ = ~new_n8460_ | ~new_n26241_;
  assign new_n26556_ = ~new_n26419_ | ~new_n26350_;
  assign new_n26557_ = ~new_n26417_ | ~new_n26349_;
  assign new_n26558_ = ~new_n8791_ | ~new_n26223_;
  assign new_n26559_ = ~new_n8461_ | ~new_n26224_;
  assign new_n26560_ = ~new_n8791_ | ~new_n26223_;
  assign new_n26561_ = ~new_n8461_ | ~new_n26224_;
  assign new_n26562_ = ~new_n26561_ | ~new_n26560_;
  assign new_n26563_ = ~new_n8788_ | ~new_n26221_;
  assign new_n26564_ = ~new_n8447_ | ~new_n26235_;
  assign new_n26565_ = ~new_n26424_ | ~new_n26243_;
  assign new_n26566_ = ~new_n26351_ | ~new_n26413_;
  assign new_n26567_ = ~new_n8785_ | ~new_n26236_;
  assign new_n26568_ = ~new_n8448_ | ~new_n26233_;
  assign new_n26569_ = ~new_n26568_ | ~new_n26567_;
  assign new_n26570_ = ~new_n8782_ | ~new_n26237_;
  assign new_n26571_ = ~new_n8444_ | ~new_n26232_;
  assign new_n26572_ = ~new_n26434_ | ~new_n26244_;
  assign new_n26573_ = ~new_n26352_ | ~new_n26426_;
  assign new_n26574_ = ~new_n8779_ | ~new_n26238_;
  assign new_n26575_ = ~new_n8437_ | ~new_n26234_;
  assign new_n26576_ = ~new_n26435_ | ~new_n26354_;
  assign new_n26577_ = ~new_n26403_ | ~new_n26353_;
  assign new_n26578_ = ~new_n8776_ | ~new_n26231_;
  assign new_n26579_ = ~new_n8441_ | ~new_n26228_;
  assign new_n26580_ = ~new_n8776_ | ~new_n26231_;
  assign new_n26581_ = ~new_n8441_ | ~new_n26228_;
  assign new_n26582_ = ~new_n26581_ | ~new_n26580_;
  assign new_n26583_ = ~new_n8773_ | ~new_n26229_;
  assign new_n26584_ = ~new_n8445_ | ~new_n26225_;
  assign new_n26585_ = ~new_n26440_ | ~new_n26245_;
  assign new_n26586_ = ~new_n26355_ | ~new_n26398_;
  assign new_n26587_ = ~new_n9286_ | ~new_n26357_;
  assign new_n26588_ = ~new_n8432_ | ~new_n26356_;
  assign new_n26589_ = ~new_n9286_ | ~new_n26357_;
  assign new_n26590_ = ~new_n8432_ | ~new_n26356_;
  assign new_n26591_ = ~new_n26590_ | ~new_n26589_;
  assign new_n26592_ = ~new_n26285_ | ~new_n8431_ | ~new_n26591_;
  assign new_n26593_ = ~new_n9277_ | ~new_n26211_ | ~new_n26286_;
  assign new_n26594_ = ~new_n9277_ | ~new_n26286_;
  assign new_n26595_ = ~new_n8431_ | ~new_n26285_;
  assign new_n26596_ = ~new_n26331_;
  assign new_n26597_ = ~new_n26504_ | ~new_n26596_;
  assign new_n26598_ = ~new_n26331_ | ~new_n26359_;
  assign new_n26599_ = ~new_n9278_ | ~new_n26284_;
  assign new_n26600_ = ~new_n8430_ | ~new_n26281_;
  assign new_n26601_ = ~new_n9278_ | ~new_n26284_;
  assign new_n26602_ = ~new_n8430_ | ~new_n26281_;
  assign new_n26603_ = ~new_n26602_ | ~new_n26601_;
  assign new_n26604_ = ~new_n9279_ | ~new_n26282_;
  assign new_n26605_ = ~new_n8434_ | ~new_n26246_;
  assign new_n26606_ = ~new_n26511_ | ~new_n26287_;
  assign new_n26607_ = ~new_n26360_ | ~new_n26499_;
  assign new_n26608_ = ~new_n9280_ | ~new_n26280_;
  assign new_n26609_ = ~new_n8435_ | ~new_n26279_;
  assign new_n26610_ = ~new_n26334_;
  assign new_n26611_ = ~new_n26495_ | ~new_n26610_;
  assign new_n26612_ = ~new_n26334_ | ~new_n26361_;
  assign new_n26613_ = ~new_n9281_ | ~new_n26278_;
  assign new_n26614_ = ~new_n8442_ | ~new_n26277_;
  assign new_n26615_ = ~new_n26335_;
  assign new_n26616_ = ~new_n26491_ | ~new_n26615_;
  assign new_n26617_ = ~new_n26335_ | ~new_n26362_;
  assign new_n26618_ = ~new_n9282_ | ~new_n26273_;
  assign new_n26619_ = ~new_n8443_ | ~new_n26270_;
  assign new_n26620_ = ~new_n26619_ | ~new_n26618_;
  assign new_n26621_ = ~new_n9283_ | ~new_n26274_;
  assign new_n26622_ = ~new_n8438_ | ~new_n26271_;
  assign new_n26623_ = ~new_n26521_ | ~new_n26288_;
  assign new_n26624_ = ~new_n26363_ | ~new_n26513_;
  assign new_n26625_ = ~new_n9284_ | ~new_n26275_;
  assign new_n26626_ = ~new_n8452_ | ~new_n26272_;
  assign new_n26627_ = ~new_n26522_ | ~new_n26365_;
  assign new_n26628_ = ~new_n26481_ | ~new_n26364_;
  assign new_n26629_ = ~new_n9285_ | ~new_n26269_;
  assign new_n26630_ = ~new_n8453_ | ~new_n26268_;
  assign new_n26631_ = ~new_n26338_;
  assign new_n26632_ = ~new_n26477_ | ~new_n26631_;
  assign new_n26633_ = ~new_n26338_ | ~new_n26366_;
  assign new_n26634_ = ~new_n8770_ | ~new_n26227_;
  assign new_n26635_ = ~new_n8455_ | ~new_n26367_;
  assign new_n26636_ = ~new_n26339_;
  assign new_n26637_ = ~new_n26396_ | ~new_n26636_;
  assign new_n26638_ = ~new_n26339_ | ~new_n26368_;
  assign new_n26639_ = ~new_n8823_ | ~new_n26267_;
  assign new_n26640_ = ~new_n8458_ | ~new_n26266_;
  assign new_n26641_ = ~new_n26340_;
  assign new_n26642_ = ~new_n26473_ | ~new_n26641_;
  assign new_n26643_ = ~new_n26340_ | ~new_n26369_;
  assign new_n26644_ = ~new_n8821_ | ~new_n26265_;
  assign new_n26645_ = ~new_n8459_ | ~new_n26370_;
  assign new_n26646_ = ~new_n26341_;
  assign new_n26647_ = ~new_n26471_ | ~new_n26646_;
  assign new_n26648_ = ~new_n26341_ | ~new_n26371_;
  assign new_n26649_ = ~new_n8818_ | ~new_n26264_;
  assign new_n26650_ = ~new_n8446_ | ~new_n26263_;
  assign new_n26651_ = ~new_n26342_;
  assign new_n26652_ = ~new_n26467_ | ~new_n26651_;
  assign new_n26653_ = ~new_n26342_ | ~new_n26372_;
  assign new_n26654_ = ~new_n8815_ | ~new_n26259_;
  assign new_n26655_ = ~new_n8450_ | ~new_n26256_;
  assign new_n26656_ = ~new_n26655_ | ~new_n26654_;
  assign new_n26657_ = ~new_n8812_ | ~new_n26260_;
  assign new_n26658_ = ~new_n8451_ | ~new_n26257_;
  assign new_n26659_ = ~new_n26532_ | ~new_n26289_;
  assign new_n26660_ = ~new_n26373_ | ~new_n26524_;
  assign new_n26661_ = ~new_n8809_ | ~new_n26261_;
  assign new_n26662_ = ~new_n8456_ | ~new_n26258_;
  assign new_n26663_ = ~new_n26533_ | ~new_n26375_;
  assign new_n26664_ = ~new_n26457_ | ~new_n26374_;
  assign new_n26665_ = ~new_n8806_ | ~new_n26255_;
  assign new_n26666_ = ~new_n8457_ | ~new_n26254_;
  assign new_n26667_ = ~new_n26345_;
  assign new_n26668_ = ~new_n26453_ | ~new_n26667_;
  assign new_n26669_ = ~new_n26345_ | ~new_n26376_;
  assign new_n26670_ = ~new_n8803_ | ~new_n26253_;
  assign new_n26671_ = ~new_n8449_ | ~new_n26252_;
  assign new_n26672_ = ~new_n26346_;
  assign new_n26673_ = ~new_n26449_ | ~new_n26672_;
  assign new_n26674_ = ~new_n26346_ | ~new_n26377_;
  assign new_n26675_ = ~new_n8800_ | ~new_n26249_;
  assign new_n26676_ = ~new_n8440_ | ~new_n26247_;
  assign new_n26677_ = ~new_n26676_ | ~new_n26675_;
  assign new_n26678_ = ~new_n8797_ | ~new_n26250_;
  assign new_n26679_ = ~new_n8439_ | ~new_n26248_;
  assign new_n26680_ = ~new_n26543_ | ~new_n26290_;
  assign new_n26681_ = ~new_n26378_ | ~new_n26535_;
  assign new_n26682_ = new_n26886_ & new_n26885_;
  assign new_n26683_ = new_n26865_ & new_n26921_;
  assign new_n26684_ = new_n26923_ & new_n26922_;
  assign new_n26685_ = new_n26866_ & new_n26938_;
  assign new_n26686_ = new_n26940_ & new_n26939_;
  assign new_n26687_ = new_n26867_ & new_n26962_;
  assign new_n26688_ = new_n26964_ & new_n26963_;
  assign new_n26689_ = new_n26889_ & new_n26884_ & new_n26870_;
  assign new_n26690_ = new_n26894_ & new_n26871_;
  assign new_n26691_ = new_n27068_ & new_n27067_;
  assign new_n26692_ = ~new_n27018_ | ~new_n27021_;
  assign new_n26693_ = ~new_n27007_ | ~new_n27010_;
  assign new_n26694_ = ~new_n26996_ | ~new_n26999_;
  assign new_n26695_ = ~new_n26988_ | ~new_n26990_;
  assign new_n26696_ = ~new_n27027_ | ~new_n26838_ | ~new_n26859_;
  assign new_n26697_ = ~new_n26917_ | ~new_n26919_;
  assign new_n26698_ = ~new_n26909_ | ~new_n26912_;
  assign new_n26699_ = ~new_n26901_ | ~new_n26903_;
  assign new_n26700_ = ~new_n26848_ | ~new_n27024_;
  assign new_n26701_ = ~new_n8447_;
  assign new_n26702_ = ~new_n8447_ | ~new_n26715_;
  assign new_n26703_ = ~new_n8461_;
  assign new_n26704_ = ~new_n8791_;
  assign new_n26705_ = ~new_n8773_;
  assign new_n26706_ = ~new_n8765_;
  assign new_n26707_ = ~new_n8455_;
  assign new_n26708_ = ~new_n8776_;
  assign new_n26709_ = ~new_n8445_;
  assign new_n26710_ = ~new_n8445_ | ~new_n26705_;
  assign new_n26711_ = ~new_n8441_;
  assign new_n26712_ = ~new_n8782_;
  assign new_n26713_ = ~new_n8785_;
  assign new_n26714_ = ~new_n8779_;
  assign new_n26715_ = ~new_n8788_;
  assign new_n26716_ = ~new_n8448_;
  assign new_n26717_ = ~new_n8444_;
  assign new_n26718_ = ~new_n8437_;
  assign new_n26719_ = ~new_n8437_ | ~new_n26714_;
  assign new_n26720_ = ~new_n26890_ | ~new_n26888_;
  assign new_n26721_ = ~new_n8794_;
  assign new_n26722_ = ~new_n8460_;
  assign new_n26723_ = ~new_n26720_ | ~new_n26891_;
  assign new_n26724_ = ~new_n26719_ | ~new_n26905_;
  assign new_n26725_ = ~new_n27025_ | ~new_n26877_ | ~new_n26861_;
  assign new_n26726_ = ~new_n9279_;
  assign new_n26727_ = ~new_n8800_;
  assign new_n26728_ = ~new_n8797_;
  assign new_n26729_ = ~new_n8440_;
  assign new_n26730_ = ~new_n8439_;
  assign new_n26731_ = ~new_n8460_ | ~new_n26721_;
  assign new_n26732_ = ~new_n8803_;
  assign new_n26733_ = ~new_n8449_;
  assign new_n26734_ = ~new_n8806_;
  assign new_n26735_ = ~new_n8457_;
  assign new_n26736_ = ~new_n8815_;
  assign new_n26737_ = ~new_n8812_;
  assign new_n26738_ = ~new_n8809_;
  assign new_n26739_ = ~new_n8450_;
  assign new_n26740_ = ~new_n8451_;
  assign new_n26741_ = ~new_n8456_;
  assign new_n26742_ = ~new_n8456_ | ~new_n26738_;
  assign new_n26743_ = ~new_n8818_;
  assign new_n26744_ = ~new_n8446_;
  assign new_n26745_ = ~new_n8459_;
  assign new_n26746_ = ~new_n8823_;
  assign new_n26747_ = ~new_n8458_;
  assign new_n26748_ = ~new_n9285_;
  assign new_n26749_ = ~new_n8453_;
  assign new_n26750_ = ~new_n9282_;
  assign new_n26751_ = ~new_n9283_;
  assign new_n26752_ = ~new_n9284_;
  assign new_n26753_ = ~new_n8443_;
  assign new_n26754_ = ~new_n8438_;
  assign new_n26755_ = ~new_n8452_;
  assign new_n26756_ = ~new_n8452_ | ~new_n26752_;
  assign new_n26757_ = ~new_n9281_;
  assign new_n26758_ = ~new_n8442_;
  assign new_n26759_ = ~new_n9280_;
  assign new_n26760_ = ~new_n8435_;
  assign new_n26761_ = ~new_n9278_;
  assign new_n26762_ = ~new_n8434_;
  assign new_n26763_ = ~new_n8434_ | ~new_n26726_;
  assign new_n26764_ = ~new_n8430_;
  assign new_n26765_ = ~new_n9277_;
  assign new_n26766_ = ~new_n8431_;
  assign new_n26767_ = ~new_n26978_ | ~new_n26977_;
  assign new_n26768_ = ~new_n26756_ | ~new_n26992_;
  assign new_n26769_ = ~new_n26742_ | ~new_n27003_;
  assign new_n26770_ = ~new_n26731_ | ~new_n27014_;
  assign new_n26771_ = ~new_n8454_;
  assign new_n26772_ = ~new_n27078_ | ~new_n27077_;
  assign new_n26773_ = ~new_n27092_ | ~new_n27091_;
  assign new_n26774_ = ~new_n27097_ | ~new_n27096_;
  assign new_n26775_ = ~new_n27113_ | ~new_n27112_;
  assign new_n26776_ = ~new_n27118_ | ~new_n27117_;
  assign new_n26777_ = ~new_n27123_ | ~new_n27122_;
  assign new_n26778_ = ~new_n27128_ | ~new_n27127_;
  assign new_n26779_ = ~new_n27133_ | ~new_n27132_;
  assign new_n26780_ = ~new_n27149_ | ~new_n27148_;
  assign new_n26781_ = ~new_n27154_ | ~new_n27153_;
  assign new_n26782_ = ~new_n27037_ | ~new_n27036_;
  assign new_n26783_ = ~new_n27046_ | ~new_n27045_;
  assign new_n26784_ = ~new_n27053_ | ~new_n27052_;
  assign new_n26785_ = ~new_n27057_ | ~new_n27056_;
  assign new_n26786_ = ~new_n27066_ | ~new_n27065_;
  assign new_n26787_ = ~new_n27087_ | ~new_n27086_;
  assign new_n26788_ = ~new_n27104_ | ~new_n27103_;
  assign new_n26789_ = ~new_n27108_ | ~new_n27107_;
  assign new_n26790_ = ~new_n27140_ | ~new_n27139_;
  assign new_n26791_ = ~new_n27144_ | ~new_n27143_;
  assign new_n26792_ = ~new_n27161_ | ~new_n27160_;
  assign new_n26793_ = new_n27028_ & new_n26869_;
  assign new_n26794_ = new_n26881_ & new_n26882_;
  assign new_n26795_ = new_n26690_ & new_n26689_;
  assign new_n26796_ = new_n27033_ & new_n27030_;
  assign new_n26797_ = new_n26702_ & new_n27039_ & new_n27038_;
  assign new_n26798_ = new_n27042_ & new_n26871_;
  assign new_n26799_ = new_n26911_ & new_n26682_;
  assign new_n26800_ = new_n27049_ & new_n26870_;
  assign new_n26801_ = new_n26710_ & new_n27059_ & new_n27058_;
  assign new_n26802_ = new_n27062_ & new_n26869_;
  assign new_n26803_ = new_n26898_ & new_n26683_;
  assign new_n26804_ = new_n26943_ & new_n26685_;
  assign new_n26805_ = new_n26967_ & new_n26687_;
  assign new_n26806_ = new_n27031_ & new_n26868_;
  assign new_n26807_ = new_n26982_ & new_n26983_;
  assign new_n26808_ = new_n26985_ & new_n27071_;
  assign new_n26809_ = new_n26982_ & new_n26983_;
  assign new_n26810_ = new_n26691_ & new_n26986_;
  assign new_n26811_ = ~new_n27075_ | ~new_n27074_;
  assign new_n26812_ = new_n26763_ & new_n27080_ & new_n27079_;
  assign new_n26813_ = new_n27083_ & new_n26868_;
  assign new_n26814_ = ~new_n27089_ | ~new_n27088_;
  assign new_n26815_ = ~new_n27094_ | ~new_n27093_;
  assign new_n26816_ = new_n26998_ & new_n26688_;
  assign new_n26817_ = new_n27100_ & new_n26867_;
  assign new_n26818_ = ~new_n27110_ | ~new_n27109_;
  assign new_n26819_ = ~new_n27115_ | ~new_n27114_;
  assign new_n26820_ = ~new_n27120_ | ~new_n27119_;
  assign new_n26821_ = ~new_n27125_ | ~new_n27124_;
  assign new_n26822_ = ~new_n27130_ | ~new_n27129_;
  assign new_n26823_ = new_n27009_ & new_n26686_;
  assign new_n26824_ = new_n27136_ & new_n26866_;
  assign new_n26825_ = ~new_n27146_ | ~new_n27145_;
  assign new_n26826_ = ~new_n27151_ | ~new_n27150_;
  assign new_n26827_ = new_n27020_ & new_n26684_;
  assign new_n26828_ = new_n27157_ & new_n26865_;
  assign new_n26829_ = new_n27035_ & new_n27034_;
  assign new_n26830_ = ~new_n26796_ | ~new_n27032_;
  assign new_n26831_ = new_n27044_ & new_n27043_;
  assign new_n26832_ = new_n27051_ & new_n27050_;
  assign new_n26833_ = new_n27055_ & new_n27054_;
  assign new_n26834_ = ~new_n26794_ | ~new_n26879_;
  assign new_n26835_ = new_n27064_ & new_n27063_;
  assign new_n26836_ = ~new_n9286_;
  assign new_n26837_ = ~new_n8432_;
  assign new_n26838_ = new_n27073_ & new_n27072_;
  assign new_n26839_ = ~new_n26807_ | ~new_n26980_;
  assign new_n26840_ = new_n27085_ & new_n27084_;
  assign new_n26841_ = ~new_n26974_ | ~new_n26973_;
  assign new_n26842_ = ~new_n26970_ | ~new_n26969_;
  assign new_n26843_ = new_n27102_ & new_n27101_;
  assign new_n26844_ = new_n27106_ & new_n27105_;
  assign new_n26845_ = ~new_n26960_ | ~new_n26959_;
  assign new_n26846_ = ~new_n26956_ | ~new_n26955_;
  assign new_n26847_ = ~new_n8770_;
  assign new_n26848_ = ~new_n8765_ | ~new_n26771_;
  assign new_n26849_ = ~new_n27026_ | ~new_n26952_ | ~new_n26860_;
  assign new_n26850_ = ~new_n8821_;
  assign new_n26851_ = ~new_n26950_ | ~new_n26949_;
  assign new_n26852_ = ~new_n26946_ | ~new_n26945_;
  assign new_n26853_ = new_n27138_ & new_n27137_;
  assign new_n26854_ = new_n27142_ & new_n27141_;
  assign new_n26855_ = ~new_n26936_ | ~new_n26935_;
  assign new_n26856_ = ~new_n26932_ | ~new_n26931_;
  assign new_n26857_ = ~new_n26928_ | ~new_n26927_;
  assign new_n26858_ = new_n27159_ & new_n27158_;
  assign new_n26859_ = ~new_n26808_ | ~new_n26839_;
  assign new_n26860_ = ~new_n26851_ | ~new_n26850_;
  assign new_n26861_ = ~new_n26848_ | ~new_n26847_;
  assign new_n26862_ = ~new_n26763_;
  assign new_n26863_ = ~new_n26710_;
  assign new_n26864_ = ~new_n26702_;
  assign new_n26865_ = ~new_n8797_ | ~new_n26730_;
  assign new_n26866_ = ~new_n8812_ | ~new_n26740_;
  assign new_n26867_ = ~new_n9283_ | ~new_n26754_;
  assign new_n26868_ = ~new_n9279_ | ~new_n26762_;
  assign new_n26869_ = ~new_n8773_ | ~new_n26709_;
  assign new_n26870_ = ~new_n8782_ | ~new_n26717_;
  assign new_n26871_ = ~new_n8788_ | ~new_n26701_;
  assign new_n26872_ = ~new_n26742_;
  assign new_n26873_ = ~new_n26756_;
  assign new_n26874_ = ~new_n26719_;
  assign new_n26875_ = ~new_n26731_;
  assign new_n26876_ = ~new_n26848_;
  assign new_n26877_ = ~new_n8455_ | ~new_n26848_;
  assign new_n26878_ = ~new_n26725_;
  assign new_n26879_ = ~new_n26793_ | ~new_n26725_;
  assign new_n26880_ = ~new_n26711_ | ~new_n26710_;
  assign new_n26881_ = ~new_n26880_ | ~new_n26708_;
  assign new_n26882_ = ~new_n8441_ | ~new_n26863_;
  assign new_n26883_ = ~new_n26834_;
  assign new_n26884_ = ~new_n8785_ | ~new_n26716_;
  assign new_n26885_ = ~new_n8448_ | ~new_n26713_;
  assign new_n26886_ = ~new_n8444_ | ~new_n26712_;
  assign new_n26887_ = ~new_n26874_ | ~new_n26870_;
  assign new_n26888_ = ~new_n26682_ | ~new_n26887_;
  assign new_n26889_ = ~new_n8779_ | ~new_n26718_;
  assign new_n26890_ = ~new_n8785_ | ~new_n26716_;
  assign new_n26891_ = ~new_n26689_ | ~new_n26834_;
  assign new_n26892_ = ~new_n26720_;
  assign new_n26893_ = ~new_n26723_;
  assign new_n26894_ = ~new_n8791_ | ~new_n26703_;
  assign new_n26895_ = ~new_n26703_ | ~new_n26702_;
  assign new_n26896_ = ~new_n8461_ | ~new_n26864_;
  assign new_n26897_ = ~new_n26830_;
  assign new_n26898_ = ~new_n8794_ | ~new_n26722_;
  assign new_n26899_ = ~new_n26898_ | ~new_n26731_;
  assign new_n26900_ = ~new_n26893_ | ~new_n26702_;
  assign new_n26901_ = ~new_n26798_ | ~new_n26900_;
  assign new_n26902_ = ~new_n26723_ | ~new_n26871_;
  assign new_n26903_ = ~new_n26797_ | ~new_n26902_;
  assign new_n26904_ = ~new_n26702_ | ~new_n26871_;
  assign new_n26905_ = ~new_n26889_ | ~new_n26834_;
  assign new_n26906_ = ~new_n26724_;
  assign new_n26907_ = ~new_n8444_ | ~new_n26712_;
  assign new_n26908_ = ~new_n26906_ | ~new_n26907_;
  assign new_n26909_ = ~new_n26800_ | ~new_n26908_;
  assign new_n26910_ = ~new_n26724_ | ~new_n26870_;
  assign new_n26911_ = ~new_n8785_ | ~new_n26716_;
  assign new_n26912_ = ~new_n26799_ | ~new_n26910_;
  assign new_n26913_ = ~new_n8444_ | ~new_n26712_;
  assign new_n26914_ = ~new_n26870_ | ~new_n26913_;
  assign new_n26915_ = ~new_n26889_ | ~new_n26719_;
  assign new_n26916_ = ~new_n26878_ | ~new_n26710_;
  assign new_n26917_ = ~new_n26802_ | ~new_n26916_;
  assign new_n26918_ = ~new_n26725_ | ~new_n26869_;
  assign new_n26919_ = ~new_n26801_ | ~new_n26918_;
  assign new_n26920_ = ~new_n26869_ | ~new_n26710_;
  assign new_n26921_ = ~new_n8800_ | ~new_n26729_;
  assign new_n26922_ = ~new_n8440_ | ~new_n26727_;
  assign new_n26923_ = ~new_n8439_ | ~new_n26728_;
  assign new_n26924_ = ~new_n26875_ | ~new_n26683_;
  assign new_n26925_ = ~new_n26684_ | ~new_n26924_;
  assign new_n26926_ = ~new_n8800_ | ~new_n26729_;
  assign new_n26927_ = ~new_n26803_ | ~new_n26830_;
  assign new_n26928_ = ~new_n26926_ | ~new_n26925_;
  assign new_n26929_ = ~new_n26857_;
  assign new_n26930_ = ~new_n8803_ | ~new_n26733_;
  assign new_n26931_ = ~new_n26930_ | ~new_n26857_;
  assign new_n26932_ = ~new_n8449_ | ~new_n26732_;
  assign new_n26933_ = ~new_n26856_;
  assign new_n26934_ = ~new_n8806_ | ~new_n26735_;
  assign new_n26935_ = ~new_n26934_ | ~new_n26856_;
  assign new_n26936_ = ~new_n8457_ | ~new_n26734_;
  assign new_n26937_ = ~new_n26855_;
  assign new_n26938_ = ~new_n8815_ | ~new_n26739_;
  assign new_n26939_ = ~new_n8450_ | ~new_n26736_;
  assign new_n26940_ = ~new_n8451_ | ~new_n26737_;
  assign new_n26941_ = ~new_n26872_ | ~new_n26685_;
  assign new_n26942_ = ~new_n26686_ | ~new_n26941_;
  assign new_n26943_ = ~new_n8809_ | ~new_n26741_;
  assign new_n26944_ = ~new_n8815_ | ~new_n26739_;
  assign new_n26945_ = ~new_n26804_ | ~new_n26855_;
  assign new_n26946_ = ~new_n26944_ | ~new_n26942_;
  assign new_n26947_ = ~new_n26852_;
  assign new_n26948_ = ~new_n8818_ | ~new_n26744_;
  assign new_n26949_ = ~new_n26948_ | ~new_n26852_;
  assign new_n26950_ = ~new_n8446_ | ~new_n26743_;
  assign new_n26951_ = ~new_n26851_;
  assign new_n26952_ = ~new_n8459_ | ~new_n26851_;
  assign new_n26953_ = ~new_n26849_;
  assign new_n26954_ = ~new_n8823_ | ~new_n26747_;
  assign new_n26955_ = ~new_n26954_ | ~new_n26849_;
  assign new_n26956_ = ~new_n8458_ | ~new_n26746_;
  assign new_n26957_ = ~new_n26846_;
  assign new_n26958_ = ~new_n9285_ | ~new_n26749_;
  assign new_n26959_ = ~new_n26958_ | ~new_n26846_;
  assign new_n26960_ = ~new_n8453_ | ~new_n26748_;
  assign new_n26961_ = ~new_n26845_;
  assign new_n26962_ = ~new_n9282_ | ~new_n26753_;
  assign new_n26963_ = ~new_n8443_ | ~new_n26750_;
  assign new_n26964_ = ~new_n8438_ | ~new_n26751_;
  assign new_n26965_ = ~new_n26873_ | ~new_n26687_;
  assign new_n26966_ = ~new_n26688_ | ~new_n26965_;
  assign new_n26967_ = ~new_n9284_ | ~new_n26755_;
  assign new_n26968_ = ~new_n9282_ | ~new_n26753_;
  assign new_n26969_ = ~new_n26805_ | ~new_n26845_;
  assign new_n26970_ = ~new_n26968_ | ~new_n26966_;
  assign new_n26971_ = ~new_n26842_;
  assign new_n26972_ = ~new_n9281_ | ~new_n26758_;
  assign new_n26973_ = ~new_n26972_ | ~new_n26842_;
  assign new_n26974_ = ~new_n8442_ | ~new_n26757_;
  assign new_n26975_ = ~new_n26841_;
  assign new_n26976_ = ~new_n9280_ | ~new_n26760_;
  assign new_n26977_ = ~new_n26976_ | ~new_n26841_;
  assign new_n26978_ = ~new_n8435_ | ~new_n26759_;
  assign new_n26979_ = ~new_n26767_;
  assign new_n26980_ = ~new_n26806_ | ~new_n26767_;
  assign new_n26981_ = ~new_n26764_ | ~new_n26763_;
  assign new_n26982_ = ~new_n26981_ | ~new_n26761_;
  assign new_n26983_ = ~new_n8430_ | ~new_n26862_;
  assign new_n26984_ = ~new_n26839_;
  assign new_n26985_ = ~new_n9277_ | ~new_n26766_;
  assign new_n26986_ = ~new_n8431_ | ~new_n26765_;
  assign new_n26987_ = ~new_n26979_ | ~new_n26763_;
  assign new_n26988_ = ~new_n26813_ | ~new_n26987_;
  assign new_n26989_ = ~new_n26767_ | ~new_n26868_;
  assign new_n26990_ = ~new_n26812_ | ~new_n26989_;
  assign new_n26991_ = ~new_n26868_ | ~new_n26763_;
  assign new_n26992_ = ~new_n26967_ | ~new_n26845_;
  assign new_n26993_ = ~new_n26768_;
  assign new_n26994_ = ~new_n8438_ | ~new_n26751_;
  assign new_n26995_ = ~new_n26993_ | ~new_n26994_;
  assign new_n26996_ = ~new_n26817_ | ~new_n26995_;
  assign new_n26997_ = ~new_n26768_ | ~new_n26867_;
  assign new_n26998_ = ~new_n9282_ | ~new_n26753_;
  assign new_n26999_ = ~new_n26816_ | ~new_n26997_;
  assign new_n27000_ = ~new_n8438_ | ~new_n26751_;
  assign new_n27001_ = ~new_n26867_ | ~new_n27000_;
  assign new_n27002_ = ~new_n26967_ | ~new_n26756_;
  assign new_n27003_ = ~new_n26943_ | ~new_n26855_;
  assign new_n27004_ = ~new_n26769_;
  assign new_n27005_ = ~new_n8451_ | ~new_n26737_;
  assign new_n27006_ = ~new_n27004_ | ~new_n27005_;
  assign new_n27007_ = ~new_n26824_ | ~new_n27006_;
  assign new_n27008_ = ~new_n26769_ | ~new_n26866_;
  assign new_n27009_ = ~new_n8815_ | ~new_n26739_;
  assign new_n27010_ = ~new_n26823_ | ~new_n27008_;
  assign new_n27011_ = ~new_n8451_ | ~new_n26737_;
  assign new_n27012_ = ~new_n26866_ | ~new_n27011_;
  assign new_n27013_ = ~new_n26943_ | ~new_n26742_;
  assign new_n27014_ = ~new_n26898_ | ~new_n26830_;
  assign new_n27015_ = ~new_n26770_;
  assign new_n27016_ = ~new_n8439_ | ~new_n26728_;
  assign new_n27017_ = ~new_n27015_ | ~new_n27016_;
  assign new_n27018_ = ~new_n26828_ | ~new_n27017_;
  assign new_n27019_ = ~new_n26770_ | ~new_n26865_;
  assign new_n27020_ = ~new_n8800_ | ~new_n26729_;
  assign new_n27021_ = ~new_n26827_ | ~new_n27019_;
  assign new_n27022_ = ~new_n8439_ | ~new_n26728_;
  assign new_n27023_ = ~new_n26865_ | ~new_n27022_;
  assign new_n27024_ = ~new_n8454_ | ~new_n26706_;
  assign new_n27025_ = ~new_n8455_ | ~new_n26847_;
  assign new_n27026_ = ~new_n8459_ | ~new_n26850_;
  assign new_n27027_ = ~new_n26810_ | ~new_n26809_ | ~new_n26980_;
  assign new_n27028_ = ~new_n8776_ | ~new_n26711_;
  assign new_n27029_ = ~new_n8791_ | ~new_n26896_;
  assign new_n27030_ = ~new_n27029_ | ~new_n26895_;
  assign new_n27031_ = ~new_n9278_ | ~new_n26764_;
  assign new_n27032_ = ~new_n26795_ | ~new_n26834_;
  assign new_n27033_ = ~new_n26892_ | ~new_n26690_;
  assign new_n27034_ = ~new_n8794_ | ~new_n26722_;
  assign new_n27035_ = ~new_n8460_ | ~new_n26721_;
  assign new_n27036_ = ~new_n26899_ | ~new_n26830_;
  assign new_n27037_ = ~new_n26897_ | ~new_n26829_;
  assign new_n27038_ = ~new_n8791_ | ~new_n26703_;
  assign new_n27039_ = ~new_n8461_ | ~new_n26704_;
  assign new_n27040_ = ~new_n8791_ | ~new_n26703_;
  assign new_n27041_ = ~new_n8461_ | ~new_n26704_;
  assign new_n27042_ = ~new_n27041_ | ~new_n27040_;
  assign new_n27043_ = ~new_n8788_ | ~new_n26701_;
  assign new_n27044_ = ~new_n8447_ | ~new_n26715_;
  assign new_n27045_ = ~new_n26904_ | ~new_n26723_;
  assign new_n27046_ = ~new_n26831_ | ~new_n26893_;
  assign new_n27047_ = ~new_n8785_ | ~new_n26716_;
  assign new_n27048_ = ~new_n8448_ | ~new_n26713_;
  assign new_n27049_ = ~new_n27048_ | ~new_n27047_;
  assign new_n27050_ = ~new_n8782_ | ~new_n26717_;
  assign new_n27051_ = ~new_n8444_ | ~new_n26712_;
  assign new_n27052_ = ~new_n26914_ | ~new_n26724_;
  assign new_n27053_ = ~new_n26832_ | ~new_n26906_;
  assign new_n27054_ = ~new_n8779_ | ~new_n26718_;
  assign new_n27055_ = ~new_n8437_ | ~new_n26714_;
  assign new_n27056_ = ~new_n26915_ | ~new_n26834_;
  assign new_n27057_ = ~new_n26883_ | ~new_n26833_;
  assign new_n27058_ = ~new_n8776_ | ~new_n26711_;
  assign new_n27059_ = ~new_n8441_ | ~new_n26708_;
  assign new_n27060_ = ~new_n8776_ | ~new_n26711_;
  assign new_n27061_ = ~new_n8441_ | ~new_n26708_;
  assign new_n27062_ = ~new_n27061_ | ~new_n27060_;
  assign new_n27063_ = ~new_n8773_ | ~new_n26709_;
  assign new_n27064_ = ~new_n8445_ | ~new_n26705_;
  assign new_n27065_ = ~new_n26920_ | ~new_n26725_;
  assign new_n27066_ = ~new_n26835_ | ~new_n26878_;
  assign new_n27067_ = ~new_n9286_ | ~new_n26837_;
  assign new_n27068_ = ~new_n8432_ | ~new_n26836_;
  assign new_n27069_ = ~new_n9286_ | ~new_n26837_;
  assign new_n27070_ = ~new_n8432_ | ~new_n26836_;
  assign new_n27071_ = ~new_n27070_ | ~new_n27069_;
  assign new_n27072_ = ~new_n26765_ | ~new_n8431_ | ~new_n27071_;
  assign new_n27073_ = ~new_n9277_ | ~new_n26691_ | ~new_n26766_;
  assign new_n27074_ = ~new_n9277_ | ~new_n26766_;
  assign new_n27075_ = ~new_n8431_ | ~new_n26765_;
  assign new_n27076_ = ~new_n26811_;
  assign new_n27077_ = ~new_n26984_ | ~new_n27076_;
  assign new_n27078_ = ~new_n26811_ | ~new_n26839_;
  assign new_n27079_ = ~new_n9278_ | ~new_n26764_;
  assign new_n27080_ = ~new_n8430_ | ~new_n26761_;
  assign new_n27081_ = ~new_n9278_ | ~new_n26764_;
  assign new_n27082_ = ~new_n8430_ | ~new_n26761_;
  assign new_n27083_ = ~new_n27082_ | ~new_n27081_;
  assign new_n27084_ = ~new_n9279_ | ~new_n26762_;
  assign new_n27085_ = ~new_n8434_ | ~new_n26726_;
  assign new_n27086_ = ~new_n26991_ | ~new_n26767_;
  assign new_n27087_ = ~new_n26840_ | ~new_n26979_;
  assign new_n27088_ = ~new_n9280_ | ~new_n26760_;
  assign new_n27089_ = ~new_n8435_ | ~new_n26759_;
  assign new_n27090_ = ~new_n26814_;
  assign new_n27091_ = ~new_n26975_ | ~new_n27090_;
  assign new_n27092_ = ~new_n26814_ | ~new_n26841_;
  assign new_n27093_ = ~new_n9281_ | ~new_n26758_;
  assign new_n27094_ = ~new_n8442_ | ~new_n26757_;
  assign new_n27095_ = ~new_n26815_;
  assign new_n27096_ = ~new_n26971_ | ~new_n27095_;
  assign new_n27097_ = ~new_n26815_ | ~new_n26842_;
  assign new_n27098_ = ~new_n9282_ | ~new_n26753_;
  assign new_n27099_ = ~new_n8443_ | ~new_n26750_;
  assign new_n27100_ = ~new_n27099_ | ~new_n27098_;
  assign new_n27101_ = ~new_n9283_ | ~new_n26754_;
  assign new_n27102_ = ~new_n8438_ | ~new_n26751_;
  assign new_n27103_ = ~new_n27001_ | ~new_n26768_;
  assign new_n27104_ = ~new_n26843_ | ~new_n26993_;
  assign new_n27105_ = ~new_n9284_ | ~new_n26755_;
  assign new_n27106_ = ~new_n8452_ | ~new_n26752_;
  assign new_n27107_ = ~new_n27002_ | ~new_n26845_;
  assign new_n27108_ = ~new_n26961_ | ~new_n26844_;
  assign new_n27109_ = ~new_n9285_ | ~new_n26749_;
  assign new_n27110_ = ~new_n8453_ | ~new_n26748_;
  assign new_n27111_ = ~new_n26818_;
  assign new_n27112_ = ~new_n26957_ | ~new_n27111_;
  assign new_n27113_ = ~new_n26818_ | ~new_n26846_;
  assign new_n27114_ = ~new_n8770_ | ~new_n26707_;
  assign new_n27115_ = ~new_n8455_ | ~new_n26847_;
  assign new_n27116_ = ~new_n26819_;
  assign new_n27117_ = ~new_n26876_ | ~new_n27116_;
  assign new_n27118_ = ~new_n26819_ | ~new_n26848_;
  assign new_n27119_ = ~new_n8823_ | ~new_n26747_;
  assign new_n27120_ = ~new_n8458_ | ~new_n26746_;
  assign new_n27121_ = ~new_n26820_;
  assign new_n27122_ = ~new_n26953_ | ~new_n27121_;
  assign new_n27123_ = ~new_n26820_ | ~new_n26849_;
  assign new_n27124_ = ~new_n8821_ | ~new_n26745_;
  assign new_n27125_ = ~new_n8459_ | ~new_n26850_;
  assign new_n27126_ = ~new_n26821_;
  assign new_n27127_ = ~new_n26951_ | ~new_n27126_;
  assign new_n27128_ = ~new_n26821_ | ~new_n26851_;
  assign new_n27129_ = ~new_n8818_ | ~new_n26744_;
  assign new_n27130_ = ~new_n8446_ | ~new_n26743_;
  assign new_n27131_ = ~new_n26822_;
  assign new_n27132_ = ~new_n26947_ | ~new_n27131_;
  assign new_n27133_ = ~new_n26822_ | ~new_n26852_;
  assign new_n27134_ = ~new_n8815_ | ~new_n26739_;
  assign new_n27135_ = ~new_n8450_ | ~new_n26736_;
  assign new_n27136_ = ~new_n27135_ | ~new_n27134_;
  assign new_n27137_ = ~new_n8812_ | ~new_n26740_;
  assign new_n27138_ = ~new_n8451_ | ~new_n26737_;
  assign new_n27139_ = ~new_n27012_ | ~new_n26769_;
  assign new_n27140_ = ~new_n26853_ | ~new_n27004_;
  assign new_n27141_ = ~new_n8809_ | ~new_n26741_;
  assign new_n27142_ = ~new_n8456_ | ~new_n26738_;
  assign new_n27143_ = ~new_n27013_ | ~new_n26855_;
  assign new_n27144_ = ~new_n26937_ | ~new_n26854_;
  assign new_n27145_ = ~new_n8806_ | ~new_n26735_;
  assign new_n27146_ = ~new_n8457_ | ~new_n26734_;
  assign new_n27147_ = ~new_n26825_;
  assign new_n27148_ = ~new_n26933_ | ~new_n27147_;
  assign new_n27149_ = ~new_n26825_ | ~new_n26856_;
  assign new_n27150_ = ~new_n8803_ | ~new_n26733_;
  assign new_n27151_ = ~new_n8449_ | ~new_n26732_;
  assign new_n27152_ = ~new_n26826_;
  assign new_n27153_ = ~new_n26929_ | ~new_n27152_;
  assign new_n27154_ = ~new_n26826_ | ~new_n26857_;
  assign new_n27155_ = ~new_n8800_ | ~new_n26729_;
  assign new_n27156_ = ~new_n8440_ | ~new_n26727_;
  assign new_n27157_ = ~new_n27156_ | ~new_n27155_;
  assign new_n27158_ = ~new_n8797_ | ~new_n26730_;
  assign new_n27159_ = ~new_n8439_ | ~new_n26728_;
  assign new_n27160_ = ~new_n27023_ | ~new_n26770_;
  assign new_n27161_ = ~new_n26858_ | ~new_n27015_;
  assign new_n27162_ = new_n27263_ & new_n27264_;
  assign new_n27163_ = new_n27274_ & new_n27273_;
  assign new_n27164_ = new_n27298_ & new_n27297_;
  assign new_n27165_ = new_n27356_ & new_n27355_;
  assign new_n27166_ = new_n27358_ & new_n27357_;
  assign new_n27167_ = ~new_n27352_ | ~new_n27166_ | ~new_n27350_;
  assign new_n27168_ = ~new_n8494_;
  assign new_n27169_ = ~new_n8472_;
  assign new_n27170_ = ~new_n8473_;
  assign new_n27171_ = ~new_n8508_;
  assign new_n27172_ = ~new_n8514_;
  assign new_n27173_ = ~new_n8513_;
  assign new_n27174_ = ~new_n8484_;
  assign new_n27175_ = ~new_n8485_;
  assign new_n27176_ = ~new_n8490_;
  assign new_n27177_ = ~new_n8491_;
  assign new_n27178_ = ~new_n8492_;
  assign new_n27179_ = ~new_n8520_;
  assign new_n27180_ = ~new_n8519_;
  assign new_n27181_ = ~new_n8524_;
  assign new_n27182_ = ~new_n8523_;
  assign new_n27183_ = ~new_n8522_;
  assign new_n27184_ = ~new_n8521_;
  assign new_n27185_ = ~new_n8489_;
  assign new_n27186_ = ~new_n8487_;
  assign new_n27187_ = ~new_n8488_;
  assign new_n27188_ = ~new_n8486_;
  assign new_n27189_ = ~new_n8518_;
  assign new_n27190_ = ~new_n8517_;
  assign new_n27191_ = ~new_n8516_;
  assign new_n27192_ = ~new_n8515_;
  assign new_n27193_ = ~new_n8479_;
  assign new_n27194_ = ~new_n8478_;
  assign new_n27195_ = ~new_n8482_;
  assign new_n27196_ = ~new_n8483_;
  assign new_n27197_ = ~new_n8481_;
  assign new_n27198_ = ~new_n8480_;
  assign new_n27199_ = ~new_n8512_;
  assign new_n27200_ = ~new_n8511_;
  assign new_n27201_ = ~new_n8510_;
  assign new_n27202_ = ~new_n8509_;
  assign new_n27203_ = ~new_n8477_;
  assign new_n27204_ = ~new_n8476_;
  assign new_n27205_ = ~new_n27313_ | ~new_n27312_;
  assign new_n27206_ = ~new_n8507_;
  assign new_n27207_ = ~new_n8474_;
  assign new_n27208_ = ~new_n8501_;
  assign new_n27209_ = ~new_n8502_;
  assign new_n27210_ = ~new_n8506_;
  assign new_n27211_ = ~new_n8505_;
  assign new_n27212_ = ~new_n8504_;
  assign new_n27213_ = ~new_n8503_;
  assign new_n27214_ = ~new_n8465_;
  assign new_n27215_ = ~new_n8467_;
  assign new_n27216_ = ~new_n8466_;
  assign new_n27217_ = ~new_n8464_;
  assign new_n27218_ = ~new_n8471_;
  assign new_n27219_ = ~new_n8470_;
  assign new_n27220_ = ~new_n8468_;
  assign new_n27221_ = ~new_n8469_;
  assign new_n27222_ = ~new_n8498_;
  assign new_n27223_ = ~new_n8497_;
  assign new_n27224_ = ~new_n27334_ | ~new_n27333_;
  assign new_n27225_ = ~new_n8499_;
  assign new_n27226_ = ~new_n8500_;
  assign new_n27227_ = ~new_n8496_;
  assign new_n27228_ = ~new_n8527_;
  assign new_n27229_ = new_n27267_ & new_n27266_;
  assign new_n27230_ = new_n27163_ & new_n27280_;
  assign new_n27231_ = new_n8489_ & new_n27184_;
  assign new_n27232_ = new_n8488_ & new_n27179_;
  assign new_n27233_ = new_n27234_ & new_n27282_ & new_n27283_;
  assign new_n27234_ = new_n27286_ & new_n27285_;
  assign new_n27235_ = new_n27162_ & new_n27236_;
  assign new_n27236_ = new_n27294_ & new_n27295_;
  assign new_n27237_ = new_n8482_ & new_n27172_;
  assign new_n27238_ = new_n8483_ & new_n27192_;
  assign new_n27239_ = new_n27241_ & new_n27299_ & new_n27300_;
  assign new_n27240_ = new_n27302_ & new_n27301_;
  assign new_n27241_ = new_n27240_ & new_n27164_;
  assign new_n27242_ = new_n8512_ & new_n27198_;
  assign new_n27243_ = new_n8511_ & new_n27193_;
  assign new_n27244_ = new_n27245_ & new_n27304_ & new_n27306_;
  assign new_n27245_ = new_n27308_ & new_n27307_;
  assign new_n27246_ = new_n27260_ & new_n27259_;
  assign new_n27247_ = new_n27318_ & new_n27317_;
  assign new_n27248_ = new_n8506_ & new_n27207_;
  assign new_n27249_ = new_n27325_ & new_n27321_ & new_n27327_ & new_n27326_;
  assign new_n27250_ = new_n27331_ & new_n27330_;
  assign new_n27251_ = new_n27328_ & new_n27332_ & new_n27252_ & new_n27329_ & new_n27250_;
  assign new_n27252_ = new_n27348_ & new_n27349_ & new_n27347_;
  assign new_n27253_ = new_n8498_ & new_n27216_;
  assign new_n27254_ = new_n27330_ & new_n27331_;
  assign new_n27255_ = new_n27354_ & new_n27342_;
  assign new_n27256_ = ~new_n8462_;
  assign new_n27257_ = ~new_n8463_;
  assign new_n27258_ = ~new_n27343_ | ~new_n27351_;
  assign new_n27259_ = ~new_n8472_ | ~new_n27212_;
  assign new_n27260_ = ~new_n8473_ | ~new_n27211_;
  assign new_n27261_ = ~new_n8508_ | ~new_n27204_;
  assign new_n27262_ = ~new_n8484_ | ~new_n27191_;
  assign new_n27263_ = ~new_n8513_ | ~new_n27197_;
  assign new_n27264_ = ~new_n8514_ | ~new_n27195_;
  assign new_n27265_ = ~new_n8485_ | ~new_n27190_;
  assign new_n27266_ = ~new_n8490_ | ~new_n27183_;
  assign new_n27267_ = ~new_n8491_ | ~new_n27182_;
  assign new_n27268_ = ~new_n8525_ | ~new_n8526_;
  assign new_n27269_ = ~new_n8493_ | ~new_n27268_;
  assign new_n27270_ = new_n8525_ | new_n8526_;
  assign new_n27271_ = ~new_n8492_ | ~new_n27181_;
  assign new_n27272_ = ~new_n27267_ | ~new_n27270_ | ~new_n27271_ | ~new_n27269_ | ~new_n27266_;
  assign new_n27273_ = ~new_n8520_ | ~new_n27187_;
  assign new_n27274_ = ~new_n8519_ | ~new_n27186_;
  assign new_n27275_ = ~new_n8524_ | ~new_n27178_;
  assign new_n27276_ = ~new_n8523_ | ~new_n27177_;
  assign new_n27277_ = ~new_n27276_ | ~new_n27275_;
  assign new_n27278_ = ~new_n27229_ | ~new_n27277_;
  assign new_n27279_ = ~new_n8522_ | ~new_n27176_;
  assign new_n27280_ = ~new_n8521_ | ~new_n27185_;
  assign new_n27281_ = ~new_n27279_ | ~new_n27230_ | ~new_n27272_ | ~new_n27278_;
  assign new_n27282_ = ~new_n27231_ | ~new_n27163_;
  assign new_n27283_ = ~new_n8487_ | ~new_n27180_;
  assign new_n27284_ = ~new_n8519_ | ~new_n27186_;
  assign new_n27285_ = ~new_n27232_ | ~new_n27284_;
  assign new_n27286_ = ~new_n8486_ | ~new_n27189_;
  assign new_n27287_ = ~new_n27281_ | ~new_n27233_;
  assign new_n27288_ = ~new_n8518_ | ~new_n27188_;
  assign new_n27289_ = ~new_n27288_ | ~new_n27287_;
  assign new_n27290_ = ~new_n27289_ | ~new_n27265_;
  assign new_n27291_ = ~new_n8517_ | ~new_n27175_;
  assign new_n27292_ = ~new_n27291_ | ~new_n27290_;
  assign new_n27293_ = ~new_n27292_ | ~new_n27262_;
  assign new_n27294_ = ~new_n8516_ | ~new_n27174_;
  assign new_n27295_ = ~new_n8515_ | ~new_n27196_;
  assign new_n27296_ = ~new_n27293_ | ~new_n27235_;
  assign new_n27297_ = ~new_n8479_ | ~new_n27200_;
  assign new_n27298_ = ~new_n8478_ | ~new_n27201_;
  assign new_n27299_ = ~new_n27237_ | ~new_n27263_;
  assign new_n27300_ = ~new_n27238_ | ~new_n27162_;
  assign new_n27301_ = ~new_n8481_ | ~new_n27173_;
  assign new_n27302_ = ~new_n8480_ | ~new_n27199_;
  assign new_n27303_ = ~new_n27296_ | ~new_n27239_;
  assign new_n27304_ = ~new_n27242_ | ~new_n27164_;
  assign new_n27305_ = ~new_n8478_ | ~new_n27201_;
  assign new_n27306_ = ~new_n27243_ | ~new_n27305_;
  assign new_n27307_ = ~new_n8510_ | ~new_n27194_;
  assign new_n27308_ = ~new_n8509_ | ~new_n27203_;
  assign new_n27309_ = ~new_n27303_ | ~new_n27244_;
  assign new_n27310_ = ~new_n8477_ | ~new_n27202_;
  assign new_n27311_ = ~new_n27310_ | ~new_n27309_;
  assign new_n27312_ = ~new_n27311_ | ~new_n27261_;
  assign new_n27313_ = ~new_n8476_ | ~new_n27171_;
  assign new_n27314_ = ~new_n27205_;
  assign new_n27315_ = ~new_n8507_ | ~new_n27314_;
  assign new_n27316_ = ~new_n8475_ | ~new_n27315_;
  assign new_n27317_ = ~new_n27205_ | ~new_n27206_;
  assign new_n27318_ = ~new_n8474_ | ~new_n27210_;
  assign new_n27319_ = ~new_n27247_ | ~new_n27246_ | ~new_n27316_;
  assign new_n27320_ = ~new_n8501_ | ~new_n27221_;
  assign new_n27321_ = ~new_n8502_ | ~new_n27219_;
  assign new_n27322_ = ~new_n27248_ | ~new_n27260_;
  assign new_n27323_ = ~new_n8505_ | ~new_n27170_;
  assign new_n27324_ = ~new_n27323_ | ~new_n27322_;
  assign new_n27325_ = ~new_n27324_ | ~new_n27259_;
  assign new_n27326_ = ~new_n8504_ | ~new_n27169_;
  assign new_n27327_ = ~new_n8503_ | ~new_n27218_;
  assign new_n27328_ = ~new_n27320_ | ~new_n27249_ | ~new_n27319_;
  assign new_n27329_ = ~new_n8465_ | ~new_n27223_;
  assign new_n27330_ = ~new_n8467_ | ~new_n27225_;
  assign new_n27331_ = ~new_n8466_ | ~new_n27222_;
  assign new_n27332_ = ~new_n8464_ | ~new_n27227_;
  assign new_n27333_ = ~new_n27253_ | ~new_n27329_;
  assign new_n27334_ = ~new_n8497_ | ~new_n27214_;
  assign new_n27335_ = ~new_n27224_;
  assign new_n27336_ = ~new_n8499_ | ~new_n27215_;
  assign new_n27337_ = ~new_n8500_ | ~new_n27220_;
  assign new_n27338_ = ~new_n27337_ | ~new_n27336_;
  assign new_n27339_ = ~new_n27335_ | ~new_n27227_;
  assign new_n27340_ = ~new_n27339_ | ~new_n27217_;
  assign new_n27341_ = ~new_n27338_ | ~new_n27332_ | ~new_n27329_ | ~new_n27254_;
  assign new_n27342_ = ~new_n8496_ | ~new_n27224_;
  assign new_n27343_ = ~new_n27165_ | ~new_n27257_;
  assign new_n27344_ = ~new_n8471_ | ~new_n27213_;
  assign new_n27345_ = ~new_n8470_ | ~new_n27209_;
  assign new_n27346_ = ~new_n27345_ | ~new_n27344_;
  assign new_n27347_ = ~new_n27320_ | ~new_n27321_ | ~new_n27346_;
  assign new_n27348_ = ~new_n8468_ | ~new_n27226_;
  assign new_n27349_ = ~new_n8469_ | ~new_n27208_;
  assign new_n27350_ = ~new_n27258_ | ~new_n27251_;
  assign new_n27351_ = ~new_n8495_ | ~new_n27165_;
  assign new_n27352_ = ~new_n27353_ | ~new_n27258_;
  assign new_n27353_ = ~new_n27255_ | ~new_n27341_ | ~new_n27340_;
  assign new_n27354_ = ~new_n8495_ | ~new_n27257_;
  assign new_n27355_ = ~new_n8462_ | ~new_n27168_;
  assign new_n27356_ = ~new_n8494_ | ~new_n27256_;
  assign new_n27357_ = ~new_n27256_ | ~new_n8494_ | ~new_n27228_;
  assign new_n27358_ = ~new_n8462_ | ~new_n8527_ | ~new_n27168_;
  assign new_n27359_ = new_n27534_ & new_n27533_;
  assign new_n27360_ = new_n27552_ & new_n27551_;
  assign new_n27361_ = new_n27592_ & new_n27591_;
  assign new_n27362_ = new_n27601_ & new_n27600_;
  assign new_n27363_ = new_n27619_ & new_n27618_;
  assign new_n27364_ = new_n27627_ & new_n27626_;
  assign new_n27365_ = new_n27706_ & new_n27703_;
  assign new_n27366_ = new_n27699_ & new_n27696_;
  assign new_n27367_ = new_n27690_ & new_n27687_;
  assign new_n27368_ = new_n27681_ & new_n27678_;
  assign new_n27369_ = new_n27675_ & new_n27673_;
  assign new_n27370_ = new_n27668_ & new_n27665_;
  assign new_n27371_ = new_n27590_ & new_n27587_;
  assign new_n27372_ = new_n27582_ & new_n27579_;
  assign new_n27373_ = new_n27568_ & new_n27565_;
  assign new_n27374_ = ~new_n8785_;
  assign new_n27375_ = ~new_n8448_;
  assign new_n27376_ = ~new_n8447_;
  assign new_n27377_ = ~new_n8448_ | ~new_n8785_;
  assign new_n27378_ = ~new_n8788_;
  assign new_n27379_ = ~new_n8779_;
  assign new_n27380_ = ~new_n8437_;
  assign new_n27381_ = ~new_n8444_;
  assign new_n27382_ = ~new_n8773_;
  assign new_n27383_ = ~new_n8445_;
  assign new_n27384_ = ~new_n8765_;
  assign new_n27385_ = ~new_n8454_;
  assign new_n27386_ = ~new_n8454_ | ~new_n8765_;
  assign new_n27387_ = ~new_n8776_;
  assign new_n27388_ = ~new_n8441_;
  assign new_n27389_ = ~new_n8437_ | ~new_n8779_;
  assign new_n27390_ = ~new_n8782_;
  assign new_n27391_ = ~new_n8791_;
  assign new_n27392_ = ~new_n8461_;
  assign new_n27393_ = ~new_n8460_;
  assign new_n27394_ = ~new_n8794_;
  assign new_n27395_ = ~new_n27416_ | ~new_n27560_;
  assign new_n27396_ = ~new_n27472_ | ~new_n27548_;
  assign new_n27397_ = ~new_n27537_ | ~new_n27538_;
  assign new_n27398_ = ~new_n8770_ | ~new_n8455_;
  assign new_n27399_ = ~new_n27477_ | ~new_n27574_;
  assign new_n27400_ = ~new_n27571_ | ~new_n27570_;
  assign new_n27401_ = ~new_n9278_;
  assign new_n27402_ = ~new_n8430_;
  assign new_n27403_ = ~new_n8434_;
  assign new_n27404_ = ~new_n9279_;
  assign new_n27405_ = ~new_n9280_;
  assign new_n27406_ = ~new_n8435_;
  assign new_n27407_ = ~new_n9281_;
  assign new_n27408_ = ~new_n8442_;
  assign new_n27409_ = ~new_n9284_;
  assign new_n27410_ = ~new_n8452_;
  assign new_n27411_ = ~new_n8815_;
  assign new_n27412_ = ~new_n8450_;
  assign new_n27413_ = ~new_n8446_;
  assign new_n27414_ = ~new_n8450_ | ~new_n8815_;
  assign new_n27415_ = ~new_n8818_;
  assign new_n27416_ = ~new_n8461_ | ~new_n8791_;
  assign new_n27417_ = ~new_n8797_;
  assign new_n27418_ = ~new_n8439_;
  assign new_n27419_ = ~new_n8803_;
  assign new_n27420_ = ~new_n8449_;
  assign new_n27421_ = ~new_n8800_;
  assign new_n27422_ = ~new_n8440_;
  assign new_n27423_ = ~new_n8440_ | ~new_n8800_;
  assign new_n27424_ = ~new_n8806_;
  assign new_n27425_ = ~new_n8457_;
  assign new_n27426_ = ~new_n8809_;
  assign new_n27427_ = ~new_n8456_;
  assign new_n27428_ = ~new_n8812_;
  assign new_n27429_ = ~new_n8451_;
  assign new_n27430_ = ~new_n8821_;
  assign new_n27431_ = ~new_n8459_;
  assign new_n27432_ = ~new_n8459_ | ~new_n8821_;
  assign new_n27433_ = ~new_n8823_;
  assign new_n27434_ = ~new_n8458_;
  assign new_n27435_ = ~new_n8458_ | ~new_n8823_;
  assign new_n27436_ = ~new_n9285_;
  assign new_n27437_ = ~new_n9283_;
  assign new_n27438_ = ~new_n8438_;
  assign new_n27439_ = ~new_n9282_;
  assign new_n27440_ = ~new_n8443_;
  assign new_n27441_ = ~new_n9279_ | ~new_n8434_;
  assign new_n27442_ = ~new_n8431_;
  assign new_n27443_ = ~new_n9277_;
  assign new_n27444_ = ~new_n27661_ | ~new_n27531_;
  assign new_n27445_ = ~new_n8453_;
  assign new_n27446_ = ~new_n27432_ | ~new_n27670_;
  assign new_n27447_ = ~new_n27616_ | ~new_n27615_;
  assign new_n27448_ = ~new_n27423_ | ~new_n27692_;
  assign new_n27449_ = ~new_n27812_ | ~new_n27811_;
  assign new_n27450_ = ~new_n27859_ | ~new_n27858_;
  assign new_n27451_ = ~new_n27730_ | ~new_n27729_;
  assign new_n27452_ = ~new_n27735_ | ~new_n27734_;
  assign new_n27453_ = ~new_n27742_ | ~new_n27741_;
  assign new_n27454_ = ~new_n27749_ | ~new_n27748_;
  assign new_n27455_ = ~new_n27754_ | ~new_n27753_;
  assign new_n27456_ = ~new_n27763_ | ~new_n27762_;
  assign new_n27457_ = ~new_n27770_ | ~new_n27769_;
  assign new_n27458_ = ~new_n27777_ | ~new_n27776_;
  assign new_n27459_ = ~new_n27784_ | ~new_n27783_;
  assign new_n27460_ = ~new_n27789_ | ~new_n27788_;
  assign new_n27461_ = ~new_n27796_ | ~new_n27795_;
  assign new_n27462_ = ~new_n27803_ | ~new_n27802_;
  assign new_n27463_ = ~new_n27817_ | ~new_n27816_;
  assign new_n27464_ = ~new_n27822_ | ~new_n27821_;
  assign new_n27465_ = ~new_n27829_ | ~new_n27828_;
  assign new_n27466_ = ~new_n27836_ | ~new_n27835_;
  assign new_n27467_ = ~new_n27843_ | ~new_n27842_;
  assign new_n27468_ = ~new_n27850_ | ~new_n27849_;
  assign new_n27469_ = ~new_n27855_ | ~new_n27854_;
  assign new_n27470_ = new_n27544_ & new_n27542_;
  assign new_n27471_ = new_n27359_ & new_n27535_;
  assign new_n27472_ = new_n27549_ & new_n27547_;
  assign new_n27473_ = new_n27556_ & new_n27555_;
  assign new_n27474_ = new_n27377_ & new_n27737_ & new_n27736_;
  assign new_n27475_ = new_n27567_ & new_n27360_;
  assign new_n27476_ = new_n27536_ & new_n27535_;
  assign new_n27477_ = new_n27575_ & new_n27573_;
  assign new_n27478_ = new_n27389_ & new_n27744_ & new_n27743_;
  assign new_n27479_ = new_n27581_ & new_n27359_;
  assign new_n27480_ = new_n27589_ & new_n27536_;
  assign new_n27481_ = new_n27559_ & new_n27361_;
  assign new_n27482_ = new_n27594_ & new_n27526_;
  assign new_n27483_ = new_n27605_ & new_n27362_;
  assign new_n27484_ = new_n27603_ & new_n27527_;
  assign new_n27485_ = new_n27623_ & new_n27622_;
  assign new_n27486_ = new_n27628_ & new_n27364_ & new_n27637_;
  assign new_n27487_ = new_n27640_ & new_n27635_;
  assign new_n27488_ = new_n27656_ & new_n27653_;
  assign new_n27489_ = new_n27723_ & new_n27657_;
  assign new_n27490_ = new_n27515_ & new_n27633_;
  assign new_n27491_ = new_n27435_ & new_n27810_ & new_n27809_;
  assign new_n27492_ = new_n27680_ & new_n27364_;
  assign new_n27493_ = new_n27414_ & new_n27824_ & new_n27823_;
  assign new_n27494_ = new_n27689_ & new_n27363_;
  assign new_n27495_ = new_n27527_ & new_n27845_ & new_n27844_;
  assign new_n27496_ = new_n27698_ & new_n27362_;
  assign new_n27497_ = new_n27526_ & new_n27857_ & new_n27856_;
  assign new_n27498_ = new_n27705_ & new_n27361_;
  assign new_n27499_ = ~new_n27473_ | ~new_n27557_;
  assign new_n27500_ = ~new_n27572_ | ~new_n27584_;
  assign new_n27501_ = ~new_n8432_;
  assign new_n27502_ = ~new_n9286_;
  assign new_n27503_ = new_n27758_ & new_n27757_;
  assign new_n27504_ = ~new_n27719_ | ~new_n27659_ | ~new_n27524_;
  assign new_n27505_ = new_n27765_ & new_n27764_;
  assign new_n27506_ = ~new_n27489_ | ~new_n27725_ | ~new_n27724_;
  assign new_n27507_ = new_n27772_ & new_n27771_;
  assign new_n27508_ = ~new_n27441_ | ~new_n27720_ | ~new_n27654_;
  assign new_n27509_ = new_n27779_ & new_n27778_;
  assign new_n27510_ = ~new_n27648_ | ~new_n27647_;
  assign new_n27511_ = new_n27791_ & new_n27790_;
  assign new_n27512_ = ~new_n27644_ | ~new_n27643_;
  assign new_n27513_ = new_n27798_ & new_n27797_;
  assign new_n27514_ = ~new_n27487_ | ~new_n27639_;
  assign new_n27515_ = new_n27805_ & new_n27804_;
  assign new_n27516_ = ~new_n27398_ | ~new_n27682_;
  assign new_n27517_ = ~new_n27485_ | ~new_n27624_;
  assign new_n27518_ = new_n27831_ & new_n27830_;
  assign new_n27519_ = ~new_n27612_ | ~new_n27611_;
  assign new_n27520_ = new_n27838_ & new_n27837_;
  assign new_n27521_ = ~new_n27608_ | ~new_n27607_;
  assign new_n27522_ = ~new_n27598_ | ~new_n27597_;
  assign new_n27523_ = ~new_n27722_ | ~new_n27721_;
  assign new_n27524_ = ~new_n8431_ | ~new_n27506_;
  assign new_n27525_ = ~new_n27389_;
  assign new_n27526_ = ~new_n8794_ | ~new_n8460_;
  assign new_n27527_ = ~new_n8449_ | ~new_n8803_;
  assign new_n27528_ = ~new_n8435_ | ~new_n9280_;
  assign new_n27529_ = ~new_n27423_;
  assign new_n27530_ = ~new_n27432_;
  assign new_n27531_ = ~new_n8442_ | ~new_n9281_;
  assign new_n27532_ = ~new_n27416_;
  assign new_n27533_ = new_n8444_ | new_n8782_;
  assign new_n27534_ = new_n8437_ | new_n8779_;
  assign new_n27535_ = new_n8776_ | new_n8441_;
  assign new_n27536_ = new_n8773_ | new_n8445_;
  assign new_n27537_ = ~new_n27386_;
  assign new_n27538_ = new_n8770_ | new_n8455_;
  assign new_n27539_ = ~new_n27397_;
  assign new_n27540_ = ~new_n27398_;
  assign new_n27541_ = ~new_n27397_ | ~new_n27398_;
  assign new_n27542_ = ~new_n8445_ | ~new_n8773_;
  assign new_n27543_ = ~new_n27541_ | ~new_n27536_;
  assign new_n27544_ = ~new_n8441_ | ~new_n8776_;
  assign new_n27545_ = ~new_n27470_ | ~new_n27543_;
  assign new_n27546_ = ~new_n27390_ | ~new_n27389_;
  assign new_n27547_ = ~new_n8444_ | ~new_n27546_;
  assign new_n27548_ = ~new_n27471_ | ~new_n27545_;
  assign new_n27549_ = ~new_n8782_ | ~new_n27525_;
  assign new_n27550_ = ~new_n27396_;
  assign new_n27551_ = new_n8447_ | new_n8788_;
  assign new_n27552_ = new_n8448_ | new_n8785_;
  assign new_n27553_ = ~new_n27377_;
  assign new_n27554_ = ~new_n27378_ | ~new_n27377_;
  assign new_n27555_ = ~new_n8447_ | ~new_n27554_;
  assign new_n27556_ = ~new_n8788_ | ~new_n27553_;
  assign new_n27557_ = ~new_n27360_ | ~new_n27396_;
  assign new_n27558_ = ~new_n27499_;
  assign new_n27559_ = new_n8791_ | new_n8461_;
  assign new_n27560_ = ~new_n27559_ | ~new_n27499_;
  assign new_n27561_ = ~new_n27395_;
  assign new_n27562_ = new_n8460_ | new_n8794_;
  assign new_n27563_ = new_n8785_ | new_n8448_;
  assign new_n27564_ = ~new_n27563_ | ~new_n27396_;
  assign new_n27565_ = ~new_n27474_ | ~new_n27564_;
  assign new_n27566_ = ~new_n27550_ | ~new_n27377_;
  assign new_n27567_ = ~new_n8788_ | ~new_n8447_;
  assign new_n27568_ = ~new_n27475_ | ~new_n27566_;
  assign new_n27569_ = new_n8448_ | new_n8785_;
  assign new_n27570_ = ~new_n27540_ | ~new_n27536_;
  assign new_n27571_ = ~new_n8445_ | ~new_n8773_;
  assign new_n27572_ = ~new_n27400_;
  assign new_n27573_ = ~new_n27476_ | ~new_n27539_;
  assign new_n27574_ = ~new_n27400_ | ~new_n27535_;
  assign new_n27575_ = ~new_n8441_ | ~new_n8776_;
  assign new_n27576_ = ~new_n27399_;
  assign new_n27577_ = new_n8779_ | new_n8437_;
  assign new_n27578_ = ~new_n27577_ | ~new_n27399_;
  assign new_n27579_ = ~new_n27478_ | ~new_n27578_;
  assign new_n27580_ = ~new_n27576_ | ~new_n27389_;
  assign new_n27581_ = ~new_n8782_ | ~new_n8444_;
  assign new_n27582_ = ~new_n27479_ | ~new_n27580_;
  assign new_n27583_ = new_n8437_ | new_n8779_;
  assign new_n27584_ = ~new_n27539_ | ~new_n27536_;
  assign new_n27585_ = ~new_n27500_;
  assign new_n27586_ = ~new_n8441_ | ~new_n8776_;
  assign new_n27587_ = ~new_n27755_ | ~new_n27397_ | ~new_n27398_ | ~new_n27756_;
  assign new_n27588_ = ~new_n27398_ | ~new_n27397_;
  assign new_n27589_ = ~new_n8445_ | ~new_n8773_;
  assign new_n27590_ = ~new_n27480_ | ~new_n27588_;
  assign new_n27591_ = new_n8460_ | new_n8794_;
  assign new_n27592_ = new_n8439_ | new_n8797_;
  assign new_n27593_ = ~new_n27532_ | ~new_n27361_;
  assign new_n27594_ = ~new_n8439_ | ~new_n8797_;
  assign new_n27595_ = ~new_n27482_ | ~new_n27593_;
  assign new_n27596_ = new_n8797_ | new_n8439_;
  assign new_n27597_ = ~new_n27481_ | ~new_n27499_;
  assign new_n27598_ = ~new_n27596_ | ~new_n27595_;
  assign new_n27599_ = ~new_n27522_;
  assign new_n27600_ = new_n8457_ | new_n8806_;
  assign new_n27601_ = new_n8449_ | new_n8803_;
  assign new_n27602_ = ~new_n27529_ | ~new_n27362_;
  assign new_n27603_ = ~new_n8457_ | ~new_n8806_;
  assign new_n27604_ = ~new_n27484_ | ~new_n27602_;
  assign new_n27605_ = new_n8800_ | new_n8440_;
  assign new_n27606_ = new_n8806_ | new_n8457_;
  assign new_n27607_ = ~new_n27483_ | ~new_n27522_;
  assign new_n27608_ = ~new_n27606_ | ~new_n27604_;
  assign new_n27609_ = ~new_n27521_;
  assign new_n27610_ = new_n8809_ | new_n8456_;
  assign new_n27611_ = ~new_n27610_ | ~new_n27521_;
  assign new_n27612_ = ~new_n8456_ | ~new_n8809_;
  assign new_n27613_ = ~new_n27519_;
  assign new_n27614_ = new_n8812_ | new_n8451_;
  assign new_n27615_ = ~new_n27614_ | ~new_n27519_;
  assign new_n27616_ = ~new_n8451_ | ~new_n8812_;
  assign new_n27617_ = ~new_n27447_;
  assign new_n27618_ = new_n8446_ | new_n8818_;
  assign new_n27619_ = new_n8450_ | new_n8815_;
  assign new_n27620_ = ~new_n27414_;
  assign new_n27621_ = ~new_n27415_ | ~new_n27414_;
  assign new_n27622_ = ~new_n8446_ | ~new_n27621_;
  assign new_n27623_ = ~new_n8818_ | ~new_n27620_;
  assign new_n27624_ = ~new_n27363_ | ~new_n27447_;
  assign new_n27625_ = ~new_n27517_;
  assign new_n27626_ = new_n8453_ | new_n9285_;
  assign new_n27627_ = new_n8458_ | new_n8823_;
  assign new_n27628_ = new_n8452_ | new_n9284_;
  assign new_n27629_ = ~new_n27435_;
  assign new_n27630_ = ~new_n9285_ | ~new_n27629_;
  assign new_n27631_ = ~new_n27630_ | ~new_n27445_;
  assign new_n27632_ = ~new_n27435_ | ~new_n27436_;
  assign new_n27633_ = ~new_n27632_ | ~new_n27631_;
  assign new_n27634_ = ~new_n27530_ | ~new_n27364_;
  assign new_n27635_ = ~new_n8452_ | ~new_n9284_;
  assign new_n27636_ = ~new_n27633_ | ~new_n27634_;
  assign new_n27637_ = new_n8821_ | new_n8459_;
  assign new_n27638_ = new_n9284_ | new_n8452_;
  assign new_n27639_ = ~new_n27517_ | ~new_n27486_;
  assign new_n27640_ = ~new_n27638_ | ~new_n27636_;
  assign new_n27641_ = ~new_n27514_;
  assign new_n27642_ = new_n9283_ | new_n8438_;
  assign new_n27643_ = ~new_n27642_ | ~new_n27514_;
  assign new_n27644_ = ~new_n8438_ | ~new_n9283_;
  assign new_n27645_ = ~new_n27512_;
  assign new_n27646_ = new_n9282_ | new_n8443_;
  assign new_n27647_ = ~new_n27646_ | ~new_n27512_;
  assign new_n27648_ = ~new_n8443_ | ~new_n9282_;
  assign new_n27649_ = ~new_n27510_;
  assign new_n27650_ = new_n8435_ | new_n9280_;
  assign new_n27651_ = ~new_n27531_ | ~new_n27528_;
  assign new_n27652_ = ~new_n27441_;
  assign new_n27653_ = new_n9281_ | new_n8442_;
  assign new_n27654_ = ~new_n27523_ | ~new_n27510_ | ~new_n27653_;
  assign new_n27655_ = ~new_n27508_;
  assign new_n27656_ = new_n9278_ | new_n8430_;
  assign new_n27657_ = ~new_n8430_ | ~new_n9278_;
  assign new_n27658_ = ~new_n27506_;
  assign new_n27659_ = ~new_n9277_ | ~new_n27506_;
  assign new_n27660_ = ~new_n27504_;
  assign new_n27661_ = ~new_n27653_ | ~new_n27510_;
  assign new_n27662_ = ~new_n27444_;
  assign new_n27663_ = new_n9280_ | new_n8435_;
  assign new_n27664_ = ~new_n27663_ | ~new_n27444_;
  assign new_n27665_ = ~new_n27509_ | ~new_n27664_ | ~new_n27528_;
  assign new_n27666_ = ~new_n27662_ | ~new_n27528_;
  assign new_n27667_ = ~new_n9279_ | ~new_n8434_;
  assign new_n27668_ = ~new_n27523_ | ~new_n27666_ | ~new_n27667_;
  assign new_n27669_ = new_n8435_ | new_n9280_;
  assign new_n27670_ = ~new_n27637_ | ~new_n27517_;
  assign new_n27671_ = ~new_n27446_;
  assign new_n27672_ = ~new_n27364_ | ~new_n27446_;
  assign new_n27673_ = ~new_n27490_ | ~new_n27672_;
  assign new_n27674_ = ~new_n27672_ | ~new_n27633_;
  assign new_n27675_ = ~new_n27808_ | ~new_n27674_;
  assign new_n27676_ = new_n8823_ | new_n8458_;
  assign new_n27677_ = ~new_n27676_ | ~new_n27446_;
  assign new_n27678_ = ~new_n27491_ | ~new_n27677_;
  assign new_n27679_ = ~new_n27671_ | ~new_n27435_;
  assign new_n27680_ = ~new_n8453_ | ~new_n9285_;
  assign new_n27681_ = ~new_n27492_ | ~new_n27679_;
  assign new_n27682_ = new_n8770_ | new_n8455_;
  assign new_n27683_ = ~new_n27516_;
  assign new_n27684_ = new_n8458_ | new_n8823_;
  assign new_n27685_ = new_n8815_ | new_n8450_;
  assign new_n27686_ = ~new_n27685_ | ~new_n27447_;
  assign new_n27687_ = ~new_n27493_ | ~new_n27686_;
  assign new_n27688_ = ~new_n27617_ | ~new_n27414_;
  assign new_n27689_ = ~new_n8818_ | ~new_n8446_;
  assign new_n27690_ = ~new_n27494_ | ~new_n27688_;
  assign new_n27691_ = new_n8450_ | new_n8815_;
  assign new_n27692_ = ~new_n27605_ | ~new_n27522_;
  assign new_n27693_ = ~new_n27448_;
  assign new_n27694_ = new_n8803_ | new_n8449_;
  assign new_n27695_ = ~new_n27694_ | ~new_n27448_;
  assign new_n27696_ = ~new_n27495_ | ~new_n27695_;
  assign new_n27697_ = ~new_n27693_ | ~new_n27527_;
  assign new_n27698_ = ~new_n8457_ | ~new_n8806_;
  assign new_n27699_ = ~new_n27496_ | ~new_n27697_;
  assign new_n27700_ = new_n8449_ | new_n8803_;
  assign new_n27701_ = new_n8794_ | new_n8460_;
  assign new_n27702_ = ~new_n27701_ | ~new_n27395_;
  assign new_n27703_ = ~new_n27497_ | ~new_n27702_;
  assign new_n27704_ = ~new_n27561_ | ~new_n27526_;
  assign new_n27705_ = ~new_n8439_ | ~new_n8797_;
  assign new_n27706_ = ~new_n27498_ | ~new_n27704_;
  assign new_n27707_ = ~new_n27562_ | ~new_n27526_;
  assign new_n27708_ = ~new_n27559_ | ~new_n27416_;
  assign new_n27709_ = ~new_n27569_ | ~new_n27377_;
  assign new_n27710_ = ~new_n27583_ | ~new_n27389_;
  assign new_n27711_ = ~new_n27586_ | ~new_n27535_;
  assign new_n27712_ = ~new_n27669_ | ~new_n27528_;
  assign new_n27713_ = ~new_n27653_ | ~new_n27531_;
  assign new_n27714_ = ~new_n27684_ | ~new_n27435_;
  assign new_n27715_ = ~new_n27637_ | ~new_n27432_;
  assign new_n27716_ = ~new_n27691_ | ~new_n27414_;
  assign new_n27717_ = ~new_n27700_ | ~new_n27527_;
  assign new_n27718_ = ~new_n27605_ | ~new_n27423_;
  assign new_n27719_ = ~new_n9277_ | ~new_n8431_;
  assign new_n27720_ = ~new_n27651_ | ~new_n27523_;
  assign new_n27721_ = ~new_n8434_ | ~new_n27650_;
  assign new_n27722_ = ~new_n9279_ | ~new_n27650_;
  assign new_n27723_ = ~new_n27656_ | ~new_n27651_ | ~new_n27523_;
  assign new_n27724_ = ~new_n27488_ | ~new_n27510_ | ~new_n27523_;
  assign new_n27725_ = ~new_n27652_ | ~new_n27656_;
  assign new_n27726_ = ~new_n8460_ | ~new_n27394_;
  assign new_n27727_ = ~new_n8794_ | ~new_n27393_;
  assign new_n27728_ = ~new_n27727_ | ~new_n27726_;
  assign new_n27729_ = ~new_n27707_ | ~new_n27395_;
  assign new_n27730_ = ~new_n27728_ | ~new_n27561_;
  assign new_n27731_ = ~new_n8461_ | ~new_n27391_;
  assign new_n27732_ = ~new_n8791_ | ~new_n27392_;
  assign new_n27733_ = ~new_n27732_ | ~new_n27731_;
  assign new_n27734_ = ~new_n27708_ | ~new_n27499_;
  assign new_n27735_ = ~new_n27558_ | ~new_n27733_;
  assign new_n27736_ = ~new_n8447_ | ~new_n27378_;
  assign new_n27737_ = ~new_n8788_ | ~new_n27376_;
  assign new_n27738_ = ~new_n8448_ | ~new_n27374_;
  assign new_n27739_ = ~new_n8785_ | ~new_n27375_;
  assign new_n27740_ = ~new_n27739_ | ~new_n27738_;
  assign new_n27741_ = ~new_n27709_ | ~new_n27396_;
  assign new_n27742_ = ~new_n27740_ | ~new_n27550_;
  assign new_n27743_ = ~new_n8444_ | ~new_n27390_;
  assign new_n27744_ = ~new_n8782_ | ~new_n27381_;
  assign new_n27745_ = ~new_n8437_ | ~new_n27379_;
  assign new_n27746_ = ~new_n8779_ | ~new_n27380_;
  assign new_n27747_ = ~new_n27746_ | ~new_n27745_;
  assign new_n27748_ = ~new_n27710_ | ~new_n27399_;
  assign new_n27749_ = ~new_n27747_ | ~new_n27576_;
  assign new_n27750_ = ~new_n8441_ | ~new_n27387_;
  assign new_n27751_ = ~new_n8776_ | ~new_n27388_;
  assign new_n27752_ = ~new_n27751_ | ~new_n27750_;
  assign new_n27753_ = ~new_n27711_ | ~new_n27500_;
  assign new_n27754_ = ~new_n27585_ | ~new_n27752_;
  assign new_n27755_ = ~new_n8445_ | ~new_n27382_;
  assign new_n27756_ = ~new_n8773_ | ~new_n27383_;
  assign new_n27757_ = ~new_n8432_ | ~new_n27502_;
  assign new_n27758_ = ~new_n9286_ | ~new_n27501_;
  assign new_n27759_ = ~new_n8432_ | ~new_n27502_;
  assign new_n27760_ = ~new_n9286_ | ~new_n27501_;
  assign new_n27761_ = ~new_n27760_ | ~new_n27759_;
  assign new_n27762_ = ~new_n27503_ | ~new_n27504_;
  assign new_n27763_ = ~new_n27660_ | ~new_n27761_;
  assign new_n27764_ = ~new_n8431_ | ~new_n27443_;
  assign new_n27765_ = ~new_n9277_ | ~new_n27442_;
  assign new_n27766_ = ~new_n8431_ | ~new_n27443_;
  assign new_n27767_ = ~new_n9277_ | ~new_n27442_;
  assign new_n27768_ = ~new_n27767_ | ~new_n27766_;
  assign new_n27769_ = ~new_n27505_ | ~new_n27506_;
  assign new_n27770_ = ~new_n27658_ | ~new_n27768_;
  assign new_n27771_ = ~new_n8430_ | ~new_n27401_;
  assign new_n27772_ = ~new_n9278_ | ~new_n27402_;
  assign new_n27773_ = ~new_n8430_ | ~new_n27401_;
  assign new_n27774_ = ~new_n9278_ | ~new_n27402_;
  assign new_n27775_ = ~new_n27774_ | ~new_n27773_;
  assign new_n27776_ = ~new_n27507_ | ~new_n27508_;
  assign new_n27777_ = ~new_n27655_ | ~new_n27775_;
  assign new_n27778_ = ~new_n8434_ | ~new_n27404_;
  assign new_n27779_ = ~new_n9279_ | ~new_n27403_;
  assign new_n27780_ = ~new_n8435_ | ~new_n27405_;
  assign new_n27781_ = ~new_n9280_ | ~new_n27406_;
  assign new_n27782_ = ~new_n27781_ | ~new_n27780_;
  assign new_n27783_ = ~new_n27712_ | ~new_n27444_;
  assign new_n27784_ = ~new_n27782_ | ~new_n27662_;
  assign new_n27785_ = ~new_n8442_ | ~new_n27407_;
  assign new_n27786_ = ~new_n9281_ | ~new_n27408_;
  assign new_n27787_ = ~new_n27786_ | ~new_n27785_;
  assign new_n27788_ = ~new_n27713_ | ~new_n27510_;
  assign new_n27789_ = ~new_n27649_ | ~new_n27787_;
  assign new_n27790_ = ~new_n8443_ | ~new_n27439_;
  assign new_n27791_ = ~new_n9282_ | ~new_n27440_;
  assign new_n27792_ = ~new_n8443_ | ~new_n27439_;
  assign new_n27793_ = ~new_n9282_ | ~new_n27440_;
  assign new_n27794_ = ~new_n27793_ | ~new_n27792_;
  assign new_n27795_ = ~new_n27511_ | ~new_n27512_;
  assign new_n27796_ = ~new_n27645_ | ~new_n27794_;
  assign new_n27797_ = ~new_n8438_ | ~new_n27437_;
  assign new_n27798_ = ~new_n9283_ | ~new_n27438_;
  assign new_n27799_ = ~new_n8438_ | ~new_n27437_;
  assign new_n27800_ = ~new_n9283_ | ~new_n27438_;
  assign new_n27801_ = ~new_n27800_ | ~new_n27799_;
  assign new_n27802_ = ~new_n27513_ | ~new_n27514_;
  assign new_n27803_ = ~new_n27641_ | ~new_n27801_;
  assign new_n27804_ = ~new_n8452_ | ~new_n27409_;
  assign new_n27805_ = ~new_n9284_ | ~new_n27410_;
  assign new_n27806_ = ~new_n8452_ | ~new_n27409_;
  assign new_n27807_ = ~new_n9284_ | ~new_n27410_;
  assign new_n27808_ = ~new_n27807_ | ~new_n27806_;
  assign new_n27809_ = ~new_n8453_ | ~new_n27436_;
  assign new_n27810_ = ~new_n9285_ | ~new_n27445_;
  assign new_n27811_ = ~new_n27537_ | ~new_n27516_;
  assign new_n27812_ = ~new_n27683_ | ~new_n27386_;
  assign new_n27813_ = ~new_n8458_ | ~new_n27433_;
  assign new_n27814_ = ~new_n8823_ | ~new_n27434_;
  assign new_n27815_ = ~new_n27814_ | ~new_n27813_;
  assign new_n27816_ = ~new_n27714_ | ~new_n27446_;
  assign new_n27817_ = ~new_n27815_ | ~new_n27671_;
  assign new_n27818_ = ~new_n8459_ | ~new_n27430_;
  assign new_n27819_ = ~new_n8821_ | ~new_n27431_;
  assign new_n27820_ = ~new_n27819_ | ~new_n27818_;
  assign new_n27821_ = ~new_n27715_ | ~new_n27517_;
  assign new_n27822_ = ~new_n27625_ | ~new_n27820_;
  assign new_n27823_ = ~new_n8446_ | ~new_n27415_;
  assign new_n27824_ = ~new_n8818_ | ~new_n27413_;
  assign new_n27825_ = ~new_n8450_ | ~new_n27411_;
  assign new_n27826_ = ~new_n8815_ | ~new_n27412_;
  assign new_n27827_ = ~new_n27826_ | ~new_n27825_;
  assign new_n27828_ = ~new_n27716_ | ~new_n27447_;
  assign new_n27829_ = ~new_n27827_ | ~new_n27617_;
  assign new_n27830_ = ~new_n8451_ | ~new_n27428_;
  assign new_n27831_ = ~new_n8812_ | ~new_n27429_;
  assign new_n27832_ = ~new_n8451_ | ~new_n27428_;
  assign new_n27833_ = ~new_n8812_ | ~new_n27429_;
  assign new_n27834_ = ~new_n27833_ | ~new_n27832_;
  assign new_n27835_ = ~new_n27518_ | ~new_n27519_;
  assign new_n27836_ = ~new_n27613_ | ~new_n27834_;
  assign new_n27837_ = ~new_n8456_ | ~new_n27426_;
  assign new_n27838_ = ~new_n8809_ | ~new_n27427_;
  assign new_n27839_ = ~new_n8456_ | ~new_n27426_;
  assign new_n27840_ = ~new_n8809_ | ~new_n27427_;
  assign new_n27841_ = ~new_n27840_ | ~new_n27839_;
  assign new_n27842_ = ~new_n27520_ | ~new_n27521_;
  assign new_n27843_ = ~new_n27609_ | ~new_n27841_;
  assign new_n27844_ = ~new_n8457_ | ~new_n27424_;
  assign new_n27845_ = ~new_n8806_ | ~new_n27425_;
  assign new_n27846_ = ~new_n8449_ | ~new_n27419_;
  assign new_n27847_ = ~new_n8803_ | ~new_n27420_;
  assign new_n27848_ = ~new_n27847_ | ~new_n27846_;
  assign new_n27849_ = ~new_n27717_ | ~new_n27448_;
  assign new_n27850_ = ~new_n27848_ | ~new_n27693_;
  assign new_n27851_ = ~new_n8440_ | ~new_n27421_;
  assign new_n27852_ = ~new_n8800_ | ~new_n27422_;
  assign new_n27853_ = ~new_n27852_ | ~new_n27851_;
  assign new_n27854_ = ~new_n27718_ | ~new_n27522_;
  assign new_n27855_ = ~new_n27599_ | ~new_n27853_;
  assign new_n27856_ = ~new_n8439_ | ~new_n27417_;
  assign new_n27857_ = ~new_n8797_ | ~new_n27418_;
  assign new_n27858_ = ~new_n8454_ | ~new_n27384_;
  assign new_n27859_ = ~new_n8765_ | ~new_n27385_;
  assign new_n27860_ = new_n8436_ & new_n27861_;
  assign new_n27861_ = ~new_n8433_;
  assign new_n27862_ = new_n28037_ & new_n28036_;
  assign new_n27863_ = new_n28055_ & new_n28054_;
  assign new_n27864_ = new_n28095_ & new_n28094_;
  assign new_n27865_ = new_n28104_ & new_n28103_;
  assign new_n27866_ = new_n28122_ & new_n28121_;
  assign new_n27867_ = new_n28130_ & new_n28129_;
  assign new_n27868_ = new_n28209_ & new_n28206_;
  assign new_n27869_ = new_n28202_ & new_n28199_;
  assign new_n27870_ = new_n28193_ & new_n28190_;
  assign new_n27871_ = new_n28184_ & new_n28181_;
  assign new_n27872_ = new_n28178_ & new_n28176_;
  assign new_n27873_ = new_n28171_ & new_n28168_;
  assign new_n27874_ = new_n28093_ & new_n28090_;
  assign new_n27875_ = new_n28085_ & new_n28082_;
  assign new_n27876_ = new_n28071_ & new_n28068_;
  assign new_n27877_ = ~new_n8785_;
  assign new_n27878_ = ~new_n8448_;
  assign new_n27879_ = ~new_n8447_;
  assign new_n27880_ = ~new_n8448_ | ~new_n8785_;
  assign new_n27881_ = ~new_n8788_;
  assign new_n27882_ = ~new_n8779_;
  assign new_n27883_ = ~new_n8437_;
  assign new_n27884_ = ~new_n8444_;
  assign new_n27885_ = ~new_n8773_;
  assign new_n27886_ = ~new_n8445_;
  assign new_n27887_ = ~new_n8765_;
  assign new_n27888_ = ~new_n8454_;
  assign new_n27889_ = ~new_n8454_ | ~new_n8765_;
  assign new_n27890_ = ~new_n8776_;
  assign new_n27891_ = ~new_n8441_;
  assign new_n27892_ = ~new_n8437_ | ~new_n8779_;
  assign new_n27893_ = ~new_n8782_;
  assign new_n27894_ = ~new_n8791_;
  assign new_n27895_ = ~new_n8461_;
  assign new_n27896_ = ~new_n8460_;
  assign new_n27897_ = ~new_n8794_;
  assign new_n27898_ = ~new_n27919_ | ~new_n28063_;
  assign new_n27899_ = ~new_n27975_ | ~new_n28051_;
  assign new_n27900_ = ~new_n28040_ | ~new_n28041_;
  assign new_n27901_ = ~new_n8770_ | ~new_n8455_;
  assign new_n27902_ = ~new_n27980_ | ~new_n28077_;
  assign new_n27903_ = ~new_n28074_ | ~new_n28073_;
  assign new_n27904_ = ~new_n9278_;
  assign new_n27905_ = ~new_n8430_;
  assign new_n27906_ = ~new_n8434_;
  assign new_n27907_ = ~new_n9279_;
  assign new_n27908_ = ~new_n9280_;
  assign new_n27909_ = ~new_n8435_;
  assign new_n27910_ = ~new_n9281_;
  assign new_n27911_ = ~new_n8442_;
  assign new_n27912_ = ~new_n9284_;
  assign new_n27913_ = ~new_n8452_;
  assign new_n27914_ = ~new_n8815_;
  assign new_n27915_ = ~new_n8450_;
  assign new_n27916_ = ~new_n8446_;
  assign new_n27917_ = ~new_n8450_ | ~new_n8815_;
  assign new_n27918_ = ~new_n8818_;
  assign new_n27919_ = ~new_n8461_ | ~new_n8791_;
  assign new_n27920_ = ~new_n8797_;
  assign new_n27921_ = ~new_n8439_;
  assign new_n27922_ = ~new_n8803_;
  assign new_n27923_ = ~new_n8449_;
  assign new_n27924_ = ~new_n8800_;
  assign new_n27925_ = ~new_n8440_;
  assign new_n27926_ = ~new_n8440_ | ~new_n8800_;
  assign new_n27927_ = ~new_n8806_;
  assign new_n27928_ = ~new_n8457_;
  assign new_n27929_ = ~new_n8809_;
  assign new_n27930_ = ~new_n8456_;
  assign new_n27931_ = ~new_n8812_;
  assign new_n27932_ = ~new_n8451_;
  assign new_n27933_ = ~new_n8821_;
  assign new_n27934_ = ~new_n8459_;
  assign new_n27935_ = ~new_n8459_ | ~new_n8821_;
  assign new_n27936_ = ~new_n8823_;
  assign new_n27937_ = ~new_n8458_;
  assign new_n27938_ = ~new_n8458_ | ~new_n8823_;
  assign new_n27939_ = ~new_n9285_;
  assign new_n27940_ = ~new_n9283_;
  assign new_n27941_ = ~new_n8438_;
  assign new_n27942_ = ~new_n9282_;
  assign new_n27943_ = ~new_n8443_;
  assign new_n27944_ = ~new_n9279_ | ~new_n8434_;
  assign new_n27945_ = ~new_n8431_;
  assign new_n27946_ = ~new_n9277_;
  assign new_n27947_ = ~new_n28164_ | ~new_n28034_;
  assign new_n27948_ = ~new_n8453_;
  assign new_n27949_ = ~new_n27935_ | ~new_n28173_;
  assign new_n27950_ = ~new_n28119_ | ~new_n28118_;
  assign new_n27951_ = ~new_n27926_ | ~new_n28195_;
  assign new_n27952_ = ~new_n28315_ | ~new_n28314_;
  assign new_n27953_ = ~new_n28362_ | ~new_n28361_;
  assign new_n27954_ = ~new_n28233_ | ~new_n28232_;
  assign new_n27955_ = ~new_n28238_ | ~new_n28237_;
  assign new_n27956_ = ~new_n28245_ | ~new_n28244_;
  assign new_n27957_ = ~new_n28252_ | ~new_n28251_;
  assign new_n27958_ = ~new_n28257_ | ~new_n28256_;
  assign new_n27959_ = ~new_n28266_ | ~new_n28265_;
  assign new_n27960_ = ~new_n28273_ | ~new_n28272_;
  assign new_n27961_ = ~new_n28280_ | ~new_n28279_;
  assign new_n27962_ = ~new_n28287_ | ~new_n28286_;
  assign new_n27963_ = ~new_n28292_ | ~new_n28291_;
  assign new_n27964_ = ~new_n28299_ | ~new_n28298_;
  assign new_n27965_ = ~new_n28306_ | ~new_n28305_;
  assign new_n27966_ = ~new_n28320_ | ~new_n28319_;
  assign new_n27967_ = ~new_n28325_ | ~new_n28324_;
  assign new_n27968_ = ~new_n28332_ | ~new_n28331_;
  assign new_n27969_ = ~new_n28339_ | ~new_n28338_;
  assign new_n27970_ = ~new_n28346_ | ~new_n28345_;
  assign new_n27971_ = ~new_n28353_ | ~new_n28352_;
  assign new_n27972_ = ~new_n28358_ | ~new_n28357_;
  assign new_n27973_ = new_n28047_ & new_n28045_;
  assign new_n27974_ = new_n27862_ & new_n28038_;
  assign new_n27975_ = new_n28052_ & new_n28050_;
  assign new_n27976_ = new_n28059_ & new_n28058_;
  assign new_n27977_ = new_n27880_ & new_n28240_ & new_n28239_;
  assign new_n27978_ = new_n28070_ & new_n27863_;
  assign new_n27979_ = new_n28039_ & new_n28038_;
  assign new_n27980_ = new_n28078_ & new_n28076_;
  assign new_n27981_ = new_n27892_ & new_n28247_ & new_n28246_;
  assign new_n27982_ = new_n28084_ & new_n27862_;
  assign new_n27983_ = new_n28092_ & new_n28039_;
  assign new_n27984_ = new_n28062_ & new_n27864_;
  assign new_n27985_ = new_n28097_ & new_n28029_;
  assign new_n27986_ = new_n28108_ & new_n27865_;
  assign new_n27987_ = new_n28106_ & new_n28030_;
  assign new_n27988_ = new_n28126_ & new_n28125_;
  assign new_n27989_ = new_n28131_ & new_n27867_ & new_n28140_;
  assign new_n27990_ = new_n28143_ & new_n28138_;
  assign new_n27991_ = new_n28159_ & new_n28156_;
  assign new_n27992_ = new_n28226_ & new_n28160_;
  assign new_n27993_ = new_n28018_ & new_n28136_;
  assign new_n27994_ = new_n27938_ & new_n28313_ & new_n28312_;
  assign new_n27995_ = new_n28183_ & new_n27867_;
  assign new_n27996_ = new_n27917_ & new_n28327_ & new_n28326_;
  assign new_n27997_ = new_n28192_ & new_n27866_;
  assign new_n27998_ = new_n28030_ & new_n28348_ & new_n28347_;
  assign new_n27999_ = new_n28201_ & new_n27865_;
  assign new_n28000_ = new_n28029_ & new_n28360_ & new_n28359_;
  assign new_n28001_ = new_n28208_ & new_n27864_;
  assign new_n28002_ = ~new_n27976_ | ~new_n28060_;
  assign new_n28003_ = ~new_n28075_ | ~new_n28087_;
  assign new_n28004_ = ~new_n8432_;
  assign new_n28005_ = ~new_n9286_;
  assign new_n28006_ = new_n28261_ & new_n28260_;
  assign new_n28007_ = ~new_n28222_ | ~new_n28162_ | ~new_n28027_;
  assign new_n28008_ = new_n28268_ & new_n28267_;
  assign new_n28009_ = ~new_n27992_ | ~new_n28228_ | ~new_n28227_;
  assign new_n28010_ = new_n28275_ & new_n28274_;
  assign new_n28011_ = ~new_n27944_ | ~new_n28223_ | ~new_n28157_;
  assign new_n28012_ = new_n28282_ & new_n28281_;
  assign new_n28013_ = ~new_n28151_ | ~new_n28150_;
  assign new_n28014_ = new_n28294_ & new_n28293_;
  assign new_n28015_ = ~new_n28147_ | ~new_n28146_;
  assign new_n28016_ = new_n28301_ & new_n28300_;
  assign new_n28017_ = ~new_n27990_ | ~new_n28142_;
  assign new_n28018_ = new_n28308_ & new_n28307_;
  assign new_n28019_ = ~new_n27901_ | ~new_n28185_;
  assign new_n28020_ = ~new_n27988_ | ~new_n28127_;
  assign new_n28021_ = new_n28334_ & new_n28333_;
  assign new_n28022_ = ~new_n28115_ | ~new_n28114_;
  assign new_n28023_ = new_n28341_ & new_n28340_;
  assign new_n28024_ = ~new_n28111_ | ~new_n28110_;
  assign new_n28025_ = ~new_n28101_ | ~new_n28100_;
  assign new_n28026_ = ~new_n28225_ | ~new_n28224_;
  assign new_n28027_ = ~new_n8431_ | ~new_n28009_;
  assign new_n28028_ = ~new_n27892_;
  assign new_n28029_ = ~new_n8794_ | ~new_n8460_;
  assign new_n28030_ = ~new_n8449_ | ~new_n8803_;
  assign new_n28031_ = ~new_n8435_ | ~new_n9280_;
  assign new_n28032_ = ~new_n27926_;
  assign new_n28033_ = ~new_n27935_;
  assign new_n28034_ = ~new_n8442_ | ~new_n9281_;
  assign new_n28035_ = ~new_n27919_;
  assign new_n28036_ = new_n8444_ | new_n8782_;
  assign new_n28037_ = new_n8437_ | new_n8779_;
  assign new_n28038_ = new_n8776_ | new_n8441_;
  assign new_n28039_ = new_n8773_ | new_n8445_;
  assign new_n28040_ = ~new_n27889_;
  assign new_n28041_ = new_n8770_ | new_n8455_;
  assign new_n28042_ = ~new_n27900_;
  assign new_n28043_ = ~new_n27901_;
  assign new_n28044_ = ~new_n27900_ | ~new_n27901_;
  assign new_n28045_ = ~new_n8445_ | ~new_n8773_;
  assign new_n28046_ = ~new_n28044_ | ~new_n28039_;
  assign new_n28047_ = ~new_n8441_ | ~new_n8776_;
  assign new_n28048_ = ~new_n27973_ | ~new_n28046_;
  assign new_n28049_ = ~new_n27893_ | ~new_n27892_;
  assign new_n28050_ = ~new_n8444_ | ~new_n28049_;
  assign new_n28051_ = ~new_n27974_ | ~new_n28048_;
  assign new_n28052_ = ~new_n8782_ | ~new_n28028_;
  assign new_n28053_ = ~new_n27899_;
  assign new_n28054_ = new_n8447_ | new_n8788_;
  assign new_n28055_ = new_n8448_ | new_n8785_;
  assign new_n28056_ = ~new_n27880_;
  assign new_n28057_ = ~new_n27881_ | ~new_n27880_;
  assign new_n28058_ = ~new_n8447_ | ~new_n28057_;
  assign new_n28059_ = ~new_n8788_ | ~new_n28056_;
  assign new_n28060_ = ~new_n27863_ | ~new_n27899_;
  assign new_n28061_ = ~new_n28002_;
  assign new_n28062_ = new_n8791_ | new_n8461_;
  assign new_n28063_ = ~new_n28062_ | ~new_n28002_;
  assign new_n28064_ = ~new_n27898_;
  assign new_n28065_ = new_n8460_ | new_n8794_;
  assign new_n28066_ = new_n8785_ | new_n8448_;
  assign new_n28067_ = ~new_n28066_ | ~new_n27899_;
  assign new_n28068_ = ~new_n27977_ | ~new_n28067_;
  assign new_n28069_ = ~new_n28053_ | ~new_n27880_;
  assign new_n28070_ = ~new_n8788_ | ~new_n8447_;
  assign new_n28071_ = ~new_n27978_ | ~new_n28069_;
  assign new_n28072_ = new_n8448_ | new_n8785_;
  assign new_n28073_ = ~new_n28043_ | ~new_n28039_;
  assign new_n28074_ = ~new_n8445_ | ~new_n8773_;
  assign new_n28075_ = ~new_n27903_;
  assign new_n28076_ = ~new_n27979_ | ~new_n28042_;
  assign new_n28077_ = ~new_n27903_ | ~new_n28038_;
  assign new_n28078_ = ~new_n8441_ | ~new_n8776_;
  assign new_n28079_ = ~new_n27902_;
  assign new_n28080_ = new_n8779_ | new_n8437_;
  assign new_n28081_ = ~new_n28080_ | ~new_n27902_;
  assign new_n28082_ = ~new_n27981_ | ~new_n28081_;
  assign new_n28083_ = ~new_n28079_ | ~new_n27892_;
  assign new_n28084_ = ~new_n8782_ | ~new_n8444_;
  assign new_n28085_ = ~new_n27982_ | ~new_n28083_;
  assign new_n28086_ = new_n8437_ | new_n8779_;
  assign new_n28087_ = ~new_n28042_ | ~new_n28039_;
  assign new_n28088_ = ~new_n28003_;
  assign new_n28089_ = ~new_n8441_ | ~new_n8776_;
  assign new_n28090_ = ~new_n28258_ | ~new_n27900_ | ~new_n27901_ | ~new_n28259_;
  assign new_n28091_ = ~new_n27901_ | ~new_n27900_;
  assign new_n28092_ = ~new_n8445_ | ~new_n8773_;
  assign new_n28093_ = ~new_n27983_ | ~new_n28091_;
  assign new_n28094_ = new_n8460_ | new_n8794_;
  assign new_n28095_ = new_n8439_ | new_n8797_;
  assign new_n28096_ = ~new_n28035_ | ~new_n27864_;
  assign new_n28097_ = ~new_n8439_ | ~new_n8797_;
  assign new_n28098_ = ~new_n27985_ | ~new_n28096_;
  assign new_n28099_ = new_n8797_ | new_n8439_;
  assign new_n28100_ = ~new_n27984_ | ~new_n28002_;
  assign new_n28101_ = ~new_n28099_ | ~new_n28098_;
  assign new_n28102_ = ~new_n28025_;
  assign new_n28103_ = new_n8457_ | new_n8806_;
  assign new_n28104_ = new_n8449_ | new_n8803_;
  assign new_n28105_ = ~new_n28032_ | ~new_n27865_;
  assign new_n28106_ = ~new_n8457_ | ~new_n8806_;
  assign new_n28107_ = ~new_n27987_ | ~new_n28105_;
  assign new_n28108_ = new_n8800_ | new_n8440_;
  assign new_n28109_ = new_n8806_ | new_n8457_;
  assign new_n28110_ = ~new_n27986_ | ~new_n28025_;
  assign new_n28111_ = ~new_n28109_ | ~new_n28107_;
  assign new_n28112_ = ~new_n28024_;
  assign new_n28113_ = new_n8809_ | new_n8456_;
  assign new_n28114_ = ~new_n28113_ | ~new_n28024_;
  assign new_n28115_ = ~new_n8456_ | ~new_n8809_;
  assign new_n28116_ = ~new_n28022_;
  assign new_n28117_ = new_n8812_ | new_n8451_;
  assign new_n28118_ = ~new_n28117_ | ~new_n28022_;
  assign new_n28119_ = ~new_n8451_ | ~new_n8812_;
  assign new_n28120_ = ~new_n27950_;
  assign new_n28121_ = new_n8446_ | new_n8818_;
  assign new_n28122_ = new_n8450_ | new_n8815_;
  assign new_n28123_ = ~new_n27917_;
  assign new_n28124_ = ~new_n27918_ | ~new_n27917_;
  assign new_n28125_ = ~new_n8446_ | ~new_n28124_;
  assign new_n28126_ = ~new_n8818_ | ~new_n28123_;
  assign new_n28127_ = ~new_n27866_ | ~new_n27950_;
  assign new_n28128_ = ~new_n28020_;
  assign new_n28129_ = new_n8453_ | new_n9285_;
  assign new_n28130_ = new_n8458_ | new_n8823_;
  assign new_n28131_ = new_n8452_ | new_n9284_;
  assign new_n28132_ = ~new_n27938_;
  assign new_n28133_ = ~new_n9285_ | ~new_n28132_;
  assign new_n28134_ = ~new_n28133_ | ~new_n27948_;
  assign new_n28135_ = ~new_n27938_ | ~new_n27939_;
  assign new_n28136_ = ~new_n28135_ | ~new_n28134_;
  assign new_n28137_ = ~new_n28033_ | ~new_n27867_;
  assign new_n28138_ = ~new_n8452_ | ~new_n9284_;
  assign new_n28139_ = ~new_n28136_ | ~new_n28137_;
  assign new_n28140_ = new_n8821_ | new_n8459_;
  assign new_n28141_ = new_n9284_ | new_n8452_;
  assign new_n28142_ = ~new_n28020_ | ~new_n27989_;
  assign new_n28143_ = ~new_n28141_ | ~new_n28139_;
  assign new_n28144_ = ~new_n28017_;
  assign new_n28145_ = new_n9283_ | new_n8438_;
  assign new_n28146_ = ~new_n28145_ | ~new_n28017_;
  assign new_n28147_ = ~new_n8438_ | ~new_n9283_;
  assign new_n28148_ = ~new_n28015_;
  assign new_n28149_ = new_n9282_ | new_n8443_;
  assign new_n28150_ = ~new_n28149_ | ~new_n28015_;
  assign new_n28151_ = ~new_n8443_ | ~new_n9282_;
  assign new_n28152_ = ~new_n28013_;
  assign new_n28153_ = new_n8435_ | new_n9280_;
  assign new_n28154_ = ~new_n28034_ | ~new_n28031_;
  assign new_n28155_ = ~new_n27944_;
  assign new_n28156_ = new_n9281_ | new_n8442_;
  assign new_n28157_ = ~new_n28026_ | ~new_n28013_ | ~new_n28156_;
  assign new_n28158_ = ~new_n28011_;
  assign new_n28159_ = new_n9278_ | new_n8430_;
  assign new_n28160_ = ~new_n8430_ | ~new_n9278_;
  assign new_n28161_ = ~new_n28009_;
  assign new_n28162_ = ~new_n9277_ | ~new_n28009_;
  assign new_n28163_ = ~new_n28007_;
  assign new_n28164_ = ~new_n28156_ | ~new_n28013_;
  assign new_n28165_ = ~new_n27947_;
  assign new_n28166_ = new_n9280_ | new_n8435_;
  assign new_n28167_ = ~new_n28166_ | ~new_n27947_;
  assign new_n28168_ = ~new_n28012_ | ~new_n28167_ | ~new_n28031_;
  assign new_n28169_ = ~new_n28165_ | ~new_n28031_;
  assign new_n28170_ = ~new_n9279_ | ~new_n8434_;
  assign new_n28171_ = ~new_n28026_ | ~new_n28169_ | ~new_n28170_;
  assign new_n28172_ = new_n8435_ | new_n9280_;
  assign new_n28173_ = ~new_n28140_ | ~new_n28020_;
  assign new_n28174_ = ~new_n27949_;
  assign new_n28175_ = ~new_n27867_ | ~new_n27949_;
  assign new_n28176_ = ~new_n27993_ | ~new_n28175_;
  assign new_n28177_ = ~new_n28175_ | ~new_n28136_;
  assign new_n28178_ = ~new_n28311_ | ~new_n28177_;
  assign new_n28179_ = new_n8823_ | new_n8458_;
  assign new_n28180_ = ~new_n28179_ | ~new_n27949_;
  assign new_n28181_ = ~new_n27994_ | ~new_n28180_;
  assign new_n28182_ = ~new_n28174_ | ~new_n27938_;
  assign new_n28183_ = ~new_n8453_ | ~new_n9285_;
  assign new_n28184_ = ~new_n27995_ | ~new_n28182_;
  assign new_n28185_ = new_n8770_ | new_n8455_;
  assign new_n28186_ = ~new_n28019_;
  assign new_n28187_ = new_n8458_ | new_n8823_;
  assign new_n28188_ = new_n8815_ | new_n8450_;
  assign new_n28189_ = ~new_n28188_ | ~new_n27950_;
  assign new_n28190_ = ~new_n27996_ | ~new_n28189_;
  assign new_n28191_ = ~new_n28120_ | ~new_n27917_;
  assign new_n28192_ = ~new_n8818_ | ~new_n8446_;
  assign new_n28193_ = ~new_n27997_ | ~new_n28191_;
  assign new_n28194_ = new_n8450_ | new_n8815_;
  assign new_n28195_ = ~new_n28108_ | ~new_n28025_;
  assign new_n28196_ = ~new_n27951_;
  assign new_n28197_ = new_n8803_ | new_n8449_;
  assign new_n28198_ = ~new_n28197_ | ~new_n27951_;
  assign new_n28199_ = ~new_n27998_ | ~new_n28198_;
  assign new_n28200_ = ~new_n28196_ | ~new_n28030_;
  assign new_n28201_ = ~new_n8457_ | ~new_n8806_;
  assign new_n28202_ = ~new_n27999_ | ~new_n28200_;
  assign new_n28203_ = new_n8449_ | new_n8803_;
  assign new_n28204_ = new_n8794_ | new_n8460_;
  assign new_n28205_ = ~new_n28204_ | ~new_n27898_;
  assign new_n28206_ = ~new_n28000_ | ~new_n28205_;
  assign new_n28207_ = ~new_n28064_ | ~new_n28029_;
  assign new_n28208_ = ~new_n8439_ | ~new_n8797_;
  assign new_n28209_ = ~new_n28001_ | ~new_n28207_;
  assign new_n28210_ = ~new_n28065_ | ~new_n28029_;
  assign new_n28211_ = ~new_n28062_ | ~new_n27919_;
  assign new_n28212_ = ~new_n28072_ | ~new_n27880_;
  assign new_n28213_ = ~new_n28086_ | ~new_n27892_;
  assign new_n28214_ = ~new_n28089_ | ~new_n28038_;
  assign new_n28215_ = ~new_n28172_ | ~new_n28031_;
  assign new_n28216_ = ~new_n28156_ | ~new_n28034_;
  assign new_n28217_ = ~new_n28187_ | ~new_n27938_;
  assign new_n28218_ = ~new_n28140_ | ~new_n27935_;
  assign new_n28219_ = ~new_n28194_ | ~new_n27917_;
  assign new_n28220_ = ~new_n28203_ | ~new_n28030_;
  assign new_n28221_ = ~new_n28108_ | ~new_n27926_;
  assign new_n28222_ = ~new_n9277_ | ~new_n8431_;
  assign new_n28223_ = ~new_n28154_ | ~new_n28026_;
  assign new_n28224_ = ~new_n8434_ | ~new_n28153_;
  assign new_n28225_ = ~new_n9279_ | ~new_n28153_;
  assign new_n28226_ = ~new_n28159_ | ~new_n28154_ | ~new_n28026_;
  assign new_n28227_ = ~new_n27991_ | ~new_n28013_ | ~new_n28026_;
  assign new_n28228_ = ~new_n28155_ | ~new_n28159_;
  assign new_n28229_ = ~new_n8460_ | ~new_n27897_;
  assign new_n28230_ = ~new_n8794_ | ~new_n27896_;
  assign new_n28231_ = ~new_n28230_ | ~new_n28229_;
  assign new_n28232_ = ~new_n28210_ | ~new_n27898_;
  assign new_n28233_ = ~new_n28231_ | ~new_n28064_;
  assign new_n28234_ = ~new_n8461_ | ~new_n27894_;
  assign new_n28235_ = ~new_n8791_ | ~new_n27895_;
  assign new_n28236_ = ~new_n28235_ | ~new_n28234_;
  assign new_n28237_ = ~new_n28211_ | ~new_n28002_;
  assign new_n28238_ = ~new_n28061_ | ~new_n28236_;
  assign new_n28239_ = ~new_n8447_ | ~new_n27881_;
  assign new_n28240_ = ~new_n8788_ | ~new_n27879_;
  assign new_n28241_ = ~new_n8448_ | ~new_n27877_;
  assign new_n28242_ = ~new_n8785_ | ~new_n27878_;
  assign new_n28243_ = ~new_n28242_ | ~new_n28241_;
  assign new_n28244_ = ~new_n28212_ | ~new_n27899_;
  assign new_n28245_ = ~new_n28243_ | ~new_n28053_;
  assign new_n28246_ = ~new_n8444_ | ~new_n27893_;
  assign new_n28247_ = ~new_n8782_ | ~new_n27884_;
  assign new_n28248_ = ~new_n8437_ | ~new_n27882_;
  assign new_n28249_ = ~new_n8779_ | ~new_n27883_;
  assign new_n28250_ = ~new_n28249_ | ~new_n28248_;
  assign new_n28251_ = ~new_n28213_ | ~new_n27902_;
  assign new_n28252_ = ~new_n28250_ | ~new_n28079_;
  assign new_n28253_ = ~new_n8441_ | ~new_n27890_;
  assign new_n28254_ = ~new_n8776_ | ~new_n27891_;
  assign new_n28255_ = ~new_n28254_ | ~new_n28253_;
  assign new_n28256_ = ~new_n28214_ | ~new_n28003_;
  assign new_n28257_ = ~new_n28088_ | ~new_n28255_;
  assign new_n28258_ = ~new_n8445_ | ~new_n27885_;
  assign new_n28259_ = ~new_n8773_ | ~new_n27886_;
  assign new_n28260_ = ~new_n8432_ | ~new_n28005_;
  assign new_n28261_ = ~new_n9286_ | ~new_n28004_;
  assign new_n28262_ = ~new_n8432_ | ~new_n28005_;
  assign new_n28263_ = ~new_n9286_ | ~new_n28004_;
  assign new_n28264_ = ~new_n28263_ | ~new_n28262_;
  assign new_n28265_ = ~new_n28006_ | ~new_n28007_;
  assign new_n28266_ = ~new_n28163_ | ~new_n28264_;
  assign new_n28267_ = ~new_n8431_ | ~new_n27946_;
  assign new_n28268_ = ~new_n9277_ | ~new_n27945_;
  assign new_n28269_ = ~new_n8431_ | ~new_n27946_;
  assign new_n28270_ = ~new_n9277_ | ~new_n27945_;
  assign new_n28271_ = ~new_n28270_ | ~new_n28269_;
  assign new_n28272_ = ~new_n28008_ | ~new_n28009_;
  assign new_n28273_ = ~new_n28161_ | ~new_n28271_;
  assign new_n28274_ = ~new_n8430_ | ~new_n27904_;
  assign new_n28275_ = ~new_n9278_ | ~new_n27905_;
  assign new_n28276_ = ~new_n8430_ | ~new_n27904_;
  assign new_n28277_ = ~new_n9278_ | ~new_n27905_;
  assign new_n28278_ = ~new_n28277_ | ~new_n28276_;
  assign new_n28279_ = ~new_n28010_ | ~new_n28011_;
  assign new_n28280_ = ~new_n28158_ | ~new_n28278_;
  assign new_n28281_ = ~new_n8434_ | ~new_n27907_;
  assign new_n28282_ = ~new_n9279_ | ~new_n27906_;
  assign new_n28283_ = ~new_n8435_ | ~new_n27908_;
  assign new_n28284_ = ~new_n9280_ | ~new_n27909_;
  assign new_n28285_ = ~new_n28284_ | ~new_n28283_;
  assign new_n28286_ = ~new_n28215_ | ~new_n27947_;
  assign new_n28287_ = ~new_n28285_ | ~new_n28165_;
  assign new_n28288_ = ~new_n8442_ | ~new_n27910_;
  assign new_n28289_ = ~new_n9281_ | ~new_n27911_;
  assign new_n28290_ = ~new_n28289_ | ~new_n28288_;
  assign new_n28291_ = ~new_n28216_ | ~new_n28013_;
  assign new_n28292_ = ~new_n28152_ | ~new_n28290_;
  assign new_n28293_ = ~new_n8443_ | ~new_n27942_;
  assign new_n28294_ = ~new_n9282_ | ~new_n27943_;
  assign new_n28295_ = ~new_n8443_ | ~new_n27942_;
  assign new_n28296_ = ~new_n9282_ | ~new_n27943_;
  assign new_n28297_ = ~new_n28296_ | ~new_n28295_;
  assign new_n28298_ = ~new_n28014_ | ~new_n28015_;
  assign new_n28299_ = ~new_n28148_ | ~new_n28297_;
  assign new_n28300_ = ~new_n8438_ | ~new_n27940_;
  assign new_n28301_ = ~new_n9283_ | ~new_n27941_;
  assign new_n28302_ = ~new_n8438_ | ~new_n27940_;
  assign new_n28303_ = ~new_n9283_ | ~new_n27941_;
  assign new_n28304_ = ~new_n28303_ | ~new_n28302_;
  assign new_n28305_ = ~new_n28016_ | ~new_n28017_;
  assign new_n28306_ = ~new_n28144_ | ~new_n28304_;
  assign new_n28307_ = ~new_n8452_ | ~new_n27912_;
  assign new_n28308_ = ~new_n9284_ | ~new_n27913_;
  assign new_n28309_ = ~new_n8452_ | ~new_n27912_;
  assign new_n28310_ = ~new_n9284_ | ~new_n27913_;
  assign new_n28311_ = ~new_n28310_ | ~new_n28309_;
  assign new_n28312_ = ~new_n8453_ | ~new_n27939_;
  assign new_n28313_ = ~new_n9285_ | ~new_n27948_;
  assign new_n28314_ = ~new_n28040_ | ~new_n28019_;
  assign new_n28315_ = ~new_n28186_ | ~new_n27889_;
  assign new_n28316_ = ~new_n8458_ | ~new_n27936_;
  assign new_n28317_ = ~new_n8823_ | ~new_n27937_;
  assign new_n28318_ = ~new_n28317_ | ~new_n28316_;
  assign new_n28319_ = ~new_n28217_ | ~new_n27949_;
  assign new_n28320_ = ~new_n28318_ | ~new_n28174_;
  assign new_n28321_ = ~new_n8459_ | ~new_n27933_;
  assign new_n28322_ = ~new_n8821_ | ~new_n27934_;
  assign new_n28323_ = ~new_n28322_ | ~new_n28321_;
  assign new_n28324_ = ~new_n28218_ | ~new_n28020_;
  assign new_n28325_ = ~new_n28128_ | ~new_n28323_;
  assign new_n28326_ = ~new_n8446_ | ~new_n27918_;
  assign new_n28327_ = ~new_n8818_ | ~new_n27916_;
  assign new_n28328_ = ~new_n8450_ | ~new_n27914_;
  assign new_n28329_ = ~new_n8815_ | ~new_n27915_;
  assign new_n28330_ = ~new_n28329_ | ~new_n28328_;
  assign new_n28331_ = ~new_n28219_ | ~new_n27950_;
  assign new_n28332_ = ~new_n28330_ | ~new_n28120_;
  assign new_n28333_ = ~new_n8451_ | ~new_n27931_;
  assign new_n28334_ = ~new_n8812_ | ~new_n27932_;
  assign new_n28335_ = ~new_n8451_ | ~new_n27931_;
  assign new_n28336_ = ~new_n8812_ | ~new_n27932_;
  assign new_n28337_ = ~new_n28336_ | ~new_n28335_;
  assign new_n28338_ = ~new_n28021_ | ~new_n28022_;
  assign new_n28339_ = ~new_n28116_ | ~new_n28337_;
  assign new_n28340_ = ~new_n8456_ | ~new_n27929_;
  assign new_n28341_ = ~new_n8809_ | ~new_n27930_;
  assign new_n28342_ = ~new_n8456_ | ~new_n27929_;
  assign new_n28343_ = ~new_n8809_ | ~new_n27930_;
  assign new_n28344_ = ~new_n28343_ | ~new_n28342_;
  assign new_n28345_ = ~new_n28023_ | ~new_n28024_;
  assign new_n28346_ = ~new_n28112_ | ~new_n28344_;
  assign new_n28347_ = ~new_n8457_ | ~new_n27927_;
  assign new_n28348_ = ~new_n8806_ | ~new_n27928_;
  assign new_n28349_ = ~new_n8449_ | ~new_n27922_;
  assign new_n28350_ = ~new_n8803_ | ~new_n27923_;
  assign new_n28351_ = ~new_n28350_ | ~new_n28349_;
  assign new_n28352_ = ~new_n28220_ | ~new_n27951_;
  assign new_n28353_ = ~new_n28351_ | ~new_n28196_;
  assign new_n28354_ = ~new_n8440_ | ~new_n27924_;
  assign new_n28355_ = ~new_n8800_ | ~new_n27925_;
  assign new_n28356_ = ~new_n28355_ | ~new_n28354_;
  assign new_n28357_ = ~new_n28221_ | ~new_n28025_;
  assign new_n28358_ = ~new_n28102_ | ~new_n28356_;
  assign new_n28359_ = ~new_n8439_ | ~new_n27920_;
  assign new_n28360_ = ~new_n8797_ | ~new_n27921_;
  assign new_n28361_ = ~new_n8454_ | ~new_n27887_;
  assign new_n28362_ = ~new_n8765_ | ~new_n27888_;
  assign new_n28363_ = new_n28538_ & new_n28537_;
  assign new_n28364_ = new_n28556_ & new_n28555_;
  assign new_n28365_ = new_n28596_ & new_n28595_;
  assign new_n28366_ = new_n28605_ & new_n28604_;
  assign new_n28367_ = new_n28623_ & new_n28622_;
  assign new_n28368_ = new_n28631_ & new_n28630_;
  assign new_n28369_ = new_n28710_ & new_n28707_;
  assign new_n28370_ = new_n28703_ & new_n28700_;
  assign new_n28371_ = new_n28694_ & new_n28691_;
  assign new_n28372_ = new_n28685_ & new_n28682_;
  assign new_n28373_ = new_n28679_ & new_n28677_;
  assign new_n28374_ = new_n28672_ & new_n28669_;
  assign new_n28375_ = new_n28594_ & new_n28591_;
  assign new_n28376_ = new_n28586_ & new_n28583_;
  assign new_n28377_ = new_n28572_ & new_n28569_;
  assign new_n28378_ = ~new_n8785_;
  assign new_n28379_ = ~new_n8448_;
  assign new_n28380_ = ~new_n8447_;
  assign new_n28381_ = ~new_n8448_ | ~new_n8785_;
  assign new_n28382_ = ~new_n8788_;
  assign new_n28383_ = ~new_n8779_;
  assign new_n28384_ = ~new_n8437_;
  assign new_n28385_ = ~new_n8444_;
  assign new_n28386_ = ~new_n8773_;
  assign new_n28387_ = ~new_n8445_;
  assign new_n28388_ = ~new_n8765_;
  assign new_n28389_ = ~new_n8454_;
  assign new_n28390_ = ~new_n8454_ | ~new_n8765_;
  assign new_n28391_ = ~new_n8776_;
  assign new_n28392_ = ~new_n8441_;
  assign new_n28393_ = ~new_n8437_ | ~new_n8779_;
  assign new_n28394_ = ~new_n8782_;
  assign new_n28395_ = ~new_n8791_;
  assign new_n28396_ = ~new_n8461_;
  assign new_n28397_ = ~new_n8460_;
  assign new_n28398_ = ~new_n8794_;
  assign new_n28399_ = ~new_n28422_ | ~new_n28564_;
  assign new_n28400_ = ~new_n28476_ | ~new_n28552_;
  assign new_n28401_ = ~new_n28541_ | ~new_n28542_;
  assign new_n28402_ = ~new_n8770_ | ~new_n8455_;
  assign new_n28403_ = ~new_n28481_ | ~new_n28578_;
  assign new_n28404_ = ~new_n28575_ | ~new_n28574_;
  assign new_n28405_ = ~new_n9278_;
  assign new_n28406_ = ~new_n8430_;
  assign new_n28407_ = ~new_n8434_;
  assign new_n28408_ = ~new_n9279_;
  assign new_n28409_ = ~new_n9280_;
  assign new_n28410_ = ~new_n8435_;
  assign new_n28411_ = ~new_n9281_;
  assign new_n28412_ = ~new_n8442_;
  assign new_n28413_ = ~new_n9284_;
  assign new_n28414_ = ~new_n8452_;
  assign new_n28415_ = ~new_n8815_;
  assign new_n28416_ = ~new_n8450_;
  assign new_n28417_ = ~new_n8446_;
  assign new_n28418_ = ~new_n8450_ | ~new_n8815_;
  assign new_n28419_ = ~new_n8818_;
  assign new_n28420_ = ~new_n8797_;
  assign new_n28421_ = ~new_n8439_;
  assign new_n28422_ = ~new_n8461_ | ~new_n8791_;
  assign new_n28423_ = ~new_n8803_;
  assign new_n28424_ = ~new_n8449_;
  assign new_n28425_ = ~new_n8800_;
  assign new_n28426_ = ~new_n8440_;
  assign new_n28427_ = ~new_n8440_ | ~new_n8800_;
  assign new_n28428_ = ~new_n8806_;
  assign new_n28429_ = ~new_n8457_;
  assign new_n28430_ = ~new_n8809_;
  assign new_n28431_ = ~new_n8456_;
  assign new_n28432_ = ~new_n8812_;
  assign new_n28433_ = ~new_n8451_;
  assign new_n28434_ = ~new_n8821_;
  assign new_n28435_ = ~new_n8459_;
  assign new_n28436_ = ~new_n8459_ | ~new_n8821_;
  assign new_n28437_ = ~new_n8823_;
  assign new_n28438_ = ~new_n8458_;
  assign new_n28439_ = ~new_n8458_ | ~new_n8823_;
  assign new_n28440_ = ~new_n9285_;
  assign new_n28441_ = ~new_n9283_;
  assign new_n28442_ = ~new_n8438_;
  assign new_n28443_ = ~new_n9282_;
  assign new_n28444_ = ~new_n8443_;
  assign new_n28445_ = ~new_n9279_ | ~new_n8434_;
  assign new_n28446_ = ~new_n8431_;
  assign new_n28447_ = ~new_n9277_;
  assign new_n28448_ = ~new_n28665_ | ~new_n28535_;
  assign new_n28449_ = ~new_n8453_;
  assign new_n28450_ = ~new_n28436_ | ~new_n28674_;
  assign new_n28451_ = ~new_n28620_ | ~new_n28619_;
  assign new_n28452_ = ~new_n28427_ | ~new_n28696_;
  assign new_n28453_ = ~new_n28816_ | ~new_n28815_;
  assign new_n28454_ = ~new_n28863_ | ~new_n28862_;
  assign new_n28455_ = ~new_n28734_ | ~new_n28733_;
  assign new_n28456_ = ~new_n28739_ | ~new_n28738_;
  assign new_n28457_ = ~new_n28746_ | ~new_n28745_;
  assign new_n28458_ = ~new_n28753_ | ~new_n28752_;
  assign new_n28459_ = ~new_n28758_ | ~new_n28757_;
  assign new_n28460_ = ~new_n28767_ | ~new_n28766_;
  assign new_n28461_ = ~new_n28774_ | ~new_n28773_;
  assign new_n28462_ = ~new_n28781_ | ~new_n28780_;
  assign new_n28463_ = ~new_n28788_ | ~new_n28787_;
  assign new_n28464_ = ~new_n28793_ | ~new_n28792_;
  assign new_n28465_ = ~new_n28800_ | ~new_n28799_;
  assign new_n28466_ = ~new_n28807_ | ~new_n28806_;
  assign new_n28467_ = ~new_n28821_ | ~new_n28820_;
  assign new_n28468_ = ~new_n28826_ | ~new_n28825_;
  assign new_n28469_ = ~new_n28833_ | ~new_n28832_;
  assign new_n28470_ = ~new_n28840_ | ~new_n28839_;
  assign new_n28471_ = ~new_n28847_ | ~new_n28846_;
  assign new_n28472_ = ~new_n28854_ | ~new_n28853_;
  assign new_n28473_ = ~new_n28859_ | ~new_n28858_;
  assign new_n28474_ = new_n28548_ & new_n28546_;
  assign new_n28475_ = new_n28363_ & new_n28539_;
  assign new_n28476_ = new_n28553_ & new_n28551_;
  assign new_n28477_ = new_n28560_ & new_n28559_;
  assign new_n28478_ = new_n28381_ & new_n28741_ & new_n28740_;
  assign new_n28479_ = new_n28571_ & new_n28364_;
  assign new_n28480_ = new_n28540_ & new_n28539_;
  assign new_n28481_ = new_n28579_ & new_n28577_;
  assign new_n28482_ = new_n28393_ & new_n28748_ & new_n28747_;
  assign new_n28483_ = new_n28585_ & new_n28363_;
  assign new_n28484_ = new_n28593_ & new_n28540_;
  assign new_n28485_ = new_n28563_ & new_n28365_;
  assign new_n28486_ = new_n28602_ & new_n28598_;
  assign new_n28487_ = new_n28609_ & new_n28366_;
  assign new_n28488_ = new_n28607_ & new_n28531_;
  assign new_n28489_ = new_n28627_ & new_n28626_;
  assign new_n28490_ = new_n28632_ & new_n28368_ & new_n28641_;
  assign new_n28491_ = new_n28644_ & new_n28639_;
  assign new_n28492_ = new_n28660_ & new_n28657_;
  assign new_n28493_ = new_n28727_ & new_n28661_;
  assign new_n28494_ = new_n28519_ & new_n28637_;
  assign new_n28495_ = new_n28439_ & new_n28814_ & new_n28813_;
  assign new_n28496_ = new_n28684_ & new_n28368_;
  assign new_n28497_ = new_n28418_ & new_n28828_ & new_n28827_;
  assign new_n28498_ = new_n28693_ & new_n28367_;
  assign new_n28499_ = new_n28531_ & new_n28849_ & new_n28848_;
  assign new_n28500_ = new_n28702_ & new_n28366_;
  assign new_n28501_ = new_n28530_ & new_n28861_ & new_n28860_;
  assign new_n28502_ = new_n28709_ & new_n28365_;
  assign new_n28503_ = ~new_n28477_ | ~new_n28561_;
  assign new_n28504_ = ~new_n28576_ | ~new_n28588_;
  assign new_n28505_ = ~new_n8432_;
  assign new_n28506_ = ~new_n9286_;
  assign new_n28507_ = new_n28762_ & new_n28761_;
  assign new_n28508_ = ~new_n28723_ | ~new_n28663_ | ~new_n28528_;
  assign new_n28509_ = new_n28769_ & new_n28768_;
  assign new_n28510_ = ~new_n28493_ | ~new_n28729_ | ~new_n28728_;
  assign new_n28511_ = new_n28776_ & new_n28775_;
  assign new_n28512_ = ~new_n28445_ | ~new_n28724_ | ~new_n28658_;
  assign new_n28513_ = new_n28783_ & new_n28782_;
  assign new_n28514_ = ~new_n28652_ | ~new_n28651_;
  assign new_n28515_ = new_n28795_ & new_n28794_;
  assign new_n28516_ = ~new_n28648_ | ~new_n28647_;
  assign new_n28517_ = new_n28802_ & new_n28801_;
  assign new_n28518_ = ~new_n28491_ | ~new_n28643_;
  assign new_n28519_ = new_n28809_ & new_n28808_;
  assign new_n28520_ = ~new_n28402_ | ~new_n28686_;
  assign new_n28521_ = ~new_n28489_ | ~new_n28628_;
  assign new_n28522_ = new_n28835_ & new_n28834_;
  assign new_n28523_ = ~new_n28616_ | ~new_n28615_;
  assign new_n28524_ = new_n28842_ & new_n28841_;
  assign new_n28525_ = ~new_n28612_ | ~new_n28611_;
  assign new_n28526_ = ~new_n28486_ | ~new_n28601_;
  assign new_n28527_ = ~new_n28726_ | ~new_n28725_;
  assign new_n28528_ = ~new_n8431_ | ~new_n28510_;
  assign new_n28529_ = ~new_n28393_;
  assign new_n28530_ = ~new_n8794_ | ~new_n8460_;
  assign new_n28531_ = ~new_n8449_ | ~new_n8803_;
  assign new_n28532_ = ~new_n8435_ | ~new_n9280_;
  assign new_n28533_ = ~new_n28427_;
  assign new_n28534_ = ~new_n28436_;
  assign new_n28535_ = ~new_n8442_ | ~new_n9281_;
  assign new_n28536_ = ~new_n28422_;
  assign new_n28537_ = new_n8444_ | new_n8782_;
  assign new_n28538_ = new_n8437_ | new_n8779_;
  assign new_n28539_ = new_n8776_ | new_n8441_;
  assign new_n28540_ = new_n8773_ | new_n8445_;
  assign new_n28541_ = ~new_n28390_;
  assign new_n28542_ = new_n8770_ | new_n8455_;
  assign new_n28543_ = ~new_n28401_;
  assign new_n28544_ = ~new_n28402_;
  assign new_n28545_ = ~new_n28401_ | ~new_n28402_;
  assign new_n28546_ = ~new_n8445_ | ~new_n8773_;
  assign new_n28547_ = ~new_n28545_ | ~new_n28540_;
  assign new_n28548_ = ~new_n8441_ | ~new_n8776_;
  assign new_n28549_ = ~new_n28474_ | ~new_n28547_;
  assign new_n28550_ = ~new_n28394_ | ~new_n28393_;
  assign new_n28551_ = ~new_n8444_ | ~new_n28550_;
  assign new_n28552_ = ~new_n28475_ | ~new_n28549_;
  assign new_n28553_ = ~new_n8782_ | ~new_n28529_;
  assign new_n28554_ = ~new_n28400_;
  assign new_n28555_ = new_n8447_ | new_n8788_;
  assign new_n28556_ = new_n8448_ | new_n8785_;
  assign new_n28557_ = ~new_n28381_;
  assign new_n28558_ = ~new_n28382_ | ~new_n28381_;
  assign new_n28559_ = ~new_n8447_ | ~new_n28558_;
  assign new_n28560_ = ~new_n8788_ | ~new_n28557_;
  assign new_n28561_ = ~new_n28364_ | ~new_n28400_;
  assign new_n28562_ = ~new_n28503_;
  assign new_n28563_ = new_n8791_ | new_n8461_;
  assign new_n28564_ = ~new_n28563_ | ~new_n28503_;
  assign new_n28565_ = ~new_n28399_;
  assign new_n28566_ = new_n8460_ | new_n8794_;
  assign new_n28567_ = new_n8785_ | new_n8448_;
  assign new_n28568_ = ~new_n28567_ | ~new_n28400_;
  assign new_n28569_ = ~new_n28478_ | ~new_n28568_;
  assign new_n28570_ = ~new_n28554_ | ~new_n28381_;
  assign new_n28571_ = ~new_n8788_ | ~new_n8447_;
  assign new_n28572_ = ~new_n28479_ | ~new_n28570_;
  assign new_n28573_ = new_n8448_ | new_n8785_;
  assign new_n28574_ = ~new_n28544_ | ~new_n28540_;
  assign new_n28575_ = ~new_n8445_ | ~new_n8773_;
  assign new_n28576_ = ~new_n28404_;
  assign new_n28577_ = ~new_n28480_ | ~new_n28543_;
  assign new_n28578_ = ~new_n28404_ | ~new_n28539_;
  assign new_n28579_ = ~new_n8441_ | ~new_n8776_;
  assign new_n28580_ = ~new_n28403_;
  assign new_n28581_ = new_n8779_ | new_n8437_;
  assign new_n28582_ = ~new_n28581_ | ~new_n28403_;
  assign new_n28583_ = ~new_n28482_ | ~new_n28582_;
  assign new_n28584_ = ~new_n28580_ | ~new_n28393_;
  assign new_n28585_ = ~new_n8782_ | ~new_n8444_;
  assign new_n28586_ = ~new_n28483_ | ~new_n28584_;
  assign new_n28587_ = new_n8437_ | new_n8779_;
  assign new_n28588_ = ~new_n28543_ | ~new_n28540_;
  assign new_n28589_ = ~new_n28504_;
  assign new_n28590_ = ~new_n8441_ | ~new_n8776_;
  assign new_n28591_ = ~new_n28759_ | ~new_n28401_ | ~new_n28402_ | ~new_n28760_;
  assign new_n28592_ = ~new_n28402_ | ~new_n28401_;
  assign new_n28593_ = ~new_n8445_ | ~new_n8773_;
  assign new_n28594_ = ~new_n28484_ | ~new_n28592_;
  assign new_n28595_ = new_n8460_ | new_n8794_;
  assign new_n28596_ = new_n8439_ | new_n8797_;
  assign new_n28597_ = ~new_n28536_ | ~new_n28365_;
  assign new_n28598_ = ~new_n8439_ | ~new_n8797_;
  assign new_n28599_ = ~new_n28530_ | ~new_n28597_;
  assign new_n28600_ = new_n8797_ | new_n8439_;
  assign new_n28601_ = ~new_n28485_ | ~new_n28503_;
  assign new_n28602_ = ~new_n28600_ | ~new_n28599_;
  assign new_n28603_ = ~new_n28526_;
  assign new_n28604_ = new_n8457_ | new_n8806_;
  assign new_n28605_ = new_n8449_ | new_n8803_;
  assign new_n28606_ = ~new_n28533_ | ~new_n28366_;
  assign new_n28607_ = ~new_n8457_ | ~new_n8806_;
  assign new_n28608_ = ~new_n28488_ | ~new_n28606_;
  assign new_n28609_ = new_n8800_ | new_n8440_;
  assign new_n28610_ = new_n8806_ | new_n8457_;
  assign new_n28611_ = ~new_n28487_ | ~new_n28526_;
  assign new_n28612_ = ~new_n28610_ | ~new_n28608_;
  assign new_n28613_ = ~new_n28525_;
  assign new_n28614_ = new_n8809_ | new_n8456_;
  assign new_n28615_ = ~new_n28614_ | ~new_n28525_;
  assign new_n28616_ = ~new_n8456_ | ~new_n8809_;
  assign new_n28617_ = ~new_n28523_;
  assign new_n28618_ = new_n8812_ | new_n8451_;
  assign new_n28619_ = ~new_n28618_ | ~new_n28523_;
  assign new_n28620_ = ~new_n8451_ | ~new_n8812_;
  assign new_n28621_ = ~new_n28451_;
  assign new_n28622_ = new_n8446_ | new_n8818_;
  assign new_n28623_ = new_n8450_ | new_n8815_;
  assign new_n28624_ = ~new_n28418_;
  assign new_n28625_ = ~new_n28419_ | ~new_n28418_;
  assign new_n28626_ = ~new_n8446_ | ~new_n28625_;
  assign new_n28627_ = ~new_n8818_ | ~new_n28624_;
  assign new_n28628_ = ~new_n28367_ | ~new_n28451_;
  assign new_n28629_ = ~new_n28521_;
  assign new_n28630_ = new_n8453_ | new_n9285_;
  assign new_n28631_ = new_n8458_ | new_n8823_;
  assign new_n28632_ = new_n8452_ | new_n9284_;
  assign new_n28633_ = ~new_n28439_;
  assign new_n28634_ = ~new_n9285_ | ~new_n28633_;
  assign new_n28635_ = ~new_n28634_ | ~new_n28449_;
  assign new_n28636_ = ~new_n28439_ | ~new_n28440_;
  assign new_n28637_ = ~new_n28636_ | ~new_n28635_;
  assign new_n28638_ = ~new_n28534_ | ~new_n28368_;
  assign new_n28639_ = ~new_n8452_ | ~new_n9284_;
  assign new_n28640_ = ~new_n28637_ | ~new_n28638_;
  assign new_n28641_ = new_n8821_ | new_n8459_;
  assign new_n28642_ = new_n9284_ | new_n8452_;
  assign new_n28643_ = ~new_n28521_ | ~new_n28490_;
  assign new_n28644_ = ~new_n28642_ | ~new_n28640_;
  assign new_n28645_ = ~new_n28518_;
  assign new_n28646_ = new_n9283_ | new_n8438_;
  assign new_n28647_ = ~new_n28646_ | ~new_n28518_;
  assign new_n28648_ = ~new_n8438_ | ~new_n9283_;
  assign new_n28649_ = ~new_n28516_;
  assign new_n28650_ = new_n9282_ | new_n8443_;
  assign new_n28651_ = ~new_n28650_ | ~new_n28516_;
  assign new_n28652_ = ~new_n8443_ | ~new_n9282_;
  assign new_n28653_ = ~new_n28514_;
  assign new_n28654_ = new_n8435_ | new_n9280_;
  assign new_n28655_ = ~new_n28535_ | ~new_n28532_;
  assign new_n28656_ = ~new_n28445_;
  assign new_n28657_ = new_n9281_ | new_n8442_;
  assign new_n28658_ = ~new_n28527_ | ~new_n28514_ | ~new_n28657_;
  assign new_n28659_ = ~new_n28512_;
  assign new_n28660_ = new_n9278_ | new_n8430_;
  assign new_n28661_ = ~new_n8430_ | ~new_n9278_;
  assign new_n28662_ = ~new_n28510_;
  assign new_n28663_ = ~new_n9277_ | ~new_n28510_;
  assign new_n28664_ = ~new_n28508_;
  assign new_n28665_ = ~new_n28657_ | ~new_n28514_;
  assign new_n28666_ = ~new_n28448_;
  assign new_n28667_ = new_n9280_ | new_n8435_;
  assign new_n28668_ = ~new_n28667_ | ~new_n28448_;
  assign new_n28669_ = ~new_n28513_ | ~new_n28668_ | ~new_n28532_;
  assign new_n28670_ = ~new_n28666_ | ~new_n28532_;
  assign new_n28671_ = ~new_n9279_ | ~new_n8434_;
  assign new_n28672_ = ~new_n28527_ | ~new_n28670_ | ~new_n28671_;
  assign new_n28673_ = new_n8435_ | new_n9280_;
  assign new_n28674_ = ~new_n28641_ | ~new_n28521_;
  assign new_n28675_ = ~new_n28450_;
  assign new_n28676_ = ~new_n28368_ | ~new_n28450_;
  assign new_n28677_ = ~new_n28494_ | ~new_n28676_;
  assign new_n28678_ = ~new_n28676_ | ~new_n28637_;
  assign new_n28679_ = ~new_n28812_ | ~new_n28678_;
  assign new_n28680_ = new_n8823_ | new_n8458_;
  assign new_n28681_ = ~new_n28680_ | ~new_n28450_;
  assign new_n28682_ = ~new_n28495_ | ~new_n28681_;
  assign new_n28683_ = ~new_n28675_ | ~new_n28439_;
  assign new_n28684_ = ~new_n8453_ | ~new_n9285_;
  assign new_n28685_ = ~new_n28496_ | ~new_n28683_;
  assign new_n28686_ = new_n8770_ | new_n8455_;
  assign new_n28687_ = ~new_n28520_;
  assign new_n28688_ = new_n8458_ | new_n8823_;
  assign new_n28689_ = new_n8815_ | new_n8450_;
  assign new_n28690_ = ~new_n28689_ | ~new_n28451_;
  assign new_n28691_ = ~new_n28497_ | ~new_n28690_;
  assign new_n28692_ = ~new_n28621_ | ~new_n28418_;
  assign new_n28693_ = ~new_n8818_ | ~new_n8446_;
  assign new_n28694_ = ~new_n28498_ | ~new_n28692_;
  assign new_n28695_ = new_n8450_ | new_n8815_;
  assign new_n28696_ = ~new_n28609_ | ~new_n28526_;
  assign new_n28697_ = ~new_n28452_;
  assign new_n28698_ = new_n8803_ | new_n8449_;
  assign new_n28699_ = ~new_n28698_ | ~new_n28452_;
  assign new_n28700_ = ~new_n28499_ | ~new_n28699_;
  assign new_n28701_ = ~new_n28697_ | ~new_n28531_;
  assign new_n28702_ = ~new_n8457_ | ~new_n8806_;
  assign new_n28703_ = ~new_n28500_ | ~new_n28701_;
  assign new_n28704_ = new_n8449_ | new_n8803_;
  assign new_n28705_ = new_n8794_ | new_n8460_;
  assign new_n28706_ = ~new_n28705_ | ~new_n28399_;
  assign new_n28707_ = ~new_n28501_ | ~new_n28706_;
  assign new_n28708_ = ~new_n28565_ | ~new_n28530_;
  assign new_n28709_ = ~new_n8439_ | ~new_n8797_;
  assign new_n28710_ = ~new_n28502_ | ~new_n28708_;
  assign new_n28711_ = ~new_n28566_ | ~new_n28530_;
  assign new_n28712_ = ~new_n28563_ | ~new_n28422_;
  assign new_n28713_ = ~new_n28573_ | ~new_n28381_;
  assign new_n28714_ = ~new_n28587_ | ~new_n28393_;
  assign new_n28715_ = ~new_n28590_ | ~new_n28539_;
  assign new_n28716_ = ~new_n28673_ | ~new_n28532_;
  assign new_n28717_ = ~new_n28657_ | ~new_n28535_;
  assign new_n28718_ = ~new_n28688_ | ~new_n28439_;
  assign new_n28719_ = ~new_n28641_ | ~new_n28436_;
  assign new_n28720_ = ~new_n28695_ | ~new_n28418_;
  assign new_n28721_ = ~new_n28704_ | ~new_n28531_;
  assign new_n28722_ = ~new_n28609_ | ~new_n28427_;
  assign new_n28723_ = ~new_n9277_ | ~new_n8431_;
  assign new_n28724_ = ~new_n28655_ | ~new_n28527_;
  assign new_n28725_ = ~new_n8434_ | ~new_n28654_;
  assign new_n28726_ = ~new_n9279_ | ~new_n28654_;
  assign new_n28727_ = ~new_n28660_ | ~new_n28655_ | ~new_n28527_;
  assign new_n28728_ = ~new_n28492_ | ~new_n28514_ | ~new_n28527_;
  assign new_n28729_ = ~new_n28656_ | ~new_n28660_;
  assign new_n28730_ = ~new_n8460_ | ~new_n28398_;
  assign new_n28731_ = ~new_n8794_ | ~new_n28397_;
  assign new_n28732_ = ~new_n28731_ | ~new_n28730_;
  assign new_n28733_ = ~new_n28711_ | ~new_n28399_;
  assign new_n28734_ = ~new_n28732_ | ~new_n28565_;
  assign new_n28735_ = ~new_n8461_ | ~new_n28395_;
  assign new_n28736_ = ~new_n8791_ | ~new_n28396_;
  assign new_n28737_ = ~new_n28736_ | ~new_n28735_;
  assign new_n28738_ = ~new_n28712_ | ~new_n28503_;
  assign new_n28739_ = ~new_n28562_ | ~new_n28737_;
  assign new_n28740_ = ~new_n8447_ | ~new_n28382_;
  assign new_n28741_ = ~new_n8788_ | ~new_n28380_;
  assign new_n28742_ = ~new_n8448_ | ~new_n28378_;
  assign new_n28743_ = ~new_n8785_ | ~new_n28379_;
  assign new_n28744_ = ~new_n28743_ | ~new_n28742_;
  assign new_n28745_ = ~new_n28713_ | ~new_n28400_;
  assign new_n28746_ = ~new_n28744_ | ~new_n28554_;
  assign new_n28747_ = ~new_n8444_ | ~new_n28394_;
  assign new_n28748_ = ~new_n8782_ | ~new_n28385_;
  assign new_n28749_ = ~new_n8437_ | ~new_n28383_;
  assign new_n28750_ = ~new_n8779_ | ~new_n28384_;
  assign new_n28751_ = ~new_n28750_ | ~new_n28749_;
  assign new_n28752_ = ~new_n28714_ | ~new_n28403_;
  assign new_n28753_ = ~new_n28751_ | ~new_n28580_;
  assign new_n28754_ = ~new_n8441_ | ~new_n28391_;
  assign new_n28755_ = ~new_n8776_ | ~new_n28392_;
  assign new_n28756_ = ~new_n28755_ | ~new_n28754_;
  assign new_n28757_ = ~new_n28715_ | ~new_n28504_;
  assign new_n28758_ = ~new_n28589_ | ~new_n28756_;
  assign new_n28759_ = ~new_n8445_ | ~new_n28386_;
  assign new_n28760_ = ~new_n8773_ | ~new_n28387_;
  assign new_n28761_ = ~new_n8432_ | ~new_n28506_;
  assign new_n28762_ = ~new_n9286_ | ~new_n28505_;
  assign new_n28763_ = ~new_n8432_ | ~new_n28506_;
  assign new_n28764_ = ~new_n9286_ | ~new_n28505_;
  assign new_n28765_ = ~new_n28764_ | ~new_n28763_;
  assign new_n28766_ = ~new_n28507_ | ~new_n28508_;
  assign new_n28767_ = ~new_n28664_ | ~new_n28765_;
  assign new_n28768_ = ~new_n8431_ | ~new_n28447_;
  assign new_n28769_ = ~new_n9277_ | ~new_n28446_;
  assign new_n28770_ = ~new_n8431_ | ~new_n28447_;
  assign new_n28771_ = ~new_n9277_ | ~new_n28446_;
  assign new_n28772_ = ~new_n28771_ | ~new_n28770_;
  assign new_n28773_ = ~new_n28509_ | ~new_n28510_;
  assign new_n28774_ = ~new_n28662_ | ~new_n28772_;
  assign new_n28775_ = ~new_n8430_ | ~new_n28405_;
  assign new_n28776_ = ~new_n9278_ | ~new_n28406_;
  assign new_n28777_ = ~new_n8430_ | ~new_n28405_;
  assign new_n28778_ = ~new_n9278_ | ~new_n28406_;
  assign new_n28779_ = ~new_n28778_ | ~new_n28777_;
  assign new_n28780_ = ~new_n28511_ | ~new_n28512_;
  assign new_n28781_ = ~new_n28659_ | ~new_n28779_;
  assign new_n28782_ = ~new_n8434_ | ~new_n28408_;
  assign new_n28783_ = ~new_n9279_ | ~new_n28407_;
  assign new_n28784_ = ~new_n8435_ | ~new_n28409_;
  assign new_n28785_ = ~new_n9280_ | ~new_n28410_;
  assign new_n28786_ = ~new_n28785_ | ~new_n28784_;
  assign new_n28787_ = ~new_n28716_ | ~new_n28448_;
  assign new_n28788_ = ~new_n28786_ | ~new_n28666_;
  assign new_n28789_ = ~new_n8442_ | ~new_n28411_;
  assign new_n28790_ = ~new_n9281_ | ~new_n28412_;
  assign new_n28791_ = ~new_n28790_ | ~new_n28789_;
  assign new_n28792_ = ~new_n28717_ | ~new_n28514_;
  assign new_n28793_ = ~new_n28653_ | ~new_n28791_;
  assign new_n28794_ = ~new_n8443_ | ~new_n28443_;
  assign new_n28795_ = ~new_n9282_ | ~new_n28444_;
  assign new_n28796_ = ~new_n8443_ | ~new_n28443_;
  assign new_n28797_ = ~new_n9282_ | ~new_n28444_;
  assign new_n28798_ = ~new_n28797_ | ~new_n28796_;
  assign new_n28799_ = ~new_n28515_ | ~new_n28516_;
  assign new_n28800_ = ~new_n28649_ | ~new_n28798_;
  assign new_n28801_ = ~new_n8438_ | ~new_n28441_;
  assign new_n28802_ = ~new_n9283_ | ~new_n28442_;
  assign new_n28803_ = ~new_n8438_ | ~new_n28441_;
  assign new_n28804_ = ~new_n9283_ | ~new_n28442_;
  assign new_n28805_ = ~new_n28804_ | ~new_n28803_;
  assign new_n28806_ = ~new_n28517_ | ~new_n28518_;
  assign new_n28807_ = ~new_n28645_ | ~new_n28805_;
  assign new_n28808_ = ~new_n8452_ | ~new_n28413_;
  assign new_n28809_ = ~new_n9284_ | ~new_n28414_;
  assign new_n28810_ = ~new_n8452_ | ~new_n28413_;
  assign new_n28811_ = ~new_n9284_ | ~new_n28414_;
  assign new_n28812_ = ~new_n28811_ | ~new_n28810_;
  assign new_n28813_ = ~new_n8453_ | ~new_n28440_;
  assign new_n28814_ = ~new_n9285_ | ~new_n28449_;
  assign new_n28815_ = ~new_n28541_ | ~new_n28520_;
  assign new_n28816_ = ~new_n28687_ | ~new_n28390_;
  assign new_n28817_ = ~new_n8458_ | ~new_n28437_;
  assign new_n28818_ = ~new_n8823_ | ~new_n28438_;
  assign new_n28819_ = ~new_n28818_ | ~new_n28817_;
  assign new_n28820_ = ~new_n28718_ | ~new_n28450_;
  assign new_n28821_ = ~new_n28819_ | ~new_n28675_;
  assign new_n28822_ = ~new_n8459_ | ~new_n28434_;
  assign new_n28823_ = ~new_n8821_ | ~new_n28435_;
  assign new_n28824_ = ~new_n28823_ | ~new_n28822_;
  assign new_n28825_ = ~new_n28719_ | ~new_n28521_;
  assign new_n28826_ = ~new_n28629_ | ~new_n28824_;
  assign new_n28827_ = ~new_n8446_ | ~new_n28419_;
  assign new_n28828_ = ~new_n8818_ | ~new_n28417_;
  assign new_n28829_ = ~new_n8450_ | ~new_n28415_;
  assign new_n28830_ = ~new_n8815_ | ~new_n28416_;
  assign new_n28831_ = ~new_n28830_ | ~new_n28829_;
  assign new_n28832_ = ~new_n28720_ | ~new_n28451_;
  assign new_n28833_ = ~new_n28831_ | ~new_n28621_;
  assign new_n28834_ = ~new_n8451_ | ~new_n28432_;
  assign new_n28835_ = ~new_n8812_ | ~new_n28433_;
  assign new_n28836_ = ~new_n8451_ | ~new_n28432_;
  assign new_n28837_ = ~new_n8812_ | ~new_n28433_;
  assign new_n28838_ = ~new_n28837_ | ~new_n28836_;
  assign new_n28839_ = ~new_n28522_ | ~new_n28523_;
  assign new_n28840_ = ~new_n28617_ | ~new_n28838_;
  assign new_n28841_ = ~new_n8456_ | ~new_n28430_;
  assign new_n28842_ = ~new_n8809_ | ~new_n28431_;
  assign new_n28843_ = ~new_n8456_ | ~new_n28430_;
  assign new_n28844_ = ~new_n8809_ | ~new_n28431_;
  assign new_n28845_ = ~new_n28844_ | ~new_n28843_;
  assign new_n28846_ = ~new_n28524_ | ~new_n28525_;
  assign new_n28847_ = ~new_n28613_ | ~new_n28845_;
  assign new_n28848_ = ~new_n8457_ | ~new_n28428_;
  assign new_n28849_ = ~new_n8806_ | ~new_n28429_;
  assign new_n28850_ = ~new_n8449_ | ~new_n28423_;
  assign new_n28851_ = ~new_n8803_ | ~new_n28424_;
  assign new_n28852_ = ~new_n28851_ | ~new_n28850_;
  assign new_n28853_ = ~new_n28721_ | ~new_n28452_;
  assign new_n28854_ = ~new_n28852_ | ~new_n28697_;
  assign new_n28855_ = ~new_n8440_ | ~new_n28425_;
  assign new_n28856_ = ~new_n8800_ | ~new_n28426_;
  assign new_n28857_ = ~new_n28856_ | ~new_n28855_;
  assign new_n28858_ = ~new_n28722_ | ~new_n28526_;
  assign new_n28859_ = ~new_n28603_ | ~new_n28857_;
  assign new_n28860_ = ~new_n8439_ | ~new_n28420_;
  assign new_n28861_ = ~new_n8797_ | ~new_n28421_;
  assign new_n28862_ = ~new_n8454_ | ~new_n28388_;
  assign new_n28863_ = ~new_n8765_ | ~new_n28389_;
  assign new_n28864_ = new_n29087_ & new_n29086_;
  assign new_n28865_ = new_n29098_ & new_n29097_;
  assign new_n28866_ = new_n29123_ & new_n29122_;
  assign new_n28867_ = new_n29137_ & new_n29136_;
  assign new_n28868_ = new_n29149_ & new_n29148_;
  assign new_n28869_ = new_n28866_ & new_n29127_;
  assign new_n28870_ = new_n28865_ & new_n29095_;
  assign new_n28871_ = new_n28869_ & new_n29120_;
  assign new_n28872_ = new_n29395_ & new_n29394_;
  assign new_n28873_ = new_n29205_ & new_n29202_;
  assign new_n28874_ = new_n29196_ & new_n29193_;
  assign new_n28875_ = new_n29189_ & new_n29186_;
  assign new_n28876_ = new_n29002_ & new_n29397_ & new_n29396_;
  assign new_n28877_ = new_n29116_ & new_n29113_;
  assign new_n28878_ = new_n29109_ & new_n29106_;
  assign new_n28879_ = ~new_n8434_ | ~new_n29166_;
  assign new_n28880_ = ~new_n8530_;
  assign new_n28881_ = ~new_n8461_;
  assign new_n28882_ = ~new_n8448_;
  assign new_n28883_ = ~new_n8448_ | ~new_n28927_;
  assign new_n28884_ = ~new_n8447_;
  assign new_n28885_ = ~new_n8444_;
  assign new_n28886_ = ~new_n8444_ | ~new_n28929_;
  assign new_n28887_ = ~new_n8445_;
  assign new_n28888_ = ~new_n8445_ | ~new_n28930_;
  assign new_n28889_ = ~new_n8441_;
  assign new_n28890_ = ~new_n8455_;
  assign new_n28891_ = ~new_n8454_;
  assign new_n28892_ = ~new_n8437_;
  assign new_n28893_ = ~new_n8460_;
  assign new_n28894_ = ~new_n29222_ | ~new_n29219_ | ~new_n29101_;
  assign new_n28895_ = ~new_n29239_ | ~new_n28886_;
  assign new_n28896_ = ~new_n29220_ | ~new_n29221_ | ~new_n29084_;
  assign new_n28897_ = ~new_n8430_;
  assign new_n28898_ = ~new_n8435_;
  assign new_n28899_ = ~new_n8442_;
  assign new_n28900_ = ~new_n8434_;
  assign new_n28901_ = ~new_n8450_;
  assign new_n28902_ = ~new_n8450_ | ~new_n28939_;
  assign new_n28903_ = ~new_n8446_;
  assign new_n28904_ = ~new_n8456_;
  assign new_n28905_ = ~new_n8449_;
  assign new_n28906_ = ~new_n8440_;
  assign new_n28907_ = ~new_n8440_ | ~new_n28944_;
  assign new_n28908_ = ~new_n8457_;
  assign new_n28909_ = ~new_n8439_;
  assign new_n28910_ = ~new_n8439_ | ~new_n28945_;
  assign new_n28911_ = ~new_n8451_;
  assign new_n28912_ = ~new_n8459_;
  assign new_n28913_ = ~new_n8453_;
  assign new_n28914_ = ~new_n8458_;
  assign new_n28915_ = ~new_n8458_ | ~new_n28948_;
  assign new_n28916_ = ~new_n8452_;
  assign new_n28917_ = ~new_n8438_;
  assign new_n28918_ = ~new_n8443_;
  assign new_n28919_ = ~new_n8435_ | ~new_n28936_;
  assign new_n28920_ = ~new_n8442_ | ~new_n28937_;
  assign new_n28921_ = ~new_n28915_ | ~new_n29182_;
  assign new_n28922_ = ~new_n29134_ | ~new_n29133_;
  assign new_n28923_ = ~new_n29225_ | ~new_n29129_;
  assign new_n28924_ = ~new_n28907_ | ~new_n29198_;
  assign new_n28925_ = ~new_n29254_ | ~new_n29253_;
  assign new_n28926_ = ~new_n29286_ | ~new_n29285_;
  assign new_n28927_ = ~new_n29283_ | ~new_n29282_;
  assign new_n28928_ = ~new_n29280_ | ~new_n29279_;
  assign new_n28929_ = ~new_n29277_ | ~new_n29276_;
  assign new_n28930_ = ~new_n29274_ | ~new_n29273_;
  assign new_n28931_ = ~new_n29271_ | ~new_n29270_;
  assign new_n28932_ = ~new_n29265_ | ~new_n29264_;
  assign new_n28933_ = ~new_n29268_ | ~new_n29267_;
  assign new_n28934_ = ~new_n29262_ | ~new_n29261_;
  assign new_n28935_ = ~new_n29326_ | ~new_n29325_;
  assign new_n28936_ = ~new_n29374_ | ~new_n29373_;
  assign new_n28937_ = ~new_n29377_ | ~new_n29376_;
  assign new_n28938_ = ~new_n29371_ | ~new_n29370_;
  assign new_n28939_ = ~new_n29350_ | ~new_n29349_;
  assign new_n28940_ = ~new_n29347_ | ~new_n29346_;
  assign new_n28941_ = ~new_n29341_ | ~new_n29340_;
  assign new_n28942_ = ~new_n29338_ | ~new_n29337_;
  assign new_n28943_ = ~new_n29335_ | ~new_n29334_;
  assign new_n28944_ = ~new_n29332_ | ~new_n29331_;
  assign new_n28945_ = ~new_n29329_ | ~new_n29328_;
  assign new_n28946_ = ~new_n29344_ | ~new_n29343_;
  assign new_n28947_ = ~new_n29353_ | ~new_n29352_;
  assign new_n28948_ = ~new_n29362_ | ~new_n29361_;
  assign new_n28949_ = ~new_n29356_ | ~new_n29355_;
  assign new_n28950_ = ~new_n29359_ | ~new_n29358_;
  assign new_n28951_ = ~new_n29365_ | ~new_n29364_;
  assign new_n28952_ = ~new_n29368_ | ~new_n29367_;
  assign new_n28953_ = ~new_n29383_ | ~new_n29382_;
  assign new_n28954_ = ~new_n29492_ | ~new_n29491_;
  assign new_n28955_ = ~new_n29289_ | ~new_n29288_;
  assign new_n28956_ = ~new_n29296_ | ~new_n29295_;
  assign new_n28957_ = ~new_n29303_ | ~new_n29302_;
  assign new_n28958_ = ~new_n29310_ | ~new_n29309_;
  assign new_n28959_ = ~new_n29317_ | ~new_n29316_;
  assign new_n28960_ = ~new_n29324_ | ~new_n29323_;
  assign new_n28961_ = ~new_n29386_ | ~new_n29385_;
  assign new_n28962_ = ~new_n29393_ | ~new_n29392_;
  assign new_n28963_ = new_n29180_ & new_n29069_;
  assign new_n28964_ = new_n29001_ & new_n28872_;
  assign new_n28965_ = ~new_n29402_ | ~new_n29401_;
  assign new_n28966_ = ~new_n29407_ | ~new_n29406_;
  assign new_n28967_ = ~new_n29414_ | ~new_n29413_;
  assign new_n28968_ = ~new_n29421_ | ~new_n29420_;
  assign new_n28969_ = ~new_n29428_ | ~new_n29427_;
  assign new_n28970_ = ~new_n29435_ | ~new_n29434_;
  assign new_n28971_ = ~new_n29440_ | ~new_n29439_;
  assign new_n28972_ = ~new_n29447_ | ~new_n29446_;
  assign new_n28973_ = ~new_n29454_ | ~new_n29453_;
  assign new_n28974_ = ~new_n29461_ | ~new_n29460_;
  assign new_n28975_ = ~new_n29468_ | ~new_n29467_;
  assign new_n28976_ = ~new_n29475_ | ~new_n29474_;
  assign new_n28977_ = ~new_n29480_ | ~new_n29479_;
  assign new_n28978_ = ~new_n29487_ | ~new_n29486_;
  assign new_n28979_ = new_n28933_ & new_n8530_;
  assign new_n28980_ = new_n29090_ & new_n29089_;
  assign new_n28981_ = new_n29102_ & new_n28870_;
  assign new_n28982_ = new_n29224_ & new_n29103_;
  assign new_n28983_ = new_n28883_ & new_n29298_ & new_n29297_;
  assign new_n28984_ = new_n29108_ & new_n28865_;
  assign new_n28985_ = new_n28888_ & new_n29319_ & new_n29318_;
  assign new_n28986_ = new_n29115_ & new_n28864_;
  assign new_n28987_ = new_n29125_ & new_n29073_;
  assign new_n28988_ = new_n29130_ & new_n28871_;
  assign new_n28989_ = new_n29233_ & new_n29131_;
  assign new_n28990_ = new_n29141_ & new_n29140_;
  assign new_n28991_ = new_n29153_ & new_n28868_;
  assign new_n28992_ = new_n29151_ & new_n29074_;
  assign new_n28993_ = new_n29174_ & new_n29236_;
  assign new_n28994_ = new_n29176_ & new_n29167_;
  assign new_n28995_ = new_n29176_ & new_n29229_;
  assign new_n28996_ = new_n29234_ & new_n29175_;
  assign new_n28997_ = ~new_n29380_ | ~new_n29379_;
  assign new_n28998_ = new_n29375_ & new_n28898_;
  assign new_n28999_ = new_n29180_ & new_n29075_;
  assign new_n29000_ = new_n29180_ & new_n29078_;
  assign new_n29001_ = new_n28920_ & new_n28919_;
  assign new_n29002_ = new_n29252_ & new_n29251_ & new_n29179_;
  assign new_n29003_ = new_n29074_ & new_n29423_ & new_n29422_;
  assign new_n29004_ = new_n29188_ & new_n28868_;
  assign new_n29005_ = new_n28902_ & new_n29449_ & new_n29448_;
  assign new_n29006_ = new_n29195_ & new_n28867_;
  assign new_n29007_ = new_n29073_ & new_n29470_ & new_n29469_;
  assign new_n29008_ = new_n29204_ & new_n28866_;
  assign new_n29009_ = ~new_n29489_ | ~new_n29488_;
  assign new_n29010_ = ~new_n8794_;
  assign new_n29011_ = new_n29257_ & new_n29256_;
  assign new_n29012_ = ~new_n8779_;
  assign new_n29013_ = ~new_n8770_;
  assign new_n29014_ = ~new_n8765_;
  assign new_n29015_ = ~new_n8776_;
  assign new_n29016_ = ~new_n8773_;
  assign new_n29017_ = ~new_n8782_;
  assign new_n29018_ = ~new_n8788_;
  assign new_n29019_ = ~new_n8785_;
  assign new_n29020_ = ~new_n8791_;
  assign new_n29021_ = ~new_n28982_ | ~new_n29243_;
  assign new_n29022_ = new_n29291_ & new_n29290_;
  assign new_n29023_ = ~new_n29223_ | ~new_n29241_;
  assign new_n29024_ = new_n29305_ & new_n29304_;
  assign new_n29025_ = ~new_n29216_ | ~new_n29093_ | ~new_n29071_;
  assign new_n29026_ = new_n29312_ & new_n29311_;
  assign new_n29027_ = ~new_n28980_ | ~new_n29091_;
  assign new_n29028_ = ~new_n9278_;
  assign new_n29029_ = ~new_n8797_;
  assign new_n29030_ = ~new_n8800_;
  assign new_n29031_ = ~new_n8806_;
  assign new_n29032_ = ~new_n8803_;
  assign new_n29033_ = ~new_n8809_;
  assign new_n29034_ = ~new_n8812_;
  assign new_n29035_ = ~new_n8818_;
  assign new_n29036_ = ~new_n8815_;
  assign new_n29037_ = ~new_n8821_;
  assign new_n29038_ = ~new_n9284_;
  assign new_n29039_ = ~new_n9285_;
  assign new_n29040_ = ~new_n8823_;
  assign new_n29041_ = ~new_n9283_;
  assign new_n29042_ = ~new_n9282_;
  assign new_n29043_ = ~new_n9279_;
  assign new_n29044_ = ~new_n9280_;
  assign new_n29045_ = ~new_n9281_;
  assign new_n29046_ = ~new_n8431_;
  assign new_n29047_ = ~new_n9277_;
  assign new_n29048_ = new_n29388_ & new_n29387_;
  assign new_n29049_ = ~new_n29171_ | ~new_n29170_;
  assign new_n29050_ = ~new_n29169_ | ~new_n29052_;
  assign new_n29051_ = ~new_n28920_ | ~new_n29050_;
  assign new_n29052_ = ~new_n29164_ | ~new_n29163_;
  assign new_n29053_ = new_n29409_ & new_n29408_;
  assign new_n29054_ = ~new_n29160_ | ~new_n29159_;
  assign new_n29055_ = new_n29416_ & new_n29415_;
  assign new_n29056_ = ~new_n29156_ | ~new_n29155_;
  assign new_n29057_ = new_n29430_ & new_n29429_;
  assign new_n29058_ = ~new_n29081_ | ~new_n29080_;
  assign new_n29059_ = ~new_n29146_ | ~new_n29145_;
  assign new_n29060_ = new_n29442_ & new_n29441_;
  assign new_n29061_ = ~new_n28990_ | ~new_n29142_;
  assign new_n29062_ = new_n29456_ & new_n29455_;
  assign new_n29063_ = ~new_n28989_ | ~new_n29249_;
  assign new_n29064_ = new_n29463_ & new_n29462_;
  assign new_n29065_ = ~new_n29232_ | ~new_n29247_;
  assign new_n29066_ = ~new_n29245_ | ~new_n28910_;
  assign new_n29067_ = new_n29482_ & new_n29481_;
  assign new_n29068_ = ~new_n29217_ | ~new_n29118_ | ~new_n29070_;
  assign new_n29069_ = ~new_n28879_ | ~new_n29227_;
  assign new_n29070_ = ~new_n28925_ | ~new_n29021_;
  assign new_n29071_ = ~new_n28934_ | ~new_n29027_;
  assign new_n29072_ = ~new_n28888_;
  assign new_n29073_ = ~new_n8449_ | ~new_n28942_;
  assign new_n29074_ = ~new_n8453_ | ~new_n28950_;
  assign new_n29075_ = ~new_n28919_;
  assign new_n29076_ = ~new_n28907_;
  assign new_n29077_ = ~new_n28915_;
  assign new_n29078_ = ~new_n28920_;
  assign new_n29079_ = ~new_n29269_ | ~new_n28880_;
  assign new_n29080_ = ~new_n8454_ | ~new_n29079_;
  assign new_n29081_ = ~new_n8530_ | ~new_n28933_;
  assign new_n29082_ = ~new_n29058_;
  assign new_n29083_ = ~new_n29266_ | ~new_n28890_;
  assign new_n29084_ = ~new_n8455_ | ~new_n28932_;
  assign new_n29085_ = ~new_n28896_;
  assign new_n29086_ = ~new_n29272_ | ~new_n28889_;
  assign new_n29087_ = ~new_n29275_ | ~new_n28887_;
  assign new_n29088_ = ~new_n28889_ | ~new_n28888_;
  assign new_n29089_ = ~new_n28931_ | ~new_n29088_;
  assign new_n29090_ = ~new_n8441_ | ~new_n29072_;
  assign new_n29091_ = ~new_n28864_ | ~new_n28896_;
  assign new_n29092_ = ~new_n29027_;
  assign new_n29093_ = ~new_n8437_ | ~new_n29027_;
  assign new_n29094_ = ~new_n29025_;
  assign new_n29095_ = ~new_n29278_ | ~new_n28885_;
  assign new_n29096_ = ~new_n28886_;
  assign new_n29097_ = ~new_n29281_ | ~new_n28884_;
  assign new_n29098_ = ~new_n29284_ | ~new_n28882_;
  assign new_n29099_ = ~new_n28883_;
  assign new_n29100_ = ~new_n28884_ | ~new_n28883_;
  assign new_n29101_ = ~new_n8447_ | ~new_n29099_;
  assign new_n29102_ = ~new_n29287_ | ~new_n28881_;
  assign new_n29103_ = ~new_n8461_ | ~new_n28926_;
  assign new_n29104_ = ~new_n29284_ | ~new_n28882_;
  assign new_n29105_ = ~new_n29104_ | ~new_n28895_;
  assign new_n29106_ = ~new_n28983_ | ~new_n29105_;
  assign new_n29107_ = ~new_n29240_ | ~new_n28883_;
  assign new_n29108_ = ~new_n8447_ | ~new_n28928_;
  assign new_n29109_ = ~new_n28984_ | ~new_n29107_;
  assign new_n29110_ = ~new_n29284_ | ~new_n28882_;
  assign new_n29111_ = ~new_n29275_ | ~new_n28887_;
  assign new_n29112_ = ~new_n29111_ | ~new_n28896_;
  assign new_n29113_ = ~new_n28985_ | ~new_n29112_;
  assign new_n29114_ = ~new_n29085_ | ~new_n28888_;
  assign new_n29115_ = ~new_n8441_ | ~new_n28931_;
  assign new_n29116_ = ~new_n28986_ | ~new_n29114_;
  assign new_n29117_ = ~new_n29275_ | ~new_n28887_;
  assign new_n29118_ = ~new_n8460_ | ~new_n29021_;
  assign new_n29119_ = ~new_n29068_;
  assign new_n29120_ = ~new_n29330_ | ~new_n28909_;
  assign new_n29121_ = ~new_n28910_;
  assign new_n29122_ = ~new_n29336_ | ~new_n28908_;
  assign new_n29123_ = ~new_n29339_ | ~new_n28905_;
  assign new_n29124_ = ~new_n29076_ | ~new_n28866_;
  assign new_n29125_ = ~new_n8457_ | ~new_n28943_;
  assign new_n29126_ = ~new_n28987_ | ~new_n29124_;
  assign new_n29127_ = ~new_n29333_ | ~new_n28906_;
  assign new_n29128_ = ~new_n29336_ | ~new_n28908_;
  assign new_n29129_ = ~new_n29128_ | ~new_n29126_;
  assign new_n29130_ = ~new_n29342_ | ~new_n28904_;
  assign new_n29131_ = ~new_n8456_ | ~new_n28941_;
  assign new_n29132_ = ~new_n29345_ | ~new_n28911_;
  assign new_n29133_ = ~new_n29132_ | ~new_n29063_;
  assign new_n29134_ = ~new_n8451_ | ~new_n28946_;
  assign new_n29135_ = ~new_n28922_;
  assign new_n29136_ = ~new_n29348_ | ~new_n28903_;
  assign new_n29137_ = ~new_n29351_ | ~new_n28901_;
  assign new_n29138_ = ~new_n28902_;
  assign new_n29139_ = ~new_n28903_ | ~new_n28902_;
  assign new_n29140_ = ~new_n28940_ | ~new_n29139_;
  assign new_n29141_ = ~new_n8446_ | ~new_n29138_;
  assign new_n29142_ = ~new_n28867_ | ~new_n28922_;
  assign new_n29143_ = ~new_n29061_;
  assign new_n29144_ = ~new_n29354_ | ~new_n28912_;
  assign new_n29145_ = ~new_n29144_ | ~new_n29061_;
  assign new_n29146_ = ~new_n8459_ | ~new_n28947_;
  assign new_n29147_ = ~new_n29059_;
  assign new_n29148_ = ~new_n29357_ | ~new_n28916_;
  assign new_n29149_ = ~new_n29360_ | ~new_n28913_;
  assign new_n29150_ = ~new_n29077_ | ~new_n28868_;
  assign new_n29151_ = ~new_n8452_ | ~new_n28949_;
  assign new_n29152_ = ~new_n28992_ | ~new_n29150_;
  assign new_n29153_ = ~new_n29363_ | ~new_n28914_;
  assign new_n29154_ = ~new_n29357_ | ~new_n28916_;
  assign new_n29155_ = ~new_n28991_ | ~new_n29059_;
  assign new_n29156_ = ~new_n29154_ | ~new_n29152_;
  assign new_n29157_ = ~new_n29056_;
  assign new_n29158_ = ~new_n29366_ | ~new_n28917_;
  assign new_n29159_ = ~new_n29158_ | ~new_n29056_;
  assign new_n29160_ = ~new_n8438_ | ~new_n28951_;
  assign new_n29161_ = ~new_n29054_;
  assign new_n29162_ = ~new_n29369_ | ~new_n28918_;
  assign new_n29163_ = ~new_n29162_ | ~new_n29054_;
  assign new_n29164_ = ~new_n8443_ | ~new_n28952_;
  assign new_n29165_ = ~new_n29052_;
  assign new_n29166_ = ~new_n29375_ | ~new_n28898_;
  assign new_n29167_ = ~new_n29168_ | ~new_n28920_ | ~new_n28919_;
  assign new_n29168_ = ~new_n8434_ | ~new_n28938_;
  assign new_n29169_ = ~new_n29378_ | ~new_n28899_;
  assign new_n29170_ = ~new_n29229_ | ~new_n29052_;
  assign new_n29171_ = ~new_n29226_ | ~new_n29167_;
  assign new_n29172_ = ~new_n29049_;
  assign new_n29173_ = ~new_n29327_ | ~new_n28897_;
  assign new_n29174_ = ~new_n8430_ | ~new_n28935_;
  assign new_n29175_ = ~new_n8430_ | ~new_n28935_;
  assign new_n29176_ = ~new_n29327_ | ~new_n28897_;
  assign new_n29177_ = ~new_n29050_;
  assign new_n29178_ = ~new_n29051_;
  assign new_n29179_ = ~new_n28998_ | ~new_n28872_;
  assign new_n29180_ = ~new_n8434_ | ~new_n28938_;
  assign new_n29181_ = ~new_n29375_ | ~new_n28898_;
  assign new_n29182_ = ~new_n29153_ | ~new_n29059_;
  assign new_n29183_ = ~new_n28921_;
  assign new_n29184_ = ~new_n29360_ | ~new_n28913_;
  assign new_n29185_ = ~new_n29184_ | ~new_n28921_;
  assign new_n29186_ = ~new_n29003_ | ~new_n29185_;
  assign new_n29187_ = ~new_n29183_ | ~new_n29074_;
  assign new_n29188_ = ~new_n8452_ | ~new_n28949_;
  assign new_n29189_ = ~new_n29004_ | ~new_n29187_;
  assign new_n29190_ = ~new_n29360_ | ~new_n28913_;
  assign new_n29191_ = ~new_n29351_ | ~new_n28901_;
  assign new_n29192_ = ~new_n29191_ | ~new_n28922_;
  assign new_n29193_ = ~new_n29005_ | ~new_n29192_;
  assign new_n29194_ = ~new_n29135_ | ~new_n28902_;
  assign new_n29195_ = ~new_n8446_ | ~new_n28940_;
  assign new_n29196_ = ~new_n29006_ | ~new_n29194_;
  assign new_n29197_ = ~new_n29351_ | ~new_n28901_;
  assign new_n29198_ = ~new_n29127_ | ~new_n29066_;
  assign new_n29199_ = ~new_n28924_;
  assign new_n29200_ = ~new_n29339_ | ~new_n28905_;
  assign new_n29201_ = ~new_n29200_ | ~new_n28924_;
  assign new_n29202_ = ~new_n29007_ | ~new_n29201_;
  assign new_n29203_ = ~new_n29199_ | ~new_n29073_;
  assign new_n29204_ = ~new_n8457_ | ~new_n28943_;
  assign new_n29205_ = ~new_n29008_ | ~new_n29203_;
  assign new_n29206_ = ~new_n29339_ | ~new_n28905_;
  assign new_n29207_ = ~new_n29110_ | ~new_n28883_;
  assign new_n29208_ = ~new_n29117_ | ~new_n28888_;
  assign new_n29209_ = ~new_n29181_ | ~new_n28919_;
  assign new_n29210_ = ~new_n29169_ | ~new_n28920_;
  assign new_n29211_ = ~new_n29190_ | ~new_n29074_;
  assign new_n29212_ = ~new_n29153_ | ~new_n28915_;
  assign new_n29213_ = ~new_n29197_ | ~new_n28902_;
  assign new_n29214_ = ~new_n29206_ | ~new_n29073_;
  assign new_n29215_ = ~new_n29127_ | ~new_n28907_;
  assign new_n29216_ = ~new_n8437_ | ~new_n28934_;
  assign new_n29217_ = ~new_n8460_ | ~new_n28925_;
  assign new_n29218_ = ~new_n28993_ | ~new_n29170_;
  assign new_n29219_ = ~new_n28928_ | ~new_n29100_;
  assign new_n29220_ = ~new_n29083_ | ~new_n8454_ | ~new_n29079_;
  assign new_n29221_ = ~new_n28979_ | ~new_n29083_;
  assign new_n29222_ = ~new_n29096_ | ~new_n28865_;
  assign new_n29223_ = ~new_n28894_;
  assign new_n29224_ = ~new_n28894_ | ~new_n29102_;
  assign new_n29225_ = ~new_n29121_ | ~new_n28869_;
  assign new_n29226_ = ~new_n28879_ | ~new_n29227_ | ~new_n29168_;
  assign new_n29227_ = ~new_n28938_ | ~new_n29166_;
  assign new_n29228_ = ~new_n28879_;
  assign new_n29229_ = ~new_n29231_ | ~new_n29230_;
  assign new_n29230_ = ~new_n28938_ | ~new_n29169_ | ~new_n29166_;
  assign new_n29231_ = ~new_n29228_ | ~new_n29169_;
  assign new_n29232_ = ~new_n28923_;
  assign new_n29233_ = ~new_n28923_ | ~new_n29130_;
  assign new_n29234_ = ~new_n28994_ | ~new_n29226_;
  assign new_n29235_ = ~new_n28995_ | ~new_n29052_;
  assign new_n29236_ = ~new_n29238_ | ~new_n29237_;
  assign new_n29237_ = ~new_n29168_ | ~new_n28920_ | ~new_n28919_;
  assign new_n29238_ = ~new_n28879_ | ~new_n29227_ | ~new_n29168_;
  assign new_n29239_ = ~new_n29095_ | ~new_n29025_;
  assign new_n29240_ = ~new_n28895_;
  assign new_n29241_ = ~new_n28870_ | ~new_n29025_;
  assign new_n29242_ = ~new_n29023_;
  assign new_n29243_ = ~new_n28981_ | ~new_n29025_;
  assign new_n29244_ = ~new_n29021_;
  assign new_n29245_ = ~new_n29120_ | ~new_n29068_;
  assign new_n29246_ = ~new_n29066_;
  assign new_n29247_ = ~new_n28871_ | ~new_n29068_;
  assign new_n29248_ = ~new_n29065_;
  assign new_n29249_ = ~new_n28988_ | ~new_n29068_;
  assign new_n29250_ = ~new_n29063_;
  assign new_n29251_ = ~new_n28999_ | ~new_n29069_;
  assign new_n29252_ = ~new_n29000_ | ~new_n29069_;
  assign new_n29253_ = ~new_n8530_ | ~new_n29010_;
  assign new_n29254_ = ~new_n8794_ | ~new_n28880_;
  assign new_n29255_ = ~new_n28925_;
  assign new_n29256_ = ~new_n29255_ | ~new_n8460_;
  assign new_n29257_ = ~new_n28925_ | ~new_n28893_;
  assign new_n29258_ = ~new_n29255_ | ~new_n8460_;
  assign new_n29259_ = ~new_n28925_ | ~new_n28893_;
  assign new_n29260_ = ~new_n29259_ | ~new_n29258_;
  assign new_n29261_ = ~new_n8530_ | ~new_n29012_;
  assign new_n29262_ = ~new_n8779_ | ~new_n28880_;
  assign new_n29263_ = ~new_n28934_;
  assign new_n29264_ = ~new_n8530_ | ~new_n29013_;
  assign new_n29265_ = ~new_n8770_ | ~new_n28880_;
  assign new_n29266_ = ~new_n28932_;
  assign new_n29267_ = ~new_n8530_ | ~new_n29014_;
  assign new_n29268_ = ~new_n8765_ | ~new_n28880_;
  assign new_n29269_ = ~new_n28933_;
  assign new_n29270_ = ~new_n8530_ | ~new_n29015_;
  assign new_n29271_ = ~new_n8776_ | ~new_n28880_;
  assign new_n29272_ = ~new_n28931_;
  assign new_n29273_ = ~new_n8530_ | ~new_n29016_;
  assign new_n29274_ = ~new_n8773_ | ~new_n28880_;
  assign new_n29275_ = ~new_n28930_;
  assign new_n29276_ = ~new_n8530_ | ~new_n29017_;
  assign new_n29277_ = ~new_n8782_ | ~new_n28880_;
  assign new_n29278_ = ~new_n28929_;
  assign new_n29279_ = ~new_n8530_ | ~new_n29018_;
  assign new_n29280_ = ~new_n8788_ | ~new_n28880_;
  assign new_n29281_ = ~new_n28928_;
  assign new_n29282_ = ~new_n8530_ | ~new_n29019_;
  assign new_n29283_ = ~new_n8785_ | ~new_n28880_;
  assign new_n29284_ = ~new_n28927_;
  assign new_n29285_ = ~new_n8530_ | ~new_n29020_;
  assign new_n29286_ = ~new_n8791_ | ~new_n28880_;
  assign new_n29287_ = ~new_n28926_;
  assign new_n29288_ = ~new_n29011_ | ~new_n29021_;
  assign new_n29289_ = ~new_n29244_ | ~new_n29260_;
  assign new_n29290_ = ~new_n29287_ | ~new_n8461_;
  assign new_n29291_ = ~new_n28926_ | ~new_n28881_;
  assign new_n29292_ = ~new_n29287_ | ~new_n8461_;
  assign new_n29293_ = ~new_n28926_ | ~new_n28881_;
  assign new_n29294_ = ~new_n29293_ | ~new_n29292_;
  assign new_n29295_ = ~new_n29022_ | ~new_n29023_;
  assign new_n29296_ = ~new_n29242_ | ~new_n29294_;
  assign new_n29297_ = ~new_n29281_ | ~new_n8447_;
  assign new_n29298_ = ~new_n28928_ | ~new_n28884_;
  assign new_n29299_ = ~new_n29284_ | ~new_n8448_;
  assign new_n29300_ = ~new_n28927_ | ~new_n28882_;
  assign new_n29301_ = ~new_n29300_ | ~new_n29299_;
  assign new_n29302_ = ~new_n28895_ | ~new_n29207_;
  assign new_n29303_ = ~new_n29301_ | ~new_n29240_;
  assign new_n29304_ = ~new_n29278_ | ~new_n8444_;
  assign new_n29305_ = ~new_n28929_ | ~new_n28885_;
  assign new_n29306_ = ~new_n29278_ | ~new_n8444_;
  assign new_n29307_ = ~new_n28929_ | ~new_n28885_;
  assign new_n29308_ = ~new_n29307_ | ~new_n29306_;
  assign new_n29309_ = ~new_n29024_ | ~new_n29025_;
  assign new_n29310_ = ~new_n29094_ | ~new_n29308_;
  assign new_n29311_ = ~new_n29263_ | ~new_n8437_;
  assign new_n29312_ = ~new_n28934_ | ~new_n28892_;
  assign new_n29313_ = ~new_n29263_ | ~new_n8437_;
  assign new_n29314_ = ~new_n28934_ | ~new_n28892_;
  assign new_n29315_ = ~new_n29314_ | ~new_n29313_;
  assign new_n29316_ = ~new_n29026_ | ~new_n29027_;
  assign new_n29317_ = ~new_n29092_ | ~new_n29315_;
  assign new_n29318_ = ~new_n29272_ | ~new_n8441_;
  assign new_n29319_ = ~new_n28931_ | ~new_n28889_;
  assign new_n29320_ = ~new_n29275_ | ~new_n8445_;
  assign new_n29321_ = ~new_n28930_ | ~new_n28887_;
  assign new_n29322_ = ~new_n29321_ | ~new_n29320_;
  assign new_n29323_ = ~new_n29208_ | ~new_n28896_;
  assign new_n29324_ = ~new_n29322_ | ~new_n29085_;
  assign new_n29325_ = ~new_n8530_ | ~new_n29028_;
  assign new_n29326_ = ~new_n9278_ | ~new_n28880_;
  assign new_n29327_ = ~new_n28935_;
  assign new_n29328_ = ~new_n8530_ | ~new_n29029_;
  assign new_n29329_ = ~new_n8797_ | ~new_n28880_;
  assign new_n29330_ = ~new_n28945_;
  assign new_n29331_ = ~new_n8530_ | ~new_n29030_;
  assign new_n29332_ = ~new_n8800_ | ~new_n28880_;
  assign new_n29333_ = ~new_n28944_;
  assign new_n29334_ = ~new_n8530_ | ~new_n29031_;
  assign new_n29335_ = ~new_n8806_ | ~new_n28880_;
  assign new_n29336_ = ~new_n28943_;
  assign new_n29337_ = ~new_n8530_ | ~new_n29032_;
  assign new_n29338_ = ~new_n8803_ | ~new_n28880_;
  assign new_n29339_ = ~new_n28942_;
  assign new_n29340_ = ~new_n8530_ | ~new_n29033_;
  assign new_n29341_ = ~new_n8809_ | ~new_n28880_;
  assign new_n29342_ = ~new_n28941_;
  assign new_n29343_ = ~new_n8530_ | ~new_n29034_;
  assign new_n29344_ = ~new_n8812_ | ~new_n28880_;
  assign new_n29345_ = ~new_n28946_;
  assign new_n29346_ = ~new_n8530_ | ~new_n29035_;
  assign new_n29347_ = ~new_n8818_ | ~new_n28880_;
  assign new_n29348_ = ~new_n28940_;
  assign new_n29349_ = ~new_n8530_ | ~new_n29036_;
  assign new_n29350_ = ~new_n8815_ | ~new_n28880_;
  assign new_n29351_ = ~new_n28939_;
  assign new_n29352_ = ~new_n8530_ | ~new_n29037_;
  assign new_n29353_ = ~new_n8821_ | ~new_n28880_;
  assign new_n29354_ = ~new_n28947_;
  assign new_n29355_ = ~new_n8530_ | ~new_n29038_;
  assign new_n29356_ = ~new_n9284_ | ~new_n28880_;
  assign new_n29357_ = ~new_n28949_;
  assign new_n29358_ = ~new_n8530_ | ~new_n29039_;
  assign new_n29359_ = ~new_n9285_ | ~new_n28880_;
  assign new_n29360_ = ~new_n28950_;
  assign new_n29361_ = ~new_n8530_ | ~new_n29040_;
  assign new_n29362_ = ~new_n8823_ | ~new_n28880_;
  assign new_n29363_ = ~new_n28948_;
  assign new_n29364_ = ~new_n8530_ | ~new_n29041_;
  assign new_n29365_ = ~new_n9283_ | ~new_n28880_;
  assign new_n29366_ = ~new_n28951_;
  assign new_n29367_ = ~new_n8530_ | ~new_n29042_;
  assign new_n29368_ = ~new_n9282_ | ~new_n28880_;
  assign new_n29369_ = ~new_n28952_;
  assign new_n29370_ = ~new_n8530_ | ~new_n29043_;
  assign new_n29371_ = ~new_n9279_ | ~new_n28880_;
  assign new_n29372_ = ~new_n28938_;
  assign new_n29373_ = ~new_n8530_ | ~new_n29044_;
  assign new_n29374_ = ~new_n9280_ | ~new_n28880_;
  assign new_n29375_ = ~new_n28936_;
  assign new_n29376_ = ~new_n8530_ | ~new_n29045_;
  assign new_n29377_ = ~new_n9281_ | ~new_n28880_;
  assign new_n29378_ = ~new_n28937_;
  assign new_n29379_ = ~new_n8530_ | ~new_n29046_;
  assign new_n29380_ = ~new_n8431_ | ~new_n28880_;
  assign new_n29381_ = ~new_n28997_;
  assign new_n29382_ = ~new_n9277_ | ~new_n29381_;
  assign new_n29383_ = ~new_n28997_ | ~new_n29047_;
  assign new_n29384_ = ~new_n28953_;
  assign new_n29385_ = ~new_n29384_ | ~new_n29218_ | ~new_n29173_;
  assign new_n29386_ = ~new_n28953_ | ~new_n28996_ | ~new_n29235_;
  assign new_n29387_ = ~new_n29327_ | ~new_n8430_;
  assign new_n29388_ = ~new_n28935_ | ~new_n28897_;
  assign new_n29389_ = ~new_n29327_ | ~new_n8430_;
  assign new_n29390_ = ~new_n28935_ | ~new_n28897_;
  assign new_n29391_ = ~new_n29390_ | ~new_n29389_;
  assign new_n29392_ = ~new_n29048_ | ~new_n29049_;
  assign new_n29393_ = ~new_n29172_ | ~new_n29391_;
  assign new_n29394_ = ~new_n29372_ | ~new_n8434_;
  assign new_n29395_ = ~new_n28938_ | ~new_n28900_;
  assign new_n29396_ = ~new_n28964_ | ~new_n29050_;
  assign new_n29397_ = ~new_n28963_ | ~new_n29177_;
  assign new_n29398_ = ~new_n29375_ | ~new_n8435_;
  assign new_n29399_ = ~new_n28936_ | ~new_n28898_;
  assign new_n29400_ = ~new_n29399_ | ~new_n29398_;
  assign new_n29401_ = ~new_n29209_ | ~new_n29051_;
  assign new_n29402_ = ~new_n29178_ | ~new_n29400_;
  assign new_n29403_ = ~new_n29378_ | ~new_n8442_;
  assign new_n29404_ = ~new_n28937_ | ~new_n28899_;
  assign new_n29405_ = ~new_n29404_ | ~new_n29403_;
  assign new_n29406_ = ~new_n29210_ | ~new_n29052_;
  assign new_n29407_ = ~new_n29165_ | ~new_n29405_;
  assign new_n29408_ = ~new_n29369_ | ~new_n8443_;
  assign new_n29409_ = ~new_n28952_ | ~new_n28918_;
  assign new_n29410_ = ~new_n29369_ | ~new_n8443_;
  assign new_n29411_ = ~new_n28952_ | ~new_n28918_;
  assign new_n29412_ = ~new_n29411_ | ~new_n29410_;
  assign new_n29413_ = ~new_n29053_ | ~new_n29054_;
  assign new_n29414_ = ~new_n29161_ | ~new_n29412_;
  assign new_n29415_ = ~new_n29366_ | ~new_n8438_;
  assign new_n29416_ = ~new_n28951_ | ~new_n28917_;
  assign new_n29417_ = ~new_n29366_ | ~new_n8438_;
  assign new_n29418_ = ~new_n28951_ | ~new_n28917_;
  assign new_n29419_ = ~new_n29418_ | ~new_n29417_;
  assign new_n29420_ = ~new_n29055_ | ~new_n29056_;
  assign new_n29421_ = ~new_n29157_ | ~new_n29419_;
  assign new_n29422_ = ~new_n29357_ | ~new_n8452_;
  assign new_n29423_ = ~new_n28949_ | ~new_n28916_;
  assign new_n29424_ = ~new_n29360_ | ~new_n8453_;
  assign new_n29425_ = ~new_n28950_ | ~new_n28913_;
  assign new_n29426_ = ~new_n29425_ | ~new_n29424_;
  assign new_n29427_ = ~new_n29211_ | ~new_n28921_;
  assign new_n29428_ = ~new_n29426_ | ~new_n29183_;
  assign new_n29429_ = ~new_n29266_ | ~new_n8455_;
  assign new_n29430_ = ~new_n28932_ | ~new_n28890_;
  assign new_n29431_ = ~new_n29266_ | ~new_n8455_;
  assign new_n29432_ = ~new_n28932_ | ~new_n28890_;
  assign new_n29433_ = ~new_n29432_ | ~new_n29431_;
  assign new_n29434_ = ~new_n29057_ | ~new_n29058_;
  assign new_n29435_ = ~new_n29082_ | ~new_n29433_;
  assign new_n29436_ = ~new_n29363_ | ~new_n8458_;
  assign new_n29437_ = ~new_n28948_ | ~new_n28914_;
  assign new_n29438_ = ~new_n29437_ | ~new_n29436_;
  assign new_n29439_ = ~new_n29212_ | ~new_n29059_;
  assign new_n29440_ = ~new_n29147_ | ~new_n29438_;
  assign new_n29441_ = ~new_n29354_ | ~new_n8459_;
  assign new_n29442_ = ~new_n28947_ | ~new_n28912_;
  assign new_n29443_ = ~new_n29354_ | ~new_n8459_;
  assign new_n29444_ = ~new_n28947_ | ~new_n28912_;
  assign new_n29445_ = ~new_n29444_ | ~new_n29443_;
  assign new_n29446_ = ~new_n29060_ | ~new_n29061_;
  assign new_n29447_ = ~new_n29143_ | ~new_n29445_;
  assign new_n29448_ = ~new_n29348_ | ~new_n8446_;
  assign new_n29449_ = ~new_n28940_ | ~new_n28903_;
  assign new_n29450_ = ~new_n29351_ | ~new_n8450_;
  assign new_n29451_ = ~new_n28939_ | ~new_n28901_;
  assign new_n29452_ = ~new_n29451_ | ~new_n29450_;
  assign new_n29453_ = ~new_n29213_ | ~new_n28922_;
  assign new_n29454_ = ~new_n29452_ | ~new_n29135_;
  assign new_n29455_ = ~new_n29345_ | ~new_n8451_;
  assign new_n29456_ = ~new_n28946_ | ~new_n28911_;
  assign new_n29457_ = ~new_n29345_ | ~new_n8451_;
  assign new_n29458_ = ~new_n28946_ | ~new_n28911_;
  assign new_n29459_ = ~new_n29458_ | ~new_n29457_;
  assign new_n29460_ = ~new_n29062_ | ~new_n29063_;
  assign new_n29461_ = ~new_n29250_ | ~new_n29459_;
  assign new_n29462_ = ~new_n29342_ | ~new_n8456_;
  assign new_n29463_ = ~new_n28941_ | ~new_n28904_;
  assign new_n29464_ = ~new_n29342_ | ~new_n8456_;
  assign new_n29465_ = ~new_n28941_ | ~new_n28904_;
  assign new_n29466_ = ~new_n29465_ | ~new_n29464_;
  assign new_n29467_ = ~new_n29064_ | ~new_n29065_;
  assign new_n29468_ = ~new_n29248_ | ~new_n29466_;
  assign new_n29469_ = ~new_n29336_ | ~new_n8457_;
  assign new_n29470_ = ~new_n28943_ | ~new_n28908_;
  assign new_n29471_ = ~new_n29339_ | ~new_n8449_;
  assign new_n29472_ = ~new_n28942_ | ~new_n28905_;
  assign new_n29473_ = ~new_n29472_ | ~new_n29471_;
  assign new_n29474_ = ~new_n29214_ | ~new_n28924_;
  assign new_n29475_ = ~new_n29473_ | ~new_n29199_;
  assign new_n29476_ = ~new_n29333_ | ~new_n8440_;
  assign new_n29477_ = ~new_n28944_ | ~new_n28906_;
  assign new_n29478_ = ~new_n29477_ | ~new_n29476_;
  assign new_n29479_ = ~new_n29066_ | ~new_n29215_;
  assign new_n29480_ = ~new_n29246_ | ~new_n29478_;
  assign new_n29481_ = ~new_n29330_ | ~new_n8439_;
  assign new_n29482_ = ~new_n28945_ | ~new_n28909_;
  assign new_n29483_ = ~new_n29330_ | ~new_n8439_;
  assign new_n29484_ = ~new_n28945_ | ~new_n28909_;
  assign new_n29485_ = ~new_n29484_ | ~new_n29483_;
  assign new_n29486_ = ~new_n29067_ | ~new_n29068_;
  assign new_n29487_ = ~new_n29119_ | ~new_n29485_;
  assign new_n29488_ = ~new_n28933_ | ~new_n28880_;
  assign new_n29489_ = ~new_n29269_ | ~new_n8530_;
  assign new_n29490_ = ~new_n29009_;
  assign new_n29491_ = ~new_n29490_ | ~new_n8454_;
  assign new_n29492_ = ~new_n29009_ | ~new_n28891_;
  assign new_n29493_ = new_n29697_ & new_n29696_;
  assign new_n29494_ = new_n29676_ & new_n29732_;
  assign new_n29495_ = new_n29734_ & new_n29733_;
  assign new_n29496_ = new_n29677_ & new_n29749_;
  assign new_n29497_ = new_n29751_ & new_n29750_;
  assign new_n29498_ = new_n29678_ & new_n29773_;
  assign new_n29499_ = new_n29775_ & new_n29774_;
  assign new_n29500_ = new_n29700_ & new_n29695_ & new_n29681_;
  assign new_n29501_ = new_n29705_ & new_n29682_;
  assign new_n29502_ = new_n29879_ & new_n29878_;
  assign new_n29503_ = ~new_n29829_ | ~new_n29832_;
  assign new_n29504_ = ~new_n29818_ | ~new_n29821_;
  assign new_n29505_ = ~new_n29807_ | ~new_n29810_;
  assign new_n29506_ = ~new_n29799_ | ~new_n29801_;
  assign new_n29507_ = ~new_n29838_ | ~new_n29649_ | ~new_n29670_;
  assign new_n29508_ = ~new_n29728_ | ~new_n29730_;
  assign new_n29509_ = ~new_n29720_ | ~new_n29723_;
  assign new_n29510_ = ~new_n29712_ | ~new_n29714_;
  assign new_n29511_ = ~new_n29659_ | ~new_n29835_;
  assign new_n29512_ = ~new_n8447_;
  assign new_n29513_ = ~new_n8447_ | ~new_n29526_;
  assign new_n29514_ = ~new_n8461_;
  assign new_n29515_ = ~new_n8791_;
  assign new_n29516_ = ~new_n8773_;
  assign new_n29517_ = ~new_n8765_;
  assign new_n29518_ = ~new_n8455_;
  assign new_n29519_ = ~new_n8776_;
  assign new_n29520_ = ~new_n8445_;
  assign new_n29521_ = ~new_n8445_ | ~new_n29516_;
  assign new_n29522_ = ~new_n8441_;
  assign new_n29523_ = ~new_n8782_;
  assign new_n29524_ = ~new_n8785_;
  assign new_n29525_ = ~new_n8779_;
  assign new_n29526_ = ~new_n8788_;
  assign new_n29527_ = ~new_n8448_;
  assign new_n29528_ = ~new_n8444_;
  assign new_n29529_ = ~new_n8437_;
  assign new_n29530_ = ~new_n8437_ | ~new_n29525_;
  assign new_n29531_ = ~new_n29701_ | ~new_n29699_;
  assign new_n29532_ = ~new_n8794_;
  assign new_n29533_ = ~new_n8460_;
  assign new_n29534_ = ~new_n29531_ | ~new_n29702_;
  assign new_n29535_ = ~new_n29530_ | ~new_n29716_;
  assign new_n29536_ = ~new_n29836_ | ~new_n29688_ | ~new_n29672_;
  assign new_n29537_ = ~new_n9279_;
  assign new_n29538_ = ~new_n8800_;
  assign new_n29539_ = ~new_n8797_;
  assign new_n29540_ = ~new_n8440_;
  assign new_n29541_ = ~new_n8439_;
  assign new_n29542_ = ~new_n8460_ | ~new_n29532_;
  assign new_n29543_ = ~new_n8803_;
  assign new_n29544_ = ~new_n8449_;
  assign new_n29545_ = ~new_n8806_;
  assign new_n29546_ = ~new_n8457_;
  assign new_n29547_ = ~new_n8815_;
  assign new_n29548_ = ~new_n8812_;
  assign new_n29549_ = ~new_n8809_;
  assign new_n29550_ = ~new_n8450_;
  assign new_n29551_ = ~new_n8451_;
  assign new_n29552_ = ~new_n8456_;
  assign new_n29553_ = ~new_n8456_ | ~new_n29549_;
  assign new_n29554_ = ~new_n8818_;
  assign new_n29555_ = ~new_n8446_;
  assign new_n29556_ = ~new_n8459_;
  assign new_n29557_ = ~new_n8823_;
  assign new_n29558_ = ~new_n8458_;
  assign new_n29559_ = ~new_n9285_;
  assign new_n29560_ = ~new_n8453_;
  assign new_n29561_ = ~new_n9282_;
  assign new_n29562_ = ~new_n9283_;
  assign new_n29563_ = ~new_n9284_;
  assign new_n29564_ = ~new_n8443_;
  assign new_n29565_ = ~new_n8438_;
  assign new_n29566_ = ~new_n8452_;
  assign new_n29567_ = ~new_n8452_ | ~new_n29563_;
  assign new_n29568_ = ~new_n9281_;
  assign new_n29569_ = ~new_n8442_;
  assign new_n29570_ = ~new_n9280_;
  assign new_n29571_ = ~new_n8435_;
  assign new_n29572_ = ~new_n9278_;
  assign new_n29573_ = ~new_n8434_;
  assign new_n29574_ = ~new_n8434_ | ~new_n29537_;
  assign new_n29575_ = ~new_n8430_;
  assign new_n29576_ = ~new_n9277_;
  assign new_n29577_ = ~new_n8431_;
  assign new_n29578_ = ~new_n29789_ | ~new_n29788_;
  assign new_n29579_ = ~new_n29567_ | ~new_n29803_;
  assign new_n29580_ = ~new_n29553_ | ~new_n29814_;
  assign new_n29581_ = ~new_n29542_ | ~new_n29825_;
  assign new_n29582_ = ~new_n8454_;
  assign new_n29583_ = ~new_n29889_ | ~new_n29888_;
  assign new_n29584_ = ~new_n29903_ | ~new_n29902_;
  assign new_n29585_ = ~new_n29908_ | ~new_n29907_;
  assign new_n29586_ = ~new_n29924_ | ~new_n29923_;
  assign new_n29587_ = ~new_n29929_ | ~new_n29928_;
  assign new_n29588_ = ~new_n29934_ | ~new_n29933_;
  assign new_n29589_ = ~new_n29939_ | ~new_n29938_;
  assign new_n29590_ = ~new_n29944_ | ~new_n29943_;
  assign new_n29591_ = ~new_n29960_ | ~new_n29959_;
  assign new_n29592_ = ~new_n29965_ | ~new_n29964_;
  assign new_n29593_ = ~new_n29848_ | ~new_n29847_;
  assign new_n29594_ = ~new_n29857_ | ~new_n29856_;
  assign new_n29595_ = ~new_n29864_ | ~new_n29863_;
  assign new_n29596_ = ~new_n29868_ | ~new_n29867_;
  assign new_n29597_ = ~new_n29877_ | ~new_n29876_;
  assign new_n29598_ = ~new_n29898_ | ~new_n29897_;
  assign new_n29599_ = ~new_n29915_ | ~new_n29914_;
  assign new_n29600_ = ~new_n29919_ | ~new_n29918_;
  assign new_n29601_ = ~new_n29951_ | ~new_n29950_;
  assign new_n29602_ = ~new_n29955_ | ~new_n29954_;
  assign new_n29603_ = ~new_n29972_ | ~new_n29971_;
  assign new_n29604_ = new_n29839_ & new_n29680_;
  assign new_n29605_ = new_n29692_ & new_n29693_;
  assign new_n29606_ = new_n29501_ & new_n29500_;
  assign new_n29607_ = new_n29844_ & new_n29841_;
  assign new_n29608_ = new_n29513_ & new_n29850_ & new_n29849_;
  assign new_n29609_ = new_n29853_ & new_n29682_;
  assign new_n29610_ = new_n29722_ & new_n29493_;
  assign new_n29611_ = new_n29860_ & new_n29681_;
  assign new_n29612_ = new_n29521_ & new_n29870_ & new_n29869_;
  assign new_n29613_ = new_n29873_ & new_n29680_;
  assign new_n29614_ = new_n29709_ & new_n29494_;
  assign new_n29615_ = new_n29754_ & new_n29496_;
  assign new_n29616_ = new_n29778_ & new_n29498_;
  assign new_n29617_ = new_n29842_ & new_n29679_;
  assign new_n29618_ = new_n29793_ & new_n29794_;
  assign new_n29619_ = new_n29796_ & new_n29882_;
  assign new_n29620_ = new_n29793_ & new_n29794_;
  assign new_n29621_ = new_n29502_ & new_n29797_;
  assign new_n29622_ = ~new_n29886_ | ~new_n29885_;
  assign new_n29623_ = new_n29574_ & new_n29891_ & new_n29890_;
  assign new_n29624_ = new_n29894_ & new_n29679_;
  assign new_n29625_ = ~new_n29900_ | ~new_n29899_;
  assign new_n29626_ = ~new_n29905_ | ~new_n29904_;
  assign new_n29627_ = new_n29809_ & new_n29499_;
  assign new_n29628_ = new_n29911_ & new_n29678_;
  assign new_n29629_ = ~new_n29921_ | ~new_n29920_;
  assign new_n29630_ = ~new_n29926_ | ~new_n29925_;
  assign new_n29631_ = ~new_n29931_ | ~new_n29930_;
  assign new_n29632_ = ~new_n29936_ | ~new_n29935_;
  assign new_n29633_ = ~new_n29941_ | ~new_n29940_;
  assign new_n29634_ = new_n29820_ & new_n29497_;
  assign new_n29635_ = new_n29947_ & new_n29677_;
  assign new_n29636_ = ~new_n29957_ | ~new_n29956_;
  assign new_n29637_ = ~new_n29962_ | ~new_n29961_;
  assign new_n29638_ = new_n29831_ & new_n29495_;
  assign new_n29639_ = new_n29968_ & new_n29676_;
  assign new_n29640_ = new_n29846_ & new_n29845_;
  assign new_n29641_ = ~new_n29607_ | ~new_n29843_;
  assign new_n29642_ = new_n29855_ & new_n29854_;
  assign new_n29643_ = new_n29862_ & new_n29861_;
  assign new_n29644_ = new_n29866_ & new_n29865_;
  assign new_n29645_ = ~new_n29605_ | ~new_n29690_;
  assign new_n29646_ = new_n29875_ & new_n29874_;
  assign new_n29647_ = ~new_n9286_;
  assign new_n29648_ = ~new_n8432_;
  assign new_n29649_ = new_n29884_ & new_n29883_;
  assign new_n29650_ = ~new_n29618_ | ~new_n29791_;
  assign new_n29651_ = new_n29896_ & new_n29895_;
  assign new_n29652_ = ~new_n29785_ | ~new_n29784_;
  assign new_n29653_ = ~new_n29781_ | ~new_n29780_;
  assign new_n29654_ = new_n29913_ & new_n29912_;
  assign new_n29655_ = new_n29917_ & new_n29916_;
  assign new_n29656_ = ~new_n29771_ | ~new_n29770_;
  assign new_n29657_ = ~new_n29767_ | ~new_n29766_;
  assign new_n29658_ = ~new_n8770_;
  assign new_n29659_ = ~new_n8765_ | ~new_n29582_;
  assign new_n29660_ = ~new_n29837_ | ~new_n29763_ | ~new_n29671_;
  assign new_n29661_ = ~new_n8821_;
  assign new_n29662_ = ~new_n29761_ | ~new_n29760_;
  assign new_n29663_ = ~new_n29757_ | ~new_n29756_;
  assign new_n29664_ = new_n29949_ & new_n29948_;
  assign new_n29665_ = new_n29953_ & new_n29952_;
  assign new_n29666_ = ~new_n29747_ | ~new_n29746_;
  assign new_n29667_ = ~new_n29743_ | ~new_n29742_;
  assign new_n29668_ = ~new_n29739_ | ~new_n29738_;
  assign new_n29669_ = new_n29970_ & new_n29969_;
  assign new_n29670_ = ~new_n29619_ | ~new_n29650_;
  assign new_n29671_ = ~new_n29662_ | ~new_n29661_;
  assign new_n29672_ = ~new_n29659_ | ~new_n29658_;
  assign new_n29673_ = ~new_n29574_;
  assign new_n29674_ = ~new_n29521_;
  assign new_n29675_ = ~new_n29513_;
  assign new_n29676_ = ~new_n8797_ | ~new_n29541_;
  assign new_n29677_ = ~new_n8812_ | ~new_n29551_;
  assign new_n29678_ = ~new_n9283_ | ~new_n29565_;
  assign new_n29679_ = ~new_n9279_ | ~new_n29573_;
  assign new_n29680_ = ~new_n8773_ | ~new_n29520_;
  assign new_n29681_ = ~new_n8782_ | ~new_n29528_;
  assign new_n29682_ = ~new_n8788_ | ~new_n29512_;
  assign new_n29683_ = ~new_n29553_;
  assign new_n29684_ = ~new_n29567_;
  assign new_n29685_ = ~new_n29530_;
  assign new_n29686_ = ~new_n29542_;
  assign new_n29687_ = ~new_n29659_;
  assign new_n29688_ = ~new_n8455_ | ~new_n29659_;
  assign new_n29689_ = ~new_n29536_;
  assign new_n29690_ = ~new_n29604_ | ~new_n29536_;
  assign new_n29691_ = ~new_n29522_ | ~new_n29521_;
  assign new_n29692_ = ~new_n29691_ | ~new_n29519_;
  assign new_n29693_ = ~new_n8441_ | ~new_n29674_;
  assign new_n29694_ = ~new_n29645_;
  assign new_n29695_ = ~new_n8785_ | ~new_n29527_;
  assign new_n29696_ = ~new_n8448_ | ~new_n29524_;
  assign new_n29697_ = ~new_n8444_ | ~new_n29523_;
  assign new_n29698_ = ~new_n29685_ | ~new_n29681_;
  assign new_n29699_ = ~new_n29493_ | ~new_n29698_;
  assign new_n29700_ = ~new_n8779_ | ~new_n29529_;
  assign new_n29701_ = ~new_n8785_ | ~new_n29527_;
  assign new_n29702_ = ~new_n29500_ | ~new_n29645_;
  assign new_n29703_ = ~new_n29531_;
  assign new_n29704_ = ~new_n29534_;
  assign new_n29705_ = ~new_n8791_ | ~new_n29514_;
  assign new_n29706_ = ~new_n29514_ | ~new_n29513_;
  assign new_n29707_ = ~new_n8461_ | ~new_n29675_;
  assign new_n29708_ = ~new_n29641_;
  assign new_n29709_ = ~new_n8794_ | ~new_n29533_;
  assign new_n29710_ = ~new_n29709_ | ~new_n29542_;
  assign new_n29711_ = ~new_n29704_ | ~new_n29513_;
  assign new_n29712_ = ~new_n29609_ | ~new_n29711_;
  assign new_n29713_ = ~new_n29534_ | ~new_n29682_;
  assign new_n29714_ = ~new_n29608_ | ~new_n29713_;
  assign new_n29715_ = ~new_n29513_ | ~new_n29682_;
  assign new_n29716_ = ~new_n29700_ | ~new_n29645_;
  assign new_n29717_ = ~new_n29535_;
  assign new_n29718_ = ~new_n8444_ | ~new_n29523_;
  assign new_n29719_ = ~new_n29717_ | ~new_n29718_;
  assign new_n29720_ = ~new_n29611_ | ~new_n29719_;
  assign new_n29721_ = ~new_n29535_ | ~new_n29681_;
  assign new_n29722_ = ~new_n8785_ | ~new_n29527_;
  assign new_n29723_ = ~new_n29610_ | ~new_n29721_;
  assign new_n29724_ = ~new_n8444_ | ~new_n29523_;
  assign new_n29725_ = ~new_n29681_ | ~new_n29724_;
  assign new_n29726_ = ~new_n29700_ | ~new_n29530_;
  assign new_n29727_ = ~new_n29689_ | ~new_n29521_;
  assign new_n29728_ = ~new_n29613_ | ~new_n29727_;
  assign new_n29729_ = ~new_n29536_ | ~new_n29680_;
  assign new_n29730_ = ~new_n29612_ | ~new_n29729_;
  assign new_n29731_ = ~new_n29680_ | ~new_n29521_;
  assign new_n29732_ = ~new_n8800_ | ~new_n29540_;
  assign new_n29733_ = ~new_n8440_ | ~new_n29538_;
  assign new_n29734_ = ~new_n8439_ | ~new_n29539_;
  assign new_n29735_ = ~new_n29686_ | ~new_n29494_;
  assign new_n29736_ = ~new_n29495_ | ~new_n29735_;
  assign new_n29737_ = ~new_n8800_ | ~new_n29540_;
  assign new_n29738_ = ~new_n29614_ | ~new_n29641_;
  assign new_n29739_ = ~new_n29737_ | ~new_n29736_;
  assign new_n29740_ = ~new_n29668_;
  assign new_n29741_ = ~new_n8803_ | ~new_n29544_;
  assign new_n29742_ = ~new_n29741_ | ~new_n29668_;
  assign new_n29743_ = ~new_n8449_ | ~new_n29543_;
  assign new_n29744_ = ~new_n29667_;
  assign new_n29745_ = ~new_n8806_ | ~new_n29546_;
  assign new_n29746_ = ~new_n29745_ | ~new_n29667_;
  assign new_n29747_ = ~new_n8457_ | ~new_n29545_;
  assign new_n29748_ = ~new_n29666_;
  assign new_n29749_ = ~new_n8815_ | ~new_n29550_;
  assign new_n29750_ = ~new_n8450_ | ~new_n29547_;
  assign new_n29751_ = ~new_n8451_ | ~new_n29548_;
  assign new_n29752_ = ~new_n29683_ | ~new_n29496_;
  assign new_n29753_ = ~new_n29497_ | ~new_n29752_;
  assign new_n29754_ = ~new_n8809_ | ~new_n29552_;
  assign new_n29755_ = ~new_n8815_ | ~new_n29550_;
  assign new_n29756_ = ~new_n29615_ | ~new_n29666_;
  assign new_n29757_ = ~new_n29755_ | ~new_n29753_;
  assign new_n29758_ = ~new_n29663_;
  assign new_n29759_ = ~new_n8818_ | ~new_n29555_;
  assign new_n29760_ = ~new_n29759_ | ~new_n29663_;
  assign new_n29761_ = ~new_n8446_ | ~new_n29554_;
  assign new_n29762_ = ~new_n29662_;
  assign new_n29763_ = ~new_n8459_ | ~new_n29662_;
  assign new_n29764_ = ~new_n29660_;
  assign new_n29765_ = ~new_n8823_ | ~new_n29558_;
  assign new_n29766_ = ~new_n29765_ | ~new_n29660_;
  assign new_n29767_ = ~new_n8458_ | ~new_n29557_;
  assign new_n29768_ = ~new_n29657_;
  assign new_n29769_ = ~new_n9285_ | ~new_n29560_;
  assign new_n29770_ = ~new_n29769_ | ~new_n29657_;
  assign new_n29771_ = ~new_n8453_ | ~new_n29559_;
  assign new_n29772_ = ~new_n29656_;
  assign new_n29773_ = ~new_n9282_ | ~new_n29564_;
  assign new_n29774_ = ~new_n8443_ | ~new_n29561_;
  assign new_n29775_ = ~new_n8438_ | ~new_n29562_;
  assign new_n29776_ = ~new_n29684_ | ~new_n29498_;
  assign new_n29777_ = ~new_n29499_ | ~new_n29776_;
  assign new_n29778_ = ~new_n9284_ | ~new_n29566_;
  assign new_n29779_ = ~new_n9282_ | ~new_n29564_;
  assign new_n29780_ = ~new_n29616_ | ~new_n29656_;
  assign new_n29781_ = ~new_n29779_ | ~new_n29777_;
  assign new_n29782_ = ~new_n29653_;
  assign new_n29783_ = ~new_n9281_ | ~new_n29569_;
  assign new_n29784_ = ~new_n29783_ | ~new_n29653_;
  assign new_n29785_ = ~new_n8442_ | ~new_n29568_;
  assign new_n29786_ = ~new_n29652_;
  assign new_n29787_ = ~new_n9280_ | ~new_n29571_;
  assign new_n29788_ = ~new_n29787_ | ~new_n29652_;
  assign new_n29789_ = ~new_n8435_ | ~new_n29570_;
  assign new_n29790_ = ~new_n29578_;
  assign new_n29791_ = ~new_n29617_ | ~new_n29578_;
  assign new_n29792_ = ~new_n29575_ | ~new_n29574_;
  assign new_n29793_ = ~new_n29792_ | ~new_n29572_;
  assign new_n29794_ = ~new_n8430_ | ~new_n29673_;
  assign new_n29795_ = ~new_n29650_;
  assign new_n29796_ = ~new_n9277_ | ~new_n29577_;
  assign new_n29797_ = ~new_n8431_ | ~new_n29576_;
  assign new_n29798_ = ~new_n29790_ | ~new_n29574_;
  assign new_n29799_ = ~new_n29624_ | ~new_n29798_;
  assign new_n29800_ = ~new_n29578_ | ~new_n29679_;
  assign new_n29801_ = ~new_n29623_ | ~new_n29800_;
  assign new_n29802_ = ~new_n29679_ | ~new_n29574_;
  assign new_n29803_ = ~new_n29778_ | ~new_n29656_;
  assign new_n29804_ = ~new_n29579_;
  assign new_n29805_ = ~new_n8438_ | ~new_n29562_;
  assign new_n29806_ = ~new_n29804_ | ~new_n29805_;
  assign new_n29807_ = ~new_n29628_ | ~new_n29806_;
  assign new_n29808_ = ~new_n29579_ | ~new_n29678_;
  assign new_n29809_ = ~new_n9282_ | ~new_n29564_;
  assign new_n29810_ = ~new_n29627_ | ~new_n29808_;
  assign new_n29811_ = ~new_n8438_ | ~new_n29562_;
  assign new_n29812_ = ~new_n29678_ | ~new_n29811_;
  assign new_n29813_ = ~new_n29778_ | ~new_n29567_;
  assign new_n29814_ = ~new_n29754_ | ~new_n29666_;
  assign new_n29815_ = ~new_n29580_;
  assign new_n29816_ = ~new_n8451_ | ~new_n29548_;
  assign new_n29817_ = ~new_n29815_ | ~new_n29816_;
  assign new_n29818_ = ~new_n29635_ | ~new_n29817_;
  assign new_n29819_ = ~new_n29580_ | ~new_n29677_;
  assign new_n29820_ = ~new_n8815_ | ~new_n29550_;
  assign new_n29821_ = ~new_n29634_ | ~new_n29819_;
  assign new_n29822_ = ~new_n8451_ | ~new_n29548_;
  assign new_n29823_ = ~new_n29677_ | ~new_n29822_;
  assign new_n29824_ = ~new_n29754_ | ~new_n29553_;
  assign new_n29825_ = ~new_n29709_ | ~new_n29641_;
  assign new_n29826_ = ~new_n29581_;
  assign new_n29827_ = ~new_n8439_ | ~new_n29539_;
  assign new_n29828_ = ~new_n29826_ | ~new_n29827_;
  assign new_n29829_ = ~new_n29639_ | ~new_n29828_;
  assign new_n29830_ = ~new_n29581_ | ~new_n29676_;
  assign new_n29831_ = ~new_n8800_ | ~new_n29540_;
  assign new_n29832_ = ~new_n29638_ | ~new_n29830_;
  assign new_n29833_ = ~new_n8439_ | ~new_n29539_;
  assign new_n29834_ = ~new_n29676_ | ~new_n29833_;
  assign new_n29835_ = ~new_n8454_ | ~new_n29517_;
  assign new_n29836_ = ~new_n8455_ | ~new_n29658_;
  assign new_n29837_ = ~new_n8459_ | ~new_n29661_;
  assign new_n29838_ = ~new_n29621_ | ~new_n29620_ | ~new_n29791_;
  assign new_n29839_ = ~new_n8776_ | ~new_n29522_;
  assign new_n29840_ = ~new_n8791_ | ~new_n29707_;
  assign new_n29841_ = ~new_n29840_ | ~new_n29706_;
  assign new_n29842_ = ~new_n9278_ | ~new_n29575_;
  assign new_n29843_ = ~new_n29606_ | ~new_n29645_;
  assign new_n29844_ = ~new_n29703_ | ~new_n29501_;
  assign new_n29845_ = ~new_n8794_ | ~new_n29533_;
  assign new_n29846_ = ~new_n8460_ | ~new_n29532_;
  assign new_n29847_ = ~new_n29710_ | ~new_n29641_;
  assign new_n29848_ = ~new_n29708_ | ~new_n29640_;
  assign new_n29849_ = ~new_n8791_ | ~new_n29514_;
  assign new_n29850_ = ~new_n8461_ | ~new_n29515_;
  assign new_n29851_ = ~new_n8791_ | ~new_n29514_;
  assign new_n29852_ = ~new_n8461_ | ~new_n29515_;
  assign new_n29853_ = ~new_n29852_ | ~new_n29851_;
  assign new_n29854_ = ~new_n8788_ | ~new_n29512_;
  assign new_n29855_ = ~new_n8447_ | ~new_n29526_;
  assign new_n29856_ = ~new_n29715_ | ~new_n29534_;
  assign new_n29857_ = ~new_n29642_ | ~new_n29704_;
  assign new_n29858_ = ~new_n8785_ | ~new_n29527_;
  assign new_n29859_ = ~new_n8448_ | ~new_n29524_;
  assign new_n29860_ = ~new_n29859_ | ~new_n29858_;
  assign new_n29861_ = ~new_n8782_ | ~new_n29528_;
  assign new_n29862_ = ~new_n8444_ | ~new_n29523_;
  assign new_n29863_ = ~new_n29725_ | ~new_n29535_;
  assign new_n29864_ = ~new_n29643_ | ~new_n29717_;
  assign new_n29865_ = ~new_n8779_ | ~new_n29529_;
  assign new_n29866_ = ~new_n8437_ | ~new_n29525_;
  assign new_n29867_ = ~new_n29726_ | ~new_n29645_;
  assign new_n29868_ = ~new_n29694_ | ~new_n29644_;
  assign new_n29869_ = ~new_n8776_ | ~new_n29522_;
  assign new_n29870_ = ~new_n8441_ | ~new_n29519_;
  assign new_n29871_ = ~new_n8776_ | ~new_n29522_;
  assign new_n29872_ = ~new_n8441_ | ~new_n29519_;
  assign new_n29873_ = ~new_n29872_ | ~new_n29871_;
  assign new_n29874_ = ~new_n8773_ | ~new_n29520_;
  assign new_n29875_ = ~new_n8445_ | ~new_n29516_;
  assign new_n29876_ = ~new_n29731_ | ~new_n29536_;
  assign new_n29877_ = ~new_n29646_ | ~new_n29689_;
  assign new_n29878_ = ~new_n9286_ | ~new_n29648_;
  assign new_n29879_ = ~new_n8432_ | ~new_n29647_;
  assign new_n29880_ = ~new_n9286_ | ~new_n29648_;
  assign new_n29881_ = ~new_n8432_ | ~new_n29647_;
  assign new_n29882_ = ~new_n29881_ | ~new_n29880_;
  assign new_n29883_ = ~new_n29576_ | ~new_n8431_ | ~new_n29882_;
  assign new_n29884_ = ~new_n9277_ | ~new_n29502_ | ~new_n29577_;
  assign new_n29885_ = ~new_n9277_ | ~new_n29577_;
  assign new_n29886_ = ~new_n8431_ | ~new_n29576_;
  assign new_n29887_ = ~new_n29622_;
  assign new_n29888_ = ~new_n29795_ | ~new_n29887_;
  assign new_n29889_ = ~new_n29622_ | ~new_n29650_;
  assign new_n29890_ = ~new_n9278_ | ~new_n29575_;
  assign new_n29891_ = ~new_n8430_ | ~new_n29572_;
  assign new_n29892_ = ~new_n9278_ | ~new_n29575_;
  assign new_n29893_ = ~new_n8430_ | ~new_n29572_;
  assign new_n29894_ = ~new_n29893_ | ~new_n29892_;
  assign new_n29895_ = ~new_n9279_ | ~new_n29573_;
  assign new_n29896_ = ~new_n8434_ | ~new_n29537_;
  assign new_n29897_ = ~new_n29802_ | ~new_n29578_;
  assign new_n29898_ = ~new_n29651_ | ~new_n29790_;
  assign new_n29899_ = ~new_n9280_ | ~new_n29571_;
  assign new_n29900_ = ~new_n8435_ | ~new_n29570_;
  assign new_n29901_ = ~new_n29625_;
  assign new_n29902_ = ~new_n29786_ | ~new_n29901_;
  assign new_n29903_ = ~new_n29625_ | ~new_n29652_;
  assign new_n29904_ = ~new_n9281_ | ~new_n29569_;
  assign new_n29905_ = ~new_n8442_ | ~new_n29568_;
  assign new_n29906_ = ~new_n29626_;
  assign new_n29907_ = ~new_n29782_ | ~new_n29906_;
  assign new_n29908_ = ~new_n29626_ | ~new_n29653_;
  assign new_n29909_ = ~new_n9282_ | ~new_n29564_;
  assign new_n29910_ = ~new_n8443_ | ~new_n29561_;
  assign new_n29911_ = ~new_n29910_ | ~new_n29909_;
  assign new_n29912_ = ~new_n9283_ | ~new_n29565_;
  assign new_n29913_ = ~new_n8438_ | ~new_n29562_;
  assign new_n29914_ = ~new_n29812_ | ~new_n29579_;
  assign new_n29915_ = ~new_n29654_ | ~new_n29804_;
  assign new_n29916_ = ~new_n9284_ | ~new_n29566_;
  assign new_n29917_ = ~new_n8452_ | ~new_n29563_;
  assign new_n29918_ = ~new_n29813_ | ~new_n29656_;
  assign new_n29919_ = ~new_n29772_ | ~new_n29655_;
  assign new_n29920_ = ~new_n9285_ | ~new_n29560_;
  assign new_n29921_ = ~new_n8453_ | ~new_n29559_;
  assign new_n29922_ = ~new_n29629_;
  assign new_n29923_ = ~new_n29768_ | ~new_n29922_;
  assign new_n29924_ = ~new_n29629_ | ~new_n29657_;
  assign new_n29925_ = ~new_n8770_ | ~new_n29518_;
  assign new_n29926_ = ~new_n8455_ | ~new_n29658_;
  assign new_n29927_ = ~new_n29630_;
  assign new_n29928_ = ~new_n29687_ | ~new_n29927_;
  assign new_n29929_ = ~new_n29630_ | ~new_n29659_;
  assign new_n29930_ = ~new_n8823_ | ~new_n29558_;
  assign new_n29931_ = ~new_n8458_ | ~new_n29557_;
  assign new_n29932_ = ~new_n29631_;
  assign new_n29933_ = ~new_n29764_ | ~new_n29932_;
  assign new_n29934_ = ~new_n29631_ | ~new_n29660_;
  assign new_n29935_ = ~new_n8821_ | ~new_n29556_;
  assign new_n29936_ = ~new_n8459_ | ~new_n29661_;
  assign new_n29937_ = ~new_n29632_;
  assign new_n29938_ = ~new_n29762_ | ~new_n29937_;
  assign new_n29939_ = ~new_n29632_ | ~new_n29662_;
  assign new_n29940_ = ~new_n8818_ | ~new_n29555_;
  assign new_n29941_ = ~new_n8446_ | ~new_n29554_;
  assign new_n29942_ = ~new_n29633_;
  assign new_n29943_ = ~new_n29758_ | ~new_n29942_;
  assign new_n29944_ = ~new_n29633_ | ~new_n29663_;
  assign new_n29945_ = ~new_n8815_ | ~new_n29550_;
  assign new_n29946_ = ~new_n8450_ | ~new_n29547_;
  assign new_n29947_ = ~new_n29946_ | ~new_n29945_;
  assign new_n29948_ = ~new_n8812_ | ~new_n29551_;
  assign new_n29949_ = ~new_n8451_ | ~new_n29548_;
  assign new_n29950_ = ~new_n29823_ | ~new_n29580_;
  assign new_n29951_ = ~new_n29664_ | ~new_n29815_;
  assign new_n29952_ = ~new_n8809_ | ~new_n29552_;
  assign new_n29953_ = ~new_n8456_ | ~new_n29549_;
  assign new_n29954_ = ~new_n29824_ | ~new_n29666_;
  assign new_n29955_ = ~new_n29748_ | ~new_n29665_;
  assign new_n29956_ = ~new_n8806_ | ~new_n29546_;
  assign new_n29957_ = ~new_n8457_ | ~new_n29545_;
  assign new_n29958_ = ~new_n29636_;
  assign new_n29959_ = ~new_n29744_ | ~new_n29958_;
  assign new_n29960_ = ~new_n29636_ | ~new_n29667_;
  assign new_n29961_ = ~new_n8803_ | ~new_n29544_;
  assign new_n29962_ = ~new_n8449_ | ~new_n29543_;
  assign new_n29963_ = ~new_n29637_;
  assign new_n29964_ = ~new_n29740_ | ~new_n29963_;
  assign new_n29965_ = ~new_n29637_ | ~new_n29668_;
  assign new_n29966_ = ~new_n8800_ | ~new_n29540_;
  assign new_n29967_ = ~new_n8440_ | ~new_n29538_;
  assign new_n29968_ = ~new_n29967_ | ~new_n29966_;
  assign new_n29969_ = ~new_n8797_ | ~new_n29541_;
  assign new_n29970_ = ~new_n8439_ | ~new_n29539_;
  assign new_n29971_ = ~new_n29834_ | ~new_n29581_;
  assign new_n29972_ = ~new_n29669_ | ~new_n29826_;
  assign new_n29973_ = new_n30069_ & new_n30085_;
  assign new_n29974_ = new_n30087_ & new_n30086_;
  assign new_n29975_ = new_n30066_ & new_n30124_;
  assign new_n29976_ = new_n30126_ & new_n30125_;
  assign new_n29977_ = new_n30067_ & new_n30141_;
  assign new_n29978_ = new_n30143_ & new_n30142_;
  assign new_n29979_ = ~new_n30174_ | ~new_n30177_;
  assign new_n29980_ = ~new_n30163_ | ~new_n30166_;
  assign new_n29981_ = ~new_n30120_ | ~new_n30122_;
  assign new_n29982_ = ~new_n30112_ | ~new_n30115_;
  assign new_n29983_ = ~new_n30104_ | ~new_n30106_;
  assign new_n29984_ = ~new_n29988_ | ~new_n30180_;
  assign new_n29985_ = ~new_n8787_;
  assign new_n29986_ = ~new_n8772_;
  assign new_n29987_ = ~new_n8764_;
  assign new_n29988_ = ~new_n8764_ | ~new_n30032_;
  assign new_n29989_ = ~new_n8951_;
  assign new_n29990_ = ~new_n8775_;
  assign new_n29991_ = ~new_n8940_;
  assign new_n29992_ = ~new_n8940_ | ~new_n29986_;
  assign new_n29993_ = ~new_n8939_;
  assign new_n29994_ = ~new_n8784_;
  assign new_n29995_ = ~new_n8781_;
  assign new_n29996_ = ~new_n8778_;
  assign new_n29997_ = ~new_n8936_;
  assign new_n29998_ = ~new_n8937_;
  assign new_n29999_ = ~new_n8938_;
  assign new_n30000_ = ~new_n8938_ | ~new_n29996_;
  assign new_n30001_ = ~new_n8790_;
  assign new_n30002_ = ~new_n8935_;
  assign new_n30003_ = ~new_n8935_ | ~new_n29985_;
  assign new_n30004_ = ~new_n8934_;
  assign new_n30005_ = ~new_n8793_;
  assign new_n30006_ = ~new_n8933_;
  assign new_n30007_ = ~new_n30093_ | ~new_n30092_;
  assign new_n30008_ = ~new_n30000_ | ~new_n30108_;
  assign new_n30009_ = ~new_n30077_ | ~new_n30076_;
  assign new_n30010_ = ~new_n8799_;
  assign new_n30011_ = ~new_n8796_;
  assign new_n30012_ = ~new_n8949_;
  assign new_n30013_ = ~new_n8950_;
  assign new_n30014_ = ~new_n8933_ | ~new_n30005_;
  assign new_n30015_ = ~new_n8802_;
  assign new_n30016_ = ~new_n8948_;
  assign new_n30017_ = ~new_n8805_;
  assign new_n30018_ = ~new_n8947_;
  assign new_n30019_ = ~new_n8814_;
  assign new_n30020_ = ~new_n8811_;
  assign new_n30021_ = ~new_n8808_;
  assign new_n30022_ = ~new_n8944_;
  assign new_n30023_ = ~new_n8945_;
  assign new_n30024_ = ~new_n8946_;
  assign new_n30025_ = ~new_n8946_ | ~new_n30021_;
  assign new_n30026_ = ~new_n8817_;
  assign new_n30027_ = ~new_n8943_;
  assign new_n30028_ = ~new_n30153_ | ~new_n30152_;
  assign new_n30029_ = ~new_n8942_;
  assign new_n30030_ = ~new_n30025_ | ~new_n30159_;
  assign new_n30031_ = ~new_n30014_ | ~new_n30170_;
  assign new_n30032_ = ~new_n8952_;
  assign new_n30033_ = ~new_n30218_ | ~new_n30217_;
  assign new_n30034_ = ~new_n30223_ | ~new_n30222_;
  assign new_n30035_ = ~new_n30228_ | ~new_n30227_;
  assign new_n30036_ = ~new_n30233_ | ~new_n30232_;
  assign new_n30037_ = ~new_n30249_ | ~new_n30248_;
  assign new_n30038_ = ~new_n30254_ | ~new_n30253_;
  assign new_n30039_ = ~new_n30184_ | ~new_n30183_;
  assign new_n30040_ = ~new_n30193_ | ~new_n30192_;
  assign new_n30041_ = ~new_n30200_ | ~new_n30199_;
  assign new_n30042_ = ~new_n30204_ | ~new_n30203_;
  assign new_n30043_ = ~new_n30213_ | ~new_n30212_;
  assign new_n30044_ = ~new_n30240_ | ~new_n30239_;
  assign new_n30045_ = ~new_n30244_ | ~new_n30243_;
  assign new_n30046_ = ~new_n30261_ | ~new_n30260_;
  assign new_n30047_ = ~new_n30215_ | ~new_n30214_;
  assign new_n30048_ = ~new_n30220_ | ~new_n30219_;
  assign new_n30049_ = ~new_n30225_ | ~new_n30224_;
  assign new_n30050_ = ~new_n30230_ | ~new_n30229_;
  assign new_n30051_ = ~new_n30246_ | ~new_n30245_;
  assign new_n30052_ = ~new_n30251_ | ~new_n30250_;
  assign new_n30053_ = ~new_n30096_ | ~new_n30098_ | ~new_n30099_;
  assign new_n30054_ = ~new_n30080_ | ~new_n30082_ | ~new_n30083_;
  assign new_n30055_ = ~new_n8769_;
  assign new_n30056_ = ~new_n8757_;
  assign new_n30057_ = ~new_n8941_;
  assign new_n30058_ = ~new_n30157_ | ~new_n30156_;
  assign new_n30059_ = ~new_n8820_;
  assign new_n30060_ = ~new_n30149_ | ~new_n30148_;
  assign new_n30061_ = ~new_n30139_ | ~new_n30138_;
  assign new_n30062_ = ~new_n30135_ | ~new_n30134_;
  assign new_n30063_ = ~new_n30131_ | ~new_n30130_;
  assign new_n30064_ = ~new_n29992_;
  assign new_n30065_ = ~new_n30003_;
  assign new_n30066_ = ~new_n8796_ | ~new_n30013_;
  assign new_n30067_ = ~new_n8811_ | ~new_n30023_;
  assign new_n30068_ = ~new_n8772_ | ~new_n29991_;
  assign new_n30069_ = ~new_n8781_ | ~new_n29998_;
  assign new_n30070_ = ~new_n8787_ | ~new_n30002_;
  assign new_n30071_ = ~new_n30025_;
  assign new_n30072_ = ~new_n30000_;
  assign new_n30073_ = ~new_n30014_;
  assign new_n30074_ = ~new_n29988_;
  assign new_n30075_ = ~new_n30074_ | ~new_n29989_;
  assign new_n30076_ = ~new_n30075_ | ~new_n30055_;
  assign new_n30077_ = ~new_n8951_ | ~new_n29988_;
  assign new_n30078_ = ~new_n30009_;
  assign new_n30079_ = ~new_n8775_ | ~new_n29993_;
  assign new_n30080_ = ~new_n30009_ | ~new_n30079_ | ~new_n30068_;
  assign new_n30081_ = ~new_n29993_ | ~new_n29992_;
  assign new_n30082_ = ~new_n30081_ | ~new_n29990_;
  assign new_n30083_ = ~new_n8939_ | ~new_n30064_;
  assign new_n30084_ = ~new_n30054_;
  assign new_n30085_ = ~new_n8784_ | ~new_n29997_;
  assign new_n30086_ = ~new_n8936_ | ~new_n29994_;
  assign new_n30087_ = ~new_n8937_ | ~new_n29995_;
  assign new_n30088_ = ~new_n30072_ | ~new_n29973_;
  assign new_n30089_ = ~new_n29974_ | ~new_n30088_;
  assign new_n30090_ = ~new_n8778_ | ~new_n29999_;
  assign new_n30091_ = ~new_n8784_ | ~new_n29997_;
  assign new_n30092_ = ~new_n30054_ | ~new_n30090_ | ~new_n29973_;
  assign new_n30093_ = ~new_n30091_ | ~new_n30089_;
  assign new_n30094_ = ~new_n30007_;
  assign new_n30095_ = ~new_n8790_ | ~new_n30004_;
  assign new_n30096_ = ~new_n30007_ | ~new_n30095_ | ~new_n30070_;
  assign new_n30097_ = ~new_n30004_ | ~new_n30003_;
  assign new_n30098_ = ~new_n30097_ | ~new_n30001_;
  assign new_n30099_ = ~new_n8934_ | ~new_n30065_;
  assign new_n30100_ = ~new_n30053_;
  assign new_n30101_ = ~new_n8793_ | ~new_n30006_;
  assign new_n30102_ = ~new_n30101_ | ~new_n30014_;
  assign new_n30103_ = ~new_n30094_ | ~new_n30003_;
  assign new_n30104_ = ~new_n30103_ | ~new_n30189_ | ~new_n30070_;
  assign new_n30105_ = ~new_n30007_ | ~new_n30070_;
  assign new_n30106_ = ~new_n30185_ | ~new_n30105_ | ~new_n30003_ | ~new_n30186_;
  assign new_n30107_ = ~new_n30003_ | ~new_n30070_;
  assign new_n30108_ = ~new_n30090_ | ~new_n30054_;
  assign new_n30109_ = ~new_n30008_;
  assign new_n30110_ = ~new_n8937_ | ~new_n29995_;
  assign new_n30111_ = ~new_n30109_ | ~new_n30110_;
  assign new_n30112_ = ~new_n30111_ | ~new_n30196_ | ~new_n30069_;
  assign new_n30113_ = ~new_n30008_ | ~new_n30069_;
  assign new_n30114_ = ~new_n8784_ | ~new_n29997_;
  assign new_n30115_ = ~new_n30113_ | ~new_n30114_ | ~new_n29974_;
  assign new_n30116_ = ~new_n8937_ | ~new_n29995_;
  assign new_n30117_ = ~new_n30069_ | ~new_n30116_;
  assign new_n30118_ = ~new_n30090_ | ~new_n30000_;
  assign new_n30119_ = ~new_n30078_ | ~new_n29992_;
  assign new_n30120_ = ~new_n30119_ | ~new_n30209_ | ~new_n30068_;
  assign new_n30121_ = ~new_n30009_ | ~new_n30068_;
  assign new_n30122_ = ~new_n30205_ | ~new_n30121_ | ~new_n29992_ | ~new_n30206_;
  assign new_n30123_ = ~new_n29992_ | ~new_n30068_;
  assign new_n30124_ = ~new_n8799_ | ~new_n30012_;
  assign new_n30125_ = ~new_n8949_ | ~new_n30010_;
  assign new_n30126_ = ~new_n8950_ | ~new_n30011_;
  assign new_n30127_ = ~new_n30073_ | ~new_n29975_;
  assign new_n30128_ = ~new_n29976_ | ~new_n30127_;
  assign new_n30129_ = ~new_n8799_ | ~new_n30012_;
  assign new_n30130_ = ~new_n30053_ | ~new_n30101_ | ~new_n29975_;
  assign new_n30131_ = ~new_n30129_ | ~new_n30128_;
  assign new_n30132_ = ~new_n30063_;
  assign new_n30133_ = ~new_n8802_ | ~new_n30016_;
  assign new_n30134_ = ~new_n30133_ | ~new_n30063_;
  assign new_n30135_ = ~new_n8948_ | ~new_n30015_;
  assign new_n30136_ = ~new_n30062_;
  assign new_n30137_ = ~new_n8805_ | ~new_n30018_;
  assign new_n30138_ = ~new_n30137_ | ~new_n30062_;
  assign new_n30139_ = ~new_n8947_ | ~new_n30017_;
  assign new_n30140_ = ~new_n30061_;
  assign new_n30141_ = ~new_n8814_ | ~new_n30022_;
  assign new_n30142_ = ~new_n8944_ | ~new_n30019_;
  assign new_n30143_ = ~new_n8945_ | ~new_n30020_;
  assign new_n30144_ = ~new_n30071_ | ~new_n29977_;
  assign new_n30145_ = ~new_n29978_ | ~new_n30144_;
  assign new_n30146_ = ~new_n8808_ | ~new_n30024_;
  assign new_n30147_ = ~new_n8814_ | ~new_n30022_;
  assign new_n30148_ = ~new_n30061_ | ~new_n30146_ | ~new_n29977_;
  assign new_n30149_ = ~new_n30147_ | ~new_n30145_;
  assign new_n30150_ = ~new_n30060_;
  assign new_n30151_ = ~new_n8817_ | ~new_n30027_;
  assign new_n30152_ = ~new_n30151_ | ~new_n30060_;
  assign new_n30153_ = ~new_n8943_ | ~new_n30026_;
  assign new_n30154_ = ~new_n30028_;
  assign new_n30155_ = ~new_n30154_ | ~new_n30029_;
  assign new_n30156_ = ~new_n30155_ | ~new_n30059_;
  assign new_n30157_ = ~new_n8942_ | ~new_n30028_;
  assign new_n30158_ = ~new_n30058_;
  assign new_n30159_ = ~new_n30146_ | ~new_n30061_;
  assign new_n30160_ = ~new_n30030_;
  assign new_n30161_ = ~new_n8945_ | ~new_n30020_;
  assign new_n30162_ = ~new_n30160_ | ~new_n30161_;
  assign new_n30163_ = ~new_n30162_ | ~new_n30236_ | ~new_n30067_;
  assign new_n30164_ = ~new_n30030_ | ~new_n30067_;
  assign new_n30165_ = ~new_n8814_ | ~new_n30022_;
  assign new_n30166_ = ~new_n30164_ | ~new_n30165_ | ~new_n29978_;
  assign new_n30167_ = ~new_n8945_ | ~new_n30020_;
  assign new_n30168_ = ~new_n30067_ | ~new_n30167_;
  assign new_n30169_ = ~new_n30146_ | ~new_n30025_;
  assign new_n30170_ = ~new_n30101_ | ~new_n30053_;
  assign new_n30171_ = ~new_n30031_;
  assign new_n30172_ = ~new_n8950_ | ~new_n30011_;
  assign new_n30173_ = ~new_n30171_ | ~new_n30172_;
  assign new_n30174_ = ~new_n30173_ | ~new_n30257_ | ~new_n30066_;
  assign new_n30175_ = ~new_n30031_ | ~new_n30066_;
  assign new_n30176_ = ~new_n8799_ | ~new_n30012_;
  assign new_n30177_ = ~new_n30175_ | ~new_n30176_ | ~new_n29976_;
  assign new_n30178_ = ~new_n8950_ | ~new_n30011_;
  assign new_n30179_ = ~new_n30066_ | ~new_n30178_;
  assign new_n30180_ = ~new_n8952_ | ~new_n29987_;
  assign new_n30181_ = ~new_n8793_ | ~new_n30006_;
  assign new_n30182_ = ~new_n8933_ | ~new_n30005_;
  assign new_n30183_ = ~new_n30102_ | ~new_n30053_;
  assign new_n30184_ = ~new_n30100_ | ~new_n30182_ | ~new_n30181_;
  assign new_n30185_ = ~new_n8790_ | ~new_n30004_;
  assign new_n30186_ = ~new_n8934_ | ~new_n30001_;
  assign new_n30187_ = ~new_n8790_ | ~new_n30004_;
  assign new_n30188_ = ~new_n8934_ | ~new_n30001_;
  assign new_n30189_ = ~new_n30188_ | ~new_n30187_;
  assign new_n30190_ = ~new_n8787_ | ~new_n30002_;
  assign new_n30191_ = ~new_n8935_ | ~new_n29985_;
  assign new_n30192_ = ~new_n30107_ | ~new_n30007_;
  assign new_n30193_ = ~new_n30094_ | ~new_n30191_ | ~new_n30190_;
  assign new_n30194_ = ~new_n8784_ | ~new_n29997_;
  assign new_n30195_ = ~new_n8936_ | ~new_n29994_;
  assign new_n30196_ = ~new_n30195_ | ~new_n30194_;
  assign new_n30197_ = ~new_n8781_ | ~new_n29998_;
  assign new_n30198_ = ~new_n8937_ | ~new_n29995_;
  assign new_n30199_ = ~new_n30117_ | ~new_n30008_;
  assign new_n30200_ = ~new_n30109_ | ~new_n30198_ | ~new_n30197_;
  assign new_n30201_ = ~new_n8778_ | ~new_n29999_;
  assign new_n30202_ = ~new_n8938_ | ~new_n29996_;
  assign new_n30203_ = ~new_n30118_ | ~new_n30054_;
  assign new_n30204_ = ~new_n30084_ | ~new_n30202_ | ~new_n30201_;
  assign new_n30205_ = ~new_n8775_ | ~new_n29993_;
  assign new_n30206_ = ~new_n8939_ | ~new_n29990_;
  assign new_n30207_ = ~new_n8775_ | ~new_n29993_;
  assign new_n30208_ = ~new_n8939_ | ~new_n29990_;
  assign new_n30209_ = ~new_n30208_ | ~new_n30207_;
  assign new_n30210_ = ~new_n8772_ | ~new_n29991_;
  assign new_n30211_ = ~new_n8940_ | ~new_n29986_;
  assign new_n30212_ = ~new_n30123_ | ~new_n30009_;
  assign new_n30213_ = ~new_n30078_ | ~new_n30211_ | ~new_n30210_;
  assign new_n30214_ = ~new_n8769_ | ~new_n29989_;
  assign new_n30215_ = ~new_n8951_ | ~new_n30055_;
  assign new_n30216_ = ~new_n30047_;
  assign new_n30217_ = ~new_n30216_ | ~new_n30074_;
  assign new_n30218_ = ~new_n30047_ | ~new_n29988_;
  assign new_n30219_ = ~new_n8757_ | ~new_n30057_;
  assign new_n30220_ = ~new_n8941_ | ~new_n30056_;
  assign new_n30221_ = ~new_n30048_;
  assign new_n30222_ = ~new_n30158_ | ~new_n30221_;
  assign new_n30223_ = ~new_n30048_ | ~new_n30058_;
  assign new_n30224_ = ~new_n8820_ | ~new_n30029_;
  assign new_n30225_ = ~new_n8942_ | ~new_n30059_;
  assign new_n30226_ = ~new_n30049_;
  assign new_n30227_ = ~new_n30226_ | ~new_n30154_;
  assign new_n30228_ = ~new_n30049_ | ~new_n30028_;
  assign new_n30229_ = ~new_n8817_ | ~new_n30027_;
  assign new_n30230_ = ~new_n8943_ | ~new_n30026_;
  assign new_n30231_ = ~new_n30050_;
  assign new_n30232_ = ~new_n30150_ | ~new_n30231_;
  assign new_n30233_ = ~new_n30050_ | ~new_n30060_;
  assign new_n30234_ = ~new_n8814_ | ~new_n30022_;
  assign new_n30235_ = ~new_n8944_ | ~new_n30019_;
  assign new_n30236_ = ~new_n30235_ | ~new_n30234_;
  assign new_n30237_ = ~new_n8811_ | ~new_n30023_;
  assign new_n30238_ = ~new_n8945_ | ~new_n30020_;
  assign new_n30239_ = ~new_n30168_ | ~new_n30030_;
  assign new_n30240_ = ~new_n30160_ | ~new_n30238_ | ~new_n30237_;
  assign new_n30241_ = ~new_n8808_ | ~new_n30024_;
  assign new_n30242_ = ~new_n8946_ | ~new_n30021_;
  assign new_n30243_ = ~new_n30169_ | ~new_n30061_;
  assign new_n30244_ = ~new_n30140_ | ~new_n30242_ | ~new_n30241_;
  assign new_n30245_ = ~new_n8805_ | ~new_n30018_;
  assign new_n30246_ = ~new_n8947_ | ~new_n30017_;
  assign new_n30247_ = ~new_n30051_;
  assign new_n30248_ = ~new_n30136_ | ~new_n30247_;
  assign new_n30249_ = ~new_n30051_ | ~new_n30062_;
  assign new_n30250_ = ~new_n8802_ | ~new_n30016_;
  assign new_n30251_ = ~new_n8948_ | ~new_n30015_;
  assign new_n30252_ = ~new_n30052_;
  assign new_n30253_ = ~new_n30132_ | ~new_n30252_;
  assign new_n30254_ = ~new_n30052_ | ~new_n30063_;
  assign new_n30255_ = ~new_n8799_ | ~new_n30012_;
  assign new_n30256_ = ~new_n8949_ | ~new_n30010_;
  assign new_n30257_ = ~new_n30256_ | ~new_n30255_;
  assign new_n30258_ = ~new_n8796_ | ~new_n30013_;
  assign new_n30259_ = ~new_n8950_ | ~new_n30011_;
  assign new_n30260_ = ~new_n30179_ | ~new_n30031_;
  assign new_n30261_ = ~new_n30171_ | ~new_n30259_ | ~new_n30258_;
  assign new_n30262_ = new_n30437_ & new_n30436_;
  assign new_n30263_ = new_n30455_ & new_n30454_;
  assign new_n30264_ = new_n30495_ & new_n30494_;
  assign new_n30265_ = new_n30504_ & new_n30503_;
  assign new_n30266_ = new_n30522_ & new_n30521_;
  assign new_n30267_ = new_n30530_ & new_n30529_;
  assign new_n30268_ = new_n30609_ & new_n30606_;
  assign new_n30269_ = new_n30602_ & new_n30599_;
  assign new_n30270_ = new_n30593_ & new_n30590_;
  assign new_n30271_ = new_n30584_ & new_n30581_;
  assign new_n30272_ = new_n30578_ & new_n30576_;
  assign new_n30273_ = new_n30571_ & new_n30568_;
  assign new_n30274_ = new_n30493_ & new_n30490_;
  assign new_n30275_ = new_n30485_ & new_n30482_;
  assign new_n30276_ = new_n30471_ & new_n30468_;
  assign new_n30277_ = ~new_n8785_;
  assign new_n30278_ = ~new_n8448_;
  assign new_n30279_ = ~new_n8447_;
  assign new_n30280_ = ~new_n8448_ | ~new_n8785_;
  assign new_n30281_ = ~new_n8788_;
  assign new_n30282_ = ~new_n8779_;
  assign new_n30283_ = ~new_n8437_;
  assign new_n30284_ = ~new_n8444_;
  assign new_n30285_ = ~new_n8773_;
  assign new_n30286_ = ~new_n8445_;
  assign new_n30287_ = ~new_n8765_;
  assign new_n30288_ = ~new_n8454_;
  assign new_n30289_ = ~new_n8454_ | ~new_n8765_;
  assign new_n30290_ = ~new_n8776_;
  assign new_n30291_ = ~new_n8441_;
  assign new_n30292_ = ~new_n8437_ | ~new_n8779_;
  assign new_n30293_ = ~new_n8782_;
  assign new_n30294_ = ~new_n8791_;
  assign new_n30295_ = ~new_n8461_;
  assign new_n30296_ = ~new_n8460_;
  assign new_n30297_ = ~new_n8794_;
  assign new_n30298_ = ~new_n30321_ | ~new_n30463_;
  assign new_n30299_ = ~new_n30375_ | ~new_n30451_;
  assign new_n30300_ = ~new_n30440_ | ~new_n30441_;
  assign new_n30301_ = ~new_n8770_ | ~new_n8455_;
  assign new_n30302_ = ~new_n30380_ | ~new_n30477_;
  assign new_n30303_ = ~new_n30474_ | ~new_n30473_;
  assign new_n30304_ = ~new_n9278_;
  assign new_n30305_ = ~new_n8430_;
  assign new_n30306_ = ~new_n8434_;
  assign new_n30307_ = ~new_n9279_;
  assign new_n30308_ = ~new_n9280_;
  assign new_n30309_ = ~new_n8435_;
  assign new_n30310_ = ~new_n9281_;
  assign new_n30311_ = ~new_n8442_;
  assign new_n30312_ = ~new_n9284_;
  assign new_n30313_ = ~new_n8452_;
  assign new_n30314_ = ~new_n8815_;
  assign new_n30315_ = ~new_n8450_;
  assign new_n30316_ = ~new_n8446_;
  assign new_n30317_ = ~new_n8450_ | ~new_n8815_;
  assign new_n30318_ = ~new_n8818_;
  assign new_n30319_ = ~new_n8797_;
  assign new_n30320_ = ~new_n8439_;
  assign new_n30321_ = ~new_n8461_ | ~new_n8791_;
  assign new_n30322_ = ~new_n8803_;
  assign new_n30323_ = ~new_n8449_;
  assign new_n30324_ = ~new_n8800_;
  assign new_n30325_ = ~new_n8440_;
  assign new_n30326_ = ~new_n8440_ | ~new_n8800_;
  assign new_n30327_ = ~new_n8806_;
  assign new_n30328_ = ~new_n8457_;
  assign new_n30329_ = ~new_n8809_;
  assign new_n30330_ = ~new_n8456_;
  assign new_n30331_ = ~new_n8812_;
  assign new_n30332_ = ~new_n8451_;
  assign new_n30333_ = ~new_n8821_;
  assign new_n30334_ = ~new_n8459_;
  assign new_n30335_ = ~new_n8459_ | ~new_n8821_;
  assign new_n30336_ = ~new_n8823_;
  assign new_n30337_ = ~new_n8458_;
  assign new_n30338_ = ~new_n8458_ | ~new_n8823_;
  assign new_n30339_ = ~new_n9285_;
  assign new_n30340_ = ~new_n9283_;
  assign new_n30341_ = ~new_n8438_;
  assign new_n30342_ = ~new_n9282_;
  assign new_n30343_ = ~new_n8443_;
  assign new_n30344_ = ~new_n9279_ | ~new_n8434_;
  assign new_n30345_ = ~new_n8431_;
  assign new_n30346_ = ~new_n9277_;
  assign new_n30347_ = ~new_n30564_ | ~new_n30434_;
  assign new_n30348_ = ~new_n8453_;
  assign new_n30349_ = ~new_n30335_ | ~new_n30573_;
  assign new_n30350_ = ~new_n30519_ | ~new_n30518_;
  assign new_n30351_ = ~new_n30326_ | ~new_n30595_;
  assign new_n30352_ = ~new_n8382_ | ~new_n8383_;
  assign new_n30353_ = ~new_n1526_ | ~new_n1527_;
  assign new_n30354_ = ~new_n30633_ | ~new_n30632_;
  assign new_n30355_ = ~new_n30638_ | ~new_n30637_;
  assign new_n30356_ = ~new_n30645_ | ~new_n30644_;
  assign new_n30357_ = ~new_n30652_ | ~new_n30651_;
  assign new_n30358_ = ~new_n30657_ | ~new_n30656_;
  assign new_n30359_ = ~new_n30666_ | ~new_n30665_;
  assign new_n30360_ = ~new_n30673_ | ~new_n30672_;
  assign new_n30361_ = ~new_n30680_ | ~new_n30679_;
  assign new_n30362_ = ~new_n30687_ | ~new_n30686_;
  assign new_n30363_ = ~new_n11441_ | ~new_n11442_;
  assign new_n30364_ = ~new_n11434_ | ~new_n11435_;
  assign new_n30365_ = ~new_n11427_ | ~new_n11428_;
  assign new_n30366_ = ~new_n8377_ | ~new_n8378_;
  assign new_n30367_ = ~new_n8372_ | ~new_n8373_;
  assign new_n30368_ = ~new_n5228_ | ~new_n5229_;
  assign new_n30369_ = ~new_n5221_ | ~new_n5222_;
  assign new_n30370_ = ~new_n5214_ | ~new_n5215_;
  assign new_n30371_ = ~new_n1935_ | ~new_n1936_;
  assign new_n30372_ = ~new_n1930_ | ~new_n1931_;
  assign new_n30373_ = new_n30447_ & new_n30445_;
  assign new_n30374_ = new_n30262_ & new_n30438_;
  assign new_n30375_ = new_n30452_ & new_n30450_;
  assign new_n30376_ = new_n30459_ & new_n30458_;
  assign new_n30377_ = new_n30280_ & new_n30640_ & new_n30639_;
  assign new_n30378_ = new_n30470_ & new_n30263_;
  assign new_n30379_ = new_n30439_ & new_n30438_;
  assign new_n30380_ = new_n30478_ & new_n30476_;
  assign new_n30381_ = new_n30292_ & new_n30647_ & new_n30646_;
  assign new_n30382_ = new_n30484_ & new_n30262_;
  assign new_n30383_ = new_n30492_ & new_n30439_;
  assign new_n30384_ = new_n30462_ & new_n30264_;
  assign new_n30385_ = new_n30501_ & new_n30497_;
  assign new_n30386_ = new_n30508_ & new_n30265_;
  assign new_n30387_ = new_n30506_ & new_n30430_;
  assign new_n30388_ = new_n30526_ & new_n30525_;
  assign new_n30389_ = new_n30531_ & new_n30267_ & new_n30540_;
  assign new_n30390_ = new_n30543_ & new_n30538_;
  assign new_n30391_ = new_n30559_ & new_n30556_;
  assign new_n30392_ = new_n30626_ & new_n30560_;
  assign new_n30393_ = new_n30418_ & new_n30536_;
  assign new_n30394_ = new_n30338_ & new_n8384_ & new_n8385_;
  assign new_n30395_ = new_n30583_ & new_n30267_;
  assign new_n30396_ = new_n30317_ & new_n5233_ & new_n8371_;
  assign new_n30397_ = new_n30592_ & new_n30266_;
  assign new_n30398_ = new_n30430_ & new_n1940_ & new_n5213_;
  assign new_n30399_ = new_n30601_ & new_n30265_;
  assign new_n30400_ = new_n30429_ & new_n1528_ & new_n1929_;
  assign new_n30401_ = new_n30608_ & new_n30264_;
  assign new_n30402_ = ~new_n30376_ | ~new_n30460_;
  assign new_n30403_ = ~new_n30475_ | ~new_n30487_;
  assign new_n30404_ = ~new_n8432_;
  assign new_n30405_ = ~new_n9286_;
  assign new_n30406_ = new_n30661_ & new_n30660_;
  assign new_n30407_ = ~new_n30622_ | ~new_n30562_ | ~new_n30427_;
  assign new_n30408_ = new_n30668_ & new_n30667_;
  assign new_n30409_ = ~new_n30392_ | ~new_n30628_ | ~new_n30627_;
  assign new_n30410_ = new_n30675_ & new_n30674_;
  assign new_n30411_ = ~new_n30344_ | ~new_n30623_ | ~new_n30557_;
  assign new_n30412_ = new_n30682_ & new_n30681_;
  assign new_n30413_ = ~new_n30551_ | ~new_n30550_;
  assign new_n30414_ = new_n11439_ & new_n11440_;
  assign new_n30415_ = ~new_n30547_ | ~new_n30546_;
  assign new_n30416_ = new_n11432_ & new_n11433_;
  assign new_n30417_ = ~new_n30390_ | ~new_n30542_;
  assign new_n30418_ = new_n8389_ & new_n8390_;
  assign new_n30419_ = ~new_n30301_ | ~new_n30585_;
  assign new_n30420_ = ~new_n30388_ | ~new_n30527_;
  assign new_n30421_ = new_n5226_ & new_n5227_;
  assign new_n30422_ = ~new_n30515_ | ~new_n30514_;
  assign new_n30423_ = new_n5219_ & new_n5220_;
  assign new_n30424_ = ~new_n30511_ | ~new_n30510_;
  assign new_n30425_ = ~new_n30385_ | ~new_n30500_;
  assign new_n30426_ = ~new_n30625_ | ~new_n30624_;
  assign new_n30427_ = ~new_n8431_ | ~new_n30409_;
  assign new_n30428_ = ~new_n30292_;
  assign new_n30429_ = ~new_n8794_ | ~new_n8460_;
  assign new_n30430_ = ~new_n8449_ | ~new_n8803_;
  assign new_n30431_ = ~new_n8435_ | ~new_n9280_;
  assign new_n30432_ = ~new_n30326_;
  assign new_n30433_ = ~new_n30335_;
  assign new_n30434_ = ~new_n8442_ | ~new_n9281_;
  assign new_n30435_ = ~new_n30321_;
  assign new_n30436_ = new_n8444_ | new_n8782_;
  assign new_n30437_ = new_n8437_ | new_n8779_;
  assign new_n30438_ = new_n8776_ | new_n8441_;
  assign new_n30439_ = new_n8773_ | new_n8445_;
  assign new_n30440_ = ~new_n30289_;
  assign new_n30441_ = new_n8770_ | new_n8455_;
  assign new_n30442_ = ~new_n30300_;
  assign new_n30443_ = ~new_n30301_;
  assign new_n30444_ = ~new_n30300_ | ~new_n30301_;
  assign new_n30445_ = ~new_n8445_ | ~new_n8773_;
  assign new_n30446_ = ~new_n30444_ | ~new_n30439_;
  assign new_n30447_ = ~new_n8441_ | ~new_n8776_;
  assign new_n30448_ = ~new_n30373_ | ~new_n30446_;
  assign new_n30449_ = ~new_n30293_ | ~new_n30292_;
  assign new_n30450_ = ~new_n8444_ | ~new_n30449_;
  assign new_n30451_ = ~new_n30374_ | ~new_n30448_;
  assign new_n30452_ = ~new_n8782_ | ~new_n30428_;
  assign new_n30453_ = ~new_n30299_;
  assign new_n30454_ = new_n8447_ | new_n8788_;
  assign new_n30455_ = new_n8448_ | new_n8785_;
  assign new_n30456_ = ~new_n30280_;
  assign new_n30457_ = ~new_n30281_ | ~new_n30280_;
  assign new_n30458_ = ~new_n8447_ | ~new_n30457_;
  assign new_n30459_ = ~new_n8788_ | ~new_n30456_;
  assign new_n30460_ = ~new_n30263_ | ~new_n30299_;
  assign new_n30461_ = ~new_n30402_;
  assign new_n30462_ = new_n8791_ | new_n8461_;
  assign new_n30463_ = ~new_n30462_ | ~new_n30402_;
  assign new_n30464_ = ~new_n30298_;
  assign new_n30465_ = new_n8460_ | new_n8794_;
  assign new_n30466_ = new_n8785_ | new_n8448_;
  assign new_n30467_ = ~new_n30466_ | ~new_n30299_;
  assign new_n30468_ = ~new_n30377_ | ~new_n30467_;
  assign new_n30469_ = ~new_n30453_ | ~new_n30280_;
  assign new_n30470_ = ~new_n8788_ | ~new_n8447_;
  assign new_n30471_ = ~new_n30378_ | ~new_n30469_;
  assign new_n30472_ = new_n8448_ | new_n8785_;
  assign new_n30473_ = ~new_n30443_ | ~new_n30439_;
  assign new_n30474_ = ~new_n8445_ | ~new_n8773_;
  assign new_n30475_ = ~new_n30303_;
  assign new_n30476_ = ~new_n30379_ | ~new_n30442_;
  assign new_n30477_ = ~new_n30303_ | ~new_n30438_;
  assign new_n30478_ = ~new_n8441_ | ~new_n8776_;
  assign new_n30479_ = ~new_n30302_;
  assign new_n30480_ = new_n8779_ | new_n8437_;
  assign new_n30481_ = ~new_n30480_ | ~new_n30302_;
  assign new_n30482_ = ~new_n30381_ | ~new_n30481_;
  assign new_n30483_ = ~new_n30479_ | ~new_n30292_;
  assign new_n30484_ = ~new_n8782_ | ~new_n8444_;
  assign new_n30485_ = ~new_n30382_ | ~new_n30483_;
  assign new_n30486_ = new_n8437_ | new_n8779_;
  assign new_n30487_ = ~new_n30442_ | ~new_n30439_;
  assign new_n30488_ = ~new_n30403_;
  assign new_n30489_ = ~new_n8441_ | ~new_n8776_;
  assign new_n30490_ = ~new_n30658_ | ~new_n30300_ | ~new_n30301_ | ~new_n30659_;
  assign new_n30491_ = ~new_n30301_ | ~new_n30300_;
  assign new_n30492_ = ~new_n8445_ | ~new_n8773_;
  assign new_n30493_ = ~new_n30383_ | ~new_n30491_;
  assign new_n30494_ = new_n8460_ | new_n8794_;
  assign new_n30495_ = new_n8439_ | new_n8797_;
  assign new_n30496_ = ~new_n30435_ | ~new_n30264_;
  assign new_n30497_ = ~new_n8439_ | ~new_n8797_;
  assign new_n30498_ = ~new_n30429_ | ~new_n30496_;
  assign new_n30499_ = new_n8797_ | new_n8439_;
  assign new_n30500_ = ~new_n30384_ | ~new_n30402_;
  assign new_n30501_ = ~new_n30499_ | ~new_n30498_;
  assign new_n30502_ = ~new_n30425_;
  assign new_n30503_ = new_n8457_ | new_n8806_;
  assign new_n30504_ = new_n8449_ | new_n8803_;
  assign new_n30505_ = ~new_n30432_ | ~new_n30265_;
  assign new_n30506_ = ~new_n8457_ | ~new_n8806_;
  assign new_n30507_ = ~new_n30387_ | ~new_n30505_;
  assign new_n30508_ = new_n8800_ | new_n8440_;
  assign new_n30509_ = new_n8806_ | new_n8457_;
  assign new_n30510_ = ~new_n30386_ | ~new_n30425_;
  assign new_n30511_ = ~new_n30509_ | ~new_n30507_;
  assign new_n30512_ = ~new_n30424_;
  assign new_n30513_ = new_n8809_ | new_n8456_;
  assign new_n30514_ = ~new_n30513_ | ~new_n30424_;
  assign new_n30515_ = ~new_n8456_ | ~new_n8809_;
  assign new_n30516_ = ~new_n30422_;
  assign new_n30517_ = new_n8812_ | new_n8451_;
  assign new_n30518_ = ~new_n30517_ | ~new_n30422_;
  assign new_n30519_ = ~new_n8451_ | ~new_n8812_;
  assign new_n30520_ = ~new_n30350_;
  assign new_n30521_ = new_n8446_ | new_n8818_;
  assign new_n30522_ = new_n8450_ | new_n8815_;
  assign new_n30523_ = ~new_n30317_;
  assign new_n30524_ = ~new_n30318_ | ~new_n30317_;
  assign new_n30525_ = ~new_n8446_ | ~new_n30524_;
  assign new_n30526_ = ~new_n8818_ | ~new_n30523_;
  assign new_n30527_ = ~new_n30266_ | ~new_n30350_;
  assign new_n30528_ = ~new_n30420_;
  assign new_n30529_ = new_n8453_ | new_n9285_;
  assign new_n30530_ = new_n8458_ | new_n8823_;
  assign new_n30531_ = new_n8452_ | new_n9284_;
  assign new_n30532_ = ~new_n30338_;
  assign new_n30533_ = ~new_n9285_ | ~new_n30532_;
  assign new_n30534_ = ~new_n30533_ | ~new_n30348_;
  assign new_n30535_ = ~new_n30338_ | ~new_n30339_;
  assign new_n30536_ = ~new_n30535_ | ~new_n30534_;
  assign new_n30537_ = ~new_n30433_ | ~new_n30267_;
  assign new_n30538_ = ~new_n8452_ | ~new_n9284_;
  assign new_n30539_ = ~new_n30536_ | ~new_n30537_;
  assign new_n30540_ = new_n8821_ | new_n8459_;
  assign new_n30541_ = new_n9284_ | new_n8452_;
  assign new_n30542_ = ~new_n30420_ | ~new_n30389_;
  assign new_n30543_ = ~new_n30541_ | ~new_n30539_;
  assign new_n30544_ = ~new_n30417_;
  assign new_n30545_ = new_n9283_ | new_n8438_;
  assign new_n30546_ = ~new_n30545_ | ~new_n30417_;
  assign new_n30547_ = ~new_n8438_ | ~new_n9283_;
  assign new_n30548_ = ~new_n30415_;
  assign new_n30549_ = new_n9282_ | new_n8443_;
  assign new_n30550_ = ~new_n30549_ | ~new_n30415_;
  assign new_n30551_ = ~new_n8443_ | ~new_n9282_;
  assign new_n30552_ = ~new_n30413_;
  assign new_n30553_ = new_n8435_ | new_n9280_;
  assign new_n30554_ = ~new_n30434_ | ~new_n30431_;
  assign new_n30555_ = ~new_n30344_;
  assign new_n30556_ = new_n9281_ | new_n8442_;
  assign new_n30557_ = ~new_n30426_ | ~new_n30413_ | ~new_n30556_;
  assign new_n30558_ = ~new_n30411_;
  assign new_n30559_ = new_n9278_ | new_n8430_;
  assign new_n30560_ = ~new_n8430_ | ~new_n9278_;
  assign new_n30561_ = ~new_n30409_;
  assign new_n30562_ = ~new_n9277_ | ~new_n30409_;
  assign new_n30563_ = ~new_n30407_;
  assign new_n30564_ = ~new_n30556_ | ~new_n30413_;
  assign new_n30565_ = ~new_n30347_;
  assign new_n30566_ = new_n9280_ | new_n8435_;
  assign new_n30567_ = ~new_n30566_ | ~new_n30347_;
  assign new_n30568_ = ~new_n30412_ | ~new_n30567_ | ~new_n30431_;
  assign new_n30569_ = ~new_n30565_ | ~new_n30431_;
  assign new_n30570_ = ~new_n9279_ | ~new_n8434_;
  assign new_n30571_ = ~new_n30426_ | ~new_n30569_ | ~new_n30570_;
  assign new_n30572_ = new_n8435_ | new_n9280_;
  assign new_n30573_ = ~new_n30540_ | ~new_n30420_;
  assign new_n30574_ = ~new_n30349_;
  assign new_n30575_ = ~new_n30267_ | ~new_n30349_;
  assign new_n30576_ = ~new_n30393_ | ~new_n30575_;
  assign new_n30577_ = ~new_n30575_ | ~new_n30536_;
  assign new_n30578_ = ~new_n8386_ | ~new_n30577_;
  assign new_n30579_ = new_n8823_ | new_n8458_;
  assign new_n30580_ = ~new_n30579_ | ~new_n30349_;
  assign new_n30581_ = ~new_n30394_ | ~new_n30580_;
  assign new_n30582_ = ~new_n30574_ | ~new_n30338_;
  assign new_n30583_ = ~new_n8453_ | ~new_n9285_;
  assign new_n30584_ = ~new_n30395_ | ~new_n30582_;
  assign new_n30585_ = new_n8770_ | new_n8455_;
  assign new_n30586_ = ~new_n30419_;
  assign new_n30587_ = new_n8458_ | new_n8823_;
  assign new_n30588_ = new_n8815_ | new_n8450_;
  assign new_n30589_ = ~new_n30588_ | ~new_n30350_;
  assign new_n30590_ = ~new_n30396_ | ~new_n30589_;
  assign new_n30591_ = ~new_n30520_ | ~new_n30317_;
  assign new_n30592_ = ~new_n8818_ | ~new_n8446_;
  assign new_n30593_ = ~new_n30397_ | ~new_n30591_;
  assign new_n30594_ = new_n8450_ | new_n8815_;
  assign new_n30595_ = ~new_n30508_ | ~new_n30425_;
  assign new_n30596_ = ~new_n30351_;
  assign new_n30597_ = new_n8803_ | new_n8449_;
  assign new_n30598_ = ~new_n30597_ | ~new_n30351_;
  assign new_n30599_ = ~new_n30398_ | ~new_n30598_;
  assign new_n30600_ = ~new_n30596_ | ~new_n30430_;
  assign new_n30601_ = ~new_n8457_ | ~new_n8806_;
  assign new_n30602_ = ~new_n30399_ | ~new_n30600_;
  assign new_n30603_ = new_n8449_ | new_n8803_;
  assign new_n30604_ = new_n8794_ | new_n8460_;
  assign new_n30605_ = ~new_n30604_ | ~new_n30298_;
  assign new_n30606_ = ~new_n30400_ | ~new_n30605_;
  assign new_n30607_ = ~new_n30464_ | ~new_n30429_;
  assign new_n30608_ = ~new_n8439_ | ~new_n8797_;
  assign new_n30609_ = ~new_n30401_ | ~new_n30607_;
  assign new_n30610_ = ~new_n30465_ | ~new_n30429_;
  assign new_n30611_ = ~new_n30462_ | ~new_n30321_;
  assign new_n30612_ = ~new_n30472_ | ~new_n30280_;
  assign new_n30613_ = ~new_n30486_ | ~new_n30292_;
  assign new_n30614_ = ~new_n30489_ | ~new_n30438_;
  assign new_n30615_ = ~new_n30572_ | ~new_n30431_;
  assign new_n30616_ = ~new_n30556_ | ~new_n30434_;
  assign new_n30617_ = ~new_n30587_ | ~new_n30338_;
  assign new_n30618_ = ~new_n30540_ | ~new_n30335_;
  assign new_n30619_ = ~new_n30594_ | ~new_n30317_;
  assign new_n30620_ = ~new_n30603_ | ~new_n30430_;
  assign new_n30621_ = ~new_n30508_ | ~new_n30326_;
  assign new_n30622_ = ~new_n9277_ | ~new_n8431_;
  assign new_n30623_ = ~new_n30554_ | ~new_n30426_;
  assign new_n30624_ = ~new_n8434_ | ~new_n30553_;
  assign new_n30625_ = ~new_n9279_ | ~new_n30553_;
  assign new_n30626_ = ~new_n30559_ | ~new_n30554_ | ~new_n30426_;
  assign new_n30627_ = ~new_n30391_ | ~new_n30413_ | ~new_n30426_;
  assign new_n30628_ = ~new_n30555_ | ~new_n30559_;
  assign new_n30629_ = ~new_n8460_ | ~new_n30297_;
  assign new_n30630_ = ~new_n8794_ | ~new_n30296_;
  assign new_n30631_ = ~new_n30630_ | ~new_n30629_;
  assign new_n30632_ = ~new_n30610_ | ~new_n30298_;
  assign new_n30633_ = ~new_n30631_ | ~new_n30464_;
  assign new_n30634_ = ~new_n8461_ | ~new_n30294_;
  assign new_n30635_ = ~new_n8791_ | ~new_n30295_;
  assign new_n30636_ = ~new_n30635_ | ~new_n30634_;
  assign new_n30637_ = ~new_n30611_ | ~new_n30402_;
  assign new_n30638_ = ~new_n30461_ | ~new_n30636_;
  assign new_n30639_ = ~new_n8447_ | ~new_n30281_;
  assign new_n30640_ = ~new_n8788_ | ~new_n30279_;
  assign new_n30641_ = ~new_n8448_ | ~new_n30277_;
  assign new_n30642_ = ~new_n8785_ | ~new_n30278_;
  assign new_n30643_ = ~new_n30642_ | ~new_n30641_;
  assign new_n30644_ = ~new_n30612_ | ~new_n30299_;
  assign new_n30645_ = ~new_n30643_ | ~new_n30453_;
  assign new_n30646_ = ~new_n8444_ | ~new_n30293_;
  assign new_n30647_ = ~new_n8782_ | ~new_n30284_;
  assign new_n30648_ = ~new_n8437_ | ~new_n30282_;
  assign new_n30649_ = ~new_n8779_ | ~new_n30283_;
  assign new_n30650_ = ~new_n30649_ | ~new_n30648_;
  assign new_n30651_ = ~new_n30613_ | ~new_n30302_;
  assign new_n30652_ = ~new_n30650_ | ~new_n30479_;
  assign new_n30653_ = ~new_n8441_ | ~new_n30290_;
  assign new_n30654_ = ~new_n8776_ | ~new_n30291_;
  assign new_n30655_ = ~new_n30654_ | ~new_n30653_;
  assign new_n30656_ = ~new_n30614_ | ~new_n30403_;
  assign new_n30657_ = ~new_n30488_ | ~new_n30655_;
  assign new_n30658_ = ~new_n8445_ | ~new_n30285_;
  assign new_n30659_ = ~new_n8773_ | ~new_n30286_;
  assign new_n30660_ = ~new_n8432_ | ~new_n30405_;
  assign new_n30661_ = ~new_n9286_ | ~new_n30404_;
  assign new_n30662_ = ~new_n8432_ | ~new_n30405_;
  assign new_n30663_ = ~new_n9286_ | ~new_n30404_;
  assign new_n30664_ = ~new_n30663_ | ~new_n30662_;
  assign new_n30665_ = ~new_n30406_ | ~new_n30407_;
  assign new_n30666_ = ~new_n30563_ | ~new_n30664_;
  assign new_n30667_ = ~new_n8431_ | ~new_n30346_;
  assign new_n30668_ = ~new_n9277_ | ~new_n30345_;
  assign new_n30669_ = ~new_n8431_ | ~new_n30346_;
  assign new_n30670_ = ~new_n9277_ | ~new_n30345_;
  assign new_n30671_ = ~new_n30670_ | ~new_n30669_;
  assign new_n30672_ = ~new_n30408_ | ~new_n30409_;
  assign new_n30673_ = ~new_n30561_ | ~new_n30671_;
  assign new_n30674_ = ~new_n8430_ | ~new_n30304_;
  assign new_n30675_ = ~new_n9278_ | ~new_n30305_;
  assign new_n30676_ = ~new_n8430_ | ~new_n30304_;
  assign new_n30677_ = ~new_n9278_ | ~new_n30305_;
  assign new_n30678_ = ~new_n30677_ | ~new_n30676_;
  assign new_n30679_ = ~new_n30410_ | ~new_n30411_;
  assign new_n30680_ = ~new_n30558_ | ~new_n30678_;
  assign new_n30681_ = ~new_n8434_ | ~new_n30307_;
  assign new_n30682_ = ~new_n9279_ | ~new_n30306_;
  assign new_n30683_ = ~new_n8435_ | ~new_n30308_;
  assign new_n30684_ = ~new_n9280_ | ~new_n30309_;
  assign new_n30685_ = ~new_n30684_ | ~new_n30683_;
  assign new_n30686_ = ~new_n30615_ | ~new_n30347_;
  assign new_n30687_ = ~new_n30685_ | ~new_n30565_;
endmodule



// Benchmark "b15" written by ABC on Sun Apr 23 00:33:20 2023

module b15 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518;
  wire new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2106_,
    new_n2107_, new_n2111_, new_n2114_, new_n2115_, new_n2123_, new_n2124_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_,
    new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_,
    new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_,
    new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_,
    new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_,
    new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_,
    new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_,
    new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_,
    new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_,
    new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_,
    new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_,
    new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_,
    new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_,
    new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_,
    new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_,
    new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_,
    new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_,
    new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_,
    new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_,
    new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_,
    new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_,
    new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_,
    new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_,
    new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_,
    new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_,
    new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_,
    new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_,
    new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_,
    new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_,
    new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_,
    new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_,
    new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_,
    new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_,
    new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_,
    new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_,
    new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_,
    new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_,
    new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_,
    new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_,
    new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_,
    new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_,
    new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_,
    new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_,
    new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_,
    new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_,
    new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_,
    new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_,
    new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_,
    new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_,
    new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_,
    new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_,
    new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_,
    new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_,
    new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_,
    new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_,
    new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_,
    new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_,
    new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_,
    new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_,
    new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_,
    new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_,
    new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_,
    new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_,
    new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_,
    new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_,
    new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_,
    new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_,
    new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_,
    new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_,
    new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_,
    new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_,
    new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_,
    new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_,
    new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_,
    new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_,
    new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_,
    new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_,
    new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_,
    new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_,
    new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_,
    new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_,
    new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_,
    new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_,
    new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_,
    new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_,
    new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_,
    new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_,
    new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_,
    new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_,
    new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_,
    new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_,
    new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_,
    new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_,
    new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_,
    new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_,
    new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_,
    new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_,
    new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_,
    new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_,
    new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8065_,
    new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_,
    new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_,
    new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_,
    new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_,
    new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_,
    new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_,
    new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_,
    new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_,
    new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_,
    new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_,
    new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_,
    new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_,
    new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_,
    new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_,
    new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_,
    new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_,
    new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_,
    new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_,
    new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_,
    new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_,
    new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_,
    new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_,
    new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_,
    new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_,
    new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_,
    new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_,
    new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_,
    new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_,
    new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_,
    new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_,
    new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_,
    new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_,
    new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_,
    new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_,
    new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_,
    new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_,
    new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_,
    new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_,
    new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_,
    new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_,
    new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_,
    new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_,
    new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_,
    new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_,
    new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_,
    new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_,
    new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_,
    new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_,
    new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_,
    new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_,
    new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_,
    new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_,
    new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8569_,
    new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_,
    new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_,
    new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_,
    new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_,
    new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_,
    new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_,
    new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_,
    new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_,
    new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_,
    new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_,
    new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_,
    new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_,
    new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_,
    new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_,
    new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_;
  assign new_n1006_ = ~new_n9322_ | ~new_n9242_;
  assign new_n1007_ = ~pi258 | ~new_n9241_;
  assign new_n1008_ = ~new_n9323_ | ~new_n9244_;
  assign new_n1009_ = ~pi478 & ~pi107;
  assign new_n1010_ = new_n2876_ & pi107;
  assign new_n1011_ = new_n2910_ & new_n3122_;
  assign new_n1012_ = new_n1878_ & new_n1107_;
  assign new_n1013_ = new_n8877_ & new_n2837_;
  assign new_n1014_ = new_n8624_ & new_n4604_ & new_n2510_;
  assign new_n1015_ = new_n1045_ & new_n2869_;
  assign new_n1016_ = pi107 & new_n2075_;
  assign new_n1017_ = pi107 & new_n2058_;
  assign new_n1018_ = new_n2869_ & pi106;
  assign new_n1019_ = new_n1016_ & new_n2853_;
  assign new_n1020_ = new_n1016_ & new_n2855_;
  assign new_n1021_ = new_n2509_ & new_n2060_;
  assign new_n1022_ = new_n2906_ & new_n2060_;
  assign new_n1023_ = new_n2074_ & new_n2075_ & pi108;
  assign new_n1024_ = new_n7786_ & pi108 & new_n2075_;
  assign new_n1025_ = new_n2880_ & pi109;
  assign new_n1026_ = new_n1019_ & new_n3142_;
  assign new_n1027_ = new_n2058_ & new_n1907_;
  assign new_n1028_ = new_n2867_ & new_n3094_;
  assign new_n1029_ = pi109 & new_n2060_;
  assign new_n1030_ = pi106 & new_n2075_;
  assign new_n1031_ = new_n1017_ & new_n2859_;
  assign new_n1032_ = new_n1017_ & new_n2861_;
  assign new_n1033_ = new_n4443_ & new_n2060_;
  assign new_n1034_ = new_n2407_ & new_n2058_;
  assign new_n1035_ = new_n1017_ & new_n4214_;
  assign new_n1036_ = new_n1020_ & new_n1924_;
  assign new_n1037_ = new_n1017_ & new_n6253_;
  assign new_n1038_ = new_n1014_ & new_n1915_;
  assign new_n1039_ = new_n1014_ & new_n3122_;
  assign new_n1040_ = new_n2867_ & new_n2035_;
  assign new_n1041_ = pi109 & new_n2061_;
  assign new_n1042_ = new_n2061_ & new_n1938_;
  assign new_n1043_ = new_n2868_ & new_n2067_;
  assign new_n1044_ = new_n2529_ & new_n2868_;
  assign new_n1045_ = pi478 & new_n2854_;
  assign new_n1046_ = new_n1109_ & new_n6139_;
  assign new_n1047_ = pi032 & new_n2869_;
  assign new_n1048_ = pi031 & new_n2869_;
  assign new_n1049_ = pi030 & new_n2869_;
  assign new_n1050_ = pi029 & new_n2869_;
  assign new_n1051_ = pi028 & new_n2869_;
  assign new_n1052_ = pi027 & new_n2869_;
  assign new_n1053_ = pi026 & new_n2869_;
  assign new_n1054_ = pi025 & new_n2869_;
  assign new_n1055_ = pi008 & new_n1015_;
  assign new_n1056_ = pi016 & new_n1015_;
  assign new_n1057_ = pi007 & new_n1015_;
  assign new_n1058_ = pi015 & new_n1015_;
  assign new_n1059_ = pi006 & new_n1015_;
  assign new_n1060_ = pi014 & new_n1015_;
  assign new_n1061_ = pi005 & new_n1015_;
  assign new_n1062_ = pi013 & new_n1015_;
  assign new_n1063_ = pi004 & new_n1015_;
  assign new_n1064_ = pi012 & new_n1015_;
  assign new_n1065_ = pi003 & new_n1015_;
  assign new_n1066_ = pi011 & new_n1015_;
  assign new_n1067_ = pi002 & new_n1015_;
  assign new_n1068_ = pi010 & new_n1015_;
  assign new_n1069_ = pi001 & new_n1015_;
  assign new_n1070_ = pi009 & new_n1015_;
  assign new_n1071_ = new_n1018_ & new_n1915_;
  assign new_n1072_ = new_n1018_ & new_n2035_;
  assign new_n1073_ = new_n1018_ & new_n1921_;
  assign new_n1074_ = new_n1018_ & new_n1928_;
  assign new_n1075_ = new_n1018_ & new_n1927_;
  assign new_n1076_ = new_n1018_ & new_n1922_;
  assign new_n1077_ = new_n1018_ & new_n2818_;
  assign new_n1078_ = new_n1018_ & new_n2816_;
  assign new_n1079_ = new_n2868_ & new_n4106_;
  assign new_n1080_ = new_n2868_ & new_n2876_;
  assign new_n1081_ = new_n1041_ & new_n1928_;
  assign new_n1082_ = new_n1025_ & new_n1105_;
  assign new_n1083_ = new_n2534_ & new_n2075_;
  assign new_n1084_ = ~pi108 & ~pi106;
  assign new_n1085_ = pi107 & pi108;
  assign new_n1086_ = new_n5011_ & new_n2075_;
  assign new_n1087_ = pi108 & new_n2031_;
  assign new_n1088_ = new_n2844_ & new_n6139_;
  assign new_n1089_ = new_n2099_ & new_n2004_;
  assign new_n1090_ = new_n3185_ & new_n2099_;
  assign new_n1091_ = new_n6341_ & new_n2004_;
  assign new_n1092_ = new_n3185_ & new_n6341_;
  assign new_n1093_ = new_n1879_ & new_n1945_;
  assign new_n1094_ = new_n3188_ & new_n1945_;
  assign new_n1095_ = new_n7959_ & new_n7942_;
  assign new_n1096_ = new_n7959_ & new_n1960_;
  assign new_n1097_ = new_n7942_ & new_n1961_;
  assign new_n1098_ = ~new_n7959_ & ~new_n7942_;
  assign new_n1099_ = new_n7950_ & new_n7951_;
  assign new_n1100_ = new_n7950_ & new_n1962_;
  assign new_n1101_ = new_n7951_ & new_n1963_;
  assign new_n1102_ = ~new_n7950_ & ~new_n7951_;
  assign new_n1103_ = pi108 & new_n2115_;
  assign new_n1104_ = new_n2222_ & new_n1109_;
  assign new_n1105_ = new_n8624_ & new_n1928_;
  assign new_n1106_ = new_n3139_ & new_n1915_;
  assign new_n1107_ = pi109 & new_n3045_;
  assign new_n1108_ = new_n2896_ & pi109;
  assign new_n1109_ = new_n2818_ & new_n2035_ & new_n3045_ & new_n1921_;
  assign new_n1110_ = pi240 & pi241 & pi239 & pi242;
  assign new_n1111_ = pi241 & new_n1910_;
  assign new_n1112_ = new_n1910_ & pi240 & pi239 & pi241;
  assign new_n1113_ = pi242 & new_n1909_;
  assign new_n1114_ = new_n1909_ & pi240 & pi239 & pi242;
  assign new_n1115_ = new_n2152_ & new_n3023_;
  assign new_n1116_ = new_n1908_ & pi241 & pi239 & pi242;
  assign new_n1117_ = pi241 & new_n1908_ & new_n1910_;
  assign new_n1118_ = new_n2151_ & new_n2150_;
  assign new_n1119_ = pi242 & new_n1908_ & new_n1909_;
  assign new_n1120_ = new_n2149_ & new_n2148_;
  assign new_n1121_ = pi239 & new_n3025_;
  assign new_n1122_ = new_n2147_ & new_n2146_;
  assign new_n1123_ = new_n2145_ & new_n2144_;
  assign new_n1124_ = new_n3023_ & pi240 & new_n1914_;
  assign new_n1125_ = new_n2143_ & new_n2142_;
  assign new_n1126_ = ~pi239 & ~pi240;
  assign new_n1127_ = new_n1126_ & pi241 & new_n1910_;
  assign new_n1128_ = new_n1126_ & pi242 & new_n1909_;
  assign new_n1129_ = new_n3025_ & new_n1914_;
  assign new_n1130_ = new_n2050_ & new_n6325_ & new_n6324_;
  assign new_n1131_ = new_n8048_ & new_n1956_;
  assign new_n1132_ = new_n2098_ & new_n2002_;
  assign new_n1133_ = new_n8007_ & new_n8048_;
  assign new_n1134_ = new_n3173_ & new_n1133_;
  assign new_n1135_ = pi245 & pi244;
  assign new_n1136_ = pi245 & new_n1947_;
  assign new_n1137_ = new_n1959_ & new_n3193_;
  assign new_n1138_ = new_n3169_ & new_n1133_;
  assign new_n1139_ = new_n1971_ & new_n3251_;
  assign new_n1140_ = new_n3170_ & new_n1133_;
  assign new_n1141_ = new_n1978_ & new_n3310_;
  assign new_n1142_ = new_n3171_ & new_n8042_;
  assign new_n1143_ = ~new_n8042_ & ~new_n8049_;
  assign new_n1144_ = new_n1143_ & new_n1133_;
  assign new_n1145_ = ~pi247 & ~pi246;
  assign new_n1146_ = new_n1982_ & new_n3367_;
  assign new_n1147_ = new_n6338_ & new_n2002_;
  assign new_n1148_ = new_n3174_ & new_n3173_;
  assign new_n1149_ = new_n1987_ & new_n3425_;
  assign new_n1150_ = new_n3174_ & new_n3169_;
  assign new_n1151_ = new_n1991_ & new_n3482_;
  assign new_n1152_ = new_n3174_ & new_n3170_;
  assign new_n1153_ = new_n1994_ & new_n3540_;
  assign new_n1154_ = new_n3174_ & new_n1143_;
  assign new_n1155_ = new_n1998_ & new_n3597_;
  assign new_n1156_ = new_n3176_ & new_n2098_;
  assign new_n1157_ = new_n2003_ & new_n2001_;
  assign new_n1158_ = new_n3169_ & new_n1131_;
  assign new_n1159_ = new_n2008_ & new_n3710_;
  assign new_n1160_ = new_n3170_ & new_n1131_;
  assign new_n1161_ = new_n2011_ & new_n3768_;
  assign new_n1162_ = new_n1143_ & new_n1131_;
  assign new_n1163_ = new_n2015_ & new_n3825_;
  assign new_n1164_ = new_n3176_ & new_n6338_;
  assign new_n1165_ = ~new_n8048_ & ~new_n8007_;
  assign new_n1166_ = new_n1165_ & new_n3173_;
  assign new_n1167_ = ~pi244 & ~pi245;
  assign new_n1168_ = new_n2018_ & new_n3883_;
  assign new_n1169_ = new_n1165_ & new_n3169_;
  assign new_n1170_ = new_n2022_ & new_n3940_;
  assign new_n1171_ = new_n1165_ & new_n3170_;
  assign new_n1172_ = new_n2025_ & new_n3998_;
  assign new_n1173_ = new_n1165_ & new_n1143_;
  assign new_n1174_ = new_n2029_ & new_n4055_;
  assign new_n1175_ = new_n4113_ & new_n6345_ & new_n6344_;
  assign new_n1176_ = new_n2389_ & new_n4144_;
  assign new_n1177_ = new_n2864_ & new_n2090_;
  assign new_n1178_ = pi242 & new_n2046_;
  assign new_n1179_ = new_n4128_ & new_n4156_;
  assign new_n1180_ = new_n1179_ & new_n1178_;
  assign new_n1181_ = new_n1910_ & new_n2046_;
  assign new_n1182_ = new_n1179_ & new_n1181_;
  assign new_n1183_ = new_n4164_ & pi242;
  assign new_n1184_ = new_n1179_ & new_n1183_;
  assign new_n1185_ = new_n4164_ & new_n1910_;
  assign new_n1186_ = new_n1179_ & new_n1185_;
  assign new_n1187_ = new_n4128_ & new_n2045_;
  assign new_n1188_ = new_n1187_ & new_n1178_;
  assign new_n1189_ = new_n1187_ & new_n1181_;
  assign new_n1190_ = new_n1187_ & new_n1183_;
  assign new_n1191_ = new_n1187_ & new_n1185_;
  assign new_n1192_ = new_n4156_ & new_n2082_;
  assign new_n1193_ = new_n1192_ & new_n1178_;
  assign new_n1194_ = new_n1192_ & new_n1181_;
  assign new_n1195_ = new_n1192_ & new_n1183_;
  assign new_n1196_ = new_n1192_ & new_n1185_;
  assign new_n1197_ = new_n2082_ & new_n2045_;
  assign new_n1198_ = new_n1178_ & new_n1197_;
  assign new_n1199_ = new_n1181_ & new_n1197_;
  assign new_n1200_ = new_n1183_ & new_n1197_;
  assign new_n1201_ = new_n1185_ & new_n1197_;
  assign new_n1202_ = new_n4125_ & new_n6365_;
  assign new_n1203_ = new_n1202_ & new_n1111_;
  assign new_n1204_ = new_n1202_ & new_n2143_;
  assign new_n1205_ = new_n1202_ & new_n3023_;
  assign new_n1206_ = new_n1202_ & new_n1113_;
  assign new_n1207_ = new_n4125_ & new_n2100_;
  assign new_n1208_ = new_n1207_ & new_n1111_;
  assign new_n1209_ = new_n1207_ & new_n2143_;
  assign new_n1210_ = new_n1207_ & new_n3023_;
  assign new_n1211_ = new_n1207_ & new_n1113_;
  assign new_n1212_ = new_n6365_ & new_n2086_;
  assign new_n1213_ = new_n1212_ & new_n1111_;
  assign new_n1214_ = new_n1212_ & new_n2143_;
  assign new_n1215_ = new_n1212_ & new_n3023_;
  assign new_n1216_ = new_n1212_ & new_n1113_;
  assign new_n1217_ = new_n2100_ & new_n2086_;
  assign new_n1218_ = new_n1217_ & new_n1111_;
  assign new_n1219_ = new_n1217_ & new_n2143_;
  assign new_n1220_ = new_n1217_ & new_n3023_;
  assign new_n1221_ = new_n1217_ & new_n1113_;
  assign new_n1222_ = new_n5710_ & new_n3024_;
  assign new_n1223_ = new_n5710_ & new_n1117_;
  assign new_n1224_ = new_n5710_ & new_n1119_;
  assign new_n1225_ = new_n5710_ & new_n3025_;
  assign new_n1226_ = new_n5710_ & pi240;
  assign new_n1227_ = new_n1226_ & new_n2143_;
  assign new_n1228_ = new_n1226_ & new_n1111_;
  assign new_n1229_ = new_n1226_ & new_n1113_;
  assign new_n1230_ = new_n1226_ & new_n3023_;
  assign new_n1231_ = new_n3024_ & new_n2089_;
  assign new_n1232_ = new_n1117_ & new_n2089_;
  assign new_n1233_ = new_n1119_ & new_n2089_;
  assign new_n1234_ = new_n3025_ & new_n2089_;
  assign new_n1235_ = pi240 & new_n2089_;
  assign new_n1236_ = new_n1235_ & new_n2143_;
  assign new_n1237_ = new_n1235_ & new_n1111_;
  assign new_n1238_ = new_n1235_ & new_n1113_;
  assign new_n1239_ = new_n1235_ & new_n3023_;
  assign new_n1240_ = new_n6435_ & new_n2829_;
  assign new_n1241_ = new_n1240_ & new_n1181_;
  assign new_n1242_ = new_n1240_ & new_n1178_;
  assign new_n1243_ = new_n1240_ & new_n1185_;
  assign new_n1244_ = new_n1240_ & new_n1183_;
  assign new_n1245_ = new_n6435_ & new_n2096_;
  assign new_n1246_ = new_n1245_ & new_n1181_;
  assign new_n1247_ = new_n1245_ & new_n1178_;
  assign new_n1248_ = new_n1245_ & new_n1185_;
  assign new_n1249_ = new_n1245_ & new_n1183_;
  assign new_n1250_ = new_n2829_ & new_n2101_;
  assign new_n1251_ = new_n1250_ & new_n1181_;
  assign new_n1252_ = new_n1250_ & new_n1178_;
  assign new_n1253_ = new_n1250_ & new_n1185_;
  assign new_n1254_ = new_n1250_ & new_n1183_;
  assign new_n1255_ = new_n2101_ & new_n2096_;
  assign new_n1256_ = new_n1255_ & new_n1181_;
  assign new_n1257_ = new_n1255_ & new_n1178_;
  assign new_n1258_ = new_n1255_ & new_n1185_;
  assign new_n1259_ = new_n1255_ & new_n1183_;
  assign new_n1260_ = pi109 & new_n2033_;
  assign new_n1261_ = pi438 & new_n1036_;
  assign new_n1262_ = new_n2175_ & new_n2176_ & new_n2177_ & new_n2178_ & new_n1264_;
  assign new_n1263_ = new_n6149_ & new_n2071_;
  assign new_n1264_ = new_n6317_ & new_n6316_;
  assign new_n1265_ = new_n6432_ & new_n6431_;
  assign new_n1266_ = ~new_n5401_ | ~new_n2650_;
  assign new_n1267_ = ~new_n5398_ | ~new_n2649_;
  assign new_n1268_ = ~new_n5395_ | ~new_n2648_;
  assign new_n1269_ = ~new_n5392_ | ~new_n2647_;
  assign new_n1270_ = ~new_n5501_ | ~new_n2671_;
  assign new_n1271_ = ~new_n5500_ | ~new_n5498_ | ~new_n5499_;
  assign new_n1272_ = ~new_n5497_ | ~new_n5495_ | ~new_n5496_;
  assign new_n1273_ = ~new_n5494_ | ~new_n5492_ | ~new_n5493_;
  assign new_n1274_ = ~new_n5491_ | ~new_n5489_ | ~new_n5490_;
  assign new_n1275_ = ~new_n5488_ | ~new_n5486_ | ~new_n5487_;
  assign new_n1276_ = ~pi259 | ~new_n9243_;
  assign new_n1277_ = new_n8144_ & new_n5391_;
  assign new_n1278_ = new_n8144_ & new_n5391_;
  assign new_n1279_ = new_n8144_ & new_n5391_;
  assign new_n1280_ = new_n8144_ & new_n5391_;
  assign new_n1281_ = new_n8144_ & new_n5391_;
  assign new_n1282_ = new_n8144_ & new_n5391_;
  assign new_n1283_ = new_n8144_ & new_n5391_;
  assign new_n1284_ = new_n8144_ & new_n5391_;
  assign new_n1285_ = new_n8144_ & new_n5391_;
  assign new_n1286_ = new_n8144_ & new_n5391_;
  assign new_n1287_ = new_n8144_ & new_n5391_;
  assign new_n1288_ = new_n8144_ & new_n5391_;
  assign new_n1289_ = new_n8144_ & new_n5391_;
  assign new_n1290_ = new_n8144_ & new_n5391_;
  assign new_n1291_ = new_n8010_ & new_n5391_;
  assign new_n1292_ = new_n8036_ & new_n5391_;
  assign new_n1293_ = new_n8037_ & new_n5391_;
  assign new_n1294_ = new_n8038_ & new_n5391_;
  assign new_n1295_ = new_n8039_ & new_n5391_;
  assign new_n1296_ = new_n8040_ & new_n5391_;
  assign new_n1297_ = new_n8041_ & new_n5391_;
  assign new_n1298_ = new_n8029_ & new_n5391_;
  assign new_n1299_ = new_n8079_ & new_n5391_;
  assign new_n1300_ = new_n8009_ & new_n5391_;
  assign new_n1301_ = new_n8008_ & new_n5391_;
  assign new_n1302_ = new_n8044_ & new_n5391_;
  assign new_n1303_ = new_n8046_ & new_n5391_;
  assign new_n1304_ = new_n8007_ & new_n5391_;
  assign new_n1305_ = ~new_n2084_ | ~new_n5514_;
  assign new_n1306_ = new_n8049_ & new_n5391_;
  assign new_n1307_ = pi107 & new_n5515_;
  assign new_n1308_ = ~new_n5415_ | ~new_n5414_ | ~new_n5413_;
  assign new_n1309_ = ~new_n5416_ | ~new_n2654_;
  assign new_n1310_ = ~new_n5425_ | ~new_n2656_;
  assign new_n1311_ = ~new_n5429_ | ~new_n2657_;
  assign new_n1312_ = ~new_n5433_ | ~new_n2658_;
  assign new_n1313_ = ~new_n5437_ | ~new_n2659_;
  assign new_n1314_ = ~new_n5441_ | ~new_n2660_;
  assign new_n1315_ = ~new_n5445_ | ~new_n2661_;
  assign new_n1316_ = ~new_n5449_ | ~new_n2662_;
  assign new_n1317_ = ~new_n5453_ | ~new_n2663_;
  assign new_n1318_ = ~new_n5457_ | ~new_n2664_;
  assign new_n1319_ = ~new_n5461_ | ~new_n2665_;
  assign new_n1320_ = ~new_n5470_ | ~new_n2667_;
  assign new_n1321_ = ~new_n5474_ | ~new_n2668_;
  assign new_n1322_ = ~new_n5478_ | ~new_n2669_;
  assign new_n1323_ = ~new_n5482_ | ~new_n2670_;
  assign new_n1324_ = ~new_n5404_ | ~new_n2651_;
  assign new_n1325_ = ~new_n5408_ | ~new_n2653_ | ~new_n5412_ | ~new_n5411_;
  assign new_n1326_ = ~new_n5420_ | ~new_n2655_ | ~new_n5424_ | ~new_n5423_;
  assign new_n1327_ = ~new_n5465_ | ~new_n2666_ | ~new_n5469_ | ~new_n5468_;
  assign new_n1328_ = ~new_n5504_ | ~new_n2672_ | ~new_n5508_ | ~new_n5507_;
  assign new_n1329_ = ~new_n5512_ | ~new_n5513_ | ~new_n5510_ | ~new_n5511_ | ~new_n5509_;
  assign new_n1330_ = ~new_n6103_ | ~new_n6102_;
  assign new_n1331_ = ~new_n6105_ | ~new_n6104_;
  assign new_n1332_ = ~new_n2813_ | ~new_n6108_;
  assign new_n1333_ = ~new_n2814_ | ~new_n6111_;
  assign new_n1334_ = ~new_n6112_ | ~new_n6439_ | ~new_n6438_;
  assign new_n1335_ = ~new_n6101_ | ~new_n1928_;
  assign new_n1336_ = ~new_n6050_ | ~new_n6049_;
  assign new_n1337_ = ~new_n6052_ | ~new_n6051_;
  assign new_n1338_ = ~new_n6056_ | ~new_n6055_;
  assign new_n1339_ = ~new_n6058_ | ~new_n6057_;
  assign new_n1340_ = ~new_n6060_ | ~new_n6059_;
  assign new_n1341_ = ~new_n6062_ | ~new_n6061_;
  assign new_n1342_ = ~new_n6064_ | ~new_n6063_;
  assign new_n1343_ = ~new_n6066_ | ~new_n6065_;
  assign new_n1344_ = ~new_n6068_ | ~new_n6067_;
  assign new_n1345_ = ~new_n6070_ | ~new_n6069_;
  assign new_n1346_ = ~new_n6072_ | ~new_n6071_;
  assign new_n1347_ = ~new_n6074_ | ~new_n6073_;
  assign new_n1348_ = ~new_n6078_ | ~new_n6077_;
  assign new_n1349_ = ~new_n6080_ | ~new_n6079_;
  assign new_n1350_ = ~new_n6082_ | ~new_n6081_;
  assign new_n1351_ = ~new_n6084_ | ~new_n6083_;
  assign new_n1352_ = ~new_n6086_ | ~new_n6085_;
  assign new_n1353_ = ~new_n6088_ | ~new_n6087_;
  assign new_n1354_ = ~new_n6090_ | ~new_n6089_;
  assign new_n1355_ = ~new_n6092_ | ~new_n6091_;
  assign new_n1356_ = ~new_n6094_ | ~new_n6093_;
  assign new_n1357_ = ~new_n6096_ | ~new_n6095_;
  assign new_n1358_ = ~new_n6038_ | ~new_n6037_;
  assign new_n1359_ = ~new_n6040_ | ~new_n6039_;
  assign new_n1360_ = ~new_n6042_ | ~new_n6041_;
  assign new_n1361_ = ~new_n6044_ | ~new_n6043_;
  assign new_n1362_ = ~new_n6046_ | ~new_n6045_;
  assign new_n1363_ = ~new_n6048_ | ~new_n6047_;
  assign new_n1364_ = ~new_n6054_ | ~new_n6053_;
  assign new_n1365_ = ~new_n6076_ | ~new_n6075_;
  assign new_n1366_ = ~new_n6098_ | ~new_n6097_;
  assign new_n1367_ = ~new_n6100_ | ~new_n6099_;
  assign new_n1368_ = ~new_n6022_ | ~new_n6021_;
  assign new_n1369_ = ~new_n6024_ | ~new_n6023_;
  assign new_n1370_ = ~new_n2810_ | ~new_n2884_;
  assign new_n1371_ = ~new_n2078_ | ~new_n2811_ | ~new_n6031_ | ~new_n6030_;
  assign new_n1372_ = ~new_n2884_ | ~new_n2812_;
  assign new_n1373_ = ~new_n6010_ | ~new_n6009_;
  assign new_n1374_ = ~new_n6012_ | ~new_n6011_;
  assign new_n1375_ = ~new_n2806_ | ~new_n6013_;
  assign new_n1376_ = ~new_n2807_ | ~new_n6015_;
  assign new_n1377_ = ~new_n2808_ | ~new_n6017_;
  assign new_n1378_ = ~new_n2809_ | ~new_n6019_;
  assign new_n1379_ = ~new_n2804_ | ~new_n2837_;
  assign new_n1380_ = new_n5881_ & new_n5728_;
  assign new_n1381_ = new_n5898_ & new_n5728_;
  assign new_n1382_ = new_n5915_ & new_n5728_;
  assign new_n1383_ = new_n6265_ & new_n5728_;
  assign new_n1384_ = new_n5947_ & new_n5728_;
  assign new_n1385_ = new_n5964_ & new_n5728_;
  assign new_n1386_ = new_n5981_ & new_n5728_;
  assign new_n1387_ = new_n5998_ & new_n5728_;
  assign new_n1388_ = ~new_n1263_ | ~new_n5999_;
  assign new_n1389_ = new_n5728_ & new_n5727_;
  assign new_n1390_ = new_n5759_ & new_n5728_;
  assign new_n1391_ = new_n5776_ & new_n5728_;
  assign new_n1392_ = new_n6263_ & new_n5728_;
  assign new_n1393_ = new_n5808_ & new_n5728_;
  assign new_n1394_ = new_n5825_ & new_n5728_;
  assign new_n1395_ = new_n5842_ & new_n5728_;
  assign new_n1396_ = new_n5859_ & new_n5728_;
  assign new_n1397_ = pi238 & new_n5708_;
  assign new_n1398_ = ~new_n2723_ | ~new_n5741_;
  assign new_n1399_ = new_n6137_ & new_n6136_;
  assign new_n1400_ = new_n6151_ & new_n6115_;
  assign new_n1401_ = new_n6124_ & new_n6123_;
  assign new_n1402_ = ~new_n5693_ | ~new_n5692_;
  assign new_n1403_ = ~new_n5695_ | ~new_n5694_;
  assign new_n1404_ = ~new_n5697_ | ~new_n5696_;
  assign new_n1405_ = ~new_n6261_ | ~new_n5698_;
  assign new_n1406_ = ~new_n5700_ | ~new_n5699_;
  assign new_n1407_ = ~new_n5702_ | ~new_n5701_;
  assign new_n1408_ = ~new_n2706_ | ~new_n5703_;
  assign new_n1409_ = ~new_n5706_ | ~new_n2707_ | ~new_n5705_;
  assign new_n1410_ = new_n5602_ & new_n5554_;
  assign new_n1411_ = new_n5619_ & new_n5554_;
  assign new_n1412_ = new_n5636_ & new_n5554_;
  assign new_n1413_ = new_n6260_ & new_n5554_;
  assign new_n1414_ = new_n5668_ & new_n5554_;
  assign new_n1415_ = new_n5685_ & new_n5554_;
  assign new_n1416_ = new_n5554_ & new_n5553_;
  assign new_n1417_ = new_n5571_ & new_n5554_;
  assign new_n1418_ = ~new_n5573_ | ~new_n5572_;
  assign new_n1419_ = ~new_n5575_ | ~new_n5574_;
  assign new_n1420_ = ~new_n5577_ | ~new_n5576_;
  assign new_n1421_ = ~new_n5579_ | ~new_n5578_;
  assign new_n1422_ = ~new_n5582_ | ~new_n5581_ | ~new_n5580_;
  assign new_n1423_ = ~new_n5585_ | ~new_n5584_ | ~new_n5583_;
  assign new_n1424_ = ~new_n5687_ | ~new_n5688_ | ~new_n5686_;
  assign new_n1425_ = ~new_n5690_ | ~new_n5691_ | ~new_n5689_;
  assign new_n1426_ = new_n8144_ & new_n2804_;
  assign new_n1427_ = new_n2804_ & new_n8144_;
  assign new_n1428_ = new_n2804_ & new_n8010_;
  assign new_n1429_ = new_n2804_ & new_n8036_;
  assign new_n1430_ = new_n2804_ & new_n8037_;
  assign new_n1431_ = new_n2804_ & new_n8038_;
  assign new_n1432_ = new_n2804_ & new_n8039_;
  assign new_n1433_ = new_n2804_ & new_n8040_;
  assign new_n1434_ = new_n2804_ & new_n8041_;
  assign new_n1435_ = new_n2804_ & new_n8029_;
  assign new_n1436_ = ~new_n5517_ | ~new_n5516_;
  assign new_n1437_ = ~new_n5519_ | ~new_n5518_;
  assign new_n1438_ = ~new_n5521_ | ~new_n5520_;
  assign new_n1439_ = ~new_n5523_ | ~new_n5522_;
  assign new_n1440_ = ~new_n5525_ | ~new_n5524_;
  assign new_n1441_ = ~new_n5527_ | ~new_n5526_;
  assign new_n1442_ = ~new_n5528_ | ~new_n5529_ | ~new_n5530_;
  assign new_n1443_ = ~new_n5531_ | ~new_n2673_ | ~new_n5532_;
  assign new_n1444_ = ~new_n5534_ | ~new_n5535_ | ~new_n5536_;
  assign po518 = ~new_n6143_ | ~new_n5262_ | ~new_n2076_;
  assign po516 = ~new_n6295_ | ~new_n5258_;
  assign po515 = ~new_n5257_ | ~new_n5256_;
  assign po513 = ~new_n2888_ | ~new_n6414_ | ~new_n6413_;
  assign po511 = ~new_n2888_ | ~new_n6410_ | ~new_n6409_;
  assign po509 = ~new_n5246_ | ~new_n2893_;
  assign po506 = ~new_n2885_ | ~new_n6402_ | ~new_n6401_;
  assign po504 = ~new_n2885_ | ~new_n6392_ | ~new_n6391_;
  assign po503 = ~new_n5240_ | ~new_n5236_ | ~new_n2594_ | ~new_n5238_ | ~new_n2593_;
  assign po502 = ~new_n5233_ | ~new_n5229_ | ~new_n2592_ | ~new_n5231_ | ~new_n2591_;
  assign po501 = ~new_n5226_ | ~new_n5222_ | ~new_n2590_ | ~new_n5224_ | ~new_n2589_;
  assign po500 = ~new_n5219_ | ~new_n5215_ | ~new_n2588_ | ~new_n5217_ | ~new_n2587_;
  assign po499 = ~new_n5212_ | ~new_n5208_ | ~new_n2586_ | ~new_n5210_ | ~new_n2585_;
  assign po498 = ~new_n5205_ | ~new_n5201_ | ~new_n2584_ | ~new_n5203_ | ~new_n2583_;
  assign po497 = ~new_n5198_ | ~new_n5194_ | ~new_n2582_ | ~new_n5196_ | ~new_n2581_;
  assign po496 = ~new_n5191_ | ~new_n5187_ | ~new_n2580_ | ~new_n5189_ | ~new_n2579_;
  assign po495 = ~new_n5184_ | ~new_n5180_ | ~new_n2578_ | ~new_n5182_ | ~new_n2577_;
  assign po494 = ~new_n5177_ | ~new_n5173_ | ~new_n2576_ | ~new_n5175_ | ~new_n2575_;
  assign po493 = ~new_n5170_ | ~new_n5166_ | ~new_n2574_ | ~new_n5168_ | ~new_n2573_;
  assign po492 = ~new_n5163_ | ~new_n5159_ | ~new_n2572_ | ~new_n5161_ | ~new_n2571_;
  assign po491 = ~new_n5156_ | ~new_n5152_ | ~new_n2570_ | ~new_n2569_ | ~new_n5154_;
  assign po490 = ~new_n5149_ | ~new_n5145_ | ~new_n2568_ | ~new_n2567_ | ~new_n5147_;
  assign po489 = ~new_n5142_ | ~new_n5138_ | ~new_n2566_ | ~new_n2565_ | ~new_n5140_;
  assign po488 = ~new_n5135_ | ~new_n2563_ | ~new_n2564_ | ~new_n5133_ | ~new_n5132_;
  assign po487 = ~new_n5128_ | ~new_n2561_ | ~new_n2562_ | ~new_n5126_ | ~new_n5125_;
  assign po486 = ~new_n5121_ | ~new_n5118_ | ~new_n2559_ | ~new_n2560_ | ~new_n5119_;
  assign po485 = ~new_n5114_ | ~new_n5111_ | ~new_n2557_ | ~new_n2558_ | ~new_n5112_;
  assign po484 = ~new_n5107_ | ~new_n5104_ | ~new_n2555_ | ~new_n2556_ | ~new_n5105_;
  assign po483 = ~new_n5100_ | ~new_n5097_ | ~new_n2553_ | ~new_n2554_ | ~new_n5098_;
  assign po482 = ~new_n5093_ | ~new_n5090_ | ~new_n2551_ | ~new_n2552_ | ~new_n5091_;
  assign po481 = ~new_n5086_ | ~new_n5083_ | ~new_n2549_ | ~new_n2550_ | ~new_n5084_;
  assign po480 = ~new_n5079_ | ~new_n5076_ | ~new_n2547_ | ~new_n2548_ | ~new_n5077_;
  assign po479 = ~new_n5072_ | ~new_n5069_ | ~new_n2545_ | ~new_n2546_ | ~new_n5070_;
  assign po478 = ~new_n5065_ | ~new_n5062_ | ~new_n2543_ | ~new_n2544_ | ~new_n5063_;
  assign po477 = ~new_n2542_ | ~new_n5055_ | ~new_n2541_ | ~new_n5054_;
  assign po476 = ~new_n5047_ | ~new_n5048_ | ~new_n2540_ | ~new_n2539_ | ~new_n5046_;
  assign po475 = ~new_n2538_ | ~new_n5039_ | ~new_n5038_ | ~new_n5037_;
  assign po474 = ~new_n2537_ | ~new_n5031_ | ~new_n5030_ | ~new_n5029_;
  assign po473 = ~new_n2536_ | ~new_n5023_ | ~new_n5022_ | ~new_n5021_;
  assign po472 = ~new_n2535_ | ~new_n5015_ | ~new_n5014_ | ~new_n5013_;
  assign po471 = ~new_n5004_ | ~new_n5003_;
  assign po470 = ~new_n5000_ | ~new_n5001_ | ~new_n5002_;
  assign po469 = ~new_n4997_ | ~new_n4998_ | ~new_n4999_;
  assign po468 = ~new_n4994_ | ~new_n4995_ | ~new_n4996_;
  assign po467 = ~new_n4991_ | ~new_n4992_ | ~new_n4993_;
  assign po466 = ~new_n4988_ | ~new_n4989_ | ~new_n4990_;
  assign po465 = ~new_n4985_ | ~new_n4986_ | ~new_n4987_;
  assign po464 = ~new_n4982_ | ~new_n4983_ | ~new_n4984_;
  assign po463 = ~new_n4979_ | ~new_n4980_ | ~new_n4981_;
  assign po462 = ~new_n4976_ | ~new_n4977_ | ~new_n4978_;
  assign po461 = ~new_n4973_ | ~new_n4974_ | ~new_n4975_;
  assign po460 = ~new_n4970_ | ~new_n4971_ | ~new_n4972_;
  assign po459 = ~new_n4967_ | ~new_n4968_ | ~new_n4969_;
  assign po458 = ~new_n4964_ | ~new_n4965_ | ~new_n4966_;
  assign po457 = ~new_n4961_ | ~new_n4962_ | ~new_n4963_;
  assign po456 = ~new_n4958_ | ~new_n4959_ | ~new_n4960_;
  assign po455 = ~new_n4955_ | ~new_n4956_ | ~new_n4957_;
  assign po454 = ~new_n4952_ | ~new_n4953_ | ~new_n4954_;
  assign po453 = ~new_n4949_ | ~new_n4950_ | ~new_n4951_;
  assign po452 = ~new_n4946_ | ~new_n4947_ | ~new_n4948_;
  assign po451 = ~new_n4943_ | ~new_n4944_ | ~new_n4945_;
  assign po450 = ~new_n4940_ | ~new_n4941_ | ~new_n4942_;
  assign po449 = ~new_n4937_ | ~new_n4938_ | ~new_n4939_;
  assign po448 = ~new_n4934_ | ~new_n4935_ | ~new_n4936_;
  assign po447 = ~new_n4931_ | ~new_n4932_ | ~new_n4933_;
  assign po446 = ~new_n4928_ | ~new_n4929_ | ~new_n4930_;
  assign po445 = ~new_n4925_ | ~new_n4926_ | ~new_n4927_;
  assign po444 = ~new_n4922_ | ~new_n4923_ | ~new_n4924_;
  assign po443 = ~new_n4919_ | ~new_n4920_ | ~new_n4921_;
  assign po442 = ~new_n4916_ | ~new_n4917_ | ~new_n4918_;
  assign po441 = ~new_n4913_ | ~new_n4914_ | ~new_n4915_;
  assign po440 = ~new_n4912_ | ~new_n4911_ | ~new_n4910_;
  assign po439 = ~new_n2821_ | ~new_n4907_;
  assign po438 = ~new_n4905_ | ~new_n4906_ | ~new_n4904_ | ~new_n4903_;
  assign po437 = ~new_n4901_ | ~new_n4902_ | ~new_n4900_ | ~new_n4899_;
  assign po436 = ~new_n4897_ | ~new_n4898_ | ~new_n4896_ | ~new_n4895_;
  assign po435 = ~new_n4893_ | ~new_n4894_ | ~new_n4892_ | ~new_n4891_;
  assign po434 = ~new_n4889_ | ~new_n4890_ | ~new_n4888_ | ~new_n4887_;
  assign po433 = ~new_n4885_ | ~new_n4886_ | ~new_n4884_ | ~new_n4883_;
  assign po432 = ~new_n4881_ | ~new_n4882_ | ~new_n4880_ | ~new_n4879_;
  assign po431 = ~new_n4877_ | ~new_n4878_ | ~new_n4876_ | ~new_n4875_;
  assign po430 = ~new_n4873_ | ~new_n4874_ | ~new_n4872_ | ~new_n4871_;
  assign po429 = ~new_n4869_ | ~new_n4870_ | ~new_n4868_ | ~new_n4867_;
  assign po428 = ~new_n4865_ | ~new_n4866_ | ~new_n4864_ | ~new_n4863_;
  assign po427 = ~new_n4861_ | ~new_n4862_ | ~new_n4860_ | ~new_n4859_;
  assign po426 = ~new_n4857_ | ~new_n4858_ | ~new_n4856_ | ~new_n4855_;
  assign po425 = ~new_n4853_ | ~new_n4854_ | ~new_n4852_ | ~new_n4851_;
  assign po424 = ~new_n4849_ | ~new_n4850_ | ~new_n4848_ | ~new_n4847_;
  assign po423 = ~new_n4845_ | ~new_n4846_ | ~new_n4844_;
  assign po422 = ~new_n4842_ | ~new_n4843_ | ~new_n4841_;
  assign po421 = ~new_n4839_ | ~new_n4840_ | ~new_n4838_;
  assign po420 = ~new_n4836_ | ~new_n4837_ | ~new_n4835_;
  assign po419 = ~new_n4833_ | ~new_n4834_ | ~new_n4832_;
  assign po418 = ~new_n4830_ | ~new_n4831_ | ~new_n4829_;
  assign po417 = ~new_n4827_ | ~new_n4828_ | ~new_n4826_;
  assign po416 = ~new_n4824_ | ~new_n4825_ | ~new_n4823_;
  assign po415 = ~new_n4821_ | ~new_n4822_ | ~new_n4820_;
  assign po414 = ~new_n4818_ | ~new_n4819_ | ~new_n4817_;
  assign po413 = ~new_n4815_ | ~new_n4816_ | ~new_n4814_;
  assign po412 = ~new_n4812_ | ~new_n4813_ | ~new_n4811_;
  assign po411 = ~new_n4809_ | ~new_n4810_ | ~new_n4808_;
  assign po410 = ~new_n4806_ | ~new_n4807_ | ~new_n4805_;
  assign po409 = ~new_n4804_ | ~new_n4803_ | ~new_n4802_;
  assign po408 = ~new_n4801_ | ~new_n4800_ | ~new_n4799_;
  assign po407 = pi374 & new_n4700_;
  assign po406 = ~new_n2527_ | ~new_n4791_;
  assign po405 = ~new_n2526_ | ~new_n4788_;
  assign po404 = ~new_n2525_ | ~new_n4785_;
  assign po403 = ~new_n2524_ | ~new_n4782_;
  assign po402 = ~new_n2523_ | ~new_n4779_;
  assign po401 = ~new_n2522_ | ~new_n4776_;
  assign po400 = ~new_n2521_ | ~new_n4773_;
  assign po399 = ~new_n2520_ | ~new_n4770_;
  assign po398 = ~new_n2519_ | ~new_n4767_;
  assign po397 = ~new_n2518_ | ~new_n4764_;
  assign po396 = ~new_n2517_ | ~new_n4761_;
  assign po395 = ~new_n2516_ | ~new_n4758_;
  assign po394 = ~new_n2515_ | ~new_n4755_;
  assign po393 = ~new_n2514_ | ~new_n4752_;
  assign po392 = ~new_n2513_ | ~new_n4749_;
  assign po391 = ~new_n4748_ | ~new_n4747_ | ~new_n4746_;
  assign po390 = ~new_n4745_ | ~new_n4744_ | ~new_n4743_;
  assign po389 = ~new_n4742_ | ~new_n4741_ | ~new_n4740_;
  assign po388 = ~new_n4739_ | ~new_n4738_ | ~new_n4737_;
  assign po387 = ~new_n4736_ | ~new_n4735_ | ~new_n4734_;
  assign po386 = ~new_n4733_ | ~new_n4732_ | ~new_n4731_;
  assign po385 = ~new_n4730_ | ~new_n4729_ | ~new_n4728_;
  assign po384 = ~new_n4727_ | ~new_n4726_ | ~new_n4725_;
  assign po383 = ~new_n4724_ | ~new_n4723_ | ~new_n4722_;
  assign po382 = ~new_n4721_ | ~new_n4720_ | ~new_n4719_;
  assign po381 = ~new_n4718_ | ~new_n4717_ | ~new_n4716_;
  assign po380 = ~new_n4715_ | ~new_n4714_ | ~new_n4713_;
  assign po379 = ~new_n4712_ | ~new_n4711_ | ~new_n4710_;
  assign po378 = ~new_n4709_ | ~new_n4708_ | ~new_n4707_;
  assign po377 = ~new_n4706_ | ~new_n4705_ | ~new_n4704_;
  assign po376 = ~new_n4703_ | ~new_n4702_ | ~new_n4701_;
  assign po375 = ~new_n6185_ | ~new_n6187_;
  assign po374 = ~new_n6184_ | ~new_n6189_;
  assign po373 = ~new_n6183_ | ~new_n6191_;
  assign po372 = ~new_n6182_ | ~new_n6193_;
  assign po371 = ~new_n6181_ | ~new_n6195_;
  assign po370 = ~new_n6180_ | ~new_n6197_;
  assign po369 = ~new_n6179_ | ~new_n6199_;
  assign po368 = ~new_n6178_ | ~new_n6201_;
  assign po367 = ~new_n6177_ | ~new_n6203_;
  assign po366 = ~new_n6176_ | ~new_n6205_;
  assign po365 = ~new_n6175_ | ~new_n6207_;
  assign po364 = ~new_n6174_ | ~new_n6209_;
  assign po363 = ~new_n6173_ | ~new_n6211_;
  assign po362 = ~new_n6172_ | ~new_n6213_;
  assign po361 = ~new_n6171_ | ~new_n6215_;
  assign po360 = ~new_n6170_ | ~new_n6217_;
  assign po359 = ~new_n6169_ | ~new_n6219_;
  assign po358 = ~new_n6168_ | ~new_n6221_;
  assign po357 = ~new_n6167_ | ~new_n6223_;
  assign po356 = ~new_n6166_ | ~new_n6225_;
  assign po355 = ~new_n6165_ | ~new_n6227_;
  assign po354 = ~new_n6164_ | ~new_n6229_;
  assign po353 = ~new_n6163_ | ~new_n6231_;
  assign po352 = ~new_n6162_ | ~new_n6233_;
  assign po351 = ~new_n6161_ | ~new_n6235_;
  assign po350 = ~new_n6160_ | ~new_n6237_;
  assign po349 = ~new_n6159_ | ~new_n6239_;
  assign po348 = ~new_n6158_ | ~new_n6241_;
  assign po347 = ~new_n6157_ | ~new_n6243_;
  assign po346 = ~new_n6156_ | ~new_n6245_;
  assign po345 = ~new_n6155_ | ~new_n6247_;
  assign po344 = ~new_n4602_ | ~new_n4600_ | ~new_n4603_ | ~new_n4601_ | ~new_n4599_;
  assign po343 = ~new_n4597_ | ~new_n4595_ | ~new_n4598_ | ~new_n4596_ | ~new_n4594_;
  assign po342 = ~new_n4592_ | ~new_n4590_ | ~new_n4593_ | ~new_n4591_ | ~new_n4589_;
  assign po341 = ~new_n4587_ | ~new_n4585_ | ~new_n4588_ | ~new_n4586_ | ~new_n4584_;
  assign po340 = ~new_n4582_ | ~new_n4580_ | ~new_n4583_ | ~new_n4581_ | ~new_n4579_;
  assign po339 = ~new_n4577_ | ~new_n4575_ | ~new_n4578_ | ~new_n4576_ | ~new_n4574_;
  assign po338 = ~new_n4572_ | ~new_n4570_ | ~new_n4573_ | ~new_n4571_ | ~new_n4569_;
  assign po337 = ~new_n4567_ | ~new_n4565_ | ~new_n4568_ | ~new_n4566_ | ~new_n4564_;
  assign po336 = ~new_n4562_ | ~new_n4560_ | ~new_n4563_ | ~new_n4561_ | ~new_n4559_;
  assign po335 = ~new_n4557_ | ~new_n4555_ | ~new_n4558_ | ~new_n4556_ | ~new_n4554_;
  assign po334 = ~new_n4552_ | ~new_n4550_ | ~new_n4553_ | ~new_n4551_ | ~new_n4549_;
  assign po333 = ~new_n4547_ | ~new_n4545_ | ~new_n4548_ | ~new_n4546_ | ~new_n4544_;
  assign po332 = ~new_n4542_ | ~new_n4540_ | ~new_n4543_ | ~new_n4541_ | ~new_n4539_;
  assign po331 = ~new_n4537_ | ~new_n4535_ | ~new_n4538_ | ~new_n4536_ | ~new_n4534_;
  assign po330 = ~new_n4532_ | ~new_n4530_ | ~new_n4533_ | ~new_n4531_ | ~new_n4529_;
  assign po329 = ~new_n4527_ | ~new_n4525_ | ~new_n4528_ | ~new_n4526_ | ~new_n4524_;
  assign po328 = ~new_n4522_ | ~new_n4520_ | ~new_n4523_ | ~new_n4521_ | ~new_n4519_;
  assign po327 = ~new_n4517_ | ~new_n4515_ | ~new_n4518_ | ~new_n4516_ | ~new_n4514_;
  assign po326 = ~new_n4512_ | ~new_n4510_ | ~new_n4513_ | ~new_n4511_ | ~new_n4509_;
  assign po325 = ~new_n4507_ | ~new_n4505_ | ~new_n4508_ | ~new_n4506_ | ~new_n4504_;
  assign po324 = ~new_n4502_ | ~new_n4500_ | ~new_n4503_ | ~new_n4501_ | ~new_n4499_;
  assign po323 = ~new_n4497_ | ~new_n4495_ | ~new_n4498_ | ~new_n4496_ | ~new_n4494_;
  assign po322 = ~new_n4492_ | ~new_n4490_ | ~new_n4493_ | ~new_n4491_ | ~new_n4489_;
  assign po321 = ~new_n4487_ | ~new_n4485_ | ~new_n4488_ | ~new_n4486_ | ~new_n4484_;
  assign po320 = ~new_n4482_ | ~new_n4483_ | ~new_n4480_ | ~new_n4481_ | ~new_n4479_;
  assign po319 = ~new_n4477_ | ~new_n4478_ | ~new_n4475_ | ~new_n4476_ | ~new_n4474_;
  assign po318 = ~new_n4472_ | ~new_n4473_ | ~new_n4470_ | ~new_n4471_ | ~new_n4469_;
  assign po317 = ~new_n4467_ | ~new_n4468_ | ~new_n4465_ | ~new_n4466_ | ~new_n4464_;
  assign po316 = ~new_n4462_ | ~new_n4463_ | ~new_n4460_ | ~new_n4461_ | ~new_n4459_;
  assign po315 = ~new_n4457_ | ~new_n4458_ | ~new_n4455_ | ~new_n4456_ | ~new_n4454_;
  assign po314 = ~new_n4452_ | ~new_n4453_ | ~new_n4451_ | ~new_n4450_ | ~new_n4449_;
  assign po313 = ~new_n4447_ | ~new_n4448_ | ~new_n4446_ | ~new_n4445_ | ~new_n4444_;
  assign po312 = ~new_n4434_ | ~new_n4432_ | ~new_n2506_ | ~new_n2504_;
  assign po311 = ~new_n4427_ | ~new_n4425_ | ~new_n2503_ | ~new_n2501_;
  assign po310 = ~new_n4420_ | ~new_n4418_ | ~new_n2500_ | ~new_n2498_;
  assign po309 = ~new_n4413_ | ~new_n4411_ | ~new_n2497_ | ~new_n2495_;
  assign po308 = ~new_n4406_ | ~new_n4404_ | ~new_n2494_ | ~new_n2492_;
  assign po307 = ~new_n4399_ | ~new_n4397_ | ~new_n2491_ | ~new_n2489_;
  assign po306 = ~new_n4392_ | ~new_n4390_ | ~new_n2488_ | ~new_n2486_;
  assign po305 = ~new_n4385_ | ~new_n4383_ | ~new_n2485_ | ~new_n2483_;
  assign po304 = ~new_n4378_ | ~new_n4376_ | ~new_n2482_ | ~new_n2480_;
  assign po303 = ~new_n4371_ | ~new_n4369_ | ~new_n2479_ | ~new_n2477_;
  assign po302 = ~new_n4364_ | ~new_n4362_ | ~new_n2476_ | ~new_n2474_;
  assign po301 = ~new_n4357_ | ~new_n4355_ | ~new_n2473_ | ~new_n2471_;
  assign po300 = ~new_n4350_ | ~new_n4348_ | ~new_n2470_ | ~new_n2468_;
  assign po299 = ~new_n4343_ | ~new_n4341_ | ~new_n2467_ | ~new_n2465_;
  assign po298 = ~new_n4336_ | ~new_n4334_ | ~new_n2464_ | ~new_n2462_;
  assign po297 = ~new_n4329_ | ~new_n4327_ | ~new_n2461_ | ~new_n2459_;
  assign po296 = ~new_n4322_ | ~new_n4320_ | ~new_n2458_ | ~new_n2456_;
  assign po295 = ~new_n4315_ | ~new_n4313_ | ~new_n2455_ | ~new_n2453_;
  assign po294 = ~new_n4308_ | ~new_n4306_ | ~new_n2452_ | ~new_n2450_;
  assign po293 = ~new_n4301_ | ~new_n2447_ | ~new_n2449_;
  assign po292 = ~new_n4294_ | ~new_n2444_ | ~new_n2446_;
  assign po291 = ~new_n4287_ | ~new_n2441_ | ~new_n2443_;
  assign po290 = ~new_n4280_ | ~new_n2438_ | ~new_n2440_;
  assign po289 = ~new_n4273_ | ~new_n2435_ | ~new_n2437_;
  assign po288 = ~new_n4266_ | ~new_n2432_ | ~new_n2434_;
  assign po287 = ~new_n4259_ | ~new_n2429_ | ~new_n2431_;
  assign po286 = ~new_n4252_ | ~new_n2426_ | ~new_n2428_;
  assign po285 = ~new_n4245_ | ~new_n2423_ | ~new_n2425_;
  assign po284 = ~new_n2420_ | ~new_n2421_;
  assign po283 = ~new_n2419_ | ~new_n2417_ | ~new_n2416_;
  assign po282 = ~new_n2415_ | ~new_n2413_ | ~new_n2412_;
  assign po281 = ~new_n2411_ | ~new_n2409_ | ~new_n2408_;
  assign po276 = pi243 & new_n4182_;
  assign po270 = ~new_n2375_ | ~new_n4105_ | ~new_n4104_;
  assign po269 = ~new_n2374_ | ~new_n4100_ | ~new_n4099_;
  assign po268 = ~new_n2373_ | ~new_n4095_ | ~new_n4094_;
  assign po267 = ~new_n2372_ | ~new_n4090_ | ~new_n4089_;
  assign po266 = ~new_n2371_ | ~new_n6257_ | ~new_n4085_;
  assign po265 = ~new_n2370_ | ~new_n4081_ | ~new_n4080_;
  assign po264 = ~new_n2369_ | ~new_n4076_ | ~new_n4075_;
  assign po263 = ~new_n2368_ | ~new_n4071_ | ~new_n4070_;
  assign po262 = ~new_n2366_ | ~new_n4049_ | ~new_n4048_;
  assign po261 = ~new_n2365_ | ~new_n4044_ | ~new_n4043_;
  assign po260 = ~new_n2364_ | ~new_n4039_ | ~new_n4038_;
  assign po259 = ~new_n2363_ | ~new_n4034_ | ~new_n4033_;
  assign po258 = ~new_n2362_ | ~new_n4029_ | ~new_n4028_;
  assign po257 = ~new_n2361_ | ~new_n4024_ | ~new_n4023_;
  assign po256 = ~new_n2360_ | ~new_n4019_ | ~new_n4018_;
  assign po255 = ~new_n2359_ | ~new_n4014_ | ~new_n4013_;
  assign po254 = ~new_n2357_ | ~new_n3991_ | ~new_n3990_;
  assign po253 = ~new_n2356_ | ~new_n3986_ | ~new_n3985_;
  assign po252 = ~new_n2355_ | ~new_n3981_ | ~new_n3980_;
  assign po251 = ~new_n2354_ | ~new_n3976_ | ~new_n3975_;
  assign po250 = ~new_n2353_ | ~new_n3971_ | ~new_n3970_;
  assign po249 = ~new_n2352_ | ~new_n3966_ | ~new_n3965_;
  assign po248 = ~new_n2351_ | ~new_n3961_ | ~new_n3960_;
  assign po247 = ~new_n2350_ | ~new_n3956_ | ~new_n3955_;
  assign po246 = ~new_n2348_ | ~new_n3934_ | ~new_n3933_;
  assign po245 = ~new_n2347_ | ~new_n3929_ | ~new_n3928_;
  assign po244 = ~new_n2346_ | ~new_n3924_ | ~new_n3923_;
  assign po243 = ~new_n2345_ | ~new_n3919_ | ~new_n3918_;
  assign po242 = ~new_n2344_ | ~new_n3914_ | ~new_n3913_;
  assign po241 = ~new_n2343_ | ~new_n3909_ | ~new_n3908_;
  assign po240 = ~new_n2342_ | ~new_n3904_ | ~new_n3903_;
  assign po239 = ~new_n2341_ | ~new_n3899_ | ~new_n3898_;
  assign po238 = ~new_n2339_ | ~new_n3876_ | ~new_n3875_;
  assign po237 = ~new_n2338_ | ~new_n3871_ | ~new_n3870_;
  assign po236 = ~new_n2337_ | ~new_n3866_ | ~new_n3865_;
  assign po235 = ~new_n2336_ | ~new_n3861_ | ~new_n3860_;
  assign po234 = ~new_n2335_ | ~new_n3856_ | ~new_n3855_;
  assign po233 = ~new_n2334_ | ~new_n3851_ | ~new_n3850_;
  assign po232 = ~new_n2333_ | ~new_n3846_ | ~new_n3845_;
  assign po231 = ~new_n2332_ | ~new_n3841_ | ~new_n3840_;
  assign po230 = ~new_n2330_ | ~new_n3819_ | ~new_n3818_;
  assign po229 = ~new_n2329_ | ~new_n3814_ | ~new_n3813_;
  assign po228 = ~new_n2328_ | ~new_n3809_ | ~new_n3808_;
  assign po227 = ~new_n2327_ | ~new_n3804_ | ~new_n3803_;
  assign po226 = ~new_n2326_ | ~new_n3799_ | ~new_n3798_;
  assign po225 = ~new_n2325_ | ~new_n3794_ | ~new_n3793_;
  assign po224 = ~new_n2324_ | ~new_n3789_ | ~new_n3788_;
  assign po223 = ~new_n2323_ | ~new_n3784_ | ~new_n3783_;
  assign po222 = ~new_n2321_ | ~new_n3761_ | ~new_n3760_;
  assign po221 = ~new_n2320_ | ~new_n3756_ | ~new_n3755_;
  assign po220 = ~new_n2319_ | ~new_n3751_ | ~new_n3750_;
  assign po219 = ~new_n2318_ | ~new_n3746_ | ~new_n3745_;
  assign po218 = ~new_n2317_ | ~new_n3741_ | ~new_n3740_;
  assign po217 = ~new_n2316_ | ~new_n3736_ | ~new_n3735_;
  assign po216 = ~new_n2315_ | ~new_n3731_ | ~new_n3730_;
  assign po215 = ~new_n2314_ | ~new_n3726_ | ~new_n3725_;
  assign po214 = ~new_n2312_ | ~new_n3704_ | ~new_n3703_;
  assign po213 = ~new_n2311_ | ~new_n3699_ | ~new_n3698_;
  assign po212 = ~new_n2310_ | ~new_n3694_ | ~new_n3693_;
  assign po211 = ~new_n2309_ | ~new_n3689_ | ~new_n3688_;
  assign po210 = ~new_n2308_ | ~new_n3684_ | ~new_n3683_;
  assign po209 = ~new_n2307_ | ~new_n3679_ | ~new_n3678_;
  assign po208 = ~new_n2306_ | ~new_n3674_ | ~new_n3673_;
  assign po207 = ~new_n2305_ | ~new_n3669_ | ~new_n3668_;
  assign po206 = ~new_n2303_ | ~new_n3648_ | ~new_n3647_;
  assign po205 = ~new_n2302_ | ~new_n3643_ | ~new_n3642_;
  assign po204 = ~new_n2301_ | ~new_n3638_ | ~new_n3637_;
  assign po203 = ~new_n2300_ | ~new_n3633_ | ~new_n3632_;
  assign po202 = ~new_n2299_ | ~new_n3628_ | ~new_n3627_;
  assign po201 = ~new_n2298_ | ~new_n3623_ | ~new_n3622_;
  assign po200 = ~new_n2297_ | ~new_n3618_ | ~new_n3617_;
  assign po199 = ~new_n2296_ | ~new_n3613_ | ~new_n3612_;
  assign po198 = ~new_n2294_ | ~new_n3591_ | ~new_n3590_;
  assign po197 = ~new_n2293_ | ~new_n3586_ | ~new_n3585_;
  assign po196 = ~new_n2292_ | ~new_n3581_ | ~new_n3580_;
  assign po195 = ~new_n2291_ | ~new_n3576_ | ~new_n3575_;
  assign po194 = ~new_n2290_ | ~new_n3571_ | ~new_n3570_;
  assign po193 = ~new_n2289_ | ~new_n3566_ | ~new_n3565_;
  assign po192 = ~new_n2288_ | ~new_n3561_ | ~new_n3560_;
  assign po191 = ~new_n2287_ | ~new_n3556_ | ~new_n3555_;
  assign po190 = ~new_n2285_ | ~new_n3533_ | ~new_n3532_;
  assign po189 = ~new_n2284_ | ~new_n3528_ | ~new_n3527_;
  assign po188 = ~new_n2283_ | ~new_n3523_ | ~new_n3522_;
  assign po187 = ~new_n2282_ | ~new_n3518_ | ~new_n3517_;
  assign po186 = ~new_n2281_ | ~new_n3513_ | ~new_n3512_;
  assign po185 = ~new_n2280_ | ~new_n3508_ | ~new_n3507_;
  assign po184 = ~new_n2279_ | ~new_n3503_ | ~new_n3502_;
  assign po183 = ~new_n2278_ | ~new_n3498_ | ~new_n3497_;
  assign po182 = ~new_n2276_ | ~new_n3476_ | ~new_n3475_;
  assign po181 = ~new_n2275_ | ~new_n3471_ | ~new_n3470_;
  assign po180 = ~new_n2274_ | ~new_n3466_ | ~new_n3465_;
  assign po179 = ~new_n2273_ | ~new_n3461_ | ~new_n3460_;
  assign po178 = ~new_n2272_ | ~new_n3456_ | ~new_n3455_;
  assign po177 = ~new_n2271_ | ~new_n3451_ | ~new_n3450_;
  assign po176 = ~new_n2270_ | ~new_n3446_ | ~new_n3445_;
  assign po175 = ~new_n2269_ | ~new_n3441_ | ~new_n3440_;
  assign po174 = ~new_n2267_ | ~new_n3418_ | ~new_n3417_;
  assign po173 = ~new_n2266_ | ~new_n3413_ | ~new_n3412_;
  assign po172 = ~new_n2265_ | ~new_n3408_ | ~new_n3407_;
  assign po171 = ~new_n2264_ | ~new_n3403_ | ~new_n3402_;
  assign po170 = ~new_n2263_ | ~new_n3398_ | ~new_n3397_;
  assign po169 = ~new_n2262_ | ~new_n3393_ | ~new_n3392_;
  assign po168 = ~new_n2261_ | ~new_n3388_ | ~new_n3387_;
  assign po167 = ~new_n2260_ | ~new_n3383_ | ~new_n3382_;
  assign po166 = ~new_n2258_ | ~new_n3361_ | ~new_n3360_;
  assign po165 = ~new_n2257_ | ~new_n3356_ | ~new_n3355_;
  assign po164 = ~new_n2256_ | ~new_n3351_ | ~new_n3350_;
  assign po163 = ~new_n2255_ | ~new_n3346_ | ~new_n3345_;
  assign po162 = ~new_n2254_ | ~new_n3341_ | ~new_n3340_;
  assign po161 = ~new_n2253_ | ~new_n3336_ | ~new_n3335_;
  assign po160 = ~new_n2252_ | ~new_n3331_ | ~new_n3330_;
  assign po159 = ~new_n2251_ | ~new_n3326_ | ~new_n3325_;
  assign po158 = ~new_n2249_ | ~new_n3302_ | ~new_n3301_;
  assign po157 = ~new_n2248_ | ~new_n3297_ | ~new_n3296_;
  assign po156 = ~new_n2247_ | ~new_n3292_ | ~new_n3291_;
  assign po155 = ~new_n2246_ | ~new_n3287_ | ~new_n3286_;
  assign po154 = ~new_n2245_ | ~new_n3282_ | ~new_n3281_;
  assign po153 = ~new_n2244_ | ~new_n3277_ | ~new_n3276_;
  assign po152 = ~new_n2243_ | ~new_n3272_ | ~new_n3271_;
  assign po151 = ~new_n2242_ | ~new_n3267_ | ~new_n3266_;
  assign po150 = ~new_n2240_ | ~new_n3244_ | ~new_n3243_;
  assign po149 = ~new_n2239_ | ~new_n3239_ | ~new_n3238_;
  assign po148 = ~new_n2238_ | ~new_n3234_ | ~new_n3233_;
  assign po147 = ~new_n2237_ | ~new_n3229_ | ~new_n3228_;
  assign po146 = ~new_n2236_ | ~new_n3224_ | ~new_n3223_;
  assign po145 = ~new_n2235_ | ~new_n3219_ | ~new_n3218_;
  assign po144 = ~new_n2234_ | ~new_n3214_ | ~new_n3213_;
  assign po143 = ~new_n2233_ | ~new_n3209_ | ~new_n3208_;
  assign po142 = ~new_n2231_ | ~new_n6335_ | ~new_n6334_;
  assign po141 = ~new_n2889_ | ~new_n3163_ | ~new_n3165_ | ~new_n3164_;
  assign po140 = ~new_n2227_ | ~new_n3161_;
  assign po138 = pi105 & new_n6295_;
  assign po137 = pi104 & new_n6295_;
  assign po136 = pi103 & new_n6295_;
  assign po135 = pi102 & new_n6295_;
  assign po134 = pi101 & new_n6295_;
  assign po133 = pi100 & new_n6295_;
  assign po132 = pi099 & new_n6295_;
  assign po131 = pi098 & new_n6295_;
  assign po130 = pi097 & new_n6295_;
  assign po129 = pi096 & new_n6295_;
  assign po128 = pi095 & new_n6295_;
  assign po127 = pi094 & new_n6295_;
  assign po126 = pi093 & new_n6295_;
  assign po125 = pi092 & new_n6295_;
  assign po124 = pi091 & new_n6295_;
  assign po123 = pi090 & new_n6295_;
  assign po122 = pi089 & new_n6295_;
  assign po121 = pi088 & new_n6295_;
  assign po120 = pi087 & new_n6295_;
  assign po119 = pi086 & new_n6295_;
  assign po118 = pi085 & new_n6295_;
  assign po117 = pi084 & new_n6295_;
  assign po116 = pi083 & new_n6295_;
  assign po115 = pi082 & new_n6295_;
  assign po114 = pi081 & new_n6295_;
  assign po113 = pi080 & new_n6295_;
  assign po112 = pi079 & new_n6295_;
  assign po111 = pi078 & new_n6295_;
  assign po110 = pi077 & new_n6295_;
  assign po109 = pi076 & new_n6295_;
  assign po106 = ~new_n3020_ | ~new_n6292_ | ~new_n6291_;
  assign po105 = ~new_n2140_ | ~new_n6290_ | ~new_n6289_;
  assign po104 = ~new_n2139_ | ~new_n3014_;
  assign po103 = ~new_n3001_ | ~new_n3000_ | ~new_n2999_;
  assign po102 = ~new_n2998_ | ~new_n2997_ | ~new_n2996_;
  assign po101 = ~new_n2995_ | ~new_n2994_ | ~new_n2993_;
  assign po100 = ~new_n2992_ | ~new_n2991_ | ~new_n2990_;
  assign po099 = ~new_n2989_ | ~new_n2988_ | ~new_n2987_;
  assign po098 = ~new_n2986_ | ~new_n2985_ | ~new_n2984_;
  assign po097 = ~new_n2983_ | ~new_n2982_ | ~new_n2981_;
  assign po096 = ~new_n2980_ | ~new_n2979_ | ~new_n2978_;
  assign po095 = ~new_n2977_ | ~new_n2976_ | ~new_n2975_;
  assign po094 = ~new_n2974_ | ~new_n2973_ | ~new_n2972_;
  assign po093 = ~new_n2971_ | ~new_n2970_ | ~new_n2969_;
  assign po092 = ~new_n2968_ | ~new_n2967_ | ~new_n2966_;
  assign po091 = ~new_n2965_ | ~new_n2964_ | ~new_n2963_;
  assign po090 = ~new_n2962_ | ~new_n2961_ | ~new_n2960_;
  assign po089 = ~new_n2959_ | ~new_n2958_ | ~new_n2957_;
  assign po088 = ~new_n2956_ | ~new_n2955_ | ~new_n2954_;
  assign po087 = ~new_n2953_ | ~new_n2952_ | ~new_n2951_;
  assign po086 = ~new_n2950_ | ~new_n2949_ | ~new_n2948_;
  assign po085 = ~new_n2947_ | ~new_n2946_ | ~new_n2945_;
  assign po084 = ~new_n2944_ | ~new_n2943_ | ~new_n2942_;
  assign po083 = ~new_n2941_ | ~new_n2940_ | ~new_n2939_;
  assign po082 = ~new_n2938_ | ~new_n2937_ | ~new_n2936_;
  assign po081 = ~new_n2935_ | ~new_n2934_ | ~new_n2933_;
  assign po080 = ~new_n2932_ | ~new_n2931_ | ~new_n2930_;
  assign po079 = ~new_n2929_ | ~new_n2928_ | ~new_n2927_;
  assign po078 = ~new_n2926_ | ~new_n2925_ | ~new_n2924_;
  assign po077 = ~new_n2923_ | ~new_n2922_ | ~new_n2921_;
  assign po076 = ~new_n2920_ | ~new_n2919_ | ~new_n2918_;
  assign po075 = ~new_n2917_ | ~new_n2916_ | ~new_n2915_;
  assign po074 = ~new_n2914_ | ~new_n2913_ | ~new_n2912_;
  assign new_n1871_ = ~new_n2643_ | ~new_n2644_ | ~new_n2646_ | ~new_n2645_;
  assign new_n1872_ = ~new_n2639_ | ~new_n2640_ | ~new_n2642_ | ~new_n2641_;
  assign new_n1873_ = ~new_n2635_ | ~new_n2636_ | ~new_n2638_ | ~new_n2637_;
  assign new_n1874_ = ~new_n2631_ | ~new_n2632_ | ~new_n2634_ | ~new_n2633_;
  assign new_n1875_ = ~new_n2627_ | ~new_n2628_ | ~new_n2630_ | ~new_n2629_;
  assign new_n1876_ = ~new_n2623_ | ~new_n2624_ | ~new_n2626_ | ~new_n2625_;
  assign new_n1877_ = ~new_n2619_ | ~new_n2620_ | ~new_n2622_ | ~new_n2621_;
  assign new_n1878_ = ~new_n2615_ | ~new_n2616_ | ~new_n2618_ | ~new_n2617_;
  assign new_n1879_ = ~new_n1973_ | ~new_n1967_;
  assign new_n1880_ = ~new_n1089_ | ~new_n1879_;
  assign new_n1881_ = ~new_n1089_ | ~new_n3188_;
  assign new_n1882_ = ~new_n1091_ | ~new_n1879_;
  assign new_n1883_ = ~new_n1091_ | ~new_n3188_;
  assign new_n1884_ = ~new_n1090_ | ~new_n1879_;
  assign new_n1885_ = ~new_n1090_ | ~new_n3188_;
  assign new_n1886_ = ~new_n1092_ | ~new_n1879_;
  assign new_n1887_ = ~new_n1092_ | ~new_n3188_;
  assign new_n1888_ = ~new_n4108_ | ~new_n2035_ | ~new_n2038_;
  assign new_n1889_ = ~new_n5731_ | ~new_n4109_;
  assign new_n1890_ = ~new_n2801_ | ~new_n2803_ | ~new_n6437_ | ~new_n6436_;
  assign new_n1891_ = ~pi479;
  assign new_n1892_ = ~pi072;
  assign new_n1893_ = ~pi072 | ~new_n1902_;
  assign new_n1894_ = ~new_n2866_ | ~new_n1895_;
  assign new_n1895_ = ~pi071;
  assign new_n1896_ = ~pi071 | ~new_n2866_;
  assign new_n1897_ = ~pi440;
  assign new_n1898_ = ~pi072 | ~new_n1895_;
  assign new_n1899_ = pi072 | pi071;
  assign new_n1900_ = ~pi036;
  assign new_n1901_ = ~pi035;
  assign new_n1902_ = ~pi073;
  assign new_n1903_ = ~pi073 | ~new_n1904_;
  assign new_n1904_ = ~pi479 | ~new_n1900_;
  assign new_n1905_ = pi036 | pi479;
  assign new_n1906_ = ~pi108;
  assign new_n1907_ = ~pi107;
  assign new_n1908_ = ~pi240;
  assign new_n1909_ = ~pi241;
  assign new_n1910_ = ~pi242;
  assign new_n1911_ = ~new_n1914_ | ~pi240 | ~pi242 | ~pi241;
  assign new_n1912_ = pi240 | pi242 | pi241;
  assign new_n1913_ = pi241 | pi242;
  assign new_n1914_ = ~pi239;
  assign new_n1915_ = ~new_n2209_ | ~new_n2210_ | ~new_n2212_ | ~new_n2211_;
  assign new_n1916_ = ~new_n3141_ | ~new_n1902_;
  assign new_n1917_ = ~new_n8624_;
  assign new_n1918_ = ~pi240 | ~new_n1914_;
  assign new_n1919_ = ~pi242 | ~pi241;
  assign new_n1920_ = ~new_n2161_ | ~new_n2162_ | ~new_n2164_ | ~new_n2163_;
  assign new_n1921_ = ~new_n2181_ | ~new_n2182_ | ~new_n2183_ | ~new_n2184_ | ~new_n2815_;
  assign new_n1922_ = ~new_n2199_ | ~new_n2200_ | ~new_n2202_ | ~new_n2201_;
  assign new_n1923_ = ~new_n2204_ | ~new_n2203_;
  assign new_n1924_ = pi478 | pi035;
  assign new_n1925_ = ~new_n8624_ | ~new_n3142_;
  assign new_n1926_ = ~new_n3122_ | ~new_n1928_;
  assign new_n1927_ = ~new_n2153_ | ~new_n2154_ | ~new_n2156_ | ~new_n2155_;
  assign new_n1928_ = ~new_n2205_ | ~new_n2206_ | ~new_n2208_ | ~new_n2207_;
  assign new_n1929_ = ~new_n1130_ | ~new_n3146_;
  assign new_n1930_ = ~new_n1046_ | ~new_n1927_;
  assign new_n1931_ = ~new_n3139_ | ~new_n3122_;
  assign new_n1932_ = ~new_n2894_ | ~new_n1104_;
  assign new_n1933_ = ~new_n1922_ | ~new_n2818_ | ~new_n3105_ | ~new_n2035_;
  assign new_n1934_ = ~new_n1915_ | ~new_n1927_;
  assign new_n1935_ = ~new_n2835_ | ~new_n1928_;
  assign new_n1936_ = ~new_n2901_ | ~new_n1088_;
  assign new_n1937_ = ~new_n8854_ | ~new_n2870_ | ~new_n6271_ | ~new_n2823_ | ~new_n3154_;
  assign new_n1938_ = ~pi109;
  assign new_n1939_ = ~pi109 | ~new_n6249_;
  assign new_n1940_ = ~pi106;
  assign new_n1941_ = ~pi107 | ~new_n1906_;
  assign new_n1942_ = pi107 | pi108;
  assign new_n1943_ = ~pi106 | ~new_n8624_;
  assign new_n1944_ = ~new_n3192_ | ~new_n1938_;
  assign new_n1945_ = ~pi247;
  assign new_n1946_ = ~pi246;
  assign new_n1947_ = ~pi244;
  assign new_n1948_ = ~pi245;
  assign new_n1949_ = ~pi246 | ~pi247;
  assign new_n1950_ = ~new_n3178_ | ~new_n1135_;
  assign new_n1951_ = pi107 | pi106;
  assign new_n1952_ = ~pi478;
  assign new_n1953_ = ~new_n8042_;
  assign new_n1954_ = ~new_n8049_;
  assign new_n1955_ = ~new_n8048_;
  assign new_n1956_ = ~new_n8007_;
  assign new_n1957_ = ~new_n8049_ | ~new_n8042_;
  assign new_n1958_ = ~new_n1976_ | ~new_n1953_;
  assign new_n1959_ = ~new_n3172_ | ~new_n1132_;
  assign new_n1960_ = ~new_n7942_;
  assign new_n1961_ = ~new_n7959_;
  assign new_n1962_ = ~new_n7951_;
  assign new_n1963_ = ~new_n7950_;
  assign new_n1964_ = ~new_n2854_ | ~new_n1952_;
  assign new_n1965_ = ~new_n1950_ | ~new_n3180_;
  assign new_n1966_ = ~new_n1950_ | ~new_n3189_;
  assign new_n1967_ = ~pi246 | ~new_n1945_;
  assign new_n1968_ = ~new_n3187_ | ~new_n1135_;
  assign new_n1969_ = ~new_n8049_ | ~new_n1953_;
  assign new_n1970_ = ~new_n8042_ | ~new_n1976_;
  assign new_n1971_ = ~new_n3245_ | ~new_n1132_;
  assign new_n1972_ = ~new_n1968_ | ~new_n3248_;
  assign new_n1973_ = ~pi247 | ~new_n1946_;
  assign new_n1974_ = ~new_n3186_ | ~new_n1135_;
  assign new_n1975_ = ~new_n8042_ | ~new_n1954_;
  assign new_n1976_ = ~new_n1969_ | ~new_n1975_;
  assign new_n1977_ = ~new_n3171_ | ~new_n1953_;
  assign new_n1978_ = ~new_n3303_ | ~new_n1132_;
  assign new_n1979_ = ~new_n1974_ | ~new_n3306_;
  assign new_n1980_ = ~new_n1974_ | ~new_n3308_;
  assign new_n1981_ = ~new_n1145_ | ~new_n1135_;
  assign new_n1982_ = ~new_n1142_ | ~new_n1132_;
  assign new_n1983_ = ~new_n1981_ | ~new_n3364_;
  assign new_n1984_ = ~pi244 | ~new_n1948_;
  assign new_n1985_ = ~new_n3183_ | ~new_n3178_;
  assign new_n1986_ = ~new_n8007_ | ~new_n1955_;
  assign new_n1987_ = ~new_n1147_ | ~new_n3172_;
  assign new_n1988_ = ~new_n1985_ | ~new_n3421_;
  assign new_n1989_ = ~new_n1985_ | ~new_n3423_;
  assign new_n1990_ = ~new_n3183_ | ~new_n3187_;
  assign new_n1991_ = ~new_n1147_ | ~new_n3245_;
  assign new_n1992_ = ~new_n1990_ | ~new_n3479_;
  assign new_n1993_ = ~new_n3183_ | ~new_n3186_;
  assign new_n1994_ = ~new_n1147_ | ~new_n3303_;
  assign new_n1995_ = ~new_n1993_ | ~new_n3536_;
  assign new_n1996_ = ~new_n1993_ | ~new_n3538_;
  assign new_n1997_ = ~new_n3183_ | ~new_n1145_;
  assign new_n1998_ = ~new_n1147_ | ~new_n1142_;
  assign new_n1999_ = ~new_n1997_ | ~new_n3594_;
  assign new_n2000_ = ~new_n1136_ | ~new_n3178_;
  assign new_n2001_ = ~new_n1131_ | ~new_n3173_;
  assign new_n2002_ = ~new_n2001_ | ~new_n1986_ | ~new_n3175_;
  assign new_n2003_ = ~new_n1156_ | ~new_n3172_;
  assign new_n2004_ = ~new_n2000_ | ~new_n1984_ | ~new_n3184_;
  assign new_n2005_ = ~new_n2000_ | ~new_n3650_;
  assign new_n2006_ = ~new_n2000_ | ~new_n3652_;
  assign new_n2007_ = ~new_n3187_ | ~new_n1136_;
  assign new_n2008_ = ~new_n1156_ | ~new_n3245_;
  assign new_n2009_ = ~new_n2007_ | ~new_n3707_;
  assign new_n2010_ = ~new_n3186_ | ~new_n1136_;
  assign new_n2011_ = ~new_n1156_ | ~new_n3303_;
  assign new_n2012_ = ~new_n2010_ | ~new_n3764_;
  assign new_n2013_ = ~new_n2010_ | ~new_n3766_;
  assign new_n2014_ = ~new_n1145_ | ~new_n1136_;
  assign new_n2015_ = ~new_n1156_ | ~new_n1142_;
  assign new_n2016_ = ~new_n2014_ | ~new_n3822_;
  assign new_n2017_ = ~new_n1167_ | ~new_n3178_;
  assign new_n2018_ = ~new_n1164_ | ~new_n3172_;
  assign new_n2019_ = ~new_n2017_ | ~new_n3879_;
  assign new_n2020_ = ~new_n2017_ | ~new_n3881_;
  assign new_n2021_ = ~new_n1167_ | ~new_n3187_;
  assign new_n2022_ = ~new_n1164_ | ~new_n3245_;
  assign new_n2023_ = ~new_n2021_ | ~new_n3937_;
  assign new_n2024_ = ~new_n1167_ | ~new_n3186_;
  assign new_n2025_ = ~new_n1164_ | ~new_n3303_;
  assign new_n2026_ = ~new_n2024_ | ~new_n3994_;
  assign new_n2027_ = ~new_n2024_ | ~new_n3996_;
  assign new_n2028_ = ~new_n1167_ | ~new_n1145_;
  assign new_n2029_ = ~new_n1164_ | ~new_n1142_;
  assign new_n2030_ = ~new_n2028_ | ~new_n4052_;
  assign new_n2031_ = ~pi476;
  assign new_n2032_ = ~new_n9223_;
  assign new_n2033_ = ~new_n1928_ | ~new_n1922_;
  assign new_n2034_ = ~new_n1928_ | ~new_n1915_;
  assign new_n2035_ = ~new_n2157_ | ~new_n2158_ | ~new_n2160_ | ~new_n2159_;
  assign new_n2036_ = ~new_n6273_ | ~new_n4135_ | ~new_n4134_;
  assign new_n2037_ = ~new_n3044_ | ~new_n1928_;
  assign new_n2038_ = ~new_n1262_ | ~new_n1921_;
  assign new_n2039_ = ~new_n3139_ | ~new_n3044_ | ~new_n6139_;
  assign new_n2040_ = ~new_n2386_ | ~new_n2892_;
  assign new_n2041_ = ~new_n3044_ | ~new_n3139_ | ~new_n1262_ | ~new_n6139_ | ~new_n3122_;
  assign new_n2042_ = ~new_n3045_ | ~new_n3094_ | ~new_n2816_ | ~new_n1262_ | ~new_n3105_;
  assign new_n2043_ = ~new_n2879_ | ~new_n2844_ | ~new_n3122_;
  assign new_n2044_ = ~new_n1106_ | ~new_n1104_;
  assign new_n2045_ = ~new_n2088_ | ~new_n4155_;
  assign new_n2046_ = ~new_n1913_ | ~new_n1919_;
  assign new_n2047_ = ~new_n8260_;
  assign new_n2048_ = ~new_n4181_ | ~new_n2887_ | ~new_n1944_;
  assign new_n2049_ = ~new_n1928_ | ~pi109 | ~new_n1922_;
  assign new_n2050_ = ~new_n1915_ | ~new_n1917_;
  assign new_n2051_ = ~new_n1921_ | ~new_n2035_;
  assign new_n2052_ = ~new_n1084_ | ~new_n1938_;
  assign new_n2053_ = ~new_n3105_ | ~new_n2035_;
  assign new_n2054_ = ~new_n2898_ | ~new_n1922_;
  assign new_n2055_ = ~new_n2835_ | ~new_n1109_;
  assign new_n2056_ = ~pi107 | ~new_n1915_;
  assign new_n2057_ = ~pi439;
  assign new_n2058_ = ~new_n2401_ | ~new_n4207_;
  assign new_n2059_ = ~new_n3045_ | ~new_n2818_;
  assign new_n2060_ = ~new_n2508_ | ~new_n2893_;
  assign new_n2061_ = ~new_n4699_ | ~new_n4698_;
  assign new_n2062_ = ~pi109 | ~new_n3139_;
  assign new_n2063_ = ~new_n3044_ | ~new_n6139_;
  assign new_n2064_ = ~new_n2851_ | ~new_n3122_;
  assign new_n2065_ = ~new_n2839_ | ~new_n1088_;
  assign new_n2066_ = ~new_n2855_ | ~pi109;
  assign new_n2067_ = ~new_n3148_ | ~new_n2035_;
  assign new_n2068_ = ~new_n2880_ | ~new_n4798_;
  assign new_n2069_ = ~pi109 | ~new_n2861_;
  assign new_n2070_ = ~new_n2880_ | ~new_n4909_;
  assign new_n2071_ = ~new_n1109_ | ~new_n2531_ | ~pi109 | ~new_n2894_;
  assign new_n2072_ = ~new_n2511_ | ~new_n1104_;
  assign new_n2073_ = ~pi438;
  assign new_n2074_ = ~new_n7786_;
  assign new_n2075_ = ~new_n2873_ | ~new_n2532_;
  assign new_n2076_ = ~new_n2854_ | ~new_n1906_;
  assign new_n2077_ = ~new_n2597_ | ~new_n2600_ | ~new_n2607_ | ~new_n2603_;
  assign new_n2078_ = ~new_n2851_ | ~new_n1915_;
  assign new_n2079_ = ~pi482;
  assign new_n2080_ = ~pi484;
  assign new_n2081_ = ~new_n1104_ | ~new_n3143_;
  assign new_n2082_ = ~new_n1911_ | ~new_n4127_;
  assign new_n2083_ = ~new_n3094_ | ~pi107;
  assign new_n2084_ = ~pi478 | ~new_n1907_;
  assign new_n2085_ = ~new_n1878_;
  assign new_n2086_ = ~new_n4124_ | ~new_n4123_;
  assign new_n2087_ = ~new_n1107_ | ~new_n2085_;
  assign new_n2088_ = ~pi242 | ~pi241 | ~new_n1908_;
  assign new_n2089_ = ~new_n1918_ | ~new_n5709_;
  assign new_n2090_ = ~new_n2842_ | ~new_n2879_;
  assign new_n2091_ = ~new_n2895_ | ~new_n2876_ | ~new_n3045_;
  assign new_n2092_ = ~new_n2895_ | ~new_n2876_ | ~new_n1922_;
  assign new_n2093_ = ~new_n3122_ | ~new_n3141_;
  assign new_n2094_ = ~new_n2722_ | ~new_n2720_ | ~new_n2719_ | ~new_n5738_;
  assign new_n2095_ = ~new_n2899_ | ~new_n2911_;
  assign new_n2096_ = ~new_n2828_ | ~new_n1912_;
  assign new_n2097_ = ~pi109 | ~new_n1262_;
  assign new_n2098_ = ~new_n6337_ | ~new_n6336_;
  assign new_n2099_ = ~new_n6340_ | ~new_n6339_;
  assign new_n2100_ = ~new_n6364_ | ~new_n6363_;
  assign new_n2101_ = ~new_n6434_ | ~new_n6433_;
  assign po070 = ~new_n6279_ | ~new_n6278_;
  assign po071 = ~new_n6281_ | ~new_n6280_;
  assign po072 = ~new_n6283_ | ~new_n6282_;
  assign po073 = ~new_n6285_ | ~new_n6284_;
  assign new_n2106_ = ~new_n6294_ | ~new_n6293_;
  assign new_n2107_ = new_n1899_ & new_n2824_;
  assign po107 = ~new_n6297_ | ~new_n6296_;
  assign po108 = ~new_n6299_ | ~new_n6298_;
  assign po139 = ~new_n6331_ | ~new_n6330_;
  assign new_n2111_ = new_n7941_ & new_n1084_ & new_n2860_;
  assign po271 = ~new_n6347_ | ~new_n6346_;
  assign po272 = ~new_n6354_ | ~new_n6353_;
  assign new_n2114_ = ~new_n6356_ | ~new_n6355_;
  assign new_n2115_ = ~new_n6359_ | ~new_n6358_;
  assign po273 = ~new_n6367_ | ~new_n6366_;
  assign po274 = ~new_n6369_ | ~new_n6368_;
  assign po275 = ~new_n6373_ | ~new_n6372_;
  assign po277 = ~new_n6375_ | ~new_n6374_;
  assign po278 = ~new_n6380_ | ~new_n6379_;
  assign po279 = ~new_n6382_ | ~new_n6381_;
  assign po280 = ~new_n6384_ | ~new_n6383_;
  assign new_n2123_ = new_n7169_ & new_n3094_;
  assign new_n2124_ = ~pi075 & ~pi440;
  assign po505 = ~new_n6400_ | ~new_n6399_;
  assign po507 = ~new_n6404_ | ~new_n6403_;
  assign po508 = ~new_n6406_ | ~new_n6405_;
  assign po510 = ~new_n6408_ | ~new_n6407_;
  assign po512 = ~new_n6412_ | ~new_n6411_;
  assign po514 = ~new_n6416_ | ~new_n6415_;
  assign po517 = ~new_n6418_ | ~new_n6417_;
  assign new_n2132_ = new_n7941_ & new_n2860_;
  assign new_n2133_ = ~new_n6420_ | ~new_n6419_;
  assign new_n2134_ = ~new_n6422_ | ~new_n6421_;
  assign new_n2135_ = ~new_n6424_ | ~new_n6423_;
  assign new_n2136_ = ~new_n6426_ | ~new_n6425_;
  assign new_n2137_ = ~new_n6428_ | ~new_n6427_;
  assign new_n2138_ = pi072 & pi035;
  assign new_n2139_ = new_n3013_ & new_n1896_;
  assign new_n2140_ = new_n3015_ & new_n1894_;
  assign new_n2141_ = pi479 & pi073;
  assign new_n2142_ = ~pi240 & ~pi239;
  assign new_n2143_ = pi242 & pi241;
  assign new_n2144_ = ~pi241 & ~pi239;
  assign new_n2145_ = pi242 & pi240;
  assign new_n2146_ = ~pi242 & ~pi239;
  assign new_n2147_ = pi241 & pi240;
  assign new_n2148_ = ~pi241 & ~pi240;
  assign new_n2149_ = pi239 & pi242;
  assign new_n2150_ = ~pi242 & ~pi240;
  assign new_n2151_ = pi239 & pi241;
  assign new_n2152_ = pi239 & pi240;
  assign new_n2153_ = new_n3028_ & new_n3029_ & new_n3031_ & new_n3030_;
  assign new_n2154_ = new_n3032_ & new_n3033_ & new_n3035_ & new_n3034_;
  assign new_n2155_ = new_n3036_ & new_n3037_ & new_n3039_ & new_n3038_;
  assign new_n2156_ = new_n3040_ & new_n3041_ & new_n3043_ & new_n3042_;
  assign new_n2157_ = new_n3078_ & new_n3079_ & new_n3081_ & new_n3080_;
  assign new_n2158_ = new_n3082_ & new_n3083_ & new_n3085_ & new_n3084_;
  assign new_n2159_ = new_n3086_ & new_n3087_ & new_n3089_ & new_n3088_;
  assign new_n2160_ = new_n3090_ & new_n3091_ & new_n3093_ & new_n3092_;
  assign new_n2161_ = new_n3061_ & new_n3062_ & new_n3064_ & new_n3063_;
  assign new_n2162_ = new_n3065_ & new_n3066_ & new_n3068_ & new_n3067_;
  assign new_n2163_ = new_n3069_ & new_n3070_ & new_n3072_ & new_n3071_;
  assign new_n2164_ = new_n3073_ & new_n3074_ & new_n3076_ & new_n3075_;
  assign new_n2165_ = ~pi241 & ~pi239;
  assign new_n2166_ = pi192 & pi242;
  assign new_n2167_ = ~pi242 & ~pi239;
  assign new_n2168_ = pi184 & pi241;
  assign new_n2169_ = pi239 & pi168;
  assign new_n2170_ = ~pi242 & ~pi240;
  assign new_n2171_ = pi152 & pi239;
  assign new_n2172_ = pi136 & pi239;
  assign new_n2173_ = ~pi241 & ~pi240;
  assign new_n2174_ = pi160 & pi242;
  assign new_n2175_ = new_n3046_ & new_n3047_ & new_n3049_ & new_n3048_;
  assign new_n2176_ = new_n3050_ & new_n3051_ & new_n3053_ & new_n3052_;
  assign new_n2177_ = new_n3054_ & new_n3055_ & new_n3057_ & new_n3056_;
  assign new_n2178_ = new_n3059_ & new_n3058_;
  assign new_n2179_ = ~pi240 & ~pi239;
  assign new_n2180_ = pi207 & pi242;
  assign new_n2181_ = new_n3095_ & new_n3096_ & new_n3098_ & new_n3097_;
  assign new_n2182_ = new_n3101_ & new_n3100_ & new_n3099_;
  assign new_n2183_ = new_n3104_ & new_n3103_ & new_n3102_;
  assign new_n2184_ = new_n6320_ & new_n6321_ & new_n6323_ & new_n6322_;
  assign new_n2185_ = ~pi240 & ~pi239;
  assign new_n2186_ = pi225 & pi242;
  assign new_n2187_ = ~pi242 & ~pi241;
  assign new_n2188_ = pi201 & pi240;
  assign new_n2189_ = ~pi242 & ~pi241;
  assign new_n2190_ = pi137 & pi240;
  assign new_n2191_ = pi242 & pi240;
  assign new_n2192_ = pi129 & pi239;
  assign new_n2193_ = ~pi242 & ~pi239;
  assign new_n2194_ = pi185 & pi240;
  assign new_n2195_ = pi241 & pi240;
  assign new_n2196_ = pi121 & pi239;
  assign new_n2197_ = ~pi241 & ~pi240;
  assign new_n2198_ = pi161 & pi239;
  assign new_n2199_ = new_n6300_ & new_n6301_ & new_n6303_ & new_n6302_;
  assign new_n2200_ = new_n6304_ & new_n6305_ & new_n6307_ & new_n6306_;
  assign new_n2201_ = new_n6308_ & new_n6309_ & new_n6311_ & new_n6310_;
  assign new_n2202_ = new_n6312_ & new_n6313_ & new_n6315_ & new_n6314_;
  assign new_n2203_ = new_n6139_ & new_n2035_ & new_n1927_;
  assign new_n2204_ = new_n3045_ & new_n3105_ & new_n1262_;
  assign new_n2205_ = new_n3123_ & new_n3124_ & new_n3126_ & new_n3125_;
  assign new_n2206_ = new_n3127_ & new_n3128_ & new_n3130_ & new_n3129_;
  assign new_n2207_ = new_n3131_ & new_n3132_ & new_n3134_ & new_n3133_;
  assign new_n2208_ = new_n3135_ & new_n3136_ & new_n3138_ & new_n3137_;
  assign new_n2209_ = new_n3106_ & new_n3107_ & new_n3109_ & new_n3108_;
  assign new_n2210_ = new_n3110_ & new_n3111_ & new_n3113_ & new_n3112_;
  assign new_n2211_ = new_n3114_ & new_n3115_ & new_n3117_ & new_n3116_;
  assign new_n2212_ = new_n3118_ & new_n3119_ & new_n3121_ & new_n3120_;
  assign new_n2213_ = new_n3022_ & new_n2853_;
  assign new_n2214_ = new_n3061_ & new_n3062_ & new_n3064_ & new_n3063_;
  assign new_n2215_ = new_n3065_ & new_n3066_ & new_n3068_ & new_n3067_;
  assign new_n2216_ = new_n3069_ & new_n3070_ & new_n3072_ & new_n3071_;
  assign new_n2217_ = new_n3073_ & new_n3074_ & new_n3076_ & new_n3075_;
  assign new_n2218_ = new_n3046_ & new_n3047_ & new_n3049_ & new_n3048_;
  assign new_n2219_ = new_n3050_ & new_n3051_ & new_n3053_ & new_n3052_;
  assign new_n2220_ = new_n3054_ & new_n3055_ & new_n3057_ & new_n3056_;
  assign new_n2221_ = new_n3059_ & new_n3058_;
  assign new_n2222_ = new_n3044_ & new_n2816_;
  assign new_n2223_ = new_n2894_ & new_n1927_;
  assign new_n2224_ = new_n6139_ & new_n3045_ & new_n1928_ & new_n1927_;
  assign new_n2225_ = new_n2862_ & new_n2044_;
  assign new_n2226_ = pi107 & new_n6248_;
  assign new_n2227_ = new_n3160_ & new_n1941_;
  assign new_n2228_ = new_n1084_ & new_n1901_;
  assign new_n2229_ = pi106 & pi109;
  assign new_n2230_ = new_n2891_ & new_n2886_;
  assign new_n2231_ = new_n2230_ & new_n3168_;
  assign new_n2232_ = new_n2869_ & new_n3197_ & new_n3198_;
  assign new_n2233_ = new_n3207_ & new_n3206_ & new_n3205_;
  assign new_n2234_ = new_n3212_ & new_n3211_ & new_n3210_;
  assign new_n2235_ = new_n3217_ & new_n3216_ & new_n3215_;
  assign new_n2236_ = new_n3222_ & new_n3221_ & new_n3220_;
  assign new_n2237_ = new_n3227_ & new_n3226_ & new_n3225_;
  assign new_n2238_ = new_n3232_ & new_n3231_ & new_n3230_;
  assign new_n2239_ = new_n3237_ & new_n3236_ & new_n3235_;
  assign new_n2240_ = new_n3242_ & new_n3241_ & new_n3240_;
  assign new_n2241_ = new_n2869_ & new_n3255_ & new_n3256_;
  assign new_n2242_ = new_n3265_ & new_n3264_ & new_n3263_;
  assign new_n2243_ = new_n3270_ & new_n3269_ & new_n3268_;
  assign new_n2244_ = new_n3275_ & new_n3274_ & new_n3273_;
  assign new_n2245_ = new_n3280_ & new_n3279_ & new_n3278_;
  assign new_n2246_ = new_n3285_ & new_n3284_ & new_n3283_;
  assign new_n2247_ = new_n3290_ & new_n3289_ & new_n3288_;
  assign new_n2248_ = new_n3295_ & new_n3294_ & new_n3293_;
  assign new_n2249_ = new_n3300_ & new_n3299_ & new_n3298_;
  assign new_n2250_ = new_n2869_ & new_n3314_ & new_n3315_;
  assign new_n2251_ = new_n3324_ & new_n3323_ & new_n3322_;
  assign new_n2252_ = new_n3329_ & new_n3328_ & new_n3327_;
  assign new_n2253_ = new_n3334_ & new_n3333_ & new_n3332_;
  assign new_n2254_ = new_n3339_ & new_n3338_ & new_n3337_;
  assign new_n2255_ = new_n3344_ & new_n3343_ & new_n3342_;
  assign new_n2256_ = new_n3349_ & new_n3348_ & new_n3347_;
  assign new_n2257_ = new_n3354_ & new_n3353_ & new_n3352_;
  assign new_n2258_ = new_n3359_ & new_n3358_ & new_n3357_;
  assign new_n2259_ = new_n2869_ & new_n3371_ & new_n3372_;
  assign new_n2260_ = new_n3381_ & new_n3380_ & new_n3379_;
  assign new_n2261_ = new_n3386_ & new_n3385_ & new_n3384_;
  assign new_n2262_ = new_n3391_ & new_n3390_ & new_n3389_;
  assign new_n2263_ = new_n3396_ & new_n3395_ & new_n3394_;
  assign new_n2264_ = new_n3401_ & new_n3400_ & new_n3399_;
  assign new_n2265_ = new_n3406_ & new_n3405_ & new_n3404_;
  assign new_n2266_ = new_n3411_ & new_n3410_ & new_n3409_;
  assign new_n2267_ = new_n3416_ & new_n3415_ & new_n3414_;
  assign new_n2268_ = new_n2869_ & new_n3429_ & new_n3430_;
  assign new_n2269_ = new_n3439_ & new_n3438_ & new_n3437_;
  assign new_n2270_ = new_n3444_ & new_n3443_ & new_n3442_;
  assign new_n2271_ = new_n3449_ & new_n3448_ & new_n3447_;
  assign new_n2272_ = new_n3454_ & new_n3453_ & new_n3452_;
  assign new_n2273_ = new_n3459_ & new_n3458_ & new_n3457_;
  assign new_n2274_ = new_n3464_ & new_n3463_ & new_n3462_;
  assign new_n2275_ = new_n3469_ & new_n3468_ & new_n3467_;
  assign new_n2276_ = new_n3474_ & new_n3473_ & new_n3472_;
  assign new_n2277_ = new_n2869_ & new_n3486_ & new_n3487_;
  assign new_n2278_ = new_n3496_ & new_n3495_ & new_n3494_;
  assign new_n2279_ = new_n3501_ & new_n3500_ & new_n3499_;
  assign new_n2280_ = new_n3506_ & new_n3505_ & new_n3504_;
  assign new_n2281_ = new_n3511_ & new_n3510_ & new_n3509_;
  assign new_n2282_ = new_n3516_ & new_n3515_ & new_n3514_;
  assign new_n2283_ = new_n3521_ & new_n3520_ & new_n3519_;
  assign new_n2284_ = new_n3526_ & new_n3525_ & new_n3524_;
  assign new_n2285_ = new_n3531_ & new_n3530_ & new_n3529_;
  assign new_n2286_ = new_n2869_ & new_n3544_ & new_n3545_;
  assign new_n2287_ = new_n3554_ & new_n3553_ & new_n3552_;
  assign new_n2288_ = new_n3559_ & new_n3558_ & new_n3557_;
  assign new_n2289_ = new_n3564_ & new_n3563_ & new_n3562_;
  assign new_n2290_ = new_n3569_ & new_n3568_ & new_n3567_;
  assign new_n2291_ = new_n3574_ & new_n3573_ & new_n3572_;
  assign new_n2292_ = new_n3579_ & new_n3578_ & new_n3577_;
  assign new_n2293_ = new_n3584_ & new_n3583_ & new_n3582_;
  assign new_n2294_ = new_n3589_ & new_n3588_ & new_n3587_;
  assign new_n2295_ = new_n2869_ & new_n3601_ & new_n3602_;
  assign new_n2296_ = new_n3611_ & new_n3610_ & new_n3609_;
  assign new_n2297_ = new_n3616_ & new_n3615_ & new_n3614_;
  assign new_n2298_ = new_n3621_ & new_n3620_ & new_n3619_;
  assign new_n2299_ = new_n3626_ & new_n3625_ & new_n3624_;
  assign new_n2300_ = new_n3631_ & new_n3630_ & new_n3629_;
  assign new_n2301_ = new_n3636_ & new_n3635_ & new_n3634_;
  assign new_n2302_ = new_n3641_ & new_n3640_ & new_n3639_;
  assign new_n2303_ = new_n3646_ & new_n3645_ & new_n3644_;
  assign new_n2304_ = new_n2869_ & new_n3657_ & new_n3658_;
  assign new_n2305_ = new_n3667_ & new_n3666_ & new_n3665_;
  assign new_n2306_ = new_n3672_ & new_n3671_ & new_n3670_;
  assign new_n2307_ = new_n3677_ & new_n3676_ & new_n3675_;
  assign new_n2308_ = new_n3682_ & new_n3681_ & new_n3680_;
  assign new_n2309_ = new_n3687_ & new_n3686_ & new_n3685_;
  assign new_n2310_ = new_n3692_ & new_n3691_ & new_n3690_;
  assign new_n2311_ = new_n3697_ & new_n3696_ & new_n3695_;
  assign new_n2312_ = new_n3702_ & new_n3701_ & new_n3700_;
  assign new_n2313_ = new_n2869_ & new_n3714_ & new_n3715_;
  assign new_n2314_ = new_n3724_ & new_n3723_ & new_n3722_;
  assign new_n2315_ = new_n3729_ & new_n3728_ & new_n3727_;
  assign new_n2316_ = new_n3734_ & new_n3733_ & new_n3732_;
  assign new_n2317_ = new_n3739_ & new_n3738_ & new_n3737_;
  assign new_n2318_ = new_n3744_ & new_n3743_ & new_n3742_;
  assign new_n2319_ = new_n3749_ & new_n3748_ & new_n3747_;
  assign new_n2320_ = new_n3754_ & new_n3753_ & new_n3752_;
  assign new_n2321_ = new_n3759_ & new_n3758_ & new_n3757_;
  assign new_n2322_ = new_n2869_ & new_n3772_ & new_n3773_;
  assign new_n2323_ = new_n3782_ & new_n3781_ & new_n3780_;
  assign new_n2324_ = new_n3787_ & new_n3786_ & new_n3785_;
  assign new_n2325_ = new_n3792_ & new_n3791_ & new_n3790_;
  assign new_n2326_ = new_n3797_ & new_n3796_ & new_n3795_;
  assign new_n2327_ = new_n3802_ & new_n3801_ & new_n3800_;
  assign new_n2328_ = new_n3807_ & new_n3806_ & new_n3805_;
  assign new_n2329_ = new_n3812_ & new_n3811_ & new_n3810_;
  assign new_n2330_ = new_n3817_ & new_n3816_ & new_n3815_;
  assign new_n2331_ = new_n2869_ & new_n3829_ & new_n3830_;
  assign new_n2332_ = new_n3839_ & new_n3838_ & new_n3837_;
  assign new_n2333_ = new_n3844_ & new_n3843_ & new_n3842_;
  assign new_n2334_ = new_n3849_ & new_n3848_ & new_n3847_;
  assign new_n2335_ = new_n3854_ & new_n3853_ & new_n3852_;
  assign new_n2336_ = new_n3859_ & new_n3858_ & new_n3857_;
  assign new_n2337_ = new_n3864_ & new_n3863_ & new_n3862_;
  assign new_n2338_ = new_n3869_ & new_n3868_ & new_n3867_;
  assign new_n2339_ = new_n3874_ & new_n3873_ & new_n3872_;
  assign new_n2340_ = new_n2869_ & new_n3887_ & new_n3888_;
  assign new_n2341_ = new_n3897_ & new_n3896_ & new_n3895_;
  assign new_n2342_ = new_n3902_ & new_n3901_ & new_n3900_;
  assign new_n2343_ = new_n3907_ & new_n3906_ & new_n3905_;
  assign new_n2344_ = new_n3912_ & new_n3911_ & new_n3910_;
  assign new_n2345_ = new_n3917_ & new_n3916_ & new_n3915_;
  assign new_n2346_ = new_n3922_ & new_n3921_ & new_n3920_;
  assign new_n2347_ = new_n3927_ & new_n3926_ & new_n3925_;
  assign new_n2348_ = new_n3932_ & new_n3931_ & new_n3930_;
  assign new_n2349_ = new_n2869_ & new_n3944_ & new_n3945_;
  assign new_n2350_ = new_n3954_ & new_n3953_ & new_n3952_;
  assign new_n2351_ = new_n3959_ & new_n3958_ & new_n3957_;
  assign new_n2352_ = new_n3964_ & new_n3963_ & new_n3962_;
  assign new_n2353_ = new_n3969_ & new_n3968_ & new_n3967_;
  assign new_n2354_ = new_n3974_ & new_n3973_ & new_n3972_;
  assign new_n2355_ = new_n3979_ & new_n3978_ & new_n3977_;
  assign new_n2356_ = new_n3984_ & new_n3983_ & new_n3982_;
  assign new_n2357_ = new_n3989_ & new_n3988_ & new_n3987_;
  assign new_n2358_ = new_n2869_ & new_n4002_ & new_n4003_;
  assign new_n2359_ = new_n4012_ & new_n4011_ & new_n4010_;
  assign new_n2360_ = new_n4017_ & new_n4016_ & new_n4015_;
  assign new_n2361_ = new_n4022_ & new_n4021_ & new_n4020_;
  assign new_n2362_ = new_n4027_ & new_n4026_ & new_n4025_;
  assign new_n2363_ = new_n4032_ & new_n4031_ & new_n4030_;
  assign new_n2364_ = new_n4037_ & new_n4036_ & new_n4035_;
  assign new_n2365_ = new_n4042_ & new_n4041_ & new_n4040_;
  assign new_n2366_ = new_n4047_ & new_n4046_ & new_n4045_;
  assign new_n2367_ = new_n2869_ & new_n4059_ & new_n4060_;
  assign new_n2368_ = new_n4069_ & new_n4068_ & new_n4067_;
  assign new_n2369_ = new_n4074_ & new_n4073_ & new_n4072_;
  assign new_n2370_ = new_n4079_ & new_n4078_ & new_n4077_;
  assign new_n2371_ = new_n4084_ & new_n4083_ & new_n4082_;
  assign new_n2372_ = new_n4088_ & new_n4087_ & new_n4086_;
  assign new_n2373_ = new_n4093_ & new_n4092_ & new_n4091_;
  assign new_n2374_ = new_n4098_ & new_n4097_ & new_n4096_;
  assign new_n2375_ = new_n4103_ & new_n4102_ & new_n4101_;
  assign new_n2376_ = pi476 & pi109;
  assign new_n2377_ = new_n3139_ & new_n3044_;
  assign new_n2378_ = new_n3142_ & new_n1901_;
  assign new_n2379_ = new_n2855_ & new_n1901_;
  assign new_n2380_ = new_n6141_ & new_n2862_;
  assign new_n2381_ = new_n4116_ & new_n4117_;
  assign new_n2382_ = new_n2381_ & new_n4115_;
  assign new_n2383_ = new_n2382_ & new_n1175_;
  assign new_n2384_ = new_n4120_ & new_n2887_;
  assign new_n2385_ = new_n4131_ & new_n4130_;
  assign new_n2386_ = new_n3094_ & new_n3045_;
  assign new_n2387_ = new_n4141_ & new_n2037_;
  assign new_n2388_ = new_n4143_ & new_n4142_;
  assign new_n2389_ = new_n2388_ & new_n2387_ & new_n4145_ & new_n6272_;
  assign new_n2390_ = new_n2908_ & new_n2041_;
  assign new_n2391_ = new_n1923_ & new_n1177_ & new_n2390_ & new_n2055_ & new_n1932_;
  assign new_n2392_ = new_n2393_ & new_n4147_;
  assign new_n2393_ = new_n4150_ & new_n4149_;
  assign new_n2394_ = new_n4158_ & new_n6362_ & new_n6361_;
  assign new_n2395_ = new_n4169_ & new_n4167_;
  assign new_n2396_ = new_n4188_ & new_n4189_;
  assign new_n2397_ = new_n4192_ & new_n4193_;
  assign new_n2398_ = new_n4197_ & new_n4198_;
  assign new_n2399_ = new_n4203_ & new_n1901_;
  assign new_n2400_ = new_n1928_ & new_n2051_;
  assign new_n2401_ = new_n4208_ & new_n4206_;
  assign new_n2402_ = new_n4212_ & new_n2042_ & new_n2043_;
  assign new_n2403_ = new_n2402_ & new_n1177_ & new_n4213_;
  assign new_n2404_ = new_n2831_ & new_n1928_;
  assign new_n2405_ = new_n2092_ & new_n1932_ & new_n2862_;
  assign new_n2406_ = new_n4211_ & new_n6152_;
  assign new_n2407_ = new_n6153_ & pi107;
  assign new_n2408_ = new_n4216_ & new_n4215_;
  assign new_n2409_ = new_n4218_ & new_n4217_;
  assign new_n2410_ = new_n4220_ & new_n4221_;
  assign new_n2411_ = new_n2410_ & new_n4219_;
  assign new_n2412_ = new_n4223_ & new_n4222_;
  assign new_n2413_ = new_n4225_ & new_n4224_;
  assign new_n2414_ = new_n4227_ & new_n4228_;
  assign new_n2415_ = new_n2414_ & new_n4226_;
  assign new_n2416_ = new_n4230_ & new_n4229_;
  assign new_n2417_ = new_n4232_ & new_n4231_;
  assign new_n2418_ = new_n4234_ & new_n4235_;
  assign new_n2419_ = new_n2418_ & new_n4233_;
  assign new_n2420_ = new_n4239_ & new_n4237_ & new_n4236_;
  assign new_n2421_ = new_n4238_ & new_n2422_ & new_n4240_;
  assign new_n2422_ = new_n4241_ & new_n4242_;
  assign new_n2423_ = new_n4246_ & new_n4244_ & new_n4243_;
  assign new_n2424_ = new_n4248_ & new_n4249_;
  assign new_n2425_ = new_n2424_ & new_n4247_;
  assign new_n2426_ = new_n4253_ & new_n4251_ & new_n4250_;
  assign new_n2427_ = new_n4255_ & new_n4256_;
  assign new_n2428_ = new_n2427_ & new_n4254_;
  assign new_n2429_ = new_n4260_ & new_n4258_ & new_n4257_;
  assign new_n2430_ = new_n4262_ & new_n4263_;
  assign new_n2431_ = new_n2430_ & new_n4261_;
  assign new_n2432_ = new_n4267_ & new_n4265_ & new_n4264_;
  assign new_n2433_ = new_n4269_ & new_n4270_;
  assign new_n2434_ = new_n2433_ & new_n4268_;
  assign new_n2435_ = new_n4274_ & new_n4272_ & new_n4271_;
  assign new_n2436_ = new_n4276_ & new_n4277_;
  assign new_n2437_ = new_n2436_ & new_n4275_;
  assign new_n2438_ = new_n4281_ & new_n4279_ & new_n4278_;
  assign new_n2439_ = new_n4283_ & new_n4284_;
  assign new_n2440_ = new_n2439_ & new_n4282_;
  assign new_n2441_ = new_n4288_ & new_n4286_ & new_n4285_;
  assign new_n2442_ = new_n4290_ & new_n4291_;
  assign new_n2443_ = new_n2442_ & new_n4289_;
  assign new_n2444_ = new_n4295_ & new_n4293_ & new_n4292_;
  assign new_n2445_ = new_n4297_ & new_n4298_;
  assign new_n2446_ = new_n2445_ & new_n4296_;
  assign new_n2447_ = new_n4302_ & new_n4300_ & new_n4299_;
  assign new_n2448_ = new_n4304_ & new_n4305_;
  assign new_n2449_ = new_n2448_ & new_n4303_;
  assign new_n2450_ = new_n4307_ & new_n4309_;
  assign new_n2451_ = new_n4311_ & new_n4312_;
  assign new_n2452_ = new_n2451_ & new_n4310_;
  assign new_n2453_ = new_n4314_ & new_n4316_;
  assign new_n2454_ = new_n4318_ & new_n4319_;
  assign new_n2455_ = new_n2454_ & new_n4317_;
  assign new_n2456_ = new_n4321_ & new_n4323_;
  assign new_n2457_ = new_n4325_ & new_n4326_;
  assign new_n2458_ = new_n2457_ & new_n4324_;
  assign new_n2459_ = new_n4328_ & new_n4330_;
  assign new_n2460_ = new_n4332_ & new_n4333_;
  assign new_n2461_ = new_n2460_ & new_n4331_;
  assign new_n2462_ = new_n4335_ & new_n4337_;
  assign new_n2463_ = new_n4339_ & new_n4340_;
  assign new_n2464_ = new_n2463_ & new_n4338_;
  assign new_n2465_ = new_n4342_ & new_n4344_;
  assign new_n2466_ = new_n4346_ & new_n4347_;
  assign new_n2467_ = new_n2466_ & new_n4345_;
  assign new_n2468_ = new_n4349_ & new_n4351_;
  assign new_n2469_ = new_n4353_ & new_n4354_;
  assign new_n2470_ = new_n2469_ & new_n4352_;
  assign new_n2471_ = new_n4356_ & new_n4358_;
  assign new_n2472_ = new_n4360_ & new_n4361_;
  assign new_n2473_ = new_n2472_ & new_n4359_;
  assign new_n2474_ = new_n4363_ & new_n4365_;
  assign new_n2475_ = new_n4367_ & new_n4368_;
  assign new_n2476_ = new_n2475_ & new_n4366_;
  assign new_n2477_ = new_n4370_ & new_n4372_;
  assign new_n2478_ = new_n4374_ & new_n4375_;
  assign new_n2479_ = new_n2478_ & new_n4373_;
  assign new_n2480_ = new_n4377_ & new_n4379_;
  assign new_n2481_ = new_n4381_ & new_n4382_;
  assign new_n2482_ = new_n2481_ & new_n4380_;
  assign new_n2483_ = new_n4384_ & new_n4386_;
  assign new_n2484_ = new_n4388_ & new_n4389_;
  assign new_n2485_ = new_n2484_ & new_n4387_;
  assign new_n2486_ = new_n4391_ & new_n4393_;
  assign new_n2487_ = new_n4395_ & new_n4396_;
  assign new_n2488_ = new_n2487_ & new_n4394_;
  assign new_n2489_ = new_n4398_ & new_n4400_;
  assign new_n2490_ = new_n4402_ & new_n4403_;
  assign new_n2491_ = new_n2490_ & new_n4401_;
  assign new_n2492_ = new_n4405_ & new_n4407_;
  assign new_n2493_ = new_n4409_ & new_n4410_;
  assign new_n2494_ = new_n2493_ & new_n4408_;
  assign new_n2495_ = new_n4412_ & new_n4414_;
  assign new_n2496_ = new_n4416_ & new_n4417_;
  assign new_n2497_ = new_n2496_ & new_n4415_;
  assign new_n2498_ = new_n4419_ & new_n4421_;
  assign new_n2499_ = new_n4423_ & new_n4424_;
  assign new_n2500_ = new_n2499_ & new_n4422_;
  assign new_n2501_ = new_n4426_ & new_n4428_;
  assign new_n2502_ = new_n4430_ & new_n4431_;
  assign new_n2503_ = new_n2502_ & new_n4429_;
  assign new_n2504_ = new_n4433_ & new_n4435_;
  assign new_n2505_ = new_n4437_ & new_n4438_;
  assign new_n2506_ = new_n2505_ & new_n4436_;
  assign new_n2507_ = new_n6139_ & new_n1927_ & new_n1906_;
  assign new_n2508_ = new_n4439_ & new_n2052_;
  assign new_n2509_ = pi108 & pi478;
  assign new_n2510_ = new_n1025_ & new_n1928_;
  assign new_n2511_ = new_n1106_ & pi109;
  assign new_n2512_ = new_n2853_ & new_n1025_;
  assign new_n2513_ = new_n4750_ & new_n4751_;
  assign new_n2514_ = new_n4753_ & new_n4754_;
  assign new_n2515_ = new_n4756_ & new_n4757_;
  assign new_n2516_ = new_n4759_ & new_n4760_;
  assign new_n2517_ = new_n4762_ & new_n4763_;
  assign new_n2518_ = new_n4765_ & new_n4766_;
  assign new_n2519_ = new_n4768_ & new_n4769_;
  assign new_n2520_ = new_n4771_ & new_n4772_;
  assign new_n2521_ = new_n4774_ & new_n4775_;
  assign new_n2522_ = new_n4777_ & new_n4778_;
  assign new_n2523_ = new_n4780_ & new_n4781_;
  assign new_n2524_ = new_n4783_ & new_n4784_;
  assign new_n2525_ = new_n4786_ & new_n4787_;
  assign new_n2526_ = new_n4789_ & new_n4790_;
  assign new_n2527_ = new_n4792_ & new_n4793_;
  assign new_n2528_ = new_n4796_ & new_n4795_;
  assign new_n2529_ = new_n1262_ & new_n2035_;
  assign new_n2530_ = new_n6139_ & pi109 & new_n1915_;
  assign new_n2531_ = new_n3044_ & new_n2816_;
  assign new_n2532_ = new_n5007_ & new_n2886_ & new_n2889_;
  assign new_n2533_ = ~pi035 & ~pi478;
  assign new_n2534_ = new_n3139_ & new_n2831_;
  assign new_n2535_ = new_n5016_ & new_n5019_ & new_n5020_ & new_n5018_ & new_n5017_;
  assign new_n2536_ = new_n5024_ & new_n5027_ & new_n5028_ & new_n5026_ & new_n5025_;
  assign new_n2537_ = new_n5032_ & new_n5035_ & new_n5036_ & new_n5034_ & new_n5033_;
  assign new_n2538_ = new_n5040_ & new_n5043_ & new_n5044_ & new_n5042_ & new_n5041_;
  assign new_n2539_ = new_n5045_ & new_n2872_;
  assign new_n2540_ = new_n5051_ & new_n5052_ & new_n5050_ & new_n5049_;
  assign new_n2541_ = new_n5053_ & new_n2872_;
  assign new_n2542_ = new_n5056_ & new_n5059_ & new_n5060_ & new_n5058_ & new_n5057_;
  assign new_n2543_ = new_n5061_ & new_n2872_;
  assign new_n2544_ = new_n5066_ & new_n5067_ & new_n5064_;
  assign new_n2545_ = new_n5068_ & new_n2872_;
  assign new_n2546_ = new_n5073_ & new_n5074_ & new_n5071_;
  assign new_n2547_ = new_n5075_ & new_n2872_;
  assign new_n2548_ = new_n5080_ & new_n5081_ & new_n5078_;
  assign new_n2549_ = new_n5082_ & new_n2872_;
  assign new_n2550_ = new_n5087_ & new_n5088_ & new_n5085_;
  assign new_n2551_ = new_n5089_ & new_n2872_;
  assign new_n2552_ = new_n5094_ & new_n5095_ & new_n5092_;
  assign new_n2553_ = new_n5096_ & new_n2872_;
  assign new_n2554_ = new_n5101_ & new_n5102_ & new_n5099_;
  assign new_n2555_ = new_n5103_ & new_n2872_;
  assign new_n2556_ = new_n5108_ & new_n5109_ & new_n5106_;
  assign new_n2557_ = new_n5110_ & new_n2872_;
  assign new_n2558_ = new_n5115_ & new_n5116_ & new_n5113_;
  assign new_n2559_ = new_n5117_ & new_n2872_;
  assign new_n2560_ = new_n5122_ & new_n5123_ & new_n5120_;
  assign new_n2561_ = new_n5124_ & new_n2872_;
  assign new_n2562_ = new_n5129_ & new_n5130_ & new_n5127_;
  assign new_n2563_ = new_n5131_ & new_n2872_;
  assign new_n2564_ = new_n5136_ & new_n5137_ & new_n5134_;
  assign new_n2565_ = new_n2872_ & new_n5139_;
  assign new_n2566_ = new_n5143_ & new_n5144_ & new_n5141_;
  assign new_n2567_ = new_n2872_ & new_n5146_;
  assign new_n2568_ = new_n5150_ & new_n5151_ & new_n5148_;
  assign new_n2569_ = new_n2872_ & new_n5153_;
  assign new_n2570_ = new_n5157_ & new_n5158_ & new_n5155_;
  assign new_n2571_ = new_n5162_ & new_n5160_;
  assign new_n2572_ = new_n5164_ & new_n5165_;
  assign new_n2573_ = new_n5169_ & new_n5167_;
  assign new_n2574_ = new_n5171_ & new_n5172_;
  assign new_n2575_ = new_n5176_ & new_n5174_;
  assign new_n2576_ = new_n5178_ & new_n5179_;
  assign new_n2577_ = new_n5183_ & new_n5181_;
  assign new_n2578_ = new_n5185_ & new_n5186_;
  assign new_n2579_ = new_n5190_ & new_n5188_;
  assign new_n2580_ = new_n5192_ & new_n5193_;
  assign new_n2581_ = new_n5197_ & new_n5195_;
  assign new_n2582_ = new_n5199_ & new_n5200_;
  assign new_n2583_ = new_n5204_ & new_n5202_;
  assign new_n2584_ = new_n5206_ & new_n5207_;
  assign new_n2585_ = new_n5211_ & new_n5209_;
  assign new_n2586_ = new_n5213_ & new_n5214_;
  assign new_n2587_ = new_n5218_ & new_n5216_;
  assign new_n2588_ = new_n5220_ & new_n5221_;
  assign new_n2589_ = new_n5225_ & new_n5223_;
  assign new_n2590_ = new_n5227_ & new_n5228_;
  assign new_n2591_ = new_n5232_ & new_n5230_;
  assign new_n2592_ = new_n5234_ & new_n5235_;
  assign new_n2593_ = new_n5239_ & new_n5237_;
  assign new_n2594_ = new_n5241_ & new_n5242_;
  assign new_n2595_ = ~pi077 & ~pi079 & ~pi078 & ~pi076;
  assign new_n2596_ = ~pi081 & ~pi083 & ~pi082 & ~pi080;
  assign new_n2597_ = new_n2596_ & new_n2595_;
  assign new_n2598_ = ~pi085 & ~pi087 & ~pi086 & ~pi084;
  assign new_n2599_ = ~pi089 & ~pi091 & ~pi090 & ~pi088;
  assign new_n2600_ = new_n2599_ & new_n2598_;
  assign new_n2601_ = ~pi093 & ~pi095 & ~pi094 & ~pi092;
  assign new_n2602_ = ~pi097 & ~pi099 & ~pi098 & ~pi096;
  assign new_n2603_ = new_n2602_ & new_n2601_;
  assign new_n2604_ = ~pi100 & ~pi101;
  assign new_n2605_ = ~pi102 & ~pi103;
  assign new_n2606_ = ~pi104 & ~pi105;
  assign new_n2607_ = new_n2604_ & new_n2605_ & new_n2606_ & new_n5243_;
  assign new_n2608_ = ~pi075 & ~pi439 & ~pi074;
  assign new_n2609_ = pi107 & new_n1901_;
  assign new_n2610_ = new_n5253_ & new_n1942_;
  assign new_n2611_ = ~pi035 & ~pi109;
  assign new_n2612_ = new_n5247_ & new_n1951_ & new_n2052_;
  assign new_n2613_ = pi107 & new_n1931_;
  assign new_n2614_ = new_n2880_ & new_n2851_;
  assign new_n2615_ = new_n5263_ & new_n5264_ & new_n5266_ & new_n5265_;
  assign new_n2616_ = new_n5267_ & new_n5268_ & new_n5270_ & new_n5269_;
  assign new_n2617_ = new_n5271_ & new_n5272_ & new_n5274_ & new_n5273_;
  assign new_n2618_ = new_n5275_ & new_n5276_ & new_n5278_ & new_n5277_;
  assign new_n2619_ = new_n5279_ & new_n5280_ & new_n5282_ & new_n5281_;
  assign new_n2620_ = new_n5283_ & new_n5284_ & new_n5286_ & new_n5285_;
  assign new_n2621_ = new_n5287_ & new_n5288_ & new_n5290_ & new_n5289_;
  assign new_n2622_ = new_n5291_ & new_n5292_ & new_n5294_ & new_n5293_;
  assign new_n2623_ = new_n5295_ & new_n5296_ & new_n5298_ & new_n5297_;
  assign new_n2624_ = new_n5299_ & new_n5300_ & new_n5302_ & new_n5301_;
  assign new_n2625_ = new_n5303_ & new_n5304_ & new_n5306_ & new_n5305_;
  assign new_n2626_ = new_n5307_ & new_n5308_ & new_n5310_ & new_n5309_;
  assign new_n2627_ = new_n5311_ & new_n5312_ & new_n5314_ & new_n5313_;
  assign new_n2628_ = new_n5315_ & new_n5316_ & new_n5318_ & new_n5317_;
  assign new_n2629_ = new_n5319_ & new_n5320_ & new_n5322_ & new_n5321_;
  assign new_n2630_ = new_n5323_ & new_n5324_ & new_n6258_ & new_n5325_;
  assign new_n2631_ = new_n5326_ & new_n5327_ & new_n5329_ & new_n5328_;
  assign new_n2632_ = new_n5330_ & new_n5331_ & new_n5333_ & new_n5332_;
  assign new_n2633_ = new_n5334_ & new_n5335_ & new_n5337_ & new_n5336_;
  assign new_n2634_ = new_n5338_ & new_n5339_ & new_n5341_ & new_n5340_;
  assign new_n2635_ = new_n5342_ & new_n5343_ & new_n5345_ & new_n5344_;
  assign new_n2636_ = new_n5346_ & new_n5347_ & new_n5349_ & new_n5348_;
  assign new_n2637_ = new_n5350_ & new_n5351_ & new_n5353_ & new_n5352_;
  assign new_n2638_ = new_n5354_ & new_n5355_ & new_n5357_ & new_n5356_;
  assign new_n2639_ = new_n5358_ & new_n5359_ & new_n5361_ & new_n5360_;
  assign new_n2640_ = new_n5362_ & new_n5363_ & new_n5365_ & new_n5364_;
  assign new_n2641_ = new_n5366_ & new_n5367_ & new_n5369_ & new_n5368_;
  assign new_n2642_ = new_n5370_ & new_n5371_ & new_n5373_ & new_n5372_;
  assign new_n2643_ = new_n5374_ & new_n5375_ & new_n5377_ & new_n5376_;
  assign new_n2644_ = new_n5378_ & new_n5379_ & new_n5381_ & new_n5380_;
  assign new_n2645_ = new_n5382_ & new_n5383_ & new_n5385_ & new_n5384_;
  assign new_n2646_ = new_n5386_ & new_n5387_ & new_n5389_ & new_n5388_;
  assign new_n2647_ = new_n5394_ & new_n5393_;
  assign new_n2648_ = new_n5397_ & new_n5396_;
  assign new_n2649_ = new_n5400_ & new_n5399_;
  assign new_n2650_ = new_n5403_ & new_n5402_;
  assign new_n2651_ = new_n5405_ & new_n2652_;
  assign new_n2652_ = new_n5407_ & new_n5406_;
  assign new_n2653_ = new_n5409_ & new_n5410_;
  assign new_n2654_ = new_n5419_ & new_n5417_ & new_n5418_;
  assign new_n2655_ = new_n5421_ & new_n5422_;
  assign new_n2656_ = new_n5428_ & new_n5426_ & new_n5427_;
  assign new_n2657_ = new_n5432_ & new_n5430_ & new_n5431_;
  assign new_n2658_ = new_n5436_ & new_n5434_ & new_n5435_;
  assign new_n2659_ = new_n5440_ & new_n5438_ & new_n5439_;
  assign new_n2660_ = new_n5444_ & new_n5442_ & new_n5443_;
  assign new_n2661_ = new_n5448_ & new_n5446_ & new_n5447_;
  assign new_n2662_ = new_n5452_ & new_n5450_ & new_n5451_;
  assign new_n2663_ = new_n5456_ & new_n5454_ & new_n5455_;
  assign new_n2664_ = new_n5460_ & new_n5458_ & new_n5459_;
  assign new_n2665_ = new_n5464_ & new_n5462_ & new_n5463_;
  assign new_n2666_ = new_n5466_ & new_n5467_;
  assign new_n2667_ = new_n5473_ & new_n5471_ & new_n5472_;
  assign new_n2668_ = new_n5477_ & new_n5475_ & new_n5476_;
  assign new_n2669_ = new_n5481_ & new_n5479_ & new_n5480_;
  assign new_n2670_ = new_n5485_ & new_n5483_ & new_n5484_;
  assign new_n2671_ = new_n5503_ & new_n5502_;
  assign new_n2672_ = new_n5505_ & new_n5506_;
  assign new_n2673_ = new_n1927_ & new_n6139_ & new_n5533_;
  assign new_n2674_ = new_n5537_ & new_n5538_ & new_n5540_ & new_n5539_;
  assign new_n2675_ = new_n5541_ & new_n5542_ & new_n5544_ & new_n5543_;
  assign new_n2676_ = new_n5545_ & new_n5546_ & new_n5548_ & new_n5547_;
  assign new_n2677_ = new_n5549_ & new_n5550_ & new_n5552_ & new_n5551_;
  assign new_n2678_ = new_n5555_ & new_n5556_ & new_n5558_ & new_n5557_;
  assign new_n2679_ = new_n5559_ & new_n5560_ & new_n5562_ & new_n5561_;
  assign new_n2680_ = new_n5563_ & new_n5564_ & new_n5566_ & new_n5565_;
  assign new_n2681_ = new_n5567_ & new_n5568_ & new_n5570_ & new_n5569_;
  assign new_n2682_ = new_n5586_ & new_n5587_ & new_n5589_ & new_n5588_;
  assign new_n2683_ = new_n5590_ & new_n5591_ & new_n5593_ & new_n5592_;
  assign new_n2684_ = new_n5594_ & new_n5595_ & new_n5597_ & new_n5596_;
  assign new_n2685_ = new_n5598_ & new_n5599_ & new_n5601_ & new_n5600_;
  assign new_n2686_ = new_n5603_ & new_n5604_ & new_n5606_ & new_n5605_;
  assign new_n2687_ = new_n5607_ & new_n5608_ & new_n5610_ & new_n5609_;
  assign new_n2688_ = new_n5611_ & new_n5612_ & new_n5614_ & new_n5613_;
  assign new_n2689_ = new_n5615_ & new_n5616_ & new_n5618_ & new_n5617_;
  assign new_n2690_ = new_n5620_ & new_n5621_ & new_n5623_ & new_n5622_;
  assign new_n2691_ = new_n5624_ & new_n5625_ & new_n5627_ & new_n5626_;
  assign new_n2692_ = new_n5628_ & new_n5629_ & new_n5631_ & new_n5630_;
  assign new_n2693_ = new_n5632_ & new_n5633_ & new_n5635_ & new_n5634_;
  assign new_n2694_ = new_n5637_ & new_n5638_ & new_n5640_ & new_n5639_;
  assign new_n2695_ = new_n5641_ & new_n5642_ & new_n5644_ & new_n5643_;
  assign new_n2696_ = new_n5645_ & new_n5646_ & new_n5648_ & new_n5647_;
  assign new_n2697_ = new_n5649_ & new_n5650_ & new_n6259_ & new_n5651_;
  assign new_n2698_ = new_n5652_ & new_n5653_ & new_n5655_ & new_n5654_;
  assign new_n2699_ = new_n5656_ & new_n5657_ & new_n5659_ & new_n5658_;
  assign new_n2700_ = new_n5660_ & new_n5661_ & new_n5663_ & new_n5662_;
  assign new_n2701_ = new_n5664_ & new_n5665_ & new_n5667_ & new_n5666_;
  assign new_n2702_ = new_n5669_ & new_n5670_ & new_n5672_ & new_n5671_;
  assign new_n2703_ = new_n5673_ & new_n5674_ & new_n5676_ & new_n5675_;
  assign new_n2704_ = new_n5677_ & new_n5678_ & new_n5680_ & new_n5679_;
  assign new_n2705_ = new_n5681_ & new_n5682_ & new_n5684_ & new_n5683_;
  assign new_n2706_ = new_n5704_ & new_n2087_;
  assign new_n2707_ = pi109 & new_n5707_;
  assign new_n2708_ = new_n5711_ & new_n5712_ & new_n5714_ & new_n5713_;
  assign new_n2709_ = new_n5715_ & new_n5716_ & new_n5718_ & new_n5717_;
  assign new_n2710_ = new_n5719_ & new_n5720_ & new_n5722_ & new_n5721_;
  assign new_n2711_ = new_n5723_ & new_n5724_ & new_n5726_ & new_n5725_;
  assign new_n2712_ = new_n2901_ & pi109;
  assign new_n2713_ = new_n3046_ & new_n3048_ & new_n3050_ & new_n3049_;
  assign new_n2714_ = new_n3053_ & new_n3052_ & new_n3051_;
  assign new_n2715_ = new_n3054_ & new_n3055_ & new_n3057_ & new_n3056_;
  assign new_n2716_ = new_n3059_ & new_n3058_;
  assign new_n2717_ = new_n3045_ & new_n2035_;
  assign new_n2718_ = pi109 & new_n1928_;
  assign new_n2719_ = new_n5735_ & new_n5734_;
  assign new_n2720_ = new_n6118_ & new_n6117_ & new_n2078_;
  assign new_n2721_ = new_n6119_ & new_n6120_ & new_n6121_;
  assign new_n2722_ = new_n2721_ & new_n1263_ & new_n6122_;
  assign new_n2723_ = new_n5742_ & new_n5740_;
  assign new_n2724_ = new_n5743_ & new_n5744_ & new_n5746_ & new_n5745_;
  assign new_n2725_ = new_n5747_ & new_n5748_ & new_n5750_ & new_n5749_;
  assign new_n2726_ = new_n5751_ & new_n5752_ & new_n5754_ & new_n5753_;
  assign new_n2727_ = new_n5755_ & new_n5756_ & new_n5758_ & new_n5757_;
  assign new_n2728_ = new_n5760_ & new_n5761_ & new_n5763_ & new_n5762_;
  assign new_n2729_ = new_n5764_ & new_n5765_ & new_n5767_ & new_n5766_;
  assign new_n2730_ = new_n5768_ & new_n5769_ & new_n5771_ & new_n5770_;
  assign new_n2731_ = new_n5772_ & new_n5773_ & new_n5775_ & new_n5774_;
  assign new_n2732_ = new_n5777_ & new_n5778_ & new_n5780_ & new_n5779_;
  assign new_n2733_ = new_n5781_ & new_n5782_ & new_n5784_ & new_n5783_;
  assign new_n2734_ = new_n5785_ & new_n5786_ & new_n5788_ & new_n5787_;
  assign new_n2735_ = new_n5790_ & new_n5789_;
  assign new_n2736_ = new_n2735_ & new_n6262_ & new_n5791_;
  assign new_n2737_ = new_n5792_ & new_n5793_ & new_n5795_ & new_n5794_;
  assign new_n2738_ = new_n5796_ & new_n5797_ & new_n5799_ & new_n5798_;
  assign new_n2739_ = new_n5800_ & new_n5801_ & new_n5803_ & new_n5802_;
  assign new_n2740_ = new_n5804_ & new_n5805_ & new_n5807_ & new_n5806_;
  assign new_n2741_ = new_n5809_ & new_n5810_ & new_n5812_ & new_n5811_;
  assign new_n2742_ = new_n5813_ & new_n5814_ & new_n5816_ & new_n5815_;
  assign new_n2743_ = new_n5817_ & new_n5818_ & new_n5820_ & new_n5819_;
  assign new_n2744_ = new_n5821_ & new_n5822_ & new_n5824_ & new_n5823_;
  assign new_n2745_ = new_n5826_ & new_n5827_ & new_n5829_ & new_n5828_;
  assign new_n2746_ = new_n5830_ & new_n5831_ & new_n5833_ & new_n5832_;
  assign new_n2747_ = new_n5834_ & new_n5835_ & new_n5837_ & new_n5836_;
  assign new_n2748_ = new_n5838_ & new_n5839_ & new_n5841_ & new_n5840_;
  assign new_n2749_ = new_n5843_ & new_n5844_ & new_n5846_ & new_n5845_;
  assign new_n2750_ = new_n5847_ & new_n5848_ & new_n5850_ & new_n5849_;
  assign new_n2751_ = new_n5851_ & new_n5852_ & new_n5854_ & new_n5853_;
  assign new_n2752_ = new_n5855_ & new_n5856_ & new_n5858_ & new_n5857_;
  assign new_n2753_ = new_n5860_ & new_n1908_;
  assign new_n2754_ = new_n5861_ & new_n5860_;
  assign new_n2755_ = new_n5862_ & new_n1909_;
  assign new_n2756_ = new_n5734_ & new_n2071_;
  assign new_n2757_ = new_n5863_ & new_n5862_;
  assign new_n2758_ = new_n6118_ & new_n2757_ & new_n6117_;
  assign new_n2759_ = new_n2758_ & new_n2756_ & new_n5735_ & new_n2078_;
  assign new_n2760_ = new_n6119_ & new_n6121_ & new_n6131_ & new_n6125_;
  assign new_n2761_ = new_n6132_ & new_n6133_ & new_n6150_ & new_n6134_;
  assign new_n2762_ = new_n5735_ & new_n5734_;
  assign new_n2763_ = new_n6118_ & new_n6117_ & new_n2078_;
  assign new_n2764_ = new_n6119_ & new_n6120_ & new_n6121_;
  assign new_n2765_ = new_n2764_ & new_n1263_ & new_n1265_ & new_n6122_;
  assign new_n2766_ = new_n5865_ & new_n5866_ & new_n5868_ & new_n5867_;
  assign new_n2767_ = new_n5869_ & new_n5870_ & new_n5872_ & new_n5871_;
  assign new_n2768_ = new_n5873_ & new_n5874_ & new_n5876_ & new_n5875_;
  assign new_n2769_ = new_n5877_ & new_n5878_ & new_n5880_ & new_n5879_;
  assign new_n2770_ = new_n5882_ & new_n5883_ & new_n5885_ & new_n5884_;
  assign new_n2771_ = new_n5886_ & new_n5887_ & new_n5889_ & new_n5888_;
  assign new_n2772_ = new_n5890_ & new_n5891_ & new_n5893_ & new_n5892_;
  assign new_n2773_ = new_n5894_ & new_n5895_ & new_n5897_ & new_n5896_;
  assign new_n2774_ = new_n5899_ & new_n5900_ & new_n5902_ & new_n5901_;
  assign new_n2775_ = new_n5903_ & new_n5904_ & new_n5906_ & new_n5905_;
  assign new_n2776_ = new_n5907_ & new_n5908_ & new_n5910_ & new_n5909_;
  assign new_n2777_ = new_n5911_ & new_n5912_ & new_n5914_ & new_n5913_;
  assign new_n2778_ = new_n5916_ & new_n5917_ & new_n5919_ & new_n5918_;
  assign new_n2779_ = new_n5920_ & new_n5921_ & new_n5923_ & new_n5922_;
  assign new_n2780_ = new_n5924_ & new_n5925_ & new_n5927_ & new_n5926_;
  assign new_n2781_ = new_n5928_ & new_n5929_ & new_n6264_ & new_n5930_;
  assign new_n2782_ = new_n5931_ & new_n5932_ & new_n5934_ & new_n5933_;
  assign new_n2783_ = new_n5935_ & new_n5936_ & new_n5938_ & new_n5937_;
  assign new_n2784_ = new_n5939_ & new_n5940_ & new_n5942_ & new_n5941_;
  assign new_n2785_ = new_n5943_ & new_n5944_ & new_n5946_ & new_n5945_;
  assign new_n2786_ = new_n5948_ & new_n5949_ & new_n5951_ & new_n5950_;
  assign new_n2787_ = new_n5952_ & new_n5953_ & new_n5955_ & new_n5954_;
  assign new_n2788_ = new_n5956_ & new_n5957_ & new_n5959_ & new_n5958_;
  assign new_n2789_ = new_n5960_ & new_n5961_ & new_n5963_ & new_n5962_;
  assign new_n2790_ = new_n5965_ & new_n5966_ & new_n5968_ & new_n5967_;
  assign new_n2791_ = new_n5969_ & new_n5970_ & new_n5972_ & new_n5971_;
  assign new_n2792_ = new_n5973_ & new_n5974_ & new_n5976_ & new_n5975_;
  assign new_n2793_ = new_n5977_ & new_n5978_ & new_n5980_ & new_n5979_;
  assign new_n2794_ = new_n5982_ & new_n5983_ & new_n5985_ & new_n5984_;
  assign new_n2795_ = new_n5986_ & new_n5987_ & new_n5989_ & new_n5988_;
  assign new_n2796_ = new_n5990_ & new_n5991_ & new_n5993_ & new_n5992_;
  assign new_n2797_ = new_n5994_ & new_n5995_ & new_n5997_ & new_n5996_;
  assign new_n2798_ = new_n1928_ & new_n2063_;
  assign new_n2799_ = new_n1927_ & new_n2035_;
  assign new_n2800_ = new_n2908_ & new_n6002_ & new_n6003_;
  assign new_n2801_ = new_n2800_ & new_n6004_;
  assign new_n2802_ = pi109 & new_n1084_;
  assign new_n2803_ = new_n2802_ & new_n6005_;
  assign new_n2804_ = new_n1915_ & new_n2818_;
  assign new_n2805_ = pi109 & new_n2818_;
  assign new_n2806_ = new_n6014_ & pi109;
  assign new_n2807_ = new_n6016_ & new_n1260_;
  assign new_n2808_ = new_n6018_ & pi109;
  assign new_n2809_ = new_n6020_ & new_n1260_;
  assign new_n2810_ = new_n6027_ & new_n6028_;
  assign new_n2811_ = new_n2097_ & new_n6029_;
  assign new_n2812_ = new_n6032_ & new_n6034_ & new_n6033_;
  assign new_n2813_ = new_n6107_ & new_n6106_;
  assign new_n2814_ = new_n6110_ & new_n6109_;
  assign new_n2815_ = new_n6319_ & new_n6318_;
  assign new_n2816_ = ~new_n2214_ | ~new_n2215_ | ~new_n2217_ | ~new_n2216_;
  assign new_n2817_ = ~new_n2384_ | ~new_n4119_;
  assign new_n2818_ = ~new_n2218_ | ~new_n2219_ | ~new_n2220_ | ~new_n2221_ | ~new_n1264_;
  assign new_n2819_ = ~pi279;
  assign new_n2820_ = new_n6371_ & new_n6370_;
  assign new_n2821_ = new_n6390_ & new_n6389_;
  assign new_n2822_ = ~new_n1025_ | ~new_n1929_;
  assign new_n2823_ = ~new_n3153_ | ~new_n2035_;
  assign new_n2824_ = ~pi034;
  assign new_n2825_ = ~new_n2612_ | ~new_n2873_;
  assign new_n2826_ = ~new_n2873_ | ~new_n2076_;
  assign new_n2827_ = ~new_n2383_ | ~new_n6343_ | ~new_n6342_;
  assign new_n2828_ = ~pi240 | ~new_n1913_;
  assign new_n2829_ = ~new_n2096_;
  assign new_n2830_ = ~pi036 | ~new_n1901_;
  assign new_n2831_ = ~new_n2056_;
  assign new_n2832_ = ~new_n2084_;
  assign new_n2833_ = ~new_n2083_;
  assign new_n2834_ = ~new_n2037_;
  assign new_n2835_ = ~new_n1934_;
  assign new_n2836_ = ~new_n2093_;
  assign new_n2837_ = ~new_n2049_;
  assign new_n2838_ = ~new_n2078_;
  assign new_n2839_ = ~new_n2064_;
  assign new_n2840_ = ~new_n2910_ | ~new_n1915_;
  assign new_n2841_ = ~new_n3105_ | ~new_n1262_;
  assign new_n2842_ = ~new_n2040_;
  assign new_n2843_ = ~new_n2069_;
  assign new_n2844_ = ~new_n1933_;
  assign new_n2845_ = ~new_n2065_;
  assign new_n2846_ = ~new_n2066_;
  assign new_n2847_ = ~new_n2072_;
  assign new_n2848_ = ~new_n2052_;
  assign new_n2849_ = ~new_n2071_;
  assign new_n2850_ = ~new_n2842_ | ~new_n2530_ | ~new_n2834_;
  assign new_n2851_ = ~new_n2062_;
  assign new_n2852_ = ~new_n2087_;
  assign new_n2853_ = ~new_n1926_;
  assign new_n2854_ = ~new_n1951_;
  assign new_n2855_ = ~new_n2034_;
  assign new_n2856_ = ~new_n2090_;
  assign new_n2857_ = ~new_n2091_;
  assign new_n2858_ = ~new_n2092_;
  assign new_n2859_ = ~new_n2044_;
  assign new_n2860_ = ~new_n1932_;
  assign new_n2861_ = ~new_n1936_;
  assign new_n2862_ = ~new_n2223_ | ~new_n1088_;
  assign new_n2863_ = ~new_n2043_;
  assign new_n2864_ = ~new_n3094_ | ~new_n1915_;
  assign new_n2865_ = ~new_n2077_;
  assign new_n2866_ = ~new_n1893_;
  assign new_n2867_ = ~new_n2070_;
  assign new_n2868_ = ~new_n2068_;
  assign new_n2869_ = ~new_n1944_;
  assign new_n2870_ = ~new_n8666_;
  assign new_n2871_ = ~new_n1964_;
  assign new_n2872_ = ~new_n2900_ | ~new_n2075_;
  assign new_n2873_ = ~new_n2880_ | ~new_n6145_;
  assign new_n2874_ = ~new_n1019_ | ~new_n1916_;
  assign new_n2875_ = ~new_n1020_ | ~new_n3022_;
  assign new_n2876_ = ~new_n2051_;
  assign new_n2877_ = ~new_n1896_;
  assign new_n2878_ = ~new_n1894_;
  assign new_n2879_ = ~new_n2039_;
  assign new_n2880_ = ~new_n1941_;
  assign new_n2881_ = ~new_n2042_;
  assign new_n2882_ = ~new_n2823_;
  assign new_n2883_ = ~new_n2001_;
  assign new_n2884_ = ~new_n3122_ | ~new_n6026_;
  assign new_n2885_ = ~new_n2608_ | ~new_n2865_;
  assign new_n2886_ = ~new_n2229_ | ~new_n2906_;
  assign new_n2887_ = ~new_n2376_ | ~new_n1085_;
  assign new_n2888_ = ~new_n3009_ | ~new_n1902_;
  assign new_n2889_ = ~new_n1009_ | ~pi108 | ~new_n1938_;
  assign new_n2890_ = ~new_n1085_ | ~new_n2047_;
  assign new_n2891_ = ~pi109 | ~pi035 | ~new_n1907_;
  assign new_n2892_ = ~new_n2038_;
  assign new_n2893_ = ~new_n1105_ | ~new_n2507_ | ~new_n1108_ | ~new_n1010_;
  assign new_n2894_ = ~new_n1931_;
  assign new_n2895_ = ~new_n2041_;
  assign new_n2896_ = ~new_n2059_;
  assign new_n2897_ = ~new_n1943_;
  assign new_n2898_ = ~new_n2053_;
  assign new_n2899_ = ~new_n2063_;
  assign new_n2900_ = ~new_n2076_;
  assign new_n2901_ = ~new_n1935_;
  assign new_n2902_ = ~new_n2033_;
  assign new_n2903_ = ~new_n1898_;
  assign new_n2904_ = ~new_n1925_;
  assign new_n2905_ = ~new_n2050_;
  assign new_n2906_ = ~new_n1942_;
  assign new_n2907_ = ~new_n1930_;
  assign new_n2908_ = ~new_n2881_ | ~new_n3044_;
  assign new_n2909_ = ~new_n2055_;
  assign new_n2910_ = ~new_n2097_;
  assign new_n2911_ = ~new_n2054_;
  assign new_n2912_ = ~pi470 | ~new_n2878_;
  assign new_n2913_ = ~pi469 | ~new_n2877_;
  assign new_n2914_ = ~pi041 | ~new_n1893_;
  assign new_n2915_ = ~pi469 | ~new_n2878_;
  assign new_n2916_ = ~pi468 | ~new_n2877_;
  assign new_n2917_ = ~pi042 | ~new_n1893_;
  assign new_n2918_ = ~pi468 | ~new_n2878_;
  assign new_n2919_ = ~pi467 | ~new_n2877_;
  assign new_n2920_ = ~pi043 | ~new_n1893_;
  assign new_n2921_ = ~pi467 | ~new_n2878_;
  assign new_n2922_ = ~pi466 | ~new_n2877_;
  assign new_n2923_ = ~pi044 | ~new_n1893_;
  assign new_n2924_ = ~pi466 | ~new_n2878_;
  assign new_n2925_ = ~pi465 | ~new_n2877_;
  assign new_n2926_ = ~pi045 | ~new_n1893_;
  assign new_n2927_ = ~pi465 | ~new_n2878_;
  assign new_n2928_ = ~pi464 | ~new_n2877_;
  assign new_n2929_ = ~pi046 | ~new_n1893_;
  assign new_n2930_ = ~pi464 | ~new_n2878_;
  assign new_n2931_ = ~pi463 | ~new_n2877_;
  assign new_n2932_ = ~pi047 | ~new_n1893_;
  assign new_n2933_ = ~pi463 | ~new_n2878_;
  assign new_n2934_ = ~pi462 | ~new_n2877_;
  assign new_n2935_ = ~pi048 | ~new_n1893_;
  assign new_n2936_ = ~pi462 | ~new_n2878_;
  assign new_n2937_ = ~pi461 | ~new_n2877_;
  assign new_n2938_ = ~pi049 | ~new_n1893_;
  assign new_n2939_ = ~pi461 | ~new_n2878_;
  assign new_n2940_ = ~pi460 | ~new_n2877_;
  assign new_n2941_ = ~pi050 | ~new_n1893_;
  assign new_n2942_ = ~pi460 | ~new_n2878_;
  assign new_n2943_ = ~pi459 | ~new_n2877_;
  assign new_n2944_ = ~pi051 | ~new_n1893_;
  assign new_n2945_ = ~pi459 | ~new_n2878_;
  assign new_n2946_ = ~pi458 | ~new_n2877_;
  assign new_n2947_ = ~pi052 | ~new_n1893_;
  assign new_n2948_ = ~pi458 | ~new_n2878_;
  assign new_n2949_ = ~pi457 | ~new_n2877_;
  assign new_n2950_ = ~pi053 | ~new_n1893_;
  assign new_n2951_ = ~pi457 | ~new_n2878_;
  assign new_n2952_ = ~pi456 | ~new_n2877_;
  assign new_n2953_ = ~pi054 | ~new_n1893_;
  assign new_n2954_ = ~pi456 | ~new_n2878_;
  assign new_n2955_ = ~pi455 | ~new_n2877_;
  assign new_n2956_ = ~pi055 | ~new_n1893_;
  assign new_n2957_ = ~pi455 | ~new_n2878_;
  assign new_n2958_ = ~pi454 | ~new_n2877_;
  assign new_n2959_ = ~pi056 | ~new_n1893_;
  assign new_n2960_ = ~pi454 | ~new_n2878_;
  assign new_n2961_ = ~pi453 | ~new_n2877_;
  assign new_n2962_ = ~pi057 | ~new_n1893_;
  assign new_n2963_ = ~pi453 | ~new_n2878_;
  assign new_n2964_ = ~pi452 | ~new_n2877_;
  assign new_n2965_ = ~pi058 | ~new_n1893_;
  assign new_n2966_ = ~pi452 | ~new_n2878_;
  assign new_n2967_ = ~pi451 | ~new_n2877_;
  assign new_n2968_ = ~pi059 | ~new_n1893_;
  assign new_n2969_ = ~pi451 | ~new_n2878_;
  assign new_n2970_ = ~pi450 | ~new_n2877_;
  assign new_n2971_ = ~pi060 | ~new_n1893_;
  assign new_n2972_ = ~pi450 | ~new_n2878_;
  assign new_n2973_ = ~pi449 | ~new_n2877_;
  assign new_n2974_ = ~pi061 | ~new_n1893_;
  assign new_n2975_ = ~pi449 | ~new_n2878_;
  assign new_n2976_ = ~pi448 | ~new_n2877_;
  assign new_n2977_ = ~pi062 | ~new_n1893_;
  assign new_n2978_ = ~pi448 | ~new_n2878_;
  assign new_n2979_ = ~pi447 | ~new_n2877_;
  assign new_n2980_ = ~pi063 | ~new_n1893_;
  assign new_n2981_ = ~pi447 | ~new_n2878_;
  assign new_n2982_ = ~pi446 | ~new_n2877_;
  assign new_n2983_ = ~pi064 | ~new_n1893_;
  assign new_n2984_ = ~pi446 | ~new_n2878_;
  assign new_n2985_ = ~pi445 | ~new_n2877_;
  assign new_n2986_ = ~pi065 | ~new_n1893_;
  assign new_n2987_ = ~pi445 | ~new_n2878_;
  assign new_n2988_ = ~pi444 | ~new_n2877_;
  assign new_n2989_ = ~pi066 | ~new_n1893_;
  assign new_n2990_ = ~pi444 | ~new_n2878_;
  assign new_n2991_ = ~pi443 | ~new_n2877_;
  assign new_n2992_ = ~pi067 | ~new_n1893_;
  assign new_n2993_ = ~pi443 | ~new_n2878_;
  assign new_n2994_ = ~pi442 | ~new_n2877_;
  assign new_n2995_ = ~pi068 | ~new_n1893_;
  assign new_n2996_ = ~pi442 | ~new_n2878_;
  assign new_n2997_ = ~pi441 | ~new_n2877_;
  assign new_n2998_ = ~pi069 | ~new_n1893_;
  assign new_n2999_ = ~pi441 | ~new_n2878_;
  assign new_n3000_ = ~pi440 | ~new_n2877_;
  assign new_n3001_ = ~pi070 | ~new_n1893_;
  assign new_n3002_ = ~new_n1904_;
  assign new_n3003_ = ~new_n3002_ | ~new_n1901_;
  assign new_n3004_ = ~pi033 | ~new_n2903_;
  assign new_n3005_ = ~new_n1905_;
  assign new_n3006_ = ~new_n3005_ | ~new_n1901_;
  assign new_n3007_ = pi073 | pi033;
  assign new_n3008_ = ~new_n6268_ | ~new_n6267_ | ~new_n3007_;
  assign new_n3009_ = ~new_n1899_;
  assign new_n3010_ = ~new_n3009_ | ~pi036 | ~new_n1891_;
  assign new_n3011_ = ~new_n2138_ | ~new_n1905_;
  assign new_n3012_ = ~new_n3011_ | ~new_n3010_;
  assign new_n3013_ = ~new_n3012_ | ~pi073 | ~new_n3004_;
  assign new_n3014_ = ~pi071 | ~new_n3008_;
  assign new_n3015_ = ~pi035 | ~new_n2866_;
  assign new_n3016_ = ~new_n2141_ | ~new_n6270_;
  assign new_n3017_ = ~pi071 | ~new_n1904_;
  assign new_n3018_ = ~pi033 | ~new_n1902_;
  assign new_n3019_ = ~new_n3018_ | ~new_n3017_;
  assign new_n3020_ = ~new_n3019_ | ~new_n1892_;
  assign new_n3021_ = ~new_n2824_ | ~new_n1899_;
  assign new_n3022_ = ~new_n1924_;
  assign new_n3023_ = ~new_n1913_;
  assign new_n3024_ = ~new_n2088_;
  assign new_n3025_ = ~new_n1912_;
  assign new_n3026_ = ~new_n1918_;
  assign new_n3027_ = ~new_n1911_;
  assign new_n3028_ = ~pi178 | ~new_n3027_;
  assign new_n3029_ = ~pi234 | ~new_n1129_;
  assign new_n3030_ = ~pi226 | ~new_n1128_;
  assign new_n3031_ = ~pi218 | ~new_n1127_;
  assign new_n3032_ = ~pi210 | ~new_n1125_;
  assign new_n3033_ = ~pi202 | ~new_n1124_;
  assign new_n3034_ = ~pi194 | ~new_n1123_;
  assign new_n3035_ = ~pi186 | ~new_n1122_;
  assign new_n3036_ = ~pi170 | ~new_n1121_;
  assign new_n3037_ = ~pi162 | ~new_n1120_;
  assign new_n3038_ = ~pi154 | ~new_n1118_;
  assign new_n3039_ = ~pi146 | ~new_n1116_;
  assign new_n3040_ = ~pi138 | ~new_n1115_;
  assign new_n3041_ = ~pi130 | ~new_n1114_;
  assign new_n3042_ = ~pi122 | ~new_n1112_;
  assign new_n3043_ = ~pi114 | ~new_n1110_;
  assign new_n3044_ = ~new_n1927_;
  assign new_n3045_ = ~new_n1922_;
  assign new_n3046_ = ~pi242 | ~pi176 | ~pi241 | ~pi240 | ~new_n1914_;
  assign new_n3047_ = ~new_n3025_ | ~pi232 | ~new_n1914_;
  assign new_n3048_ = ~new_n1909_ | ~pi242 | ~pi224 | ~new_n1126_;
  assign new_n3049_ = ~new_n1910_ | ~pi241 | ~pi216 | ~new_n1126_;
  assign new_n3050_ = ~new_n1914_ | ~pi240 | ~pi200 | ~new_n3023_;
  assign new_n3051_ = ~new_n2166_ | ~new_n2165_ | ~pi240;
  assign new_n3052_ = ~new_n2168_ | ~new_n2167_ | ~pi240;
  assign new_n3053_ = ~new_n2169_ | ~new_n3025_;
  assign new_n3054_ = ~new_n2171_ | ~new_n2170_ | ~pi241;
  assign new_n3055_ = ~pi239 | ~pi144 | ~pi242 | ~pi241 | ~new_n1908_;
  assign new_n3056_ = ~new_n2172_ | ~new_n3023_ | ~pi240;
  assign new_n3057_ = ~pi239 | ~pi128 | ~pi242 | ~pi240 | ~new_n1909_;
  assign new_n3058_ = ~pi239 | ~pi120 | ~pi241 | ~pi240 | ~new_n1910_;
  assign new_n3059_ = ~pi239 | ~pi112 | ~pi242 | ~pi241 | ~pi240;
  assign new_n3060_ = ~new_n2818_;
  assign new_n3061_ = ~pi179 | ~new_n3027_;
  assign new_n3062_ = ~pi235 | ~new_n1129_;
  assign new_n3063_ = ~pi227 | ~new_n1128_;
  assign new_n3064_ = ~pi219 | ~new_n1127_;
  assign new_n3065_ = ~pi211 | ~new_n1125_;
  assign new_n3066_ = ~pi203 | ~new_n1124_;
  assign new_n3067_ = ~pi195 | ~new_n1123_;
  assign new_n3068_ = ~pi187 | ~new_n1122_;
  assign new_n3069_ = ~pi171 | ~new_n1121_;
  assign new_n3070_ = ~pi163 | ~new_n1120_;
  assign new_n3071_ = ~pi155 | ~new_n1118_;
  assign new_n3072_ = ~pi147 | ~new_n1116_;
  assign new_n3073_ = ~pi139 | ~new_n1115_;
  assign new_n3074_ = ~pi131 | ~new_n1114_;
  assign new_n3075_ = ~pi123 | ~new_n1112_;
  assign new_n3076_ = ~pi115 | ~new_n1110_;
  assign new_n3077_ = ~new_n2816_;
  assign new_n3078_ = ~pi174 | ~new_n3027_;
  assign new_n3079_ = ~pi230 | ~new_n1129_;
  assign new_n3080_ = ~pi222 | ~new_n1128_;
  assign new_n3081_ = ~pi214 | ~new_n1127_;
  assign new_n3082_ = ~pi206 | ~new_n1125_;
  assign new_n3083_ = ~pi198 | ~new_n1124_;
  assign new_n3084_ = ~pi190 | ~new_n1123_;
  assign new_n3085_ = ~pi182 | ~new_n1122_;
  assign new_n3086_ = ~pi166 | ~new_n1121_;
  assign new_n3087_ = ~pi158 | ~new_n1120_;
  assign new_n3088_ = ~pi150 | ~new_n1118_;
  assign new_n3089_ = ~pi142 | ~new_n1116_;
  assign new_n3090_ = ~pi134 | ~new_n1115_;
  assign new_n3091_ = ~pi126 | ~new_n1114_;
  assign new_n3092_ = ~pi118 | ~new_n1112_;
  assign new_n3093_ = ~pi110 | ~new_n1110_;
  assign new_n3094_ = ~new_n2035_;
  assign new_n3095_ = ~pi175 | ~new_n2143_ | ~new_n3026_;
  assign new_n3096_ = ~new_n1113_ | ~pi223 | ~new_n1126_;
  assign new_n3097_ = ~new_n1111_ | ~pi215 | ~new_n1126_;
  assign new_n3098_ = ~new_n3026_ | ~pi199 | ~new_n3023_;
  assign new_n3099_ = ~pi191 | ~new_n1113_ | ~new_n3026_;
  assign new_n3100_ = ~pi183 | ~new_n1111_ | ~new_n3026_;
  assign new_n3101_ = ~new_n2152_ | ~pi135 | ~new_n3023_;
  assign new_n3102_ = ~pi127 | ~new_n2152_ | ~new_n1113_;
  assign new_n3103_ = ~pi119 | ~new_n2152_ | ~new_n1111_;
  assign new_n3104_ = ~pi111 | ~new_n2152_ | ~new_n2143_;
  assign new_n3105_ = ~new_n1921_;
  assign new_n3106_ = ~pi180 | ~new_n3027_;
  assign new_n3107_ = ~pi236 | ~new_n1129_;
  assign new_n3108_ = ~pi228 | ~new_n1128_;
  assign new_n3109_ = ~pi220 | ~new_n1127_;
  assign new_n3110_ = ~pi212 | ~new_n1125_;
  assign new_n3111_ = ~pi204 | ~new_n1124_;
  assign new_n3112_ = ~pi196 | ~new_n1123_;
  assign new_n3113_ = ~pi188 | ~new_n1122_;
  assign new_n3114_ = ~pi172 | ~new_n1121_;
  assign new_n3115_ = ~pi164 | ~new_n1120_;
  assign new_n3116_ = ~pi156 | ~new_n1118_;
  assign new_n3117_ = ~pi148 | ~new_n1116_;
  assign new_n3118_ = ~pi140 | ~new_n1115_;
  assign new_n3119_ = ~pi132 | ~new_n1114_;
  assign new_n3120_ = ~pi124 | ~new_n1112_;
  assign new_n3121_ = ~pi116 | ~new_n1110_;
  assign new_n3122_ = ~new_n1915_;
  assign new_n3123_ = ~pi181 | ~new_n3027_;
  assign new_n3124_ = ~pi237 | ~new_n1129_;
  assign new_n3125_ = ~pi229 | ~new_n1128_;
  assign new_n3126_ = ~pi221 | ~new_n1127_;
  assign new_n3127_ = ~pi213 | ~new_n1125_;
  assign new_n3128_ = ~pi205 | ~new_n1124_;
  assign new_n3129_ = ~pi197 | ~new_n1123_;
  assign new_n3130_ = ~pi189 | ~new_n1122_;
  assign new_n3131_ = ~pi173 | ~new_n1121_;
  assign new_n3132_ = ~pi165 | ~new_n1120_;
  assign new_n3133_ = ~pi157 | ~new_n1118_;
  assign new_n3134_ = ~pi149 | ~new_n1116_;
  assign new_n3135_ = ~pi141 | ~new_n1115_;
  assign new_n3136_ = ~pi133 | ~new_n1114_;
  assign new_n3137_ = ~pi125 | ~new_n1112_;
  assign new_n3138_ = ~pi117 | ~new_n1110_;
  assign new_n3139_ = ~new_n1928_;
  assign new_n3140_ = ~pi071 | ~new_n1892_;
  assign new_n3141_ = ~new_n1898_ | ~new_n3140_;
  assign new_n3142_ = ~new_n1916_;
  assign new_n3143_ = ~new_n3122_ | ~new_n2032_;
  assign new_n3144_ = ~new_n2081_;
  assign new_n3145_ = ~new_n1931_ | ~new_n1916_ | ~new_n2034_;
  assign new_n3146_ = ~new_n3145_ | ~new_n1901_;
  assign new_n3147_ = ~new_n1929_;
  assign new_n3148_ = ~new_n3105_ | ~new_n2818_;
  assign new_n3149_ = ~new_n2841_ | ~new_n1930_;
  assign new_n3150_ = ~new_n3149_ | ~new_n2224_;
  assign new_n3151_ = ~new_n2225_ | ~new_n3150_;
  assign new_n3152_ = ~new_n2860_ | ~new_n2032_;
  assign new_n3153_ = ~new_n3152_ | ~new_n6327_ | ~new_n6326_;
  assign new_n3154_ = ~new_n1105_ | ~new_n2907_;
  assign new_n3155_ = pi477 | pi476;
  assign new_n3156_ = ~new_n1937_;
  assign new_n3157_ = ~new_n3156_ | ~new_n1906_;
  assign new_n3158_ = ~pi108 | ~pi035;
  assign new_n3159_ = ~new_n1939_;
  assign new_n3160_ = ~pi108 | ~new_n6333_ | ~new_n6332_;
  assign new_n3161_ = ~pi107 | ~new_n1939_;
  assign new_n3162_ = ~new_n6249_ | ~new_n2891_;
  assign new_n3163_ = ~new_n2228_ | ~new_n3159_;
  assign new_n3164_ = ~pi108 | ~new_n3162_;
  assign new_n3165_ = ~new_n1025_ | ~new_n6249_;
  assign new_n3166_ = ~new_n2897_ | ~new_n2906_;
  assign new_n3167_ = ~new_n6249_ | ~new_n2890_;
  assign new_n3168_ = ~new_n1025_ | ~new_n1937_;
  assign new_n3169_ = ~new_n1969_;
  assign new_n3170_ = ~new_n1975_;
  assign new_n3171_ = ~new_n1976_;
  assign new_n3172_ = ~new_n1958_;
  assign new_n3173_ = ~new_n1957_;
  assign new_n3174_ = ~new_n1986_;
  assign new_n3175_ = ~new_n8007_ | ~new_n1957_;
  assign new_n3176_ = ~new_n2002_;
  assign new_n3177_ = ~new_n1959_;
  assign new_n3178_ = ~new_n1949_;
  assign new_n3179_ = ~new_n1950_;
  assign new_n3180_ = ~new_n1095_ | ~new_n1099_;
  assign new_n3181_ = ~new_n1965_;
  assign new_n3182_ = ~new_n2000_;
  assign new_n3183_ = ~new_n1984_;
  assign new_n3184_ = ~pi244 | ~new_n1949_;
  assign new_n3185_ = ~new_n2004_;
  assign new_n3186_ = ~new_n1973_;
  assign new_n3187_ = ~new_n1967_;
  assign new_n3188_ = ~new_n1879_;
  assign new_n3189_ = ~new_n1089_ | ~new_n1093_;
  assign new_n3190_ = ~new_n1966_;
  assign new_n3191_ = ~pi108 | ~new_n1907_;
  assign new_n3192_ = ~new_n1943_ | ~new_n3191_ | ~new_n1941_;
  assign new_n3193_ = ~new_n3173_ | ~new_n1133_;
  assign new_n3194_ = ~new_n1137_ | ~new_n1015_;
  assign new_n3195_ = ~new_n1964_ | ~new_n3194_;
  assign new_n3196_ = ~new_n3181_ | ~new_n3195_;
  assign new_n3197_ = ~pi106 | ~new_n1950_;
  assign new_n3198_ = ~new_n3190_ | ~pi107;
  assign new_n3199_ = ~new_n3196_ | ~new_n2232_;
  assign new_n3200_ = ~new_n1137_ | ~new_n1045_;
  assign new_n3201_ = ~new_n1964_ | ~new_n3200_;
  assign new_n3202_ = ~new_n3201_ | ~new_n1965_;
  assign new_n3203_ = ~pi107 | ~new_n1966_;
  assign new_n3204_ = ~new_n3203_ | ~new_n3202_;
  assign new_n3205_ = ~new_n1072_ | ~new_n3179_;
  assign new_n3206_ = ~new_n1070_ | ~new_n1134_;
  assign new_n3207_ = ~new_n1069_ | ~new_n3177_;
  assign new_n3208_ = ~new_n1054_ | ~new_n3204_;
  assign new_n3209_ = ~pi110 | ~new_n3199_;
  assign new_n3210_ = ~new_n1073_ | ~new_n3179_;
  assign new_n3211_ = ~new_n1068_ | ~new_n1134_;
  assign new_n3212_ = ~new_n1067_ | ~new_n3177_;
  assign new_n3213_ = ~new_n1053_ | ~new_n3204_;
  assign new_n3214_ = ~pi111 | ~new_n3199_;
  assign new_n3215_ = ~new_n1077_ | ~new_n3179_;
  assign new_n3216_ = ~new_n1066_ | ~new_n1134_;
  assign new_n3217_ = ~new_n1065_ | ~new_n3177_;
  assign new_n3218_ = ~new_n1052_ | ~new_n3204_;
  assign new_n3219_ = ~pi112 | ~new_n3199_;
  assign new_n3220_ = ~new_n1076_ | ~new_n3179_;
  assign new_n3221_ = ~new_n1064_ | ~new_n1134_;
  assign new_n3222_ = ~new_n1063_ | ~new_n3177_;
  assign new_n3223_ = ~new_n1051_ | ~new_n3204_;
  assign new_n3224_ = ~pi113 | ~new_n3199_;
  assign new_n3225_ = ~new_n1075_ | ~new_n3179_;
  assign new_n3226_ = ~new_n1062_ | ~new_n1134_;
  assign new_n3227_ = ~new_n1061_ | ~new_n3177_;
  assign new_n3228_ = ~new_n1050_ | ~new_n3204_;
  assign new_n3229_ = ~pi114 | ~new_n3199_;
  assign new_n3230_ = ~new_n1078_ | ~new_n3179_;
  assign new_n3231_ = ~new_n1060_ | ~new_n1134_;
  assign new_n3232_ = ~new_n1059_ | ~new_n3177_;
  assign new_n3233_ = ~new_n1049_ | ~new_n3204_;
  assign new_n3234_ = ~pi115 | ~new_n3199_;
  assign new_n3235_ = ~new_n1071_ | ~new_n3179_;
  assign new_n3236_ = ~new_n1058_ | ~new_n1134_;
  assign new_n3237_ = ~new_n1057_ | ~new_n3177_;
  assign new_n3238_ = ~new_n1048_ | ~new_n3204_;
  assign new_n3239_ = ~pi116 | ~new_n3199_;
  assign new_n3240_ = ~new_n1074_ | ~new_n3179_;
  assign new_n3241_ = ~new_n1056_ | ~new_n1134_;
  assign new_n3242_ = ~new_n1055_ | ~new_n3177_;
  assign new_n3243_ = ~new_n1047_ | ~new_n3204_;
  assign new_n3244_ = ~pi117 | ~new_n3199_;
  assign new_n3245_ = ~new_n1970_;
  assign new_n3246_ = ~new_n1971_;
  assign new_n3247_ = ~new_n1968_;
  assign new_n3248_ = ~new_n1100_ | ~new_n1095_;
  assign new_n3249_ = ~new_n1972_;
  assign new_n3250_ = ~new_n1880_;
  assign new_n3251_ = ~new_n3169_ | ~new_n1133_;
  assign new_n3252_ = ~new_n1139_ | ~new_n1015_;
  assign new_n3253_ = ~new_n1964_ | ~new_n3252_;
  assign new_n3254_ = ~new_n3249_ | ~new_n3253_;
  assign new_n3255_ = ~pi106 | ~new_n1968_;
  assign new_n3256_ = ~pi107 | ~new_n1880_;
  assign new_n3257_ = ~new_n3254_ | ~new_n2241_;
  assign new_n3258_ = ~new_n1139_ | ~new_n1045_;
  assign new_n3259_ = ~new_n1964_ | ~new_n3258_;
  assign new_n3260_ = ~new_n3259_ | ~new_n1972_;
  assign new_n3261_ = ~pi107 | ~new_n3250_;
  assign new_n3262_ = ~new_n3261_ | ~new_n3260_;
  assign new_n3263_ = ~new_n3247_ | ~new_n1072_;
  assign new_n3264_ = ~new_n1138_ | ~new_n1070_;
  assign new_n3265_ = ~new_n3246_ | ~new_n1069_;
  assign new_n3266_ = ~new_n1054_ | ~new_n3262_;
  assign new_n3267_ = ~pi118 | ~new_n3257_;
  assign new_n3268_ = ~new_n3247_ | ~new_n1073_;
  assign new_n3269_ = ~new_n1138_ | ~new_n1068_;
  assign new_n3270_ = ~new_n3246_ | ~new_n1067_;
  assign new_n3271_ = ~new_n1053_ | ~new_n3262_;
  assign new_n3272_ = ~pi119 | ~new_n3257_;
  assign new_n3273_ = ~new_n3247_ | ~new_n1077_;
  assign new_n3274_ = ~new_n1138_ | ~new_n1066_;
  assign new_n3275_ = ~new_n3246_ | ~new_n1065_;
  assign new_n3276_ = ~new_n1052_ | ~new_n3262_;
  assign new_n3277_ = ~pi120 | ~new_n3257_;
  assign new_n3278_ = ~new_n3247_ | ~new_n1076_;
  assign new_n3279_ = ~new_n1138_ | ~new_n1064_;
  assign new_n3280_ = ~new_n3246_ | ~new_n1063_;
  assign new_n3281_ = ~new_n1051_ | ~new_n3262_;
  assign new_n3282_ = ~pi121 | ~new_n3257_;
  assign new_n3283_ = ~new_n3247_ | ~new_n1075_;
  assign new_n3284_ = ~new_n1138_ | ~new_n1062_;
  assign new_n3285_ = ~new_n3246_ | ~new_n1061_;
  assign new_n3286_ = ~new_n1050_ | ~new_n3262_;
  assign new_n3287_ = ~pi122 | ~new_n3257_;
  assign new_n3288_ = ~new_n3247_ | ~new_n1078_;
  assign new_n3289_ = ~new_n1138_ | ~new_n1060_;
  assign new_n3290_ = ~new_n3246_ | ~new_n1059_;
  assign new_n3291_ = ~new_n1049_ | ~new_n3262_;
  assign new_n3292_ = ~pi123 | ~new_n3257_;
  assign new_n3293_ = ~new_n3247_ | ~new_n1071_;
  assign new_n3294_ = ~new_n1138_ | ~new_n1058_;
  assign new_n3295_ = ~new_n3246_ | ~new_n1057_;
  assign new_n3296_ = ~new_n1048_ | ~new_n3262_;
  assign new_n3297_ = ~pi124 | ~new_n3257_;
  assign new_n3298_ = ~new_n3247_ | ~new_n1074_;
  assign new_n3299_ = ~new_n1138_ | ~new_n1056_;
  assign new_n3300_ = ~new_n3246_ | ~new_n1055_;
  assign new_n3301_ = ~new_n1047_ | ~new_n3262_;
  assign new_n3302_ = ~pi125 | ~new_n3257_;
  assign new_n3303_ = ~new_n1977_;
  assign new_n3304_ = ~new_n1978_;
  assign new_n3305_ = ~new_n1974_;
  assign new_n3306_ = ~new_n1101_ | ~new_n1095_;
  assign new_n3307_ = ~new_n1979_;
  assign new_n3308_ = ~new_n1094_ | ~new_n1089_;
  assign new_n3309_ = ~new_n1980_;
  assign new_n3310_ = ~new_n3170_ | ~new_n1133_;
  assign new_n3311_ = ~new_n1141_ | ~new_n1015_;
  assign new_n3312_ = ~new_n1964_ | ~new_n3311_;
  assign new_n3313_ = ~new_n3307_ | ~new_n3312_;
  assign new_n3314_ = ~pi106 | ~new_n1974_;
  assign new_n3315_ = ~new_n3309_ | ~pi107;
  assign new_n3316_ = ~new_n3313_ | ~new_n2250_;
  assign new_n3317_ = ~new_n1141_ | ~new_n1045_;
  assign new_n3318_ = ~new_n1964_ | ~new_n3317_;
  assign new_n3319_ = ~new_n3318_ | ~new_n1979_;
  assign new_n3320_ = ~pi107 | ~new_n1980_;
  assign new_n3321_ = ~new_n3320_ | ~new_n3319_;
  assign new_n3322_ = ~new_n3305_ | ~new_n1072_;
  assign new_n3323_ = ~new_n1140_ | ~new_n1070_;
  assign new_n3324_ = ~new_n3304_ | ~new_n1069_;
  assign new_n3325_ = ~new_n1054_ | ~new_n3321_;
  assign new_n3326_ = ~pi126 | ~new_n3316_;
  assign new_n3327_ = ~new_n3305_ | ~new_n1073_;
  assign new_n3328_ = ~new_n1140_ | ~new_n1068_;
  assign new_n3329_ = ~new_n3304_ | ~new_n1067_;
  assign new_n3330_ = ~new_n1053_ | ~new_n3321_;
  assign new_n3331_ = ~pi127 | ~new_n3316_;
  assign new_n3332_ = ~new_n3305_ | ~new_n1077_;
  assign new_n3333_ = ~new_n1140_ | ~new_n1066_;
  assign new_n3334_ = ~new_n3304_ | ~new_n1065_;
  assign new_n3335_ = ~new_n1052_ | ~new_n3321_;
  assign new_n3336_ = ~pi128 | ~new_n3316_;
  assign new_n3337_ = ~new_n3305_ | ~new_n1076_;
  assign new_n3338_ = ~new_n1140_ | ~new_n1064_;
  assign new_n3339_ = ~new_n3304_ | ~new_n1063_;
  assign new_n3340_ = ~new_n1051_ | ~new_n3321_;
  assign new_n3341_ = ~pi129 | ~new_n3316_;
  assign new_n3342_ = ~new_n3305_ | ~new_n1075_;
  assign new_n3343_ = ~new_n1140_ | ~new_n1062_;
  assign new_n3344_ = ~new_n3304_ | ~new_n1061_;
  assign new_n3345_ = ~new_n1050_ | ~new_n3321_;
  assign new_n3346_ = ~pi130 | ~new_n3316_;
  assign new_n3347_ = ~new_n3305_ | ~new_n1078_;
  assign new_n3348_ = ~new_n1140_ | ~new_n1060_;
  assign new_n3349_ = ~new_n3304_ | ~new_n1059_;
  assign new_n3350_ = ~new_n1049_ | ~new_n3321_;
  assign new_n3351_ = ~pi131 | ~new_n3316_;
  assign new_n3352_ = ~new_n3305_ | ~new_n1071_;
  assign new_n3353_ = ~new_n1140_ | ~new_n1058_;
  assign new_n3354_ = ~new_n3304_ | ~new_n1057_;
  assign new_n3355_ = ~new_n1048_ | ~new_n3321_;
  assign new_n3356_ = ~pi132 | ~new_n3316_;
  assign new_n3357_ = ~new_n3305_ | ~new_n1074_;
  assign new_n3358_ = ~new_n1140_ | ~new_n1056_;
  assign new_n3359_ = ~new_n3304_ | ~new_n1055_;
  assign new_n3360_ = ~new_n1047_ | ~new_n3321_;
  assign new_n3361_ = ~pi133 | ~new_n3316_;
  assign new_n3362_ = ~new_n1982_;
  assign new_n3363_ = ~new_n1981_;
  assign new_n3364_ = ~new_n1102_ | ~new_n1095_;
  assign new_n3365_ = ~new_n1983_;
  assign new_n3366_ = ~new_n1881_;
  assign new_n3367_ = ~new_n1143_ | ~new_n1133_;
  assign new_n3368_ = ~new_n1146_ | ~new_n1015_;
  assign new_n3369_ = ~new_n1964_ | ~new_n3368_;
  assign new_n3370_ = ~new_n3365_ | ~new_n3369_;
  assign new_n3371_ = ~pi106 | ~new_n1981_;
  assign new_n3372_ = ~pi107 | ~new_n1881_;
  assign new_n3373_ = ~new_n3370_ | ~new_n2259_;
  assign new_n3374_ = ~new_n1146_ | ~new_n1045_;
  assign new_n3375_ = ~new_n1964_ | ~new_n3374_;
  assign new_n3376_ = ~new_n3375_ | ~new_n1983_;
  assign new_n3377_ = ~pi107 | ~new_n3366_;
  assign new_n3378_ = ~new_n3377_ | ~new_n3376_;
  assign new_n3379_ = ~new_n3363_ | ~new_n1072_;
  assign new_n3380_ = ~new_n1144_ | ~new_n1070_;
  assign new_n3381_ = ~new_n3362_ | ~new_n1069_;
  assign new_n3382_ = ~new_n1054_ | ~new_n3378_;
  assign new_n3383_ = ~pi134 | ~new_n3373_;
  assign new_n3384_ = ~new_n3363_ | ~new_n1073_;
  assign new_n3385_ = ~new_n1144_ | ~new_n1068_;
  assign new_n3386_ = ~new_n3362_ | ~new_n1067_;
  assign new_n3387_ = ~new_n1053_ | ~new_n3378_;
  assign new_n3388_ = ~pi135 | ~new_n3373_;
  assign new_n3389_ = ~new_n3363_ | ~new_n1077_;
  assign new_n3390_ = ~new_n1144_ | ~new_n1066_;
  assign new_n3391_ = ~new_n3362_ | ~new_n1065_;
  assign new_n3392_ = ~new_n1052_ | ~new_n3378_;
  assign new_n3393_ = ~pi136 | ~new_n3373_;
  assign new_n3394_ = ~new_n3363_ | ~new_n1076_;
  assign new_n3395_ = ~new_n1144_ | ~new_n1064_;
  assign new_n3396_ = ~new_n3362_ | ~new_n1063_;
  assign new_n3397_ = ~new_n1051_ | ~new_n3378_;
  assign new_n3398_ = ~pi137 | ~new_n3373_;
  assign new_n3399_ = ~new_n3363_ | ~new_n1075_;
  assign new_n3400_ = ~new_n1144_ | ~new_n1062_;
  assign new_n3401_ = ~new_n3362_ | ~new_n1061_;
  assign new_n3402_ = ~new_n1050_ | ~new_n3378_;
  assign new_n3403_ = ~pi138 | ~new_n3373_;
  assign new_n3404_ = ~new_n3363_ | ~new_n1078_;
  assign new_n3405_ = ~new_n1144_ | ~new_n1060_;
  assign new_n3406_ = ~new_n3362_ | ~new_n1059_;
  assign new_n3407_ = ~new_n1049_ | ~new_n3378_;
  assign new_n3408_ = ~pi139 | ~new_n3373_;
  assign new_n3409_ = ~new_n3363_ | ~new_n1071_;
  assign new_n3410_ = ~new_n1144_ | ~new_n1058_;
  assign new_n3411_ = ~new_n3362_ | ~new_n1057_;
  assign new_n3412_ = ~new_n1048_ | ~new_n3378_;
  assign new_n3413_ = ~pi140 | ~new_n3373_;
  assign new_n3414_ = ~new_n3363_ | ~new_n1074_;
  assign new_n3415_ = ~new_n1144_ | ~new_n1056_;
  assign new_n3416_ = ~new_n3362_ | ~new_n1055_;
  assign new_n3417_ = ~new_n1047_ | ~new_n3378_;
  assign new_n3418_ = ~pi141 | ~new_n3373_;
  assign new_n3419_ = ~new_n1987_;
  assign new_n3420_ = ~new_n1985_;
  assign new_n3421_ = ~new_n1097_ | ~new_n1099_;
  assign new_n3422_ = ~new_n1988_;
  assign new_n3423_ = ~new_n1091_ | ~new_n1093_;
  assign new_n3424_ = ~new_n1989_;
  assign new_n3425_ = ~new_n3174_ | ~new_n3173_;
  assign new_n3426_ = ~new_n1149_ | ~new_n1015_;
  assign new_n3427_ = ~new_n1964_ | ~new_n3426_;
  assign new_n3428_ = ~new_n3422_ | ~new_n3427_;
  assign new_n3429_ = ~pi106 | ~new_n1985_;
  assign new_n3430_ = ~new_n3424_ | ~pi107;
  assign new_n3431_ = ~new_n3428_ | ~new_n2268_;
  assign new_n3432_ = ~new_n1149_ | ~new_n1045_;
  assign new_n3433_ = ~new_n1964_ | ~new_n3432_;
  assign new_n3434_ = ~new_n3433_ | ~new_n1988_;
  assign new_n3435_ = ~pi107 | ~new_n1989_;
  assign new_n3436_ = ~new_n3435_ | ~new_n3434_;
  assign new_n3437_ = ~new_n3420_ | ~new_n1072_;
  assign new_n3438_ = ~new_n1148_ | ~new_n1070_;
  assign new_n3439_ = ~new_n3419_ | ~new_n1069_;
  assign new_n3440_ = ~new_n1054_ | ~new_n3436_;
  assign new_n3441_ = ~pi142 | ~new_n3431_;
  assign new_n3442_ = ~new_n3420_ | ~new_n1073_;
  assign new_n3443_ = ~new_n1148_ | ~new_n1068_;
  assign new_n3444_ = ~new_n3419_ | ~new_n1067_;
  assign new_n3445_ = ~new_n1053_ | ~new_n3436_;
  assign new_n3446_ = ~pi143 | ~new_n3431_;
  assign new_n3447_ = ~new_n3420_ | ~new_n1077_;
  assign new_n3448_ = ~new_n1148_ | ~new_n1066_;
  assign new_n3449_ = ~new_n3419_ | ~new_n1065_;
  assign new_n3450_ = ~new_n1052_ | ~new_n3436_;
  assign new_n3451_ = ~pi144 | ~new_n3431_;
  assign new_n3452_ = ~new_n3420_ | ~new_n1076_;
  assign new_n3453_ = ~new_n1148_ | ~new_n1064_;
  assign new_n3454_ = ~new_n3419_ | ~new_n1063_;
  assign new_n3455_ = ~new_n1051_ | ~new_n3436_;
  assign new_n3456_ = ~pi145 | ~new_n3431_;
  assign new_n3457_ = ~new_n3420_ | ~new_n1075_;
  assign new_n3458_ = ~new_n1148_ | ~new_n1062_;
  assign new_n3459_ = ~new_n3419_ | ~new_n1061_;
  assign new_n3460_ = ~new_n1050_ | ~new_n3436_;
  assign new_n3461_ = ~pi146 | ~new_n3431_;
  assign new_n3462_ = ~new_n3420_ | ~new_n1078_;
  assign new_n3463_ = ~new_n1148_ | ~new_n1060_;
  assign new_n3464_ = ~new_n3419_ | ~new_n1059_;
  assign new_n3465_ = ~new_n1049_ | ~new_n3436_;
  assign new_n3466_ = ~pi147 | ~new_n3431_;
  assign new_n3467_ = ~new_n3420_ | ~new_n1071_;
  assign new_n3468_ = ~new_n1148_ | ~new_n1058_;
  assign new_n3469_ = ~new_n3419_ | ~new_n1057_;
  assign new_n3470_ = ~new_n1048_ | ~new_n3436_;
  assign new_n3471_ = ~pi148 | ~new_n3431_;
  assign new_n3472_ = ~new_n3420_ | ~new_n1074_;
  assign new_n3473_ = ~new_n1148_ | ~new_n1056_;
  assign new_n3474_ = ~new_n3419_ | ~new_n1055_;
  assign new_n3475_ = ~new_n1047_ | ~new_n3436_;
  assign new_n3476_ = ~pi149 | ~new_n3431_;
  assign new_n3477_ = ~new_n1991_;
  assign new_n3478_ = ~new_n1990_;
  assign new_n3479_ = ~new_n1097_ | ~new_n1100_;
  assign new_n3480_ = ~new_n1992_;
  assign new_n3481_ = ~new_n1882_;
  assign new_n3482_ = ~new_n3174_ | ~new_n3169_;
  assign new_n3483_ = ~new_n1151_ | ~new_n1015_;
  assign new_n3484_ = ~new_n1964_ | ~new_n3483_;
  assign new_n3485_ = ~new_n3480_ | ~new_n3484_;
  assign new_n3486_ = ~pi106 | ~new_n1990_;
  assign new_n3487_ = ~pi107 | ~new_n1882_;
  assign new_n3488_ = ~new_n3485_ | ~new_n2277_;
  assign new_n3489_ = ~new_n1151_ | ~new_n1045_;
  assign new_n3490_ = ~new_n1964_ | ~new_n3489_;
  assign new_n3491_ = ~new_n3490_ | ~new_n1992_;
  assign new_n3492_ = ~pi107 | ~new_n3481_;
  assign new_n3493_ = ~new_n3492_ | ~new_n3491_;
  assign new_n3494_ = ~new_n3478_ | ~new_n1072_;
  assign new_n3495_ = ~new_n1150_ | ~new_n1070_;
  assign new_n3496_ = ~new_n3477_ | ~new_n1069_;
  assign new_n3497_ = ~new_n1054_ | ~new_n3493_;
  assign new_n3498_ = ~pi150 | ~new_n3488_;
  assign new_n3499_ = ~new_n3478_ | ~new_n1073_;
  assign new_n3500_ = ~new_n1150_ | ~new_n1068_;
  assign new_n3501_ = ~new_n3477_ | ~new_n1067_;
  assign new_n3502_ = ~new_n1053_ | ~new_n3493_;
  assign new_n3503_ = ~pi151 | ~new_n3488_;
  assign new_n3504_ = ~new_n3478_ | ~new_n1077_;
  assign new_n3505_ = ~new_n1150_ | ~new_n1066_;
  assign new_n3506_ = ~new_n3477_ | ~new_n1065_;
  assign new_n3507_ = ~new_n1052_ | ~new_n3493_;
  assign new_n3508_ = ~pi152 | ~new_n3488_;
  assign new_n3509_ = ~new_n3478_ | ~new_n1076_;
  assign new_n3510_ = ~new_n1150_ | ~new_n1064_;
  assign new_n3511_ = ~new_n3477_ | ~new_n1063_;
  assign new_n3512_ = ~new_n1051_ | ~new_n3493_;
  assign new_n3513_ = ~pi153 | ~new_n3488_;
  assign new_n3514_ = ~new_n3478_ | ~new_n1075_;
  assign new_n3515_ = ~new_n1150_ | ~new_n1062_;
  assign new_n3516_ = ~new_n3477_ | ~new_n1061_;
  assign new_n3517_ = ~new_n1050_ | ~new_n3493_;
  assign new_n3518_ = ~pi154 | ~new_n3488_;
  assign new_n3519_ = ~new_n3478_ | ~new_n1078_;
  assign new_n3520_ = ~new_n1150_ | ~new_n1060_;
  assign new_n3521_ = ~new_n3477_ | ~new_n1059_;
  assign new_n3522_ = ~new_n1049_ | ~new_n3493_;
  assign new_n3523_ = ~pi155 | ~new_n3488_;
  assign new_n3524_ = ~new_n3478_ | ~new_n1071_;
  assign new_n3525_ = ~new_n1150_ | ~new_n1058_;
  assign new_n3526_ = ~new_n3477_ | ~new_n1057_;
  assign new_n3527_ = ~new_n1048_ | ~new_n3493_;
  assign new_n3528_ = ~pi156 | ~new_n3488_;
  assign new_n3529_ = ~new_n3478_ | ~new_n1074_;
  assign new_n3530_ = ~new_n1150_ | ~new_n1056_;
  assign new_n3531_ = ~new_n3477_ | ~new_n1055_;
  assign new_n3532_ = ~new_n1047_ | ~new_n3493_;
  assign new_n3533_ = ~pi157 | ~new_n3488_;
  assign new_n3534_ = ~new_n1994_;
  assign new_n3535_ = ~new_n1993_;
  assign new_n3536_ = ~new_n1097_ | ~new_n1101_;
  assign new_n3537_ = ~new_n1995_;
  assign new_n3538_ = ~new_n1091_ | ~new_n1094_;
  assign new_n3539_ = ~new_n1996_;
  assign new_n3540_ = ~new_n3174_ | ~new_n3170_;
  assign new_n3541_ = ~new_n1153_ | ~new_n1015_;
  assign new_n3542_ = ~new_n1964_ | ~new_n3541_;
  assign new_n3543_ = ~new_n3537_ | ~new_n3542_;
  assign new_n3544_ = ~pi106 | ~new_n1993_;
  assign new_n3545_ = ~new_n3539_ | ~pi107;
  assign new_n3546_ = ~new_n3543_ | ~new_n2286_;
  assign new_n3547_ = ~new_n1153_ | ~new_n1045_;
  assign new_n3548_ = ~new_n1964_ | ~new_n3547_;
  assign new_n3549_ = ~new_n3548_ | ~new_n1995_;
  assign new_n3550_ = ~pi107 | ~new_n1996_;
  assign new_n3551_ = ~new_n3550_ | ~new_n3549_;
  assign new_n3552_ = ~new_n3535_ | ~new_n1072_;
  assign new_n3553_ = ~new_n1152_ | ~new_n1070_;
  assign new_n3554_ = ~new_n3534_ | ~new_n1069_;
  assign new_n3555_ = ~new_n1054_ | ~new_n3551_;
  assign new_n3556_ = ~pi158 | ~new_n3546_;
  assign new_n3557_ = ~new_n3535_ | ~new_n1073_;
  assign new_n3558_ = ~new_n1152_ | ~new_n1068_;
  assign new_n3559_ = ~new_n3534_ | ~new_n1067_;
  assign new_n3560_ = ~new_n1053_ | ~new_n3551_;
  assign new_n3561_ = ~pi159 | ~new_n3546_;
  assign new_n3562_ = ~new_n3535_ | ~new_n1077_;
  assign new_n3563_ = ~new_n1152_ | ~new_n1066_;
  assign new_n3564_ = ~new_n3534_ | ~new_n1065_;
  assign new_n3565_ = ~new_n1052_ | ~new_n3551_;
  assign new_n3566_ = ~pi160 | ~new_n3546_;
  assign new_n3567_ = ~new_n3535_ | ~new_n1076_;
  assign new_n3568_ = ~new_n1152_ | ~new_n1064_;
  assign new_n3569_ = ~new_n3534_ | ~new_n1063_;
  assign new_n3570_ = ~new_n1051_ | ~new_n3551_;
  assign new_n3571_ = ~pi161 | ~new_n3546_;
  assign new_n3572_ = ~new_n3535_ | ~new_n1075_;
  assign new_n3573_ = ~new_n1152_ | ~new_n1062_;
  assign new_n3574_ = ~new_n3534_ | ~new_n1061_;
  assign new_n3575_ = ~new_n1050_ | ~new_n3551_;
  assign new_n3576_ = ~pi162 | ~new_n3546_;
  assign new_n3577_ = ~new_n3535_ | ~new_n1078_;
  assign new_n3578_ = ~new_n1152_ | ~new_n1060_;
  assign new_n3579_ = ~new_n3534_ | ~new_n1059_;
  assign new_n3580_ = ~new_n1049_ | ~new_n3551_;
  assign new_n3581_ = ~pi163 | ~new_n3546_;
  assign new_n3582_ = ~new_n3535_ | ~new_n1071_;
  assign new_n3583_ = ~new_n1152_ | ~new_n1058_;
  assign new_n3584_ = ~new_n3534_ | ~new_n1057_;
  assign new_n3585_ = ~new_n1048_ | ~new_n3551_;
  assign new_n3586_ = ~pi164 | ~new_n3546_;
  assign new_n3587_ = ~new_n3535_ | ~new_n1074_;
  assign new_n3588_ = ~new_n1152_ | ~new_n1056_;
  assign new_n3589_ = ~new_n3534_ | ~new_n1055_;
  assign new_n3590_ = ~new_n1047_ | ~new_n3551_;
  assign new_n3591_ = ~pi165 | ~new_n3546_;
  assign new_n3592_ = ~new_n1998_;
  assign new_n3593_ = ~new_n1997_;
  assign new_n3594_ = ~new_n1097_ | ~new_n1102_;
  assign new_n3595_ = ~new_n1999_;
  assign new_n3596_ = ~new_n1883_;
  assign new_n3597_ = ~new_n3174_ | ~new_n1143_;
  assign new_n3598_ = ~new_n1155_ | ~new_n1015_;
  assign new_n3599_ = ~new_n1964_ | ~new_n3598_;
  assign new_n3600_ = ~new_n3595_ | ~new_n3599_;
  assign new_n3601_ = ~pi106 | ~new_n1997_;
  assign new_n3602_ = ~pi107 | ~new_n1883_;
  assign new_n3603_ = ~new_n3600_ | ~new_n2295_;
  assign new_n3604_ = ~new_n1155_ | ~new_n1045_;
  assign new_n3605_ = ~new_n1964_ | ~new_n3604_;
  assign new_n3606_ = ~new_n3605_ | ~new_n1999_;
  assign new_n3607_ = ~pi107 | ~new_n3596_;
  assign new_n3608_ = ~new_n3607_ | ~new_n3606_;
  assign new_n3609_ = ~new_n3593_ | ~new_n1072_;
  assign new_n3610_ = ~new_n1154_ | ~new_n1070_;
  assign new_n3611_ = ~new_n3592_ | ~new_n1069_;
  assign new_n3612_ = ~new_n1054_ | ~new_n3608_;
  assign new_n3613_ = ~pi166 | ~new_n3603_;
  assign new_n3614_ = ~new_n3593_ | ~new_n1073_;
  assign new_n3615_ = ~new_n1154_ | ~new_n1068_;
  assign new_n3616_ = ~new_n3592_ | ~new_n1067_;
  assign new_n3617_ = ~new_n1053_ | ~new_n3608_;
  assign new_n3618_ = ~pi167 | ~new_n3603_;
  assign new_n3619_ = ~new_n3593_ | ~new_n1077_;
  assign new_n3620_ = ~new_n1154_ | ~new_n1066_;
  assign new_n3621_ = ~new_n3592_ | ~new_n1065_;
  assign new_n3622_ = ~new_n1052_ | ~new_n3608_;
  assign new_n3623_ = ~pi168 | ~new_n3603_;
  assign new_n3624_ = ~new_n3593_ | ~new_n1076_;
  assign new_n3625_ = ~new_n1154_ | ~new_n1064_;
  assign new_n3626_ = ~new_n3592_ | ~new_n1063_;
  assign new_n3627_ = ~new_n1051_ | ~new_n3608_;
  assign new_n3628_ = ~pi169 | ~new_n3603_;
  assign new_n3629_ = ~new_n3593_ | ~new_n1075_;
  assign new_n3630_ = ~new_n1154_ | ~new_n1062_;
  assign new_n3631_ = ~new_n3592_ | ~new_n1061_;
  assign new_n3632_ = ~new_n1050_ | ~new_n3608_;
  assign new_n3633_ = ~pi170 | ~new_n3603_;
  assign new_n3634_ = ~new_n3593_ | ~new_n1078_;
  assign new_n3635_ = ~new_n1154_ | ~new_n1060_;
  assign new_n3636_ = ~new_n3592_ | ~new_n1059_;
  assign new_n3637_ = ~new_n1049_ | ~new_n3608_;
  assign new_n3638_ = ~pi171 | ~new_n3603_;
  assign new_n3639_ = ~new_n3593_ | ~new_n1071_;
  assign new_n3640_ = ~new_n1154_ | ~new_n1058_;
  assign new_n3641_ = ~new_n3592_ | ~new_n1057_;
  assign new_n3642_ = ~new_n1048_ | ~new_n3608_;
  assign new_n3643_ = ~pi172 | ~new_n3603_;
  assign new_n3644_ = ~new_n3593_ | ~new_n1074_;
  assign new_n3645_ = ~new_n1154_ | ~new_n1056_;
  assign new_n3646_ = ~new_n3592_ | ~new_n1055_;
  assign new_n3647_ = ~new_n1047_ | ~new_n3608_;
  assign new_n3648_ = ~pi173 | ~new_n3603_;
  assign new_n3649_ = ~new_n2003_;
  assign new_n3650_ = ~new_n1096_ | ~new_n1099_;
  assign new_n3651_ = ~new_n2005_;
  assign new_n3652_ = ~new_n1090_ | ~new_n1093_;
  assign new_n3653_ = ~new_n2006_;
  assign new_n3654_ = ~new_n1157_ | ~new_n1015_;
  assign new_n3655_ = ~new_n1964_ | ~new_n3654_;
  assign new_n3656_ = ~new_n3651_ | ~new_n3655_;
  assign new_n3657_ = ~pi106 | ~new_n2000_;
  assign new_n3658_ = ~new_n3653_ | ~pi107;
  assign new_n3659_ = ~new_n3656_ | ~new_n2304_;
  assign new_n3660_ = ~new_n1157_ | ~new_n1045_;
  assign new_n3661_ = ~new_n1964_ | ~new_n3660_;
  assign new_n3662_ = ~new_n3661_ | ~new_n2005_;
  assign new_n3663_ = ~pi107 | ~new_n2006_;
  assign new_n3664_ = ~new_n3663_ | ~new_n3662_;
  assign new_n3665_ = ~new_n3182_ | ~new_n1072_;
  assign new_n3666_ = ~new_n2883_ | ~new_n1070_;
  assign new_n3667_ = ~new_n3649_ | ~new_n1069_;
  assign new_n3668_ = ~new_n1054_ | ~new_n3664_;
  assign new_n3669_ = ~pi174 | ~new_n3659_;
  assign new_n3670_ = ~new_n3182_ | ~new_n1073_;
  assign new_n3671_ = ~new_n2883_ | ~new_n1068_;
  assign new_n3672_ = ~new_n3649_ | ~new_n1067_;
  assign new_n3673_ = ~new_n1053_ | ~new_n3664_;
  assign new_n3674_ = ~pi175 | ~new_n3659_;
  assign new_n3675_ = ~new_n3182_ | ~new_n1077_;
  assign new_n3676_ = ~new_n2883_ | ~new_n1066_;
  assign new_n3677_ = ~new_n3649_ | ~new_n1065_;
  assign new_n3678_ = ~new_n1052_ | ~new_n3664_;
  assign new_n3679_ = ~pi176 | ~new_n3659_;
  assign new_n3680_ = ~new_n3182_ | ~new_n1076_;
  assign new_n3681_ = ~new_n2883_ | ~new_n1064_;
  assign new_n3682_ = ~new_n3649_ | ~new_n1063_;
  assign new_n3683_ = ~new_n1051_ | ~new_n3664_;
  assign new_n3684_ = ~pi177 | ~new_n3659_;
  assign new_n3685_ = ~new_n3182_ | ~new_n1075_;
  assign new_n3686_ = ~new_n2883_ | ~new_n1062_;
  assign new_n3687_ = ~new_n3649_ | ~new_n1061_;
  assign new_n3688_ = ~new_n1050_ | ~new_n3664_;
  assign new_n3689_ = ~pi178 | ~new_n3659_;
  assign new_n3690_ = ~new_n3182_ | ~new_n1078_;
  assign new_n3691_ = ~new_n2883_ | ~new_n1060_;
  assign new_n3692_ = ~new_n3649_ | ~new_n1059_;
  assign new_n3693_ = ~new_n1049_ | ~new_n3664_;
  assign new_n3694_ = ~pi179 | ~new_n3659_;
  assign new_n3695_ = ~new_n3182_ | ~new_n1071_;
  assign new_n3696_ = ~new_n2883_ | ~new_n1058_;
  assign new_n3697_ = ~new_n3649_ | ~new_n1057_;
  assign new_n3698_ = ~new_n1048_ | ~new_n3664_;
  assign new_n3699_ = ~pi180 | ~new_n3659_;
  assign new_n3700_ = ~new_n3182_ | ~new_n1074_;
  assign new_n3701_ = ~new_n2883_ | ~new_n1056_;
  assign new_n3702_ = ~new_n3649_ | ~new_n1055_;
  assign new_n3703_ = ~new_n1047_ | ~new_n3664_;
  assign new_n3704_ = ~pi181 | ~new_n3659_;
  assign new_n3705_ = ~new_n2008_;
  assign new_n3706_ = ~new_n2007_;
  assign new_n3707_ = ~new_n1096_ | ~new_n1100_;
  assign new_n3708_ = ~new_n2009_;
  assign new_n3709_ = ~new_n1884_;
  assign new_n3710_ = ~new_n3169_ | ~new_n1131_;
  assign new_n3711_ = ~new_n1159_ | ~new_n1015_;
  assign new_n3712_ = ~new_n1964_ | ~new_n3711_;
  assign new_n3713_ = ~new_n3708_ | ~new_n3712_;
  assign new_n3714_ = ~pi106 | ~new_n2007_;
  assign new_n3715_ = ~pi107 | ~new_n1884_;
  assign new_n3716_ = ~new_n3713_ | ~new_n2313_;
  assign new_n3717_ = ~new_n1159_ | ~new_n1045_;
  assign new_n3718_ = ~new_n1964_ | ~new_n3717_;
  assign new_n3719_ = ~new_n3718_ | ~new_n2009_;
  assign new_n3720_ = ~pi107 | ~new_n3709_;
  assign new_n3721_ = ~new_n3720_ | ~new_n3719_;
  assign new_n3722_ = ~new_n3706_ | ~new_n1072_;
  assign new_n3723_ = ~new_n1158_ | ~new_n1070_;
  assign new_n3724_ = ~new_n3705_ | ~new_n1069_;
  assign new_n3725_ = ~new_n1054_ | ~new_n3721_;
  assign new_n3726_ = ~pi182 | ~new_n3716_;
  assign new_n3727_ = ~new_n3706_ | ~new_n1073_;
  assign new_n3728_ = ~new_n1158_ | ~new_n1068_;
  assign new_n3729_ = ~new_n3705_ | ~new_n1067_;
  assign new_n3730_ = ~new_n1053_ | ~new_n3721_;
  assign new_n3731_ = ~pi183 | ~new_n3716_;
  assign new_n3732_ = ~new_n3706_ | ~new_n1077_;
  assign new_n3733_ = ~new_n1158_ | ~new_n1066_;
  assign new_n3734_ = ~new_n3705_ | ~new_n1065_;
  assign new_n3735_ = ~new_n1052_ | ~new_n3721_;
  assign new_n3736_ = ~pi184 | ~new_n3716_;
  assign new_n3737_ = ~new_n3706_ | ~new_n1076_;
  assign new_n3738_ = ~new_n1158_ | ~new_n1064_;
  assign new_n3739_ = ~new_n3705_ | ~new_n1063_;
  assign new_n3740_ = ~new_n1051_ | ~new_n3721_;
  assign new_n3741_ = ~pi185 | ~new_n3716_;
  assign new_n3742_ = ~new_n3706_ | ~new_n1075_;
  assign new_n3743_ = ~new_n1158_ | ~new_n1062_;
  assign new_n3744_ = ~new_n3705_ | ~new_n1061_;
  assign new_n3745_ = ~new_n1050_ | ~new_n3721_;
  assign new_n3746_ = ~pi186 | ~new_n3716_;
  assign new_n3747_ = ~new_n3706_ | ~new_n1078_;
  assign new_n3748_ = ~new_n1158_ | ~new_n1060_;
  assign new_n3749_ = ~new_n3705_ | ~new_n1059_;
  assign new_n3750_ = ~new_n1049_ | ~new_n3721_;
  assign new_n3751_ = ~pi187 | ~new_n3716_;
  assign new_n3752_ = ~new_n3706_ | ~new_n1071_;
  assign new_n3753_ = ~new_n1158_ | ~new_n1058_;
  assign new_n3754_ = ~new_n3705_ | ~new_n1057_;
  assign new_n3755_ = ~new_n1048_ | ~new_n3721_;
  assign new_n3756_ = ~pi188 | ~new_n3716_;
  assign new_n3757_ = ~new_n3706_ | ~new_n1074_;
  assign new_n3758_ = ~new_n1158_ | ~new_n1056_;
  assign new_n3759_ = ~new_n3705_ | ~new_n1055_;
  assign new_n3760_ = ~new_n1047_ | ~new_n3721_;
  assign new_n3761_ = ~pi189 | ~new_n3716_;
  assign new_n3762_ = ~new_n2011_;
  assign new_n3763_ = ~new_n2010_;
  assign new_n3764_ = ~new_n1096_ | ~new_n1101_;
  assign new_n3765_ = ~new_n2012_;
  assign new_n3766_ = ~new_n1090_ | ~new_n1094_;
  assign new_n3767_ = ~new_n2013_;
  assign new_n3768_ = ~new_n3170_ | ~new_n1131_;
  assign new_n3769_ = ~new_n1161_ | ~new_n1015_;
  assign new_n3770_ = ~new_n1964_ | ~new_n3769_;
  assign new_n3771_ = ~new_n3765_ | ~new_n3770_;
  assign new_n3772_ = ~pi106 | ~new_n2010_;
  assign new_n3773_ = ~new_n3767_ | ~pi107;
  assign new_n3774_ = ~new_n3771_ | ~new_n2322_;
  assign new_n3775_ = ~new_n1161_ | ~new_n1045_;
  assign new_n3776_ = ~new_n1964_ | ~new_n3775_;
  assign new_n3777_ = ~new_n3776_ | ~new_n2012_;
  assign new_n3778_ = ~pi107 | ~new_n2013_;
  assign new_n3779_ = ~new_n3778_ | ~new_n3777_;
  assign new_n3780_ = ~new_n3763_ | ~new_n1072_;
  assign new_n3781_ = ~new_n1160_ | ~new_n1070_;
  assign new_n3782_ = ~new_n3762_ | ~new_n1069_;
  assign new_n3783_ = ~new_n1054_ | ~new_n3779_;
  assign new_n3784_ = ~pi190 | ~new_n3774_;
  assign new_n3785_ = ~new_n3763_ | ~new_n1073_;
  assign new_n3786_ = ~new_n1160_ | ~new_n1068_;
  assign new_n3787_ = ~new_n3762_ | ~new_n1067_;
  assign new_n3788_ = ~new_n1053_ | ~new_n3779_;
  assign new_n3789_ = ~pi191 | ~new_n3774_;
  assign new_n3790_ = ~new_n3763_ | ~new_n1077_;
  assign new_n3791_ = ~new_n1160_ | ~new_n1066_;
  assign new_n3792_ = ~new_n3762_ | ~new_n1065_;
  assign new_n3793_ = ~new_n1052_ | ~new_n3779_;
  assign new_n3794_ = ~pi192 | ~new_n3774_;
  assign new_n3795_ = ~new_n3763_ | ~new_n1076_;
  assign new_n3796_ = ~new_n1160_ | ~new_n1064_;
  assign new_n3797_ = ~new_n3762_ | ~new_n1063_;
  assign new_n3798_ = ~new_n1051_ | ~new_n3779_;
  assign new_n3799_ = ~pi193 | ~new_n3774_;
  assign new_n3800_ = ~new_n3763_ | ~new_n1075_;
  assign new_n3801_ = ~new_n1160_ | ~new_n1062_;
  assign new_n3802_ = ~new_n3762_ | ~new_n1061_;
  assign new_n3803_ = ~new_n1050_ | ~new_n3779_;
  assign new_n3804_ = ~pi194 | ~new_n3774_;
  assign new_n3805_ = ~new_n3763_ | ~new_n1078_;
  assign new_n3806_ = ~new_n1160_ | ~new_n1060_;
  assign new_n3807_ = ~new_n3762_ | ~new_n1059_;
  assign new_n3808_ = ~new_n1049_ | ~new_n3779_;
  assign new_n3809_ = ~pi195 | ~new_n3774_;
  assign new_n3810_ = ~new_n3763_ | ~new_n1071_;
  assign new_n3811_ = ~new_n1160_ | ~new_n1058_;
  assign new_n3812_ = ~new_n3762_ | ~new_n1057_;
  assign new_n3813_ = ~new_n1048_ | ~new_n3779_;
  assign new_n3814_ = ~pi196 | ~new_n3774_;
  assign new_n3815_ = ~new_n3763_ | ~new_n1074_;
  assign new_n3816_ = ~new_n1160_ | ~new_n1056_;
  assign new_n3817_ = ~new_n3762_ | ~new_n1055_;
  assign new_n3818_ = ~new_n1047_ | ~new_n3779_;
  assign new_n3819_ = ~pi197 | ~new_n3774_;
  assign new_n3820_ = ~new_n2015_;
  assign new_n3821_ = ~new_n2014_;
  assign new_n3822_ = ~new_n1096_ | ~new_n1102_;
  assign new_n3823_ = ~new_n2016_;
  assign new_n3824_ = ~new_n1885_;
  assign new_n3825_ = ~new_n1143_ | ~new_n1131_;
  assign new_n3826_ = ~new_n1163_ | ~new_n1015_;
  assign new_n3827_ = ~new_n1964_ | ~new_n3826_;
  assign new_n3828_ = ~new_n3823_ | ~new_n3827_;
  assign new_n3829_ = ~pi106 | ~new_n2014_;
  assign new_n3830_ = ~pi107 | ~new_n1885_;
  assign new_n3831_ = ~new_n3828_ | ~new_n2331_;
  assign new_n3832_ = ~new_n1163_ | ~new_n1045_;
  assign new_n3833_ = ~new_n1964_ | ~new_n3832_;
  assign new_n3834_ = ~new_n3833_ | ~new_n2016_;
  assign new_n3835_ = ~pi107 | ~new_n3824_;
  assign new_n3836_ = ~new_n3835_ | ~new_n3834_;
  assign new_n3837_ = ~new_n3821_ | ~new_n1072_;
  assign new_n3838_ = ~new_n1162_ | ~new_n1070_;
  assign new_n3839_ = ~new_n3820_ | ~new_n1069_;
  assign new_n3840_ = ~new_n1054_ | ~new_n3836_;
  assign new_n3841_ = ~pi198 | ~new_n3831_;
  assign new_n3842_ = ~new_n3821_ | ~new_n1073_;
  assign new_n3843_ = ~new_n1162_ | ~new_n1068_;
  assign new_n3844_ = ~new_n3820_ | ~new_n1067_;
  assign new_n3845_ = ~new_n1053_ | ~new_n3836_;
  assign new_n3846_ = ~pi199 | ~new_n3831_;
  assign new_n3847_ = ~new_n3821_ | ~new_n1077_;
  assign new_n3848_ = ~new_n1162_ | ~new_n1066_;
  assign new_n3849_ = ~new_n3820_ | ~new_n1065_;
  assign new_n3850_ = ~new_n1052_ | ~new_n3836_;
  assign new_n3851_ = ~pi200 | ~new_n3831_;
  assign new_n3852_ = ~new_n3821_ | ~new_n1076_;
  assign new_n3853_ = ~new_n1162_ | ~new_n1064_;
  assign new_n3854_ = ~new_n3820_ | ~new_n1063_;
  assign new_n3855_ = ~new_n1051_ | ~new_n3836_;
  assign new_n3856_ = ~pi201 | ~new_n3831_;
  assign new_n3857_ = ~new_n3821_ | ~new_n1075_;
  assign new_n3858_ = ~new_n1162_ | ~new_n1062_;
  assign new_n3859_ = ~new_n3820_ | ~new_n1061_;
  assign new_n3860_ = ~new_n1050_ | ~new_n3836_;
  assign new_n3861_ = ~pi202 | ~new_n3831_;
  assign new_n3862_ = ~new_n3821_ | ~new_n1078_;
  assign new_n3863_ = ~new_n1162_ | ~new_n1060_;
  assign new_n3864_ = ~new_n3820_ | ~new_n1059_;
  assign new_n3865_ = ~new_n1049_ | ~new_n3836_;
  assign new_n3866_ = ~pi203 | ~new_n3831_;
  assign new_n3867_ = ~new_n3821_ | ~new_n1071_;
  assign new_n3868_ = ~new_n1162_ | ~new_n1058_;
  assign new_n3869_ = ~new_n3820_ | ~new_n1057_;
  assign new_n3870_ = ~new_n1048_ | ~new_n3836_;
  assign new_n3871_ = ~pi204 | ~new_n3831_;
  assign new_n3872_ = ~new_n3821_ | ~new_n1074_;
  assign new_n3873_ = ~new_n1162_ | ~new_n1056_;
  assign new_n3874_ = ~new_n3820_ | ~new_n1055_;
  assign new_n3875_ = ~new_n1047_ | ~new_n3836_;
  assign new_n3876_ = ~pi205 | ~new_n3831_;
  assign new_n3877_ = ~new_n2018_;
  assign new_n3878_ = ~new_n2017_;
  assign new_n3879_ = ~new_n1098_ | ~new_n1099_;
  assign new_n3880_ = ~new_n2019_;
  assign new_n3881_ = ~new_n1092_ | ~new_n1093_;
  assign new_n3882_ = ~new_n2020_;
  assign new_n3883_ = ~new_n1165_ | ~new_n3173_;
  assign new_n3884_ = ~new_n1168_ | ~new_n1015_;
  assign new_n3885_ = ~new_n1964_ | ~new_n3884_;
  assign new_n3886_ = ~new_n3880_ | ~new_n3885_;
  assign new_n3887_ = ~pi106 | ~new_n2017_;
  assign new_n3888_ = ~new_n3882_ | ~pi107;
  assign new_n3889_ = ~new_n3886_ | ~new_n2340_;
  assign new_n3890_ = ~new_n1168_ | ~new_n1045_;
  assign new_n3891_ = ~new_n1964_ | ~new_n3890_;
  assign new_n3892_ = ~new_n3891_ | ~new_n2019_;
  assign new_n3893_ = ~pi107 | ~new_n2020_;
  assign new_n3894_ = ~new_n3893_ | ~new_n3892_;
  assign new_n3895_ = ~new_n3878_ | ~new_n1072_;
  assign new_n3896_ = ~new_n1166_ | ~new_n1070_;
  assign new_n3897_ = ~new_n3877_ | ~new_n1069_;
  assign new_n3898_ = ~new_n1054_ | ~new_n3894_;
  assign new_n3899_ = ~pi206 | ~new_n3889_;
  assign new_n3900_ = ~new_n3878_ | ~new_n1073_;
  assign new_n3901_ = ~new_n1166_ | ~new_n1068_;
  assign new_n3902_ = ~new_n3877_ | ~new_n1067_;
  assign new_n3903_ = ~new_n1053_ | ~new_n3894_;
  assign new_n3904_ = ~pi207 | ~new_n3889_;
  assign new_n3905_ = ~new_n3878_ | ~new_n1077_;
  assign new_n3906_ = ~new_n1166_ | ~new_n1066_;
  assign new_n3907_ = ~new_n3877_ | ~new_n1065_;
  assign new_n3908_ = ~new_n1052_ | ~new_n3894_;
  assign new_n3909_ = ~pi208 | ~new_n3889_;
  assign new_n3910_ = ~new_n3878_ | ~new_n1076_;
  assign new_n3911_ = ~new_n1166_ | ~new_n1064_;
  assign new_n3912_ = ~new_n3877_ | ~new_n1063_;
  assign new_n3913_ = ~new_n1051_ | ~new_n3894_;
  assign new_n3914_ = ~pi209 | ~new_n3889_;
  assign new_n3915_ = ~new_n3878_ | ~new_n1075_;
  assign new_n3916_ = ~new_n1166_ | ~new_n1062_;
  assign new_n3917_ = ~new_n3877_ | ~new_n1061_;
  assign new_n3918_ = ~new_n1050_ | ~new_n3894_;
  assign new_n3919_ = ~pi210 | ~new_n3889_;
  assign new_n3920_ = ~new_n3878_ | ~new_n1078_;
  assign new_n3921_ = ~new_n1166_ | ~new_n1060_;
  assign new_n3922_ = ~new_n3877_ | ~new_n1059_;
  assign new_n3923_ = ~new_n1049_ | ~new_n3894_;
  assign new_n3924_ = ~pi211 | ~new_n3889_;
  assign new_n3925_ = ~new_n3878_ | ~new_n1071_;
  assign new_n3926_ = ~new_n1166_ | ~new_n1058_;
  assign new_n3927_ = ~new_n3877_ | ~new_n1057_;
  assign new_n3928_ = ~new_n1048_ | ~new_n3894_;
  assign new_n3929_ = ~pi212 | ~new_n3889_;
  assign new_n3930_ = ~new_n3878_ | ~new_n1074_;
  assign new_n3931_ = ~new_n1166_ | ~new_n1056_;
  assign new_n3932_ = ~new_n3877_ | ~new_n1055_;
  assign new_n3933_ = ~new_n1047_ | ~new_n3894_;
  assign new_n3934_ = ~pi213 | ~new_n3889_;
  assign new_n3935_ = ~new_n2022_;
  assign new_n3936_ = ~new_n2021_;
  assign new_n3937_ = ~new_n1098_ | ~new_n1100_;
  assign new_n3938_ = ~new_n2023_;
  assign new_n3939_ = ~new_n1886_;
  assign new_n3940_ = ~new_n1165_ | ~new_n3169_;
  assign new_n3941_ = ~new_n1170_ | ~new_n1015_;
  assign new_n3942_ = ~new_n1964_ | ~new_n3941_;
  assign new_n3943_ = ~new_n3938_ | ~new_n3942_;
  assign new_n3944_ = ~pi106 | ~new_n2021_;
  assign new_n3945_ = ~pi107 | ~new_n1886_;
  assign new_n3946_ = ~new_n3943_ | ~new_n2349_;
  assign new_n3947_ = ~new_n1170_ | ~new_n1045_;
  assign new_n3948_ = ~new_n1964_ | ~new_n3947_;
  assign new_n3949_ = ~new_n3948_ | ~new_n2023_;
  assign new_n3950_ = ~pi107 | ~new_n3939_;
  assign new_n3951_ = ~new_n3950_ | ~new_n3949_;
  assign new_n3952_ = ~new_n3936_ | ~new_n1072_;
  assign new_n3953_ = ~new_n1169_ | ~new_n1070_;
  assign new_n3954_ = ~new_n3935_ | ~new_n1069_;
  assign new_n3955_ = ~new_n1054_ | ~new_n3951_;
  assign new_n3956_ = ~pi214 | ~new_n3946_;
  assign new_n3957_ = ~new_n3936_ | ~new_n1073_;
  assign new_n3958_ = ~new_n1169_ | ~new_n1068_;
  assign new_n3959_ = ~new_n3935_ | ~new_n1067_;
  assign new_n3960_ = ~new_n1053_ | ~new_n3951_;
  assign new_n3961_ = ~pi215 | ~new_n3946_;
  assign new_n3962_ = ~new_n3936_ | ~new_n1077_;
  assign new_n3963_ = ~new_n1169_ | ~new_n1066_;
  assign new_n3964_ = ~new_n3935_ | ~new_n1065_;
  assign new_n3965_ = ~new_n1052_ | ~new_n3951_;
  assign new_n3966_ = ~pi216 | ~new_n3946_;
  assign new_n3967_ = ~new_n3936_ | ~new_n1076_;
  assign new_n3968_ = ~new_n1169_ | ~new_n1064_;
  assign new_n3969_ = ~new_n3935_ | ~new_n1063_;
  assign new_n3970_ = ~new_n1051_ | ~new_n3951_;
  assign new_n3971_ = ~pi217 | ~new_n3946_;
  assign new_n3972_ = ~new_n3936_ | ~new_n1075_;
  assign new_n3973_ = ~new_n1169_ | ~new_n1062_;
  assign new_n3974_ = ~new_n3935_ | ~new_n1061_;
  assign new_n3975_ = ~new_n1050_ | ~new_n3951_;
  assign new_n3976_ = ~pi218 | ~new_n3946_;
  assign new_n3977_ = ~new_n3936_ | ~new_n1078_;
  assign new_n3978_ = ~new_n1169_ | ~new_n1060_;
  assign new_n3979_ = ~new_n3935_ | ~new_n1059_;
  assign new_n3980_ = ~new_n1049_ | ~new_n3951_;
  assign new_n3981_ = ~pi219 | ~new_n3946_;
  assign new_n3982_ = ~new_n3936_ | ~new_n1071_;
  assign new_n3983_ = ~new_n1169_ | ~new_n1058_;
  assign new_n3984_ = ~new_n3935_ | ~new_n1057_;
  assign new_n3985_ = ~new_n1048_ | ~new_n3951_;
  assign new_n3986_ = ~pi220 | ~new_n3946_;
  assign new_n3987_ = ~new_n3936_ | ~new_n1074_;
  assign new_n3988_ = ~new_n1169_ | ~new_n1056_;
  assign new_n3989_ = ~new_n3935_ | ~new_n1055_;
  assign new_n3990_ = ~new_n1047_ | ~new_n3951_;
  assign new_n3991_ = ~pi221 | ~new_n3946_;
  assign new_n3992_ = ~new_n2025_;
  assign new_n3993_ = ~new_n2024_;
  assign new_n3994_ = ~new_n1098_ | ~new_n1101_;
  assign new_n3995_ = ~new_n2026_;
  assign new_n3996_ = ~new_n1092_ | ~new_n1094_;
  assign new_n3997_ = ~new_n2027_;
  assign new_n3998_ = ~new_n1165_ | ~new_n3170_;
  assign new_n3999_ = ~new_n1172_ | ~new_n1015_;
  assign new_n4000_ = ~new_n1964_ | ~new_n3999_;
  assign new_n4001_ = ~new_n3995_ | ~new_n4000_;
  assign new_n4002_ = ~pi106 | ~new_n2024_;
  assign new_n4003_ = ~new_n3997_ | ~pi107;
  assign new_n4004_ = ~new_n4001_ | ~new_n2358_;
  assign new_n4005_ = ~new_n1172_ | ~new_n1045_;
  assign new_n4006_ = ~new_n1964_ | ~new_n4005_;
  assign new_n4007_ = ~new_n4006_ | ~new_n2026_;
  assign new_n4008_ = ~pi107 | ~new_n2027_;
  assign new_n4009_ = ~new_n4008_ | ~new_n4007_;
  assign new_n4010_ = ~new_n3993_ | ~new_n1072_;
  assign new_n4011_ = ~new_n1171_ | ~new_n1070_;
  assign new_n4012_ = ~new_n3992_ | ~new_n1069_;
  assign new_n4013_ = ~new_n1054_ | ~new_n4009_;
  assign new_n4014_ = ~pi222 | ~new_n4004_;
  assign new_n4015_ = ~new_n3993_ | ~new_n1073_;
  assign new_n4016_ = ~new_n1171_ | ~new_n1068_;
  assign new_n4017_ = ~new_n3992_ | ~new_n1067_;
  assign new_n4018_ = ~new_n1053_ | ~new_n4009_;
  assign new_n4019_ = ~pi223 | ~new_n4004_;
  assign new_n4020_ = ~new_n3993_ | ~new_n1077_;
  assign new_n4021_ = ~new_n1171_ | ~new_n1066_;
  assign new_n4022_ = ~new_n3992_ | ~new_n1065_;
  assign new_n4023_ = ~new_n1052_ | ~new_n4009_;
  assign new_n4024_ = ~pi224 | ~new_n4004_;
  assign new_n4025_ = ~new_n3993_ | ~new_n1076_;
  assign new_n4026_ = ~new_n1171_ | ~new_n1064_;
  assign new_n4027_ = ~new_n3992_ | ~new_n1063_;
  assign new_n4028_ = ~new_n1051_ | ~new_n4009_;
  assign new_n4029_ = ~pi225 | ~new_n4004_;
  assign new_n4030_ = ~new_n3993_ | ~new_n1075_;
  assign new_n4031_ = ~new_n1171_ | ~new_n1062_;
  assign new_n4032_ = ~new_n3992_ | ~new_n1061_;
  assign new_n4033_ = ~new_n1050_ | ~new_n4009_;
  assign new_n4034_ = ~pi226 | ~new_n4004_;
  assign new_n4035_ = ~new_n3993_ | ~new_n1078_;
  assign new_n4036_ = ~new_n1171_ | ~new_n1060_;
  assign new_n4037_ = ~new_n3992_ | ~new_n1059_;
  assign new_n4038_ = ~new_n1049_ | ~new_n4009_;
  assign new_n4039_ = ~pi227 | ~new_n4004_;
  assign new_n4040_ = ~new_n3993_ | ~new_n1071_;
  assign new_n4041_ = ~new_n1171_ | ~new_n1058_;
  assign new_n4042_ = ~new_n3992_ | ~new_n1057_;
  assign new_n4043_ = ~new_n1048_ | ~new_n4009_;
  assign new_n4044_ = ~pi228 | ~new_n4004_;
  assign new_n4045_ = ~new_n3993_ | ~new_n1074_;
  assign new_n4046_ = ~new_n1171_ | ~new_n1056_;
  assign new_n4047_ = ~new_n3992_ | ~new_n1055_;
  assign new_n4048_ = ~new_n1047_ | ~new_n4009_;
  assign new_n4049_ = ~pi229 | ~new_n4004_;
  assign new_n4050_ = ~new_n2029_;
  assign new_n4051_ = ~new_n2028_;
  assign new_n4052_ = ~new_n1098_ | ~new_n1102_;
  assign new_n4053_ = ~new_n2030_;
  assign new_n4054_ = ~new_n1887_;
  assign new_n4055_ = ~new_n1165_ | ~new_n1143_;
  assign new_n4056_ = ~new_n1174_ | ~new_n1015_;
  assign new_n4057_ = ~new_n1964_ | ~new_n4056_;
  assign new_n4058_ = ~new_n4053_ | ~new_n4057_;
  assign new_n4059_ = ~pi106 | ~new_n2028_;
  assign new_n4060_ = ~pi107 | ~new_n1887_;
  assign new_n4061_ = ~new_n4058_ | ~new_n2367_;
  assign new_n4062_ = ~new_n1174_ | ~new_n1045_;
  assign new_n4063_ = ~new_n1964_ | ~new_n4062_;
  assign new_n4064_ = ~new_n4063_ | ~new_n2030_;
  assign new_n4065_ = ~pi107 | ~new_n4054_;
  assign new_n4066_ = ~new_n4065_ | ~new_n4064_;
  assign new_n4067_ = ~new_n4051_ | ~new_n1072_;
  assign new_n4068_ = ~new_n1173_ | ~new_n1070_;
  assign new_n4069_ = ~new_n4050_ | ~new_n1069_;
  assign new_n4070_ = ~new_n1054_ | ~new_n4066_;
  assign new_n4071_ = ~pi230 | ~new_n4061_;
  assign new_n4072_ = ~new_n4051_ | ~new_n1073_;
  assign new_n4073_ = ~new_n1173_ | ~new_n1068_;
  assign new_n4074_ = ~new_n4050_ | ~new_n1067_;
  assign new_n4075_ = ~new_n1053_ | ~new_n4066_;
  assign new_n4076_ = ~pi231 | ~new_n4061_;
  assign new_n4077_ = ~new_n4051_ | ~new_n1077_;
  assign new_n4078_ = ~new_n1173_ | ~new_n1066_;
  assign new_n4079_ = ~new_n4050_ | ~new_n1065_;
  assign new_n4080_ = ~new_n1052_ | ~new_n4066_;
  assign new_n4081_ = ~pi232 | ~new_n4061_;
  assign new_n4082_ = ~new_n4051_ | ~new_n1076_;
  assign new_n4083_ = ~new_n1173_ | ~new_n1064_;
  assign new_n4084_ = ~new_n4050_ | ~new_n1063_;
  assign new_n4085_ = ~new_n1051_ | ~new_n4066_;
  assign new_n4086_ = ~new_n4051_ | ~new_n1075_;
  assign new_n4087_ = ~new_n1173_ | ~new_n1062_;
  assign new_n4088_ = ~new_n4050_ | ~new_n1061_;
  assign new_n4089_ = ~new_n1050_ | ~new_n4066_;
  assign new_n4090_ = ~pi234 | ~new_n4061_;
  assign new_n4091_ = ~new_n4051_ | ~new_n1078_;
  assign new_n4092_ = ~new_n1173_ | ~new_n1060_;
  assign new_n4093_ = ~new_n4050_ | ~new_n1059_;
  assign new_n4094_ = ~new_n1049_ | ~new_n4066_;
  assign new_n4095_ = ~pi235 | ~new_n4061_;
  assign new_n4096_ = ~new_n4051_ | ~new_n1071_;
  assign new_n4097_ = ~new_n1173_ | ~new_n1058_;
  assign new_n4098_ = ~new_n4050_ | ~new_n1057_;
  assign new_n4099_ = ~new_n1048_ | ~new_n4066_;
  assign new_n4100_ = ~pi236 | ~new_n4061_;
  assign new_n4101_ = ~new_n4051_ | ~new_n1074_;
  assign new_n4102_ = ~new_n1173_ | ~new_n1056_;
  assign new_n4103_ = ~new_n4050_ | ~new_n1055_;
  assign new_n4104_ = ~new_n1047_ | ~new_n4066_;
  assign new_n4105_ = ~pi237 | ~new_n4061_;
  assign new_n4106_ = ~new_n2067_;
  assign new_n4107_ = ~new_n3148_ | ~new_n2035_ | ~new_n2038_;
  assign new_n4108_ = ~new_n3105_ | ~new_n3045_ | ~new_n2818_;
  assign new_n4109_ = ~new_n1888_;
  assign new_n4110_ = ~new_n3139_ | ~new_n1933_;
  assign new_n4111_ = ~new_n4109_ | ~new_n4110_ | ~new_n1927_;
  assign new_n4112_ = ~new_n2377_ | ~new_n1109_;
  assign new_n4113_ = ~new_n2853_ | ~new_n4107_;
  assign new_n4114_ = ~new_n2378_ | ~new_n6254_;
  assign new_n4115_ = ~new_n9223_ | ~new_n2860_ | ~new_n1901_;
  assign new_n4116_ = ~new_n1106_ | ~new_n6139_;
  assign new_n4117_ = ~new_n2902_ | ~new_n3148_;
  assign new_n4118_ = ~new_n2827_;
  assign new_n4119_ = ~new_n1025_ | ~new_n2827_;
  assign new_n4120_ = ~pi106 | ~new_n1938_;
  assign new_n4121_ = ~new_n2817_;
  assign new_n4122_ = ~pi241 | ~pi240;
  assign new_n4123_ = ~pi239 | ~new_n4122_;
  assign new_n4124_ = ~new_n3026_ | ~pi241;
  assign new_n4125_ = ~new_n2086_;
  assign new_n4126_ = ~new_n2143_ | ~pi240;
  assign new_n4127_ = ~pi239 | ~new_n4126_;
  assign new_n4128_ = ~new_n2082_;
  assign new_n4129_ = ~new_n1919_ | ~new_n1908_;
  assign new_n4130_ = ~pi239 | ~new_n4129_;
  assign new_n4131_ = ~new_n1126_ | ~new_n1919_;
  assign new_n4132_ = ~new_n3139_ | ~new_n1934_;
  assign new_n4133_ = ~new_n3045_ | ~new_n1262_;
  assign new_n4134_ = ~new_n6139_ | ~new_n6349_ | ~new_n6348_;
  assign new_n4135_ = ~new_n3094_ | ~new_n4133_;
  assign new_n4136_ = ~new_n2053_ | ~new_n3045_ | ~new_n2038_;
  assign new_n4137_ = ~new_n4136_ | ~new_n2816_;
  assign new_n4138_ = ~new_n6274_ | ~new_n4137_;
  assign new_n4139_ = ~new_n3105_ | ~new_n2816_;
  assign new_n4140_ = ~new_n2039_ | ~new_n4139_;
  assign new_n4141_ = ~new_n2853_ | ~new_n4107_;
  assign new_n4142_ = ~new_n2902_ | ~new_n3148_;
  assign new_n4143_ = ~new_n4140_ | ~new_n1915_;
  assign new_n4144_ = ~new_n3139_ | ~new_n6352_;
  assign new_n4145_ = ~new_n2835_ | ~new_n1888_;
  assign new_n4146_ = ~new_n1936_ | ~new_n2862_;
  assign new_n4147_ = ~new_n2385_ | ~new_n4146_;
  assign new_n4148_ = ~new_n7942_ | ~new_n6154_;
  assign new_n4149_ = ~new_n2863_ | ~new_n2082_;
  assign new_n4150_ = ~new_n2859_ | ~new_n2086_;
  assign new_n4151_ = ~new_n4148_ | ~new_n2392_;
  assign new_n4152_ = ~new_n2897_ | ~new_n2082_;
  assign new_n4153_ = ~new_n1084_ | ~new_n4151_;
  assign new_n4154_ = ~new_n4153_ | ~new_n4152_;
  assign new_n4155_ = ~pi240 | ~new_n1919_;
  assign new_n4156_ = ~new_n2045_;
  assign new_n4157_ = ~new_n7959_ | ~new_n6154_;
  assign new_n4158_ = ~new_n2859_ | ~new_n2100_;
  assign new_n4159_ = ~new_n2394_ | ~new_n4157_;
  assign new_n4160_ = ~new_n1103_ | ~new_n2114_;
  assign new_n4161_ = ~new_n2897_ | ~new_n2045_;
  assign new_n4162_ = ~new_n1084_ | ~new_n4159_;
  assign new_n4163_ = ~new_n4161_ | ~new_n4162_ | ~new_n4160_;
  assign new_n4164_ = ~new_n2046_;
  assign new_n4165_ = ~new_n1088_ | ~new_n2894_;
  assign new_n4166_ = ~new_n1936_ | ~new_n4165_;
  assign new_n4167_ = ~new_n4164_ | ~new_n4166_;
  assign new_n4168_ = ~new_n7950_ | ~new_n6154_;
  assign new_n4169_ = ~new_n2859_ | ~new_n1909_;
  assign new_n4170_ = ~new_n2395_ | ~new_n4168_;
  assign new_n4171_ = ~new_n6357_ | ~new_n1103_;
  assign new_n4172_ = ~new_n4164_ | ~new_n2897_;
  assign new_n4173_ = ~new_n1084_ | ~new_n4170_;
  assign new_n4174_ = ~new_n4172_ | ~new_n4173_ | ~new_n4171_;
  assign new_n4175_ = ~new_n7951_ | ~new_n6154_;
  assign new_n4176_ = ~new_n2820_ | ~new_n4175_;
  assign new_n4177_ = ~new_n2897_ | ~new_n1910_;
  assign new_n4178_ = ~new_n1084_ | ~new_n4176_;
  assign new_n4179_ = ~new_n6360_ | ~pi108;
  assign new_n4180_ = ~new_n4177_ | ~new_n4178_ | ~new_n4179_;
  assign new_n4181_ = ~new_n8260_ | ~new_n1085_ | ~pi109;
  assign new_n4182_ = ~new_n2048_;
  assign new_n4183_ = ~pi108 | ~new_n1940_;
  assign new_n4184_ = ~new_n3172_ | ~new_n2098_;
  assign new_n4185_ = ~new_n2002_ | ~new_n4184_;
  assign new_n4186_ = ~new_n2003_ | ~new_n4185_;
  assign new_n4187_ = ~new_n1045_ | ~new_n4186_;
  assign new_n4188_ = ~new_n7942_ | ~new_n4183_;
  assign new_n4189_ = ~new_n2871_ | ~new_n8007_;
  assign new_n4190_ = ~new_n2396_ | ~new_n4187_;
  assign new_n4191_ = ~new_n1045_ | ~new_n6378_;
  assign new_n4192_ = ~new_n7959_ | ~new_n4183_;
  assign new_n4193_ = ~new_n2871_ | ~new_n8048_;
  assign new_n4194_ = ~new_n2397_ | ~new_n4191_;
  assign new_n4195_ = ~new_n1970_ | ~new_n1977_;
  assign new_n4196_ = ~new_n1045_ | ~new_n4195_;
  assign new_n4197_ = ~new_n7950_ | ~new_n4183_;
  assign new_n4198_ = ~new_n2871_ | ~new_n8049_;
  assign new_n4199_ = ~new_n2398_ | ~new_n4196_;
  assign new_n4200_ = ~new_n7951_ | ~new_n4183_;
  assign new_n4201_ = ~new_n8042_ | ~new_n2854_;
  assign new_n4202_ = ~new_n2890_ | ~new_n4200_ | ~new_n4201_;
  assign new_n4203_ = ~new_n3122_ | ~new_n1916_;
  assign new_n4204_ = ~new_n2905_ | ~new_n1088_;
  assign new_n4205_ = ~new_n6387_ | ~new_n6388_ | ~new_n1175_ | ~new_n4204_;
  assign new_n4206_ = ~new_n2837_ | ~new_n2880_ | ~new_n3148_;
  assign new_n4207_ = ~new_n1025_ | ~new_n4205_;
  assign new_n4208_ = ~new_n2848_ | ~new_n1907_;
  assign new_n4209_ = ~new_n2058_;
  assign new_n4210_ = ~new_n2907_ | ~new_n2853_;
  assign new_n4211_ = ~new_n2901_ | ~new_n1046_;
  assign new_n4212_ = ~new_n2911_ | ~new_n2895_;
  assign new_n4213_ = ~new_n2909_ | ~new_n3139_;
  assign new_n4214_ = ~new_n2403_ | ~new_n1176_;
  assign new_n4215_ = ~new_n8349_ | ~new_n1037_;
  assign new_n4216_ = ~new_n6467_ | ~new_n1035_;
  assign new_n4217_ = ~new_n6677_ | ~new_n1034_;
  assign new_n4218_ = ~new_n9040_ | ~new_n1032_;
  assign new_n4219_ = ~pi248 | ~new_n1031_;
  assign new_n4220_ = ~pi439 | ~new_n1027_;
  assign new_n4221_ = ~new_n4209_ | ~pi248;
  assign new_n4222_ = ~new_n8350_ | ~new_n1037_;
  assign new_n4223_ = ~new_n6533_ | ~new_n1035_;
  assign new_n4224_ = ~new_n6702_ | ~new_n1034_;
  assign new_n4225_ = ~new_n9117_ | ~new_n1032_;
  assign new_n4226_ = ~new_n9225_ | ~new_n1031_;
  assign new_n4227_ = ~new_n1027_ | ~pi440;
  assign new_n4228_ = ~new_n4209_ | ~pi249;
  assign new_n4229_ = ~new_n8401_ | ~new_n1037_;
  assign new_n4230_ = ~new_n6522_ | ~new_n1035_;
  assign new_n4231_ = ~new_n6761_ | ~new_n1034_;
  assign new_n4232_ = ~new_n9041_ | ~new_n1032_;
  assign new_n4233_ = ~new_n9292_ | ~new_n1031_;
  assign new_n4234_ = ~new_n1027_ | ~pi441;
  assign new_n4235_ = ~pi250 | ~new_n4209_;
  assign new_n4236_ = ~new_n8305_ | ~new_n1037_;
  assign new_n4237_ = ~new_n6519_ | ~new_n1035_;
  assign new_n4238_ = ~new_n6752_ | ~new_n1034_;
  assign new_n4239_ = ~new_n9129_ | ~new_n1032_;
  assign new_n4240_ = ~new_n9289_ | ~new_n1031_;
  assign new_n4241_ = ~new_n1027_ | ~pi442;
  assign new_n4242_ = ~pi251 | ~new_n4209_;
  assign new_n4243_ = ~new_n8304_ | ~new_n1037_;
  assign new_n4244_ = ~new_n6518_ | ~new_n1035_;
  assign new_n4245_ = ~new_n6749_ | ~new_n1034_;
  assign new_n4246_ = ~new_n9104_ | ~new_n1032_;
  assign new_n4247_ = ~new_n9288_ | ~new_n1031_;
  assign new_n4248_ = ~new_n1027_ | ~pi443;
  assign new_n4249_ = ~pi252 | ~new_n4209_;
  assign new_n4250_ = ~new_n8303_ | ~new_n1037_;
  assign new_n4251_ = ~new_n6517_ | ~new_n1035_;
  assign new_n4252_ = ~new_n6746_ | ~new_n1034_;
  assign new_n4253_ = ~new_n9103_ | ~new_n1032_;
  assign new_n4254_ = ~new_n9287_ | ~new_n1031_;
  assign new_n4255_ = ~new_n1027_ | ~pi444;
  assign new_n4256_ = ~pi253 | ~new_n4209_;
  assign new_n4257_ = ~new_n8302_ | ~new_n1037_;
  assign new_n4258_ = ~new_n6516_ | ~new_n1035_;
  assign new_n4259_ = ~new_n6743_ | ~new_n1034_;
  assign new_n4260_ = ~new_n9102_ | ~new_n1032_;
  assign new_n4261_ = ~new_n9286_ | ~new_n1031_;
  assign new_n4262_ = ~new_n1027_ | ~pi445;
  assign new_n4263_ = ~pi254 | ~new_n4209_;
  assign new_n4264_ = ~new_n8301_ | ~new_n1037_;
  assign new_n4265_ = ~new_n6515_ | ~new_n1035_;
  assign new_n4266_ = ~new_n6740_ | ~new_n1034_;
  assign new_n4267_ = ~new_n9101_ | ~new_n1032_;
  assign new_n4268_ = ~new_n9285_ | ~new_n1031_;
  assign new_n4269_ = ~new_n1027_ | ~pi446;
  assign new_n4270_ = ~pi255 | ~new_n4209_;
  assign new_n4271_ = ~new_n8300_ | ~new_n1037_;
  assign new_n4272_ = ~new_n6514_ | ~new_n1035_;
  assign new_n4273_ = ~new_n6737_ | ~new_n1034_;
  assign new_n4274_ = ~new_n9100_ | ~new_n1032_;
  assign new_n4275_ = ~new_n9284_ | ~new_n1031_;
  assign new_n4276_ = ~new_n1027_ | ~pi447;
  assign new_n4277_ = ~pi256 | ~new_n4209_;
  assign new_n4278_ = ~new_n8299_ | ~new_n1037_;
  assign new_n4279_ = ~new_n6513_ | ~new_n1035_;
  assign new_n4280_ = ~new_n6734_ | ~new_n1034_;
  assign new_n4281_ = ~new_n9099_ | ~new_n1032_;
  assign new_n4282_ = ~new_n9283_ | ~new_n1031_;
  assign new_n4283_ = ~new_n1027_ | ~pi448;
  assign new_n4284_ = ~pi257 | ~new_n4209_;
  assign new_n4285_ = ~new_n8348_ | ~new_n1037_;
  assign new_n4286_ = ~new_n6543_ | ~new_n1035_;
  assign new_n4287_ = ~new_n6820_ | ~new_n1034_;
  assign new_n4288_ = ~new_n9127_ | ~new_n1032_;
  assign new_n4289_ = ~new_n9312_ | ~new_n1031_;
  assign new_n4290_ = ~new_n1027_ | ~pi449;
  assign new_n4291_ = ~pi258 | ~new_n4209_;
  assign new_n4292_ = ~new_n8347_ | ~new_n1037_;
  assign new_n4293_ = ~new_n6542_ | ~new_n1035_;
  assign new_n4294_ = ~new_n6817_ | ~new_n1034_;
  assign new_n4295_ = ~new_n9126_ | ~new_n1032_;
  assign new_n4296_ = ~new_n9311_ | ~new_n1031_;
  assign new_n4297_ = ~new_n1027_ | ~pi450;
  assign new_n4298_ = ~pi259 | ~new_n4209_;
  assign new_n4299_ = ~new_n8346_ | ~new_n1037_;
  assign new_n4300_ = ~new_n6541_ | ~new_n1035_;
  assign new_n4301_ = ~new_n6814_ | ~new_n1034_;
  assign new_n4302_ = ~new_n9125_ | ~new_n1032_;
  assign new_n4303_ = ~new_n9310_ | ~new_n1031_;
  assign new_n4304_ = ~new_n1027_ | ~pi451;
  assign new_n4305_ = ~pi260 | ~new_n4209_;
  assign new_n4306_ = ~new_n8345_ | ~new_n1037_;
  assign new_n4307_ = ~new_n6540_ | ~new_n1035_;
  assign new_n4308_ = ~new_n6811_ | ~new_n1034_;
  assign new_n4309_ = ~new_n9124_ | ~new_n1032_;
  assign new_n4310_ = ~new_n9309_ | ~new_n1031_;
  assign new_n4311_ = ~new_n1027_ | ~pi452;
  assign new_n4312_ = ~pi261 | ~new_n4209_;
  assign new_n4313_ = ~new_n8344_ | ~new_n1037_;
  assign new_n4314_ = ~new_n6539_ | ~new_n1035_;
  assign new_n4315_ = ~new_n6808_ | ~new_n1034_;
  assign new_n4316_ = ~new_n9123_ | ~new_n1032_;
  assign new_n4317_ = ~new_n9308_ | ~new_n1031_;
  assign new_n4318_ = ~new_n1027_ | ~pi453;
  assign new_n4319_ = ~pi262 | ~new_n4209_;
  assign new_n4320_ = ~new_n8343_ | ~new_n1037_;
  assign new_n4321_ = ~new_n6538_ | ~new_n1035_;
  assign new_n4322_ = ~new_n6805_ | ~new_n1034_;
  assign new_n4323_ = ~new_n9122_ | ~new_n1032_;
  assign new_n4324_ = ~new_n9307_ | ~new_n1031_;
  assign new_n4325_ = ~new_n1027_ | ~pi454;
  assign new_n4326_ = ~pi263 | ~new_n4209_;
  assign new_n4327_ = ~new_n8342_ | ~new_n1037_;
  assign new_n4328_ = ~new_n6537_ | ~new_n1035_;
  assign new_n4329_ = ~new_n6802_ | ~new_n1034_;
  assign new_n4330_ = ~new_n9121_ | ~new_n1032_;
  assign new_n4331_ = ~new_n9306_ | ~new_n1031_;
  assign new_n4332_ = ~new_n1027_ | ~pi455;
  assign new_n4333_ = ~pi264 | ~new_n4209_;
  assign new_n4334_ = ~new_n8341_ | ~new_n1037_;
  assign new_n4335_ = ~new_n6536_ | ~new_n1035_;
  assign new_n4336_ = ~new_n6799_ | ~new_n1034_;
  assign new_n4337_ = ~new_n9120_ | ~new_n1032_;
  assign new_n4338_ = ~new_n9305_ | ~new_n1031_;
  assign new_n4339_ = ~new_n1027_ | ~pi456;
  assign new_n4340_ = ~pi265 | ~new_n4209_;
  assign new_n4341_ = ~new_n8340_ | ~new_n1037_;
  assign new_n4342_ = ~new_n6535_ | ~new_n1035_;
  assign new_n4343_ = ~new_n6796_ | ~new_n1034_;
  assign new_n4344_ = ~new_n9119_ | ~new_n1032_;
  assign new_n4345_ = ~new_n9304_ | ~new_n1031_;
  assign new_n4346_ = ~new_n1027_ | ~pi457;
  assign new_n4347_ = ~pi266 | ~new_n4209_;
  assign new_n4348_ = ~new_n8339_ | ~new_n1037_;
  assign new_n4349_ = ~new_n6534_ | ~new_n1035_;
  assign new_n4350_ = ~new_n6793_ | ~new_n1034_;
  assign new_n4351_ = ~new_n9118_ | ~new_n1032_;
  assign new_n4352_ = ~new_n9303_ | ~new_n1031_;
  assign new_n4353_ = ~new_n1027_ | ~pi458;
  assign new_n4354_ = ~pi267 | ~new_n4209_;
  assign new_n4355_ = ~new_n8338_ | ~new_n1037_;
  assign new_n4356_ = ~new_n6532_ | ~new_n1035_;
  assign new_n4357_ = ~new_n6789_ | ~new_n1034_;
  assign new_n4358_ = ~new_n9116_ | ~new_n1032_;
  assign new_n4359_ = ~new_n9302_ | ~new_n1031_;
  assign new_n4360_ = ~new_n1027_ | ~pi459;
  assign new_n4361_ = ~pi268 | ~new_n4209_;
  assign new_n4362_ = ~new_n8337_ | ~new_n1037_;
  assign new_n4363_ = ~new_n6531_ | ~new_n1035_;
  assign new_n4364_ = ~new_n6786_ | ~new_n1034_;
  assign new_n4365_ = ~new_n9115_ | ~new_n1032_;
  assign new_n4366_ = ~new_n9301_ | ~new_n1031_;
  assign new_n4367_ = ~new_n1027_ | ~pi460;
  assign new_n4368_ = ~pi269 | ~new_n4209_;
  assign new_n4369_ = ~new_n8336_ | ~new_n1037_;
  assign new_n4370_ = ~new_n6530_ | ~new_n1035_;
  assign new_n4371_ = ~new_n6783_ | ~new_n1034_;
  assign new_n4372_ = ~new_n9114_ | ~new_n1032_;
  assign new_n4373_ = ~new_n9300_ | ~new_n1031_;
  assign new_n4374_ = ~new_n1027_ | ~pi461;
  assign new_n4375_ = ~pi270 | ~new_n4209_;
  assign new_n4376_ = ~new_n8335_ | ~new_n1037_;
  assign new_n4377_ = ~new_n6529_ | ~new_n1035_;
  assign new_n4378_ = ~new_n6780_ | ~new_n1034_;
  assign new_n4379_ = ~new_n9113_ | ~new_n1032_;
  assign new_n4380_ = ~new_n9299_ | ~new_n1031_;
  assign new_n4381_ = ~new_n1027_ | ~pi462;
  assign new_n4382_ = ~pi271 | ~new_n4209_;
  assign new_n4383_ = ~new_n8334_ | ~new_n1037_;
  assign new_n4384_ = ~new_n6528_ | ~new_n1035_;
  assign new_n4385_ = ~new_n6777_ | ~new_n1034_;
  assign new_n4386_ = ~new_n9112_ | ~new_n1032_;
  assign new_n4387_ = ~new_n9298_ | ~new_n1031_;
  assign new_n4388_ = ~new_n1027_ | ~pi463;
  assign new_n4389_ = ~pi272 | ~new_n4209_;
  assign new_n4390_ = ~new_n8333_ | ~new_n1037_;
  assign new_n4391_ = ~new_n6527_ | ~new_n1035_;
  assign new_n4392_ = ~new_n6774_ | ~new_n1034_;
  assign new_n4393_ = ~new_n9111_ | ~new_n1032_;
  assign new_n4394_ = ~new_n9297_ | ~new_n1031_;
  assign new_n4395_ = ~new_n1027_ | ~pi464;
  assign new_n4396_ = ~pi273 | ~new_n4209_;
  assign new_n4397_ = ~new_n8332_ | ~new_n1037_;
  assign new_n4398_ = ~new_n6526_ | ~new_n1035_;
  assign new_n4399_ = ~new_n6771_ | ~new_n1034_;
  assign new_n4400_ = ~new_n9110_ | ~new_n1032_;
  assign new_n4401_ = ~new_n9296_ | ~new_n1031_;
  assign new_n4402_ = ~new_n1027_ | ~pi465;
  assign new_n4403_ = ~pi274 | ~new_n4209_;
  assign new_n4404_ = ~new_n8331_ | ~new_n1037_;
  assign new_n4405_ = ~new_n6525_ | ~new_n1035_;
  assign new_n4406_ = ~new_n6768_ | ~new_n1034_;
  assign new_n4407_ = ~new_n9109_ | ~new_n1032_;
  assign new_n4408_ = ~new_n9295_ | ~new_n1031_;
  assign new_n4409_ = ~new_n1027_ | ~pi466;
  assign new_n4410_ = ~pi275 | ~new_n4209_;
  assign new_n4411_ = ~new_n8330_ | ~new_n1037_;
  assign new_n4412_ = ~new_n6524_ | ~new_n1035_;
  assign new_n4413_ = ~new_n6765_ | ~new_n1034_;
  assign new_n4414_ = ~new_n9108_ | ~new_n1032_;
  assign new_n4415_ = ~new_n9294_ | ~new_n1031_;
  assign new_n4416_ = ~new_n1027_ | ~pi467;
  assign new_n4417_ = ~pi276 | ~new_n4209_;
  assign new_n4418_ = ~new_n8329_ | ~new_n1037_;
  assign new_n4419_ = ~new_n6523_ | ~new_n1035_;
  assign new_n4420_ = ~new_n6763_ | ~new_n1034_;
  assign new_n4421_ = ~new_n9107_ | ~new_n1032_;
  assign new_n4422_ = ~new_n9293_ | ~new_n1031_;
  assign new_n4423_ = ~new_n1027_ | ~pi468;
  assign new_n4424_ = ~pi277 | ~new_n4209_;
  assign new_n4425_ = ~new_n8328_ | ~new_n1037_;
  assign new_n4426_ = ~new_n6521_ | ~new_n1035_;
  assign new_n4427_ = ~new_n6758_ | ~new_n1034_;
  assign new_n4428_ = ~new_n9106_ | ~new_n1032_;
  assign new_n4429_ = ~new_n9291_ | ~new_n1031_;
  assign new_n4430_ = ~new_n1027_ | ~pi469;
  assign new_n4431_ = ~pi278 | ~new_n4209_;
  assign new_n4432_ = ~new_n8327_ | ~new_n1037_;
  assign new_n4433_ = ~new_n6520_ | ~new_n1035_;
  assign new_n4434_ = ~new_n6756_ | ~new_n1034_;
  assign new_n4435_ = ~new_n9105_ | ~new_n1032_;
  assign new_n4436_ = ~new_n9290_ | ~new_n1031_;
  assign new_n4437_ = ~new_n1027_ | ~pi470;
  assign new_n4438_ = ~pi279 | ~new_n4209_;
  assign new_n4439_ = ~new_n2854_ | ~new_n1938_;
  assign new_n4440_ = ~new_n2060_;
  assign new_n4441_ = ~pi107 | ~new_n1938_;
  assign new_n4442_ = ~pi108 | ~new_n1952_;
  assign new_n4443_ = ~new_n4442_ | ~new_n4441_;
  assign new_n4444_ = ~pi280 | ~new_n1033_;
  assign new_n4445_ = ~new_n1029_ | ~new_n6677_;
  assign new_n4446_ = ~new_n1022_ | ~pi439;
  assign new_n4447_ = ~new_n7160_ | ~new_n1021_;
  assign new_n4448_ = ~pi280 | ~new_n4440_;
  assign new_n4449_ = ~new_n7733_ | ~new_n1033_;
  assign new_n4450_ = ~new_n1029_ | ~new_n6702_;
  assign new_n4451_ = ~new_n1022_ | ~pi440;
  assign new_n4452_ = ~new_n7190_ | ~new_n1021_;
  assign new_n4453_ = ~pi281 | ~new_n4440_;
  assign new_n4454_ = ~new_n7788_ | ~new_n1033_;
  assign new_n4455_ = ~new_n1029_ | ~new_n6761_;
  assign new_n4456_ = ~new_n1022_ | ~pi441;
  assign new_n4457_ = ~new_n7097_ | ~new_n1021_;
  assign new_n4458_ = ~pi282 | ~new_n4440_;
  assign new_n4459_ = ~new_n7785_ | ~new_n1033_;
  assign new_n4460_ = ~new_n1029_ | ~new_n6752_;
  assign new_n4461_ = ~new_n1022_ | ~pi442;
  assign new_n4462_ = ~new_n7098_ | ~new_n1021_;
  assign new_n4463_ = ~pi283 | ~new_n4440_;
  assign new_n4464_ = ~new_n7784_ | ~new_n1033_;
  assign new_n4465_ = ~new_n1029_ | ~new_n6749_;
  assign new_n4466_ = ~new_n1022_ | ~pi443;
  assign new_n4467_ = ~new_n7168_ | ~new_n1021_;
  assign new_n4468_ = ~pi284 | ~new_n4440_;
  assign new_n4469_ = ~new_n7783_ | ~new_n1033_;
  assign new_n4470_ = ~new_n1029_ | ~new_n6746_;
  assign new_n4471_ = ~new_n1022_ | ~pi444;
  assign new_n4472_ = ~new_n7166_ | ~new_n1021_;
  assign new_n4473_ = ~pi285 | ~new_n4440_;
  assign new_n4474_ = ~new_n7782_ | ~new_n1033_;
  assign new_n4475_ = ~new_n1029_ | ~new_n6743_;
  assign new_n4476_ = ~new_n1022_ | ~pi445;
  assign new_n4477_ = ~new_n7164_ | ~new_n1021_;
  assign new_n4478_ = ~pi286 | ~new_n4440_;
  assign new_n4479_ = ~new_n7781_ | ~new_n1033_;
  assign new_n4480_ = ~new_n1029_ | ~new_n6740_;
  assign new_n4481_ = ~new_n1022_ | ~pi446;
  assign new_n4482_ = ~new_n7099_ | ~new_n1021_;
  assign new_n4483_ = ~pi287 | ~new_n4440_;
  assign new_n4484_ = ~new_n7780_ | ~new_n1033_;
  assign new_n4485_ = ~new_n1029_ | ~new_n6737_;
  assign new_n4486_ = ~new_n1022_ | ~pi447;
  assign new_n4487_ = ~new_n7163_ | ~new_n1021_;
  assign new_n4488_ = ~pi288 | ~new_n4440_;
  assign new_n4489_ = ~new_n7779_ | ~new_n1033_;
  assign new_n4490_ = ~new_n1029_ | ~new_n6734_;
  assign new_n4491_ = ~new_n1022_ | ~pi448;
  assign new_n4492_ = ~new_n7161_ | ~new_n1021_;
  assign new_n4493_ = ~pi289 | ~new_n4440_;
  assign new_n4494_ = ~new_n7808_ | ~new_n1033_;
  assign new_n4495_ = ~new_n1029_ | ~new_n6820_;
  assign new_n4496_ = ~new_n1022_ | ~pi449;
  assign new_n4497_ = ~new_n7092_ | ~new_n1021_;
  assign new_n4498_ = ~pi290 | ~new_n4440_;
  assign new_n4499_ = ~new_n7807_ | ~new_n1033_;
  assign new_n4500_ = ~new_n1029_ | ~new_n6817_;
  assign new_n4501_ = ~new_n1022_ | ~pi450;
  assign new_n4502_ = ~new_n7093_ | ~new_n1021_;
  assign new_n4503_ = ~pi291 | ~new_n4440_;
  assign new_n4504_ = ~new_n7806_ | ~new_n1033_;
  assign new_n4505_ = ~new_n1029_ | ~new_n6814_;
  assign new_n4506_ = ~new_n1022_ | ~pi451;
  assign new_n4507_ = ~new_n7200_ | ~new_n1021_;
  assign new_n4508_ = ~pi292 | ~new_n4440_;
  assign new_n4509_ = ~new_n7805_ | ~new_n1033_;
  assign new_n4510_ = ~new_n1029_ | ~new_n6811_;
  assign new_n4511_ = ~new_n1022_ | ~pi452;
  assign new_n4512_ = ~new_n7198_ | ~new_n1021_;
  assign new_n4513_ = ~pi293 | ~new_n4440_;
  assign new_n4514_ = ~new_n7804_ | ~new_n1033_;
  assign new_n4515_ = ~new_n1029_ | ~new_n6808_;
  assign new_n4516_ = ~new_n1022_ | ~pi453;
  assign new_n4517_ = ~new_n7197_ | ~new_n1021_;
  assign new_n4518_ = ~pi294 | ~new_n4440_;
  assign new_n4519_ = ~new_n7803_ | ~new_n1033_;
  assign new_n4520_ = ~new_n1029_ | ~new_n6805_;
  assign new_n4521_ = ~new_n1022_ | ~pi454;
  assign new_n4522_ = ~new_n7094_ | ~new_n1021_;
  assign new_n4523_ = ~pi295 | ~new_n4440_;
  assign new_n4524_ = ~new_n7802_ | ~new_n1033_;
  assign new_n4525_ = ~new_n1029_ | ~new_n6802_;
  assign new_n4526_ = ~new_n1022_ | ~pi455;
  assign new_n4527_ = ~new_n7095_ | ~new_n1021_;
  assign new_n4528_ = ~pi296 | ~new_n4440_;
  assign new_n4529_ = ~new_n7801_ | ~new_n1033_;
  assign new_n4530_ = ~new_n1029_ | ~new_n6799_;
  assign new_n4531_ = ~new_n1022_ | ~pi456;
  assign new_n4532_ = ~new_n7196_ | ~new_n1021_;
  assign new_n4533_ = ~pi297 | ~new_n4440_;
  assign new_n4534_ = ~new_n7800_ | ~new_n1033_;
  assign new_n4535_ = ~new_n1029_ | ~new_n6796_;
  assign new_n4536_ = ~new_n1022_ | ~pi457;
  assign new_n4537_ = ~new_n7194_ | ~new_n1021_;
  assign new_n4538_ = ~pi298 | ~new_n4440_;
  assign new_n4539_ = ~new_n7799_ | ~new_n1033_;
  assign new_n4540_ = ~new_n1029_ | ~new_n6793_;
  assign new_n4541_ = ~new_n1022_ | ~pi458;
  assign new_n4542_ = ~new_n7192_ | ~new_n1021_;
  assign new_n4543_ = ~pi299 | ~new_n4440_;
  assign new_n4544_ = ~new_n7798_ | ~new_n1033_;
  assign new_n4545_ = ~new_n1029_ | ~new_n6789_;
  assign new_n4546_ = ~new_n1022_ | ~pi459;
  assign new_n4547_ = ~new_n7188_ | ~new_n1021_;
  assign new_n4548_ = ~pi300 | ~new_n4440_;
  assign new_n4549_ = ~new_n7797_ | ~new_n1033_;
  assign new_n4550_ = ~new_n1029_ | ~new_n6786_;
  assign new_n4551_ = ~new_n1022_ | ~pi460;
  assign new_n4552_ = ~new_n7096_ | ~new_n1021_;
  assign new_n4553_ = ~pi301 | ~new_n4440_;
  assign new_n4554_ = ~new_n7796_ | ~new_n1033_;
  assign new_n4555_ = ~new_n1029_ | ~new_n6783_;
  assign new_n4556_ = ~new_n1022_ | ~pi461;
  assign new_n4557_ = ~new_n7187_ | ~new_n1021_;
  assign new_n4558_ = ~pi302 | ~new_n4440_;
  assign new_n4559_ = ~new_n7795_ | ~new_n1033_;
  assign new_n4560_ = ~new_n1029_ | ~new_n6780_;
  assign new_n4561_ = ~new_n1022_ | ~pi462;
  assign new_n4562_ = ~new_n7185_ | ~new_n1021_;
  assign new_n4563_ = ~pi303 | ~new_n4440_;
  assign new_n4564_ = ~new_n7794_ | ~new_n1033_;
  assign new_n4565_ = ~new_n1029_ | ~new_n6777_;
  assign new_n4566_ = ~new_n1022_ | ~pi463;
  assign new_n4567_ = ~new_n7183_ | ~new_n1021_;
  assign new_n4568_ = ~pi304 | ~new_n4440_;
  assign new_n4569_ = ~new_n7793_ | ~new_n1033_;
  assign new_n4570_ = ~new_n1029_ | ~new_n6774_;
  assign new_n4571_ = ~new_n1022_ | ~pi464;
  assign new_n4572_ = ~new_n7181_ | ~new_n1021_;
  assign new_n4573_ = ~pi305 | ~new_n4440_;
  assign new_n4574_ = ~new_n7792_ | ~new_n1033_;
  assign new_n4575_ = ~new_n1029_ | ~new_n6771_;
  assign new_n4576_ = ~new_n1022_ | ~pi465;
  assign new_n4577_ = ~new_n7179_ | ~new_n1021_;
  assign new_n4578_ = ~pi306 | ~new_n4440_;
  assign new_n4579_ = ~new_n7791_ | ~new_n1033_;
  assign new_n4580_ = ~new_n1029_ | ~new_n6768_;
  assign new_n4581_ = ~new_n1022_ | ~pi466;
  assign new_n4582_ = ~new_n7177_ | ~new_n1021_;
  assign new_n4583_ = ~pi307 | ~new_n4440_;
  assign new_n4584_ = ~new_n7790_ | ~new_n1033_;
  assign new_n4585_ = ~new_n1029_ | ~new_n6765_;
  assign new_n4586_ = ~new_n1022_ | ~pi467;
  assign new_n4587_ = ~new_n7175_ | ~new_n1021_;
  assign new_n4588_ = ~pi308 | ~new_n4440_;
  assign new_n4589_ = ~new_n7789_ | ~new_n1033_;
  assign new_n4590_ = ~new_n1029_ | ~new_n6763_;
  assign new_n4591_ = ~new_n1022_ | ~pi468;
  assign new_n4592_ = ~new_n7173_ | ~new_n1021_;
  assign new_n4593_ = ~pi309 | ~new_n4440_;
  assign new_n4594_ = ~new_n7787_ | ~new_n1033_;
  assign new_n4595_ = ~new_n1029_ | ~new_n6758_;
  assign new_n4596_ = ~new_n1022_ | ~pi469;
  assign new_n4597_ = ~new_n7171_ | ~new_n1021_;
  assign new_n4598_ = ~pi310 | ~new_n4440_;
  assign new_n4599_ = ~new_n7786_ | ~new_n1033_;
  assign new_n4600_ = ~new_n1029_ | ~new_n6756_;
  assign new_n4601_ = ~new_n1022_ | ~pi470;
  assign new_n4602_ = ~new_n7169_ | ~new_n1021_;
  assign new_n4603_ = ~pi311 | ~new_n4440_;
  assign new_n4604_ = ~pi035 | ~new_n1926_;
  assign new_n4605_ = ~pi390 | ~new_n1039_;
  assign new_n4606_ = ~pi017 | ~new_n1038_;
  assign new_n4607_ = ~new_n4606_ | ~new_n4605_;
  assign new_n4608_ = ~pi389 | ~new_n1039_;
  assign new_n4609_ = ~pi018 | ~new_n1038_;
  assign new_n4610_ = ~new_n4609_ | ~new_n4608_;
  assign new_n4611_ = ~pi388 | ~new_n1039_;
  assign new_n4612_ = ~pi019 | ~new_n1038_;
  assign new_n4613_ = ~new_n4612_ | ~new_n4611_;
  assign new_n4614_ = ~pi387 | ~new_n1039_;
  assign new_n4615_ = ~pi020 | ~new_n1038_;
  assign new_n4616_ = ~new_n4615_ | ~new_n4614_;
  assign new_n4617_ = ~pi386 | ~new_n1039_;
  assign new_n4618_ = ~pi021 | ~new_n1038_;
  assign new_n4619_ = ~new_n4618_ | ~new_n4617_;
  assign new_n4620_ = ~pi385 | ~new_n1039_;
  assign new_n4621_ = ~pi022 | ~new_n1038_;
  assign new_n4622_ = ~new_n4621_ | ~new_n4620_;
  assign new_n4623_ = ~pi384 | ~new_n1039_;
  assign new_n4624_ = ~pi023 | ~new_n1038_;
  assign new_n4625_ = ~new_n4624_ | ~new_n4623_;
  assign new_n4626_ = ~pi383 | ~new_n1039_;
  assign new_n4627_ = ~pi024 | ~new_n1038_;
  assign new_n4628_ = ~new_n4627_ | ~new_n4626_;
  assign new_n4629_ = ~pi382 | ~new_n1039_;
  assign new_n4630_ = ~new_n1038_ | ~pi025;
  assign new_n4631_ = ~new_n4630_ | ~new_n4629_;
  assign new_n4632_ = ~pi381 | ~new_n1039_;
  assign new_n4633_ = ~new_n1038_ | ~pi026;
  assign new_n4634_ = ~new_n4633_ | ~new_n4632_;
  assign new_n4635_ = ~pi380 | ~new_n1039_;
  assign new_n4636_ = ~new_n1038_ | ~pi027;
  assign new_n4637_ = ~new_n4636_ | ~new_n4635_;
  assign new_n4638_ = ~pi379 | ~new_n1039_;
  assign new_n4639_ = ~new_n1038_ | ~pi028;
  assign new_n4640_ = ~new_n4639_ | ~new_n4638_;
  assign new_n4641_ = ~pi378 | ~new_n1039_;
  assign new_n4642_ = ~new_n1038_ | ~pi029;
  assign new_n4643_ = ~new_n4642_ | ~new_n4641_;
  assign new_n4644_ = ~pi377 | ~new_n1039_;
  assign new_n4645_ = ~new_n1038_ | ~pi030;
  assign new_n4646_ = ~new_n4645_ | ~new_n4644_;
  assign new_n4647_ = ~pi376 | ~new_n1039_;
  assign new_n4648_ = ~new_n1038_ | ~pi031;
  assign new_n4649_ = ~new_n4648_ | ~new_n4647_;
  assign new_n4650_ = ~pi375 | ~new_n1039_;
  assign new_n4651_ = ~new_n1038_ | ~pi032;
  assign new_n4652_ = ~new_n4651_ | ~new_n4650_;
  assign new_n4653_ = ~pi405 | ~new_n1039_;
  assign new_n4654_ = ~pi018 | ~new_n1038_;
  assign new_n4655_ = ~new_n4654_ | ~new_n4653_;
  assign new_n4656_ = ~pi404 | ~new_n1039_;
  assign new_n4657_ = ~pi019 | ~new_n1038_;
  assign new_n4658_ = ~new_n4657_ | ~new_n4656_;
  assign new_n4659_ = ~pi403 | ~new_n1039_;
  assign new_n4660_ = ~pi020 | ~new_n1038_;
  assign new_n4661_ = ~new_n4660_ | ~new_n4659_;
  assign new_n4662_ = ~pi402 | ~new_n1039_;
  assign new_n4663_ = ~pi021 | ~new_n1038_;
  assign new_n4664_ = ~new_n4663_ | ~new_n4662_;
  assign new_n4665_ = ~pi401 | ~new_n1039_;
  assign new_n4666_ = ~pi022 | ~new_n1038_;
  assign new_n4667_ = ~new_n4666_ | ~new_n4665_;
  assign new_n4668_ = ~pi400 | ~new_n1039_;
  assign new_n4669_ = ~pi023 | ~new_n1038_;
  assign new_n4670_ = ~new_n4669_ | ~new_n4668_;
  assign new_n4671_ = ~pi399 | ~new_n1039_;
  assign new_n4672_ = ~pi024 | ~new_n1038_;
  assign new_n4673_ = ~new_n4672_ | ~new_n4671_;
  assign new_n4674_ = ~pi398 | ~new_n1039_;
  assign new_n4675_ = ~new_n1038_ | ~pi025;
  assign new_n4676_ = ~new_n4675_ | ~new_n4674_;
  assign new_n4677_ = ~pi397 | ~new_n1039_;
  assign new_n4678_ = ~new_n1038_ | ~pi026;
  assign new_n4679_ = ~new_n4678_ | ~new_n4677_;
  assign new_n4680_ = ~pi396 | ~new_n1039_;
  assign new_n4681_ = ~new_n1038_ | ~pi027;
  assign new_n4682_ = ~new_n4681_ | ~new_n4680_;
  assign new_n4683_ = ~pi395 | ~new_n1039_;
  assign new_n4684_ = ~new_n1038_ | ~pi028;
  assign new_n4685_ = ~new_n4684_ | ~new_n4683_;
  assign new_n4686_ = ~pi394 | ~new_n1039_;
  assign new_n4687_ = ~new_n1038_ | ~pi029;
  assign new_n4688_ = ~new_n4687_ | ~new_n4686_;
  assign new_n4689_ = ~pi393 | ~new_n1039_;
  assign new_n4690_ = ~new_n1038_ | ~pi030;
  assign new_n4691_ = ~new_n4690_ | ~new_n4689_;
  assign new_n4692_ = ~pi392 | ~new_n1039_;
  assign new_n4693_ = ~new_n1038_ | ~pi031;
  assign new_n4694_ = ~new_n4693_ | ~new_n4692_;
  assign new_n4695_ = ~pi391 | ~new_n1039_;
  assign new_n4696_ = ~new_n1038_ | ~pi032;
  assign new_n4697_ = ~new_n4696_ | ~new_n4695_;
  assign new_n4698_ = ~new_n2904_ | ~new_n2880_ | ~new_n6251_;
  assign new_n4699_ = ~new_n1085_ | ~new_n1938_;
  assign new_n4700_ = ~new_n2061_;
  assign new_n4701_ = ~new_n1042_ | ~pi327;
  assign new_n4702_ = ~new_n1041_ | ~pi375;
  assign new_n4703_ = ~pi343 | ~new_n4700_;
  assign new_n4704_ = ~new_n1042_ | ~pi326;
  assign new_n4705_ = ~new_n1041_ | ~pi376;
  assign new_n4706_ = ~pi344 | ~new_n4700_;
  assign new_n4707_ = ~new_n1042_ | ~pi325;
  assign new_n4708_ = ~new_n1041_ | ~pi377;
  assign new_n4709_ = ~pi345 | ~new_n4700_;
  assign new_n4710_ = ~new_n1042_ | ~pi324;
  assign new_n4711_ = ~new_n1041_ | ~pi378;
  assign new_n4712_ = ~pi346 | ~new_n4700_;
  assign new_n4713_ = ~new_n1042_ | ~pi323;
  assign new_n4714_ = ~new_n1041_ | ~pi379;
  assign new_n4715_ = ~pi347 | ~new_n4700_;
  assign new_n4716_ = ~new_n1042_ | ~pi322;
  assign new_n4717_ = ~new_n1041_ | ~pi380;
  assign new_n4718_ = ~pi348 | ~new_n4700_;
  assign new_n4719_ = ~new_n1042_ | ~pi321;
  assign new_n4720_ = ~new_n1041_ | ~pi381;
  assign new_n4721_ = ~pi349 | ~new_n4700_;
  assign new_n4722_ = ~new_n1042_ | ~pi320;
  assign new_n4723_ = ~new_n1041_ | ~pi382;
  assign new_n4724_ = ~pi350 | ~new_n4700_;
  assign new_n4725_ = ~new_n1042_ | ~pi319;
  assign new_n4726_ = ~new_n1041_ | ~pi383;
  assign new_n4727_ = ~pi351 | ~new_n4700_;
  assign new_n4728_ = ~new_n1042_ | ~pi318;
  assign new_n4729_ = ~new_n1041_ | ~pi384;
  assign new_n4730_ = ~pi352 | ~new_n4700_;
  assign new_n4731_ = ~new_n1042_ | ~pi317;
  assign new_n4732_ = ~new_n1041_ | ~pi385;
  assign new_n4733_ = ~pi353 | ~new_n4700_;
  assign new_n4734_ = ~new_n1042_ | ~pi316;
  assign new_n4735_ = ~new_n1041_ | ~pi386;
  assign new_n4736_ = ~pi354 | ~new_n4700_;
  assign new_n4737_ = ~new_n1042_ | ~pi315;
  assign new_n4738_ = ~new_n1041_ | ~pi387;
  assign new_n4739_ = ~pi355 | ~new_n4700_;
  assign new_n4740_ = ~new_n1042_ | ~pi314;
  assign new_n4741_ = ~new_n1041_ | ~pi388;
  assign new_n4742_ = ~pi356 | ~new_n4700_;
  assign new_n4743_ = ~new_n1042_ | ~pi313;
  assign new_n4744_ = ~new_n1041_ | ~pi389;
  assign new_n4745_ = ~pi357 | ~new_n4700_;
  assign new_n4746_ = ~new_n1042_ | ~pi312;
  assign new_n4747_ = ~new_n1041_ | ~pi390;
  assign new_n4748_ = ~pi358 | ~new_n4700_;
  assign new_n4749_ = ~new_n1081_ | ~pi391;
  assign new_n4750_ = ~new_n1042_ | ~pi342;
  assign new_n4751_ = ~pi359 | ~new_n4700_;
  assign new_n4752_ = ~new_n1081_ | ~pi392;
  assign new_n4753_ = ~new_n1042_ | ~pi341;
  assign new_n4754_ = ~pi360 | ~new_n4700_;
  assign new_n4755_ = ~new_n1081_ | ~pi393;
  assign new_n4756_ = ~new_n1042_ | ~pi340;
  assign new_n4757_ = ~pi361 | ~new_n4700_;
  assign new_n4758_ = ~new_n1081_ | ~pi394;
  assign new_n4759_ = ~new_n1042_ | ~pi339;
  assign new_n4760_ = ~pi362 | ~new_n4700_;
  assign new_n4761_ = ~new_n1081_ | ~pi395;
  assign new_n4762_ = ~new_n1042_ | ~pi338;
  assign new_n4763_ = ~pi363 | ~new_n4700_;
  assign new_n4764_ = ~new_n1081_ | ~pi396;
  assign new_n4765_ = ~new_n1042_ | ~pi337;
  assign new_n4766_ = ~pi364 | ~new_n4700_;
  assign new_n4767_ = ~new_n1081_ | ~pi397;
  assign new_n4768_ = ~new_n1042_ | ~pi336;
  assign new_n4769_ = ~pi365 | ~new_n4700_;
  assign new_n4770_ = ~new_n1081_ | ~pi398;
  assign new_n4771_ = ~new_n1042_ | ~pi335;
  assign new_n4772_ = ~pi366 | ~new_n4700_;
  assign new_n4773_ = ~new_n1081_ | ~pi399;
  assign new_n4774_ = ~new_n1042_ | ~pi334;
  assign new_n4775_ = ~pi367 | ~new_n4700_;
  assign new_n4776_ = ~new_n1081_ | ~pi400;
  assign new_n4777_ = ~new_n1042_ | ~pi333;
  assign new_n4778_ = ~pi368 | ~new_n4700_;
  assign new_n4779_ = ~new_n1081_ | ~pi401;
  assign new_n4780_ = ~new_n1042_ | ~pi332;
  assign new_n4781_ = ~pi369 | ~new_n4700_;
  assign new_n4782_ = ~new_n1081_ | ~pi402;
  assign new_n4783_ = ~new_n1042_ | ~pi331;
  assign new_n4784_ = ~pi370 | ~new_n4700_;
  assign new_n4785_ = ~new_n1081_ | ~pi403;
  assign new_n4786_ = ~new_n1042_ | ~pi330;
  assign new_n4787_ = ~pi371 | ~new_n4700_;
  assign new_n4788_ = ~new_n1081_ | ~pi404;
  assign new_n4789_ = ~new_n1042_ | ~pi329;
  assign new_n4790_ = ~pi372 | ~new_n4700_;
  assign new_n4791_ = ~new_n1081_ | ~pi405;
  assign new_n4792_ = ~new_n1042_ | ~pi328;
  assign new_n4793_ = ~pi373 | ~new_n4700_;
  assign new_n4794_ = ~new_n9223_ | ~new_n2839_ | ~new_n1104_;
  assign new_n4795_ = ~new_n2839_ | ~new_n2899_ | ~new_n2842_;
  assign new_n4796_ = ~new_n8624_ | ~new_n2845_ | ~new_n1927_;
  assign new_n4797_ = ~new_n6148_ | ~new_n1901_;
  assign new_n4798_ = ~new_n2528_ | ~new_n4797_;
  assign new_n4799_ = ~new_n1079_ | ~pi032;
  assign new_n4800_ = ~new_n1043_ | ~new_n7160_;
  assign new_n4801_ = ~pi375 | ~new_n2068_;
  assign new_n4802_ = ~new_n1079_ | ~pi031;
  assign new_n4803_ = ~new_n1043_ | ~new_n7190_;
  assign new_n4804_ = ~pi376 | ~new_n2068_;
  assign new_n4805_ = ~new_n1079_ | ~pi030;
  assign new_n4806_ = ~new_n1043_ | ~new_n7097_;
  assign new_n4807_ = ~pi377 | ~new_n2068_;
  assign new_n4808_ = ~new_n1079_ | ~pi029;
  assign new_n4809_ = ~new_n1043_ | ~new_n7098_;
  assign new_n4810_ = ~pi378 | ~new_n2068_;
  assign new_n4811_ = ~new_n1079_ | ~pi028;
  assign new_n4812_ = ~new_n1043_ | ~new_n7168_;
  assign new_n4813_ = ~pi379 | ~new_n2068_;
  assign new_n4814_ = ~new_n1079_ | ~pi027;
  assign new_n4815_ = ~new_n1043_ | ~new_n7166_;
  assign new_n4816_ = ~pi380 | ~new_n2068_;
  assign new_n4817_ = ~new_n1079_ | ~pi026;
  assign new_n4818_ = ~new_n1043_ | ~new_n7164_;
  assign new_n4819_ = ~pi381 | ~new_n2068_;
  assign new_n4820_ = ~new_n1079_ | ~pi025;
  assign new_n4821_ = ~new_n1043_ | ~new_n7099_;
  assign new_n4822_ = ~pi382 | ~new_n2068_;
  assign new_n4823_ = ~new_n1079_ | ~pi024;
  assign new_n4824_ = ~new_n1043_ | ~new_n7163_;
  assign new_n4825_ = ~pi383 | ~new_n2068_;
  assign new_n4826_ = ~new_n1079_ | ~pi023;
  assign new_n4827_ = ~new_n1043_ | ~new_n7161_;
  assign new_n4828_ = ~pi384 | ~new_n2068_;
  assign new_n4829_ = ~new_n1079_ | ~pi022;
  assign new_n4830_ = ~new_n1043_ | ~new_n7092_;
  assign new_n4831_ = ~pi385 | ~new_n2068_;
  assign new_n4832_ = ~new_n1079_ | ~pi021;
  assign new_n4833_ = ~new_n1043_ | ~new_n7093_;
  assign new_n4834_ = ~pi386 | ~new_n2068_;
  assign new_n4835_ = ~new_n1079_ | ~pi020;
  assign new_n4836_ = ~new_n1043_ | ~new_n7200_;
  assign new_n4837_ = ~pi387 | ~new_n2068_;
  assign new_n4838_ = ~new_n1079_ | ~pi019;
  assign new_n4839_ = ~new_n1043_ | ~new_n7198_;
  assign new_n4840_ = ~pi388 | ~new_n2068_;
  assign new_n4841_ = ~new_n1079_ | ~pi018;
  assign new_n4842_ = ~new_n1043_ | ~new_n7197_;
  assign new_n4843_ = ~pi389 | ~new_n2068_;
  assign new_n4844_ = ~new_n1079_ | ~pi017;
  assign new_n4845_ = ~new_n1043_ | ~new_n7094_;
  assign new_n4846_ = ~pi390 | ~new_n2068_;
  assign new_n4847_ = ~new_n1080_ | ~pi016;
  assign new_n4848_ = ~new_n1044_ | ~pi032;
  assign new_n4849_ = ~new_n1043_ | ~new_n7095_;
  assign new_n4850_ = ~pi391 | ~new_n2068_;
  assign new_n4851_ = ~new_n1080_ | ~pi015;
  assign new_n4852_ = ~new_n1044_ | ~pi031;
  assign new_n4853_ = ~new_n1043_ | ~new_n7196_;
  assign new_n4854_ = ~pi392 | ~new_n2068_;
  assign new_n4855_ = ~new_n1080_ | ~pi014;
  assign new_n4856_ = ~new_n1044_ | ~pi030;
  assign new_n4857_ = ~new_n1043_ | ~new_n7194_;
  assign new_n4858_ = ~pi393 | ~new_n2068_;
  assign new_n4859_ = ~new_n1080_ | ~pi013;
  assign new_n4860_ = ~new_n1044_ | ~pi029;
  assign new_n4861_ = ~new_n1043_ | ~new_n7192_;
  assign new_n4862_ = ~pi394 | ~new_n2068_;
  assign new_n4863_ = ~new_n1080_ | ~pi012;
  assign new_n4864_ = ~new_n1044_ | ~pi028;
  assign new_n4865_ = ~new_n1043_ | ~new_n7188_;
  assign new_n4866_ = ~pi395 | ~new_n2068_;
  assign new_n4867_ = ~new_n1080_ | ~pi011;
  assign new_n4868_ = ~new_n1044_ | ~pi027;
  assign new_n4869_ = ~new_n1043_ | ~new_n7096_;
  assign new_n4870_ = ~pi396 | ~new_n2068_;
  assign new_n4871_ = ~new_n1080_ | ~pi010;
  assign new_n4872_ = ~new_n1044_ | ~pi026;
  assign new_n4873_ = ~new_n1043_ | ~new_n7187_;
  assign new_n4874_ = ~pi397 | ~new_n2068_;
  assign new_n4875_ = ~new_n1080_ | ~pi009;
  assign new_n4876_ = ~new_n1044_ | ~pi025;
  assign new_n4877_ = ~new_n1043_ | ~new_n7185_;
  assign new_n4878_ = ~pi398 | ~new_n2068_;
  assign new_n4879_ = ~new_n1080_ | ~pi008;
  assign new_n4880_ = ~new_n1044_ | ~pi024;
  assign new_n4881_ = ~new_n1043_ | ~new_n7183_;
  assign new_n4882_ = ~pi399 | ~new_n2068_;
  assign new_n4883_ = ~new_n1080_ | ~pi007;
  assign new_n4884_ = ~new_n1044_ | ~pi023;
  assign new_n4885_ = ~new_n1043_ | ~new_n7181_;
  assign new_n4886_ = ~pi400 | ~new_n2068_;
  assign new_n4887_ = ~new_n1080_ | ~pi006;
  assign new_n4888_ = ~new_n1044_ | ~pi022;
  assign new_n4889_ = ~new_n1043_ | ~new_n7179_;
  assign new_n4890_ = ~pi401 | ~new_n2068_;
  assign new_n4891_ = ~new_n1080_ | ~pi005;
  assign new_n4892_ = ~new_n1044_ | ~pi021;
  assign new_n4893_ = ~new_n1043_ | ~new_n7177_;
  assign new_n4894_ = ~pi402 | ~new_n2068_;
  assign new_n4895_ = ~new_n1080_ | ~pi004;
  assign new_n4896_ = ~new_n1044_ | ~pi020;
  assign new_n4897_ = ~new_n1043_ | ~new_n7175_;
  assign new_n4898_ = ~pi403 | ~new_n2068_;
  assign new_n4899_ = ~new_n1080_ | ~pi003;
  assign new_n4900_ = ~new_n1044_ | ~pi019;
  assign new_n4901_ = ~new_n1043_ | ~new_n7173_;
  assign new_n4902_ = ~pi404 | ~new_n2068_;
  assign new_n4903_ = ~new_n1080_ | ~pi002;
  assign new_n4904_ = ~new_n1044_ | ~pi018;
  assign new_n4905_ = ~new_n1043_ | ~new_n7171_;
  assign new_n4906_ = ~pi405 | ~new_n2068_;
  assign new_n4907_ = ~new_n1080_ | ~pi001;
  assign new_n4908_ = ~new_n2843_ | ~new_n1917_;
  assign new_n4909_ = ~new_n2850_ | ~new_n4908_;
  assign new_n4910_ = ~new_n1040_ | ~new_n7160_;
  assign new_n4911_ = ~new_n1028_ | ~new_n8349_;
  assign new_n4912_ = ~pi407 | ~new_n2070_;
  assign new_n4913_ = ~new_n1040_ | ~new_n7190_;
  assign new_n4914_ = ~new_n1028_ | ~new_n8350_;
  assign new_n4915_ = ~pi408 | ~new_n2070_;
  assign new_n4916_ = ~new_n1040_ | ~new_n7097_;
  assign new_n4917_ = ~new_n1028_ | ~new_n8401_;
  assign new_n4918_ = ~pi409 | ~new_n2070_;
  assign new_n4919_ = ~new_n1040_ | ~new_n7098_;
  assign new_n4920_ = ~new_n1028_ | ~new_n8305_;
  assign new_n4921_ = ~pi410 | ~new_n2070_;
  assign new_n4922_ = ~new_n1040_ | ~new_n7168_;
  assign new_n4923_ = ~new_n1028_ | ~new_n8304_;
  assign new_n4924_ = ~pi411 | ~new_n2070_;
  assign new_n4925_ = ~new_n1040_ | ~new_n7166_;
  assign new_n4926_ = ~new_n1028_ | ~new_n8303_;
  assign new_n4927_ = ~pi412 | ~new_n2070_;
  assign new_n4928_ = ~new_n1040_ | ~new_n7164_;
  assign new_n4929_ = ~new_n1028_ | ~new_n8302_;
  assign new_n4930_ = ~pi413 | ~new_n2070_;
  assign new_n4931_ = ~new_n1040_ | ~new_n7099_;
  assign new_n4932_ = ~new_n1028_ | ~new_n8301_;
  assign new_n4933_ = ~pi414 | ~new_n2070_;
  assign new_n4934_ = ~new_n1040_ | ~new_n7163_;
  assign new_n4935_ = ~new_n1028_ | ~new_n8300_;
  assign new_n4936_ = ~pi415 | ~new_n2070_;
  assign new_n4937_ = ~new_n1040_ | ~new_n7161_;
  assign new_n4938_ = ~new_n1028_ | ~new_n8299_;
  assign new_n4939_ = ~pi416 | ~new_n2070_;
  assign new_n4940_ = ~new_n1040_ | ~new_n7092_;
  assign new_n4941_ = ~new_n1028_ | ~new_n8348_;
  assign new_n4942_ = ~pi417 | ~new_n2070_;
  assign new_n4943_ = ~new_n1040_ | ~new_n7093_;
  assign new_n4944_ = ~new_n1028_ | ~new_n8347_;
  assign new_n4945_ = ~pi418 | ~new_n2070_;
  assign new_n4946_ = ~new_n1040_ | ~new_n7200_;
  assign new_n4947_ = ~new_n1028_ | ~new_n8346_;
  assign new_n4948_ = ~pi419 | ~new_n2070_;
  assign new_n4949_ = ~new_n1040_ | ~new_n7198_;
  assign new_n4950_ = ~new_n1028_ | ~new_n8345_;
  assign new_n4951_ = ~pi420 | ~new_n2070_;
  assign new_n4952_ = ~new_n1040_ | ~new_n7197_;
  assign new_n4953_ = ~new_n1028_ | ~new_n8344_;
  assign new_n4954_ = ~pi421 | ~new_n2070_;
  assign new_n4955_ = ~new_n1040_ | ~new_n7094_;
  assign new_n4956_ = ~new_n1028_ | ~new_n8343_;
  assign new_n4957_ = ~pi422 | ~new_n2070_;
  assign new_n4958_ = ~new_n1040_ | ~new_n7095_;
  assign new_n4959_ = ~new_n1028_ | ~new_n8342_;
  assign new_n4960_ = ~pi423 | ~new_n2070_;
  assign new_n4961_ = ~new_n1040_ | ~new_n7196_;
  assign new_n4962_ = ~new_n1028_ | ~new_n8341_;
  assign new_n4963_ = ~pi424 | ~new_n2070_;
  assign new_n4964_ = ~new_n1040_ | ~new_n7194_;
  assign new_n4965_ = ~new_n1028_ | ~new_n8340_;
  assign new_n4966_ = ~pi425 | ~new_n2070_;
  assign new_n4967_ = ~new_n1040_ | ~new_n7192_;
  assign new_n4968_ = ~new_n1028_ | ~new_n8339_;
  assign new_n4969_ = ~pi426 | ~new_n2070_;
  assign new_n4970_ = ~new_n1040_ | ~new_n7188_;
  assign new_n4971_ = ~new_n1028_ | ~new_n8338_;
  assign new_n4972_ = ~pi427 | ~new_n2070_;
  assign new_n4973_ = ~new_n1040_ | ~new_n7096_;
  assign new_n4974_ = ~new_n1028_ | ~new_n8337_;
  assign new_n4975_ = ~pi428 | ~new_n2070_;
  assign new_n4976_ = ~new_n1040_ | ~new_n7187_;
  assign new_n4977_ = ~new_n1028_ | ~new_n8336_;
  assign new_n4978_ = ~pi429 | ~new_n2070_;
  assign new_n4979_ = ~new_n1040_ | ~new_n7185_;
  assign new_n4980_ = ~new_n1028_ | ~new_n8335_;
  assign new_n4981_ = ~pi430 | ~new_n2070_;
  assign new_n4982_ = ~new_n1040_ | ~new_n7183_;
  assign new_n4983_ = ~new_n1028_ | ~new_n8334_;
  assign new_n4984_ = ~pi431 | ~new_n2070_;
  assign new_n4985_ = ~new_n1040_ | ~new_n7181_;
  assign new_n4986_ = ~new_n1028_ | ~new_n8333_;
  assign new_n4987_ = ~pi432 | ~new_n2070_;
  assign new_n4988_ = ~new_n1040_ | ~new_n7179_;
  assign new_n4989_ = ~new_n1028_ | ~new_n8332_;
  assign new_n4990_ = ~pi433 | ~new_n2070_;
  assign new_n4991_ = ~new_n1040_ | ~new_n7177_;
  assign new_n4992_ = ~new_n1028_ | ~new_n8331_;
  assign new_n4993_ = ~pi434 | ~new_n2070_;
  assign new_n4994_ = ~new_n1040_ | ~new_n7175_;
  assign new_n4995_ = ~new_n1028_ | ~new_n8330_;
  assign new_n4996_ = ~pi435 | ~new_n2070_;
  assign new_n4997_ = ~new_n1040_ | ~new_n7173_;
  assign new_n4998_ = ~new_n1028_ | ~new_n8329_;
  assign new_n4999_ = ~pi436 | ~new_n2070_;
  assign new_n5000_ = ~new_n1040_ | ~new_n7171_;
  assign new_n5001_ = ~new_n1028_ | ~new_n8328_;
  assign new_n5002_ = ~pi437 | ~new_n2070_;
  assign new_n5003_ = ~new_n1028_ | ~new_n8327_;
  assign new_n5004_ = ~pi438 | ~new_n2070_;
  assign new_n5005_ = ~new_n2849_ | ~new_n9223_;
  assign new_n5006_ = ~new_n2847_ | ~new_n8624_;
  assign new_n5007_ = ~new_n2848_ | ~new_n1907_;
  assign new_n5008_ = ~new_n2075_;
  assign new_n5009_ = ~new_n2894_ | ~pi107;
  assign new_n5010_ = ~new_n7786_ | ~pi108;
  assign new_n5011_ = ~new_n5010_ | ~new_n5009_;
  assign new_n5012_ = pi478 | pi035;
  assign new_n5013_ = ~new_n1261_ | ~new_n8349_;
  assign new_n5014_ = ~pi439 | ~new_n6130_;
  assign new_n5015_ = ~pi407 | ~new_n6129_;
  assign new_n5016_ = ~new_n1086_ | ~new_n7160_;
  assign new_n5017_ = ~new_n1083_ | ~new_n7951_;
  assign new_n5018_ = ~new_n1030_ | ~pi280;
  assign new_n5019_ = ~new_n1023_ | ~pi280;
  assign new_n5020_ = ~new_n5008_ | ~pi439;
  assign new_n5021_ = ~new_n1261_ | ~new_n8350_;
  assign new_n5022_ = ~new_n8675_ | ~new_n6130_;
  assign new_n5023_ = ~pi408 | ~new_n6129_;
  assign new_n5024_ = ~new_n1086_ | ~new_n7190_;
  assign new_n5025_ = ~new_n1083_ | ~new_n7950_;
  assign new_n5026_ = ~new_n1030_ | ~pi281;
  assign new_n5027_ = ~new_n1023_ | ~new_n7733_;
  assign new_n5028_ = ~new_n5008_ | ~pi440;
  assign new_n5029_ = ~new_n1261_ | ~new_n8401_;
  assign new_n5030_ = ~new_n8742_ | ~new_n6130_;
  assign new_n5031_ = ~pi409 | ~new_n6129_;
  assign new_n5032_ = ~new_n1086_ | ~new_n7097_;
  assign new_n5033_ = ~new_n1083_ | ~new_n7959_;
  assign new_n5034_ = ~new_n1030_ | ~pi282;
  assign new_n5035_ = ~new_n1023_ | ~new_n7788_;
  assign new_n5036_ = ~new_n5008_ | ~pi441;
  assign new_n5037_ = ~new_n1261_ | ~new_n8305_;
  assign new_n5038_ = ~new_n8739_ | ~new_n6130_;
  assign new_n5039_ = ~pi410 | ~new_n6129_;
  assign new_n5040_ = ~new_n1086_ | ~new_n7098_;
  assign new_n5041_ = ~new_n1083_ | ~new_n7942_;
  assign new_n5042_ = ~new_n1030_ | ~pi283;
  assign new_n5043_ = ~new_n1023_ | ~new_n7785_;
  assign new_n5044_ = ~new_n5008_ | ~pi442;
  assign new_n5045_ = ~new_n1261_ | ~new_n8304_;
  assign new_n5046_ = ~new_n8738_ | ~new_n6130_;
  assign new_n5047_ = ~pi411 | ~new_n6129_;
  assign new_n5048_ = ~new_n1086_ | ~new_n7168_;
  assign new_n5049_ = ~new_n1083_ | ~new_n7941_;
  assign new_n5050_ = ~new_n1030_ | ~pi284;
  assign new_n5051_ = ~new_n1023_ | ~new_n7784_;
  assign new_n5052_ = ~new_n5008_ | ~pi443;
  assign new_n5053_ = ~new_n1261_ | ~new_n8303_;
  assign new_n5054_ = ~new_n8737_ | ~new_n6130_;
  assign new_n5055_ = ~pi412 | ~new_n6129_;
  assign new_n5056_ = ~new_n1086_ | ~new_n7166_;
  assign new_n5057_ = ~new_n7922_ | ~new_n1083_;
  assign new_n5058_ = ~new_n1030_ | ~pi285;
  assign new_n5059_ = ~new_n1023_ | ~new_n7783_;
  assign new_n5060_ = ~new_n5008_ | ~pi444;
  assign new_n5061_ = ~new_n1261_ | ~new_n8302_;
  assign new_n5062_ = ~new_n8736_ | ~new_n6130_;
  assign new_n5063_ = ~pi413 | ~new_n6129_;
  assign new_n5064_ = ~new_n1030_ | ~pi286;
  assign new_n5065_ = ~new_n1024_ | ~new_n7164_;
  assign new_n5066_ = ~new_n1023_ | ~new_n7782_;
  assign new_n5067_ = ~new_n5008_ | ~pi445;
  assign new_n5068_ = ~new_n1261_ | ~new_n8301_;
  assign new_n5069_ = ~new_n8735_ | ~new_n6130_;
  assign new_n5070_ = ~pi414 | ~new_n6129_;
  assign new_n5071_ = ~new_n1030_ | ~pi287;
  assign new_n5072_ = ~new_n1024_ | ~new_n7099_;
  assign new_n5073_ = ~new_n1023_ | ~new_n7781_;
  assign new_n5074_ = ~new_n5008_ | ~pi446;
  assign new_n5075_ = ~new_n1261_ | ~new_n8300_;
  assign new_n5076_ = ~new_n8734_ | ~new_n6130_;
  assign new_n5077_ = ~pi415 | ~new_n6129_;
  assign new_n5078_ = ~new_n1030_ | ~pi288;
  assign new_n5079_ = ~new_n1024_ | ~new_n7163_;
  assign new_n5080_ = ~new_n1023_ | ~new_n7780_;
  assign new_n5081_ = ~new_n5008_ | ~pi447;
  assign new_n5082_ = ~new_n1261_ | ~new_n8299_;
  assign new_n5083_ = ~new_n8733_ | ~new_n6130_;
  assign new_n5084_ = ~pi416 | ~new_n6129_;
  assign new_n5085_ = ~new_n1030_ | ~pi289;
  assign new_n5086_ = ~new_n1024_ | ~new_n7161_;
  assign new_n5087_ = ~new_n1023_ | ~new_n7779_;
  assign new_n5088_ = ~new_n5008_ | ~pi448;
  assign new_n5089_ = ~new_n1261_ | ~new_n8348_;
  assign new_n5090_ = ~new_n8762_ | ~new_n6130_;
  assign new_n5091_ = ~pi417 | ~new_n6129_;
  assign new_n5092_ = ~new_n1030_ | ~pi290;
  assign new_n5093_ = ~new_n1024_ | ~new_n7092_;
  assign new_n5094_ = ~new_n1023_ | ~new_n7808_;
  assign new_n5095_ = ~new_n5008_ | ~pi449;
  assign new_n5096_ = ~new_n1261_ | ~new_n8347_;
  assign new_n5097_ = ~new_n8761_ | ~new_n6130_;
  assign new_n5098_ = ~pi418 | ~new_n6129_;
  assign new_n5099_ = ~new_n1030_ | ~pi291;
  assign new_n5100_ = ~new_n1024_ | ~new_n7093_;
  assign new_n5101_ = ~new_n1023_ | ~new_n7807_;
  assign new_n5102_ = ~new_n5008_ | ~pi450;
  assign new_n5103_ = ~new_n1261_ | ~new_n8346_;
  assign new_n5104_ = ~new_n8760_ | ~new_n6130_;
  assign new_n5105_ = ~pi419 | ~new_n6129_;
  assign new_n5106_ = ~new_n1030_ | ~pi292;
  assign new_n5107_ = ~new_n1024_ | ~new_n7200_;
  assign new_n5108_ = ~new_n1023_ | ~new_n7806_;
  assign new_n5109_ = ~new_n5008_ | ~pi451;
  assign new_n5110_ = ~new_n1261_ | ~new_n8345_;
  assign new_n5111_ = ~new_n8759_ | ~new_n6130_;
  assign new_n5112_ = ~pi420 | ~new_n6129_;
  assign new_n5113_ = ~new_n1030_ | ~pi293;
  assign new_n5114_ = ~new_n1024_ | ~new_n7198_;
  assign new_n5115_ = ~new_n1023_ | ~new_n7805_;
  assign new_n5116_ = ~new_n5008_ | ~pi452;
  assign new_n5117_ = ~new_n1261_ | ~new_n8344_;
  assign new_n5118_ = ~new_n8758_ | ~new_n6130_;
  assign new_n5119_ = ~pi421 | ~new_n6129_;
  assign new_n5120_ = ~new_n1030_ | ~pi294;
  assign new_n5121_ = ~new_n1024_ | ~new_n7197_;
  assign new_n5122_ = ~new_n1023_ | ~new_n7804_;
  assign new_n5123_ = ~new_n5008_ | ~pi453;
  assign new_n5124_ = ~new_n1261_ | ~new_n8343_;
  assign new_n5125_ = ~new_n8757_ | ~new_n6130_;
  assign new_n5126_ = ~pi422 | ~new_n6129_;
  assign new_n5127_ = ~new_n1030_ | ~pi295;
  assign new_n5128_ = ~new_n1024_ | ~new_n7094_;
  assign new_n5129_ = ~new_n1023_ | ~new_n7803_;
  assign new_n5130_ = ~new_n5008_ | ~pi454;
  assign new_n5131_ = ~new_n1261_ | ~new_n8342_;
  assign new_n5132_ = ~new_n8756_ | ~new_n6130_;
  assign new_n5133_ = ~pi423 | ~new_n6129_;
  assign new_n5134_ = ~new_n1030_ | ~pi296;
  assign new_n5135_ = ~new_n1024_ | ~new_n7095_;
  assign new_n5136_ = ~new_n1023_ | ~new_n7802_;
  assign new_n5137_ = ~new_n5008_ | ~pi455;
  assign new_n5138_ = ~new_n1261_ | ~new_n8341_;
  assign new_n5139_ = ~new_n8755_ | ~new_n6130_;
  assign new_n5140_ = ~pi424 | ~new_n6129_;
  assign new_n5141_ = ~new_n1030_ | ~pi297;
  assign new_n5142_ = ~new_n1024_ | ~new_n7196_;
  assign new_n5143_ = ~new_n1023_ | ~new_n7801_;
  assign new_n5144_ = ~new_n5008_ | ~pi456;
  assign new_n5145_ = ~new_n1261_ | ~new_n8340_;
  assign new_n5146_ = ~new_n8754_ | ~new_n6130_;
  assign new_n5147_ = ~pi425 | ~new_n6129_;
  assign new_n5148_ = ~new_n1030_ | ~pi298;
  assign new_n5149_ = ~new_n1024_ | ~new_n7194_;
  assign new_n5150_ = ~new_n1023_ | ~new_n7800_;
  assign new_n5151_ = ~new_n5008_ | ~pi457;
  assign new_n5152_ = ~new_n1261_ | ~new_n8339_;
  assign new_n5153_ = ~new_n8753_ | ~new_n6130_;
  assign new_n5154_ = ~pi426 | ~new_n6129_;
  assign new_n5155_ = ~new_n1030_ | ~pi299;
  assign new_n5156_ = ~new_n1024_ | ~new_n7192_;
  assign new_n5157_ = ~new_n1023_ | ~new_n7799_;
  assign new_n5158_ = ~new_n5008_ | ~pi458;
  assign new_n5159_ = ~new_n1261_ | ~new_n8338_;
  assign new_n5160_ = ~new_n8752_ | ~new_n6130_;
  assign new_n5161_ = ~pi427 | ~new_n6129_;
  assign new_n5162_ = ~new_n1030_ | ~pi300;
  assign new_n5163_ = ~new_n1024_ | ~new_n7188_;
  assign new_n5164_ = ~new_n1023_ | ~new_n7798_;
  assign new_n5165_ = ~new_n5008_ | ~pi459;
  assign new_n5166_ = ~new_n1261_ | ~new_n8337_;
  assign new_n5167_ = ~new_n8751_ | ~new_n6130_;
  assign new_n5168_ = ~pi428 | ~new_n6129_;
  assign new_n5169_ = ~new_n1030_ | ~pi301;
  assign new_n5170_ = ~new_n1024_ | ~new_n7096_;
  assign new_n5171_ = ~new_n1023_ | ~new_n7797_;
  assign new_n5172_ = ~new_n5008_ | ~pi460;
  assign new_n5173_ = ~new_n1261_ | ~new_n8336_;
  assign new_n5174_ = ~new_n8750_ | ~new_n6130_;
  assign new_n5175_ = ~pi429 | ~new_n6129_;
  assign new_n5176_ = ~new_n1030_ | ~pi302;
  assign new_n5177_ = ~new_n1024_ | ~new_n7187_;
  assign new_n5178_ = ~new_n1023_ | ~new_n7796_;
  assign new_n5179_ = ~new_n5008_ | ~pi461;
  assign new_n5180_ = ~new_n1261_ | ~new_n8335_;
  assign new_n5181_ = ~new_n8749_ | ~new_n6130_;
  assign new_n5182_ = ~pi430 | ~new_n6129_;
  assign new_n5183_ = ~new_n1030_ | ~pi303;
  assign new_n5184_ = ~new_n1024_ | ~new_n7185_;
  assign new_n5185_ = ~new_n1023_ | ~new_n7795_;
  assign new_n5186_ = ~new_n5008_ | ~pi462;
  assign new_n5187_ = ~new_n1261_ | ~new_n8334_;
  assign new_n5188_ = ~new_n8748_ | ~new_n6130_;
  assign new_n5189_ = ~pi431 | ~new_n6129_;
  assign new_n5190_ = ~new_n1030_ | ~pi304;
  assign new_n5191_ = ~new_n1024_ | ~new_n7183_;
  assign new_n5192_ = ~new_n1023_ | ~new_n7794_;
  assign new_n5193_ = ~new_n5008_ | ~pi463;
  assign new_n5194_ = ~new_n1261_ | ~new_n8333_;
  assign new_n5195_ = ~new_n8747_ | ~new_n6130_;
  assign new_n5196_ = ~pi432 | ~new_n6129_;
  assign new_n5197_ = ~new_n1030_ | ~pi305;
  assign new_n5198_ = ~new_n1024_ | ~new_n7181_;
  assign new_n5199_ = ~new_n1023_ | ~new_n7793_;
  assign new_n5200_ = ~new_n5008_ | ~pi464;
  assign new_n5201_ = ~new_n1261_ | ~new_n8332_;
  assign new_n5202_ = ~new_n8746_ | ~new_n6130_;
  assign new_n5203_ = ~pi433 | ~new_n6129_;
  assign new_n5204_ = ~new_n1030_ | ~pi306;
  assign new_n5205_ = ~new_n1024_ | ~new_n7179_;
  assign new_n5206_ = ~new_n1023_ | ~new_n7792_;
  assign new_n5207_ = ~new_n5008_ | ~pi465;
  assign new_n5208_ = ~new_n1261_ | ~new_n8331_;
  assign new_n5209_ = ~new_n8745_ | ~new_n6130_;
  assign new_n5210_ = ~pi434 | ~new_n6129_;
  assign new_n5211_ = ~new_n1030_ | ~pi307;
  assign new_n5212_ = ~new_n1024_ | ~new_n7177_;
  assign new_n5213_ = ~new_n1023_ | ~new_n7791_;
  assign new_n5214_ = ~new_n5008_ | ~pi466;
  assign new_n5215_ = ~new_n1261_ | ~new_n8330_;
  assign new_n5216_ = ~new_n8744_ | ~new_n6130_;
  assign new_n5217_ = ~pi435 | ~new_n6129_;
  assign new_n5218_ = ~new_n1030_ | ~pi308;
  assign new_n5219_ = ~new_n1024_ | ~new_n7175_;
  assign new_n5220_ = ~new_n1023_ | ~new_n7790_;
  assign new_n5221_ = ~new_n5008_ | ~pi467;
  assign new_n5222_ = ~new_n1261_ | ~new_n8329_;
  assign new_n5223_ = ~new_n8743_ | ~new_n6130_;
  assign new_n5224_ = ~pi436 | ~new_n6129_;
  assign new_n5225_ = ~new_n1030_ | ~pi309;
  assign new_n5226_ = ~new_n1024_ | ~new_n7173_;
  assign new_n5227_ = ~new_n1023_ | ~new_n7789_;
  assign new_n5228_ = ~new_n5008_ | ~pi468;
  assign new_n5229_ = ~new_n1261_ | ~new_n8328_;
  assign new_n5230_ = ~new_n8741_ | ~new_n6130_;
  assign new_n5231_ = ~pi437 | ~new_n6129_;
  assign new_n5232_ = ~new_n1030_ | ~pi310;
  assign new_n5233_ = ~new_n1024_ | ~new_n7171_;
  assign new_n5234_ = ~new_n1023_ | ~new_n7787_;
  assign new_n5235_ = ~new_n5008_ | ~pi469;
  assign new_n5236_ = ~new_n1261_ | ~new_n8327_;
  assign new_n5237_ = ~new_n8740_ | ~new_n6130_;
  assign new_n5238_ = ~pi438 | ~new_n6129_;
  assign new_n5239_ = ~new_n1030_ | ~pi311;
  assign new_n5240_ = ~new_n1024_ | ~new_n7169_;
  assign new_n5241_ = ~new_n1023_ | ~new_n7786_;
  assign new_n5242_ = ~new_n5008_ | ~pi470;
  assign new_n5243_ = ~pi075 | ~pi074;
  assign new_n5244_ = pi440 | pi439;
  assign new_n5245_ = ~new_n2822_;
  assign new_n5246_ = ~pi476 | ~new_n2822_;
  assign new_n5247_ = ~new_n2611_ | ~new_n1085_;
  assign new_n5248_ = ~new_n2825_;
  assign new_n5249_ = ~pi478 | ~new_n3142_;
  assign new_n5250_ = ~new_n2853_ | ~new_n5249_;
  assign new_n5251_ = ~new_n2609_ | ~new_n5250_;
  assign new_n5252_ = ~pi109 | ~new_n5251_;
  assign new_n5253_ = ~new_n2838_ | ~new_n1916_;
  assign new_n5254_ = ~new_n2610_ | ~new_n5252_;
  assign new_n5255_ = ~new_n1025_ | ~new_n1130_;
  assign new_n5256_ = ~pi482 | ~new_n5255_;
  assign new_n5257_ = ~new_n2900_ | ~pi109;
  assign new_n5258_ = ~pi483 | ~pi073;
  assign new_n5259_ = ~new_n2826_;
  assign new_n5260_ = ~new_n2613_ | ~new_n1935_;
  assign new_n5261_ = ~new_n2050_ | ~new_n3144_ | ~new_n2614_;
  assign new_n5262_ = ~pi485 | ~new_n5261_;
  assign new_n5263_ = ~new_n1201_ | ~pi110;
  assign new_n5264_ = ~new_n1200_ | ~pi118;
  assign new_n5265_ = ~new_n1199_ | ~pi126;
  assign new_n5266_ = ~new_n1198_ | ~pi134;
  assign new_n5267_ = ~new_n1196_ | ~pi142;
  assign new_n5268_ = ~new_n1195_ | ~pi150;
  assign new_n5269_ = ~new_n1194_ | ~pi158;
  assign new_n5270_ = ~new_n1193_ | ~pi166;
  assign new_n5271_ = ~new_n1191_ | ~pi174;
  assign new_n5272_ = ~new_n1190_ | ~pi182;
  assign new_n5273_ = ~new_n1189_ | ~pi190;
  assign new_n5274_ = ~new_n1188_ | ~pi198;
  assign new_n5275_ = ~new_n1186_ | ~pi206;
  assign new_n5276_ = ~new_n1184_ | ~pi214;
  assign new_n5277_ = ~new_n1182_ | ~pi222;
  assign new_n5278_ = ~new_n1180_ | ~pi230;
  assign new_n5279_ = ~new_n1201_ | ~pi111;
  assign new_n5280_ = ~new_n1200_ | ~pi119;
  assign new_n5281_ = ~new_n1199_ | ~pi127;
  assign new_n5282_ = ~new_n1198_ | ~pi135;
  assign new_n5283_ = ~new_n1196_ | ~pi143;
  assign new_n5284_ = ~new_n1195_ | ~pi151;
  assign new_n5285_ = ~new_n1194_ | ~pi159;
  assign new_n5286_ = ~new_n1193_ | ~pi167;
  assign new_n5287_ = ~new_n1191_ | ~pi175;
  assign new_n5288_ = ~new_n1190_ | ~pi183;
  assign new_n5289_ = ~new_n1189_ | ~pi191;
  assign new_n5290_ = ~new_n1188_ | ~pi199;
  assign new_n5291_ = ~new_n1186_ | ~pi207;
  assign new_n5292_ = ~new_n1184_ | ~pi215;
  assign new_n5293_ = ~new_n1182_ | ~pi223;
  assign new_n5294_ = ~new_n1180_ | ~pi231;
  assign new_n5295_ = ~new_n1201_ | ~pi112;
  assign new_n5296_ = ~new_n1200_ | ~pi120;
  assign new_n5297_ = ~new_n1199_ | ~pi128;
  assign new_n5298_ = ~new_n1198_ | ~pi136;
  assign new_n5299_ = ~new_n1196_ | ~pi144;
  assign new_n5300_ = ~new_n1195_ | ~pi152;
  assign new_n5301_ = ~new_n1194_ | ~pi160;
  assign new_n5302_ = ~new_n1193_ | ~pi168;
  assign new_n5303_ = ~new_n1191_ | ~pi176;
  assign new_n5304_ = ~new_n1190_ | ~pi184;
  assign new_n5305_ = ~new_n1189_ | ~pi192;
  assign new_n5306_ = ~new_n1188_ | ~pi200;
  assign new_n5307_ = ~new_n1186_ | ~pi208;
  assign new_n5308_ = ~new_n1184_ | ~pi216;
  assign new_n5309_ = ~new_n1182_ | ~pi224;
  assign new_n5310_ = ~new_n1180_ | ~pi232;
  assign new_n5311_ = ~new_n1201_ | ~pi113;
  assign new_n5312_ = ~new_n1200_ | ~pi121;
  assign new_n5313_ = ~new_n1199_ | ~pi129;
  assign new_n5314_ = ~new_n1198_ | ~pi137;
  assign new_n5315_ = ~new_n1196_ | ~pi145;
  assign new_n5316_ = ~new_n1195_ | ~pi153;
  assign new_n5317_ = ~new_n1194_ | ~pi161;
  assign new_n5318_ = ~new_n1193_ | ~pi169;
  assign new_n5319_ = ~new_n1191_ | ~pi177;
  assign new_n5320_ = ~new_n1190_ | ~pi185;
  assign new_n5321_ = ~new_n1189_ | ~pi193;
  assign new_n5322_ = ~new_n1188_ | ~pi201;
  assign new_n5323_ = ~new_n1186_ | ~pi209;
  assign new_n5324_ = ~new_n1184_ | ~pi217;
  assign new_n5325_ = ~new_n1182_ | ~pi225;
  assign new_n5326_ = ~new_n1201_ | ~pi114;
  assign new_n5327_ = ~new_n1200_ | ~pi122;
  assign new_n5328_ = ~new_n1199_ | ~pi130;
  assign new_n5329_ = ~new_n1198_ | ~pi138;
  assign new_n5330_ = ~new_n1196_ | ~pi146;
  assign new_n5331_ = ~new_n1195_ | ~pi154;
  assign new_n5332_ = ~new_n1194_ | ~pi162;
  assign new_n5333_ = ~new_n1193_ | ~pi170;
  assign new_n5334_ = ~new_n1191_ | ~pi178;
  assign new_n5335_ = ~new_n1190_ | ~pi186;
  assign new_n5336_ = ~new_n1189_ | ~pi194;
  assign new_n5337_ = ~new_n1188_ | ~pi202;
  assign new_n5338_ = ~new_n1186_ | ~pi210;
  assign new_n5339_ = ~new_n1184_ | ~pi218;
  assign new_n5340_ = ~new_n1182_ | ~pi226;
  assign new_n5341_ = ~new_n1180_ | ~pi234;
  assign new_n5342_ = ~new_n1201_ | ~pi115;
  assign new_n5343_ = ~new_n1200_ | ~pi123;
  assign new_n5344_ = ~new_n1199_ | ~pi131;
  assign new_n5345_ = ~new_n1198_ | ~pi139;
  assign new_n5346_ = ~new_n1196_ | ~pi147;
  assign new_n5347_ = ~new_n1195_ | ~pi155;
  assign new_n5348_ = ~new_n1194_ | ~pi163;
  assign new_n5349_ = ~new_n1193_ | ~pi171;
  assign new_n5350_ = ~new_n1191_ | ~pi179;
  assign new_n5351_ = ~new_n1190_ | ~pi187;
  assign new_n5352_ = ~new_n1189_ | ~pi195;
  assign new_n5353_ = ~new_n1188_ | ~pi203;
  assign new_n5354_ = ~new_n1186_ | ~pi211;
  assign new_n5355_ = ~new_n1184_ | ~pi219;
  assign new_n5356_ = ~new_n1182_ | ~pi227;
  assign new_n5357_ = ~new_n1180_ | ~pi235;
  assign new_n5358_ = ~new_n1201_ | ~pi116;
  assign new_n5359_ = ~new_n1200_ | ~pi124;
  assign new_n5360_ = ~new_n1199_ | ~pi132;
  assign new_n5361_ = ~new_n1198_ | ~pi140;
  assign new_n5362_ = ~new_n1196_ | ~pi148;
  assign new_n5363_ = ~new_n1195_ | ~pi156;
  assign new_n5364_ = ~new_n1194_ | ~pi164;
  assign new_n5365_ = ~new_n1193_ | ~pi172;
  assign new_n5366_ = ~new_n1191_ | ~pi180;
  assign new_n5367_ = ~new_n1190_ | ~pi188;
  assign new_n5368_ = ~new_n1189_ | ~pi196;
  assign new_n5369_ = ~new_n1188_ | ~pi204;
  assign new_n5370_ = ~new_n1186_ | ~pi212;
  assign new_n5371_ = ~new_n1184_ | ~pi220;
  assign new_n5372_ = ~new_n1182_ | ~pi228;
  assign new_n5373_ = ~new_n1180_ | ~pi236;
  assign new_n5374_ = ~new_n1201_ | ~pi117;
  assign new_n5375_ = ~new_n1200_ | ~pi125;
  assign new_n5376_ = ~new_n1199_ | ~pi133;
  assign new_n5377_ = ~new_n1198_ | ~pi141;
  assign new_n5378_ = ~new_n1196_ | ~pi149;
  assign new_n5379_ = ~new_n1195_ | ~pi157;
  assign new_n5380_ = ~new_n1194_ | ~pi165;
  assign new_n5381_ = ~new_n1193_ | ~pi173;
  assign new_n5382_ = ~new_n1191_ | ~pi181;
  assign new_n5383_ = ~new_n1190_ | ~pi189;
  assign new_n5384_ = ~new_n1189_ | ~pi197;
  assign new_n5385_ = ~new_n1188_ | ~pi205;
  assign new_n5386_ = ~new_n1186_ | ~pi213;
  assign new_n5387_ = ~new_n1184_ | ~pi221;
  assign new_n5388_ = ~new_n1182_ | ~pi229;
  assign new_n5389_ = ~new_n1180_ | ~pi237;
  assign new_n5390_ = ~new_n3105_ | ~pi107;
  assign new_n5391_ = ~new_n2056_ | ~new_n5390_;
  assign new_n5392_ = ~new_n2833_ | ~pi384;
  assign new_n5393_ = ~new_n2832_ | ~pi289;
  assign new_n5394_ = ~new_n7779_ | ~new_n1009_;
  assign new_n5395_ = ~new_n2833_ | ~pi383;
  assign new_n5396_ = ~new_n2832_ | ~pi288;
  assign new_n5397_ = ~new_n7780_ | ~new_n1009_;
  assign new_n5398_ = ~new_n2833_ | ~pi382;
  assign new_n5399_ = ~new_n2832_ | ~pi287;
  assign new_n5400_ = ~new_n7781_ | ~new_n1009_;
  assign new_n5401_ = ~new_n2833_ | ~pi381;
  assign new_n5402_ = ~new_n2832_ | ~pi286;
  assign new_n5403_ = ~new_n7782_ | ~new_n1009_;
  assign new_n5404_ = ~new_n7922_ | ~new_n5391_;
  assign new_n5405_ = ~new_n2833_ | ~pi380;
  assign new_n5406_ = ~new_n2832_ | ~pi285;
  assign new_n5407_ = ~new_n7783_ | ~new_n1009_;
  assign new_n5408_ = ~new_n7941_ | ~new_n5391_;
  assign new_n5409_ = ~new_n2833_ | ~pi379;
  assign new_n5410_ = ~new_n2832_ | ~pi284;
  assign new_n5411_ = ~new_n7784_ | ~new_n1009_;
  assign new_n5412_ = ~new_n1010_ | ~pi238;
  assign new_n5413_ = ~new_n2833_ | ~pi406;
  assign new_n5414_ = ~new_n2832_ | ~pi311;
  assign new_n5415_ = ~new_n7786_ | ~new_n1009_;
  assign new_n5416_ = ~new_n7943_ | ~new_n5391_;
  assign new_n5417_ = ~new_n2833_ | ~pi405;
  assign new_n5418_ = ~new_n2832_ | ~pi310;
  assign new_n5419_ = ~new_n7787_ | ~new_n1009_;
  assign new_n5420_ = ~new_n7942_ | ~new_n5391_;
  assign new_n5421_ = ~new_n2833_ | ~pi378;
  assign new_n5422_ = ~new_n2832_ | ~pi283;
  assign new_n5423_ = ~new_n7785_ | ~new_n1009_;
  assign new_n5424_ = ~new_n1010_ | ~pi239;
  assign new_n5425_ = ~new_n7944_ | ~new_n5391_;
  assign new_n5426_ = ~new_n2833_ | ~pi404;
  assign new_n5427_ = ~new_n2832_ | ~pi309;
  assign new_n5428_ = ~new_n7789_ | ~new_n1009_;
  assign new_n5429_ = ~new_n7945_ | ~new_n5391_;
  assign new_n5430_ = ~new_n2833_ | ~pi403;
  assign new_n5431_ = ~new_n2832_ | ~pi308;
  assign new_n5432_ = ~new_n7790_ | ~new_n1009_;
  assign new_n5433_ = ~new_n7946_ | ~new_n5391_;
  assign new_n5434_ = ~new_n2833_ | ~pi402;
  assign new_n5435_ = ~new_n2832_ | ~pi307;
  assign new_n5436_ = ~new_n7791_ | ~new_n1009_;
  assign new_n5437_ = ~new_n7947_ | ~new_n5391_;
  assign new_n5438_ = ~new_n2833_ | ~pi401;
  assign new_n5439_ = ~new_n2832_ | ~pi306;
  assign new_n5440_ = ~new_n7792_ | ~new_n1009_;
  assign new_n5441_ = ~new_n7948_ | ~new_n5391_;
  assign new_n5442_ = ~new_n2833_ | ~pi400;
  assign new_n5443_ = ~new_n2832_ | ~pi305;
  assign new_n5444_ = ~new_n7793_ | ~new_n1009_;
  assign new_n5445_ = ~new_n7949_ | ~new_n5391_;
  assign new_n5446_ = ~new_n2833_ | ~pi399;
  assign new_n5447_ = ~new_n2832_ | ~pi304;
  assign new_n5448_ = ~new_n7794_ | ~new_n1009_;
  assign new_n5449_ = ~new_n7923_ | ~new_n5391_;
  assign new_n5450_ = ~new_n2833_ | ~pi398;
  assign new_n5451_ = ~new_n2832_ | ~pi303;
  assign new_n5452_ = ~new_n7795_ | ~new_n1009_;
  assign new_n5453_ = ~new_n1381_ | ~new_n5391_;
  assign new_n5454_ = ~new_n2833_ | ~pi397;
  assign new_n5455_ = ~new_n2832_ | ~pi302;
  assign new_n5456_ = ~new_n7796_ | ~new_n1009_;
  assign new_n5457_ = ~new_n1382_ | ~new_n5391_;
  assign new_n5458_ = ~new_n2833_ | ~pi396;
  assign new_n5459_ = ~new_n2832_ | ~pi301;
  assign new_n5460_ = ~new_n7797_ | ~new_n1009_;
  assign new_n5461_ = ~new_n1383_ | ~new_n5391_;
  assign new_n5462_ = ~new_n2833_ | ~pi395;
  assign new_n5463_ = ~new_n2832_ | ~pi300;
  assign new_n5464_ = ~new_n7798_ | ~new_n1009_;
  assign new_n5465_ = ~new_n7959_ | ~new_n5391_;
  assign new_n5466_ = ~new_n2833_ | ~pi377;
  assign new_n5467_ = ~new_n2832_ | ~pi282;
  assign new_n5468_ = ~new_n7788_ | ~new_n1009_;
  assign new_n5469_ = ~new_n1010_ | ~pi240;
  assign new_n5470_ = ~new_n1384_ | ~new_n5391_;
  assign new_n5471_ = ~new_n2833_ | ~pi394;
  assign new_n5472_ = ~new_n2832_ | ~pi299;
  assign new_n5473_ = ~new_n7799_ | ~new_n1009_;
  assign new_n5474_ = ~new_n1385_ | ~new_n5391_;
  assign new_n5475_ = ~new_n2833_ | ~pi393;
  assign new_n5476_ = ~new_n2832_ | ~pi298;
  assign new_n5477_ = ~new_n7800_ | ~new_n1009_;
  assign new_n5478_ = ~new_n1386_ | ~new_n5391_;
  assign new_n5479_ = ~new_n2833_ | ~pi392;
  assign new_n5480_ = ~new_n2832_ | ~pi297;
  assign new_n5481_ = ~new_n7801_ | ~new_n1009_;
  assign new_n5482_ = ~new_n1387_ | ~new_n5391_;
  assign new_n5483_ = ~new_n2833_ | ~pi391;
  assign new_n5484_ = ~new_n2832_ | ~pi296;
  assign new_n5485_ = ~new_n7802_ | ~new_n1009_;
  assign new_n5486_ = ~new_n2833_ | ~pi390;
  assign new_n5487_ = ~new_n2832_ | ~pi295;
  assign new_n5488_ = ~new_n7803_ | ~new_n1009_;
  assign new_n5489_ = ~new_n2833_ | ~pi389;
  assign new_n5490_ = ~new_n2832_ | ~pi294;
  assign new_n5491_ = ~new_n7804_ | ~new_n1009_;
  assign new_n5492_ = ~new_n2833_ | ~pi388;
  assign new_n5493_ = ~new_n2832_ | ~pi293;
  assign new_n5494_ = ~new_n7805_ | ~new_n1009_;
  assign new_n5495_ = ~new_n2833_ | ~pi387;
  assign new_n5496_ = ~new_n2832_ | ~pi292;
  assign new_n5497_ = ~new_n7806_ | ~new_n1009_;
  assign new_n5498_ = ~new_n2833_ | ~pi386;
  assign new_n5499_ = ~new_n2832_ | ~pi291;
  assign new_n5500_ = ~new_n7807_ | ~new_n1009_;
  assign new_n5501_ = ~new_n2833_ | ~pi385;
  assign new_n5502_ = ~new_n2832_ | ~pi290;
  assign new_n5503_ = ~new_n7808_ | ~new_n1009_;
  assign new_n5504_ = ~new_n7950_ | ~new_n5391_;
  assign new_n5505_ = ~new_n2833_ | ~pi376;
  assign new_n5506_ = ~new_n2832_ | ~pi281;
  assign new_n5507_ = ~new_n7733_ | ~new_n1009_;
  assign new_n5508_ = ~new_n1010_ | ~pi241;
  assign new_n5509_ = ~new_n7951_ | ~new_n5391_;
  assign new_n5510_ = ~new_n2833_ | ~pi375;
  assign new_n5511_ = ~new_n2832_ | ~pi280;
  assign new_n5512_ = ~pi280 | ~new_n1009_;
  assign new_n5513_ = ~new_n1010_ | ~pi242;
  assign new_n5514_ = ~new_n8048_ | ~new_n5391_;
  assign new_n5515_ = ~new_n1953_ | ~new_n2083_ | ~new_n3105_;
  assign new_n5516_ = ~new_n2804_ | ~new_n8079_;
  assign new_n5517_ = ~new_n9001_ | ~new_n2853_;
  assign new_n5518_ = ~new_n2804_ | ~new_n8009_;
  assign new_n5519_ = ~new_n9012_ | ~new_n2853_;
  assign new_n5520_ = ~new_n2804_ | ~new_n8008_;
  assign new_n5521_ = ~new_n9013_ | ~new_n2853_;
  assign new_n5522_ = ~new_n2804_ | ~new_n8044_;
  assign new_n5523_ = ~new_n9014_ | ~new_n2853_;
  assign new_n5524_ = ~new_n2804_ | ~new_n8046_;
  assign new_n5525_ = ~new_n9015_ | ~new_n2853_;
  assign new_n5526_ = ~new_n2804_ | ~new_n8007_;
  assign new_n5527_ = ~new_n9020_ | ~new_n2853_;
  assign new_n5528_ = ~new_n2804_ | ~new_n8048_;
  assign new_n5529_ = ~new_n9000_ | ~new_n2853_;
  assign new_n5530_ = ~new_n3139_ | ~new_n1927_;
  assign new_n5531_ = ~new_n2804_ | ~new_n8049_;
  assign new_n5532_ = ~new_n9016_ | ~new_n2853_;
  assign new_n5533_ = ~new_n1262_ | ~new_n1928_;
  assign new_n5534_ = ~new_n2804_ | ~new_n8042_;
  assign new_n5535_ = ~new_n8999_ | ~new_n2853_;
  assign new_n5536_ = ~new_n3139_ | ~new_n1927_;
  assign new_n5537_ = ~new_n1221_ | ~pi116;
  assign new_n5538_ = ~new_n1220_ | ~pi124;
  assign new_n5539_ = ~new_n1219_ | ~pi132;
  assign new_n5540_ = ~new_n1218_ | ~pi140;
  assign new_n5541_ = ~new_n1216_ | ~pi148;
  assign new_n5542_ = ~new_n1215_ | ~pi156;
  assign new_n5543_ = ~new_n1214_ | ~pi164;
  assign new_n5544_ = ~new_n1213_ | ~pi172;
  assign new_n5545_ = ~new_n1211_ | ~pi180;
  assign new_n5546_ = ~new_n1210_ | ~pi188;
  assign new_n5547_ = ~new_n1209_ | ~pi196;
  assign new_n5548_ = ~new_n1208_ | ~pi204;
  assign new_n5549_ = ~new_n1206_ | ~pi212;
  assign new_n5550_ = ~new_n1205_ | ~pi220;
  assign new_n5551_ = ~new_n1204_ | ~pi228;
  assign new_n5552_ = ~new_n1203_ | ~pi236;
  assign new_n5553_ = ~new_n2674_ | ~new_n2675_ | ~new_n2677_ | ~new_n2676_;
  assign new_n5554_ = ~new_n2049_ | ~new_n2062_;
  assign new_n5555_ = ~new_n1221_ | ~pi117;
  assign new_n5556_ = ~new_n1220_ | ~pi125;
  assign new_n5557_ = ~new_n1219_ | ~pi133;
  assign new_n5558_ = ~new_n1218_ | ~pi141;
  assign new_n5559_ = ~new_n1216_ | ~pi149;
  assign new_n5560_ = ~new_n1215_ | ~pi157;
  assign new_n5561_ = ~new_n1214_ | ~pi165;
  assign new_n5562_ = ~new_n1213_ | ~pi173;
  assign new_n5563_ = ~new_n1211_ | ~pi181;
  assign new_n5564_ = ~new_n1210_ | ~pi189;
  assign new_n5565_ = ~new_n1209_ | ~pi197;
  assign new_n5566_ = ~new_n1208_ | ~pi205;
  assign new_n5567_ = ~new_n1206_ | ~pi213;
  assign new_n5568_ = ~new_n1205_ | ~pi221;
  assign new_n5569_ = ~new_n1204_ | ~pi229;
  assign new_n5570_ = ~new_n1203_ | ~pi237;
  assign new_n5571_ = ~new_n2678_ | ~new_n2679_ | ~new_n2681_ | ~new_n2680_;
  assign new_n5572_ = ~new_n2852_ | ~new_n1878_;
  assign new_n5573_ = ~new_n1012_ | ~new_n8660_;
  assign new_n5574_ = ~new_n2852_ | ~new_n1877_;
  assign new_n5575_ = ~new_n8658_ | ~new_n1012_;
  assign new_n5576_ = ~new_n2852_ | ~new_n1876_;
  assign new_n5577_ = ~new_n8661_ | ~new_n1012_;
  assign new_n5578_ = ~new_n2852_ | ~new_n1875_;
  assign new_n5579_ = ~new_n8665_ | ~new_n1012_;
  assign new_n5580_ = ~new_n2852_ | ~new_n1874_;
  assign new_n5581_ = ~new_n8663_ | ~new_n1012_;
  assign new_n5582_ = ~new_n7942_ | ~new_n1938_;
  assign new_n5583_ = ~new_n2852_ | ~new_n1873_;
  assign new_n5584_ = ~new_n8664_ | ~new_n1012_;
  assign new_n5585_ = ~new_n7959_ | ~new_n1938_;
  assign new_n5586_ = ~new_n1221_ | ~pi110;
  assign new_n5587_ = ~new_n1220_ | ~pi118;
  assign new_n5588_ = ~new_n1219_ | ~pi126;
  assign new_n5589_ = ~new_n1218_ | ~pi134;
  assign new_n5590_ = ~new_n1216_ | ~pi142;
  assign new_n5591_ = ~new_n1215_ | ~pi150;
  assign new_n5592_ = ~new_n1214_ | ~pi158;
  assign new_n5593_ = ~new_n1213_ | ~pi166;
  assign new_n5594_ = ~new_n1211_ | ~pi174;
  assign new_n5595_ = ~new_n1210_ | ~pi182;
  assign new_n5596_ = ~new_n1209_ | ~pi190;
  assign new_n5597_ = ~new_n1208_ | ~pi198;
  assign new_n5598_ = ~new_n1206_ | ~pi206;
  assign new_n5599_ = ~new_n1205_ | ~pi214;
  assign new_n5600_ = ~new_n1204_ | ~pi222;
  assign new_n5601_ = ~new_n1203_ | ~pi230;
  assign new_n5602_ = ~new_n2682_ | ~new_n2683_ | ~new_n2685_ | ~new_n2684_;
  assign new_n5603_ = ~new_n1221_ | ~pi111;
  assign new_n5604_ = ~new_n1220_ | ~pi119;
  assign new_n5605_ = ~new_n1219_ | ~pi127;
  assign new_n5606_ = ~new_n1218_ | ~pi135;
  assign new_n5607_ = ~new_n1216_ | ~pi143;
  assign new_n5608_ = ~new_n1215_ | ~pi151;
  assign new_n5609_ = ~new_n1214_ | ~pi159;
  assign new_n5610_ = ~new_n1213_ | ~pi167;
  assign new_n5611_ = ~new_n1211_ | ~pi175;
  assign new_n5612_ = ~new_n1210_ | ~pi183;
  assign new_n5613_ = ~new_n1209_ | ~pi191;
  assign new_n5614_ = ~new_n1208_ | ~pi199;
  assign new_n5615_ = ~new_n1206_ | ~pi207;
  assign new_n5616_ = ~new_n1205_ | ~pi215;
  assign new_n5617_ = ~new_n1204_ | ~pi223;
  assign new_n5618_ = ~new_n1203_ | ~pi231;
  assign new_n5619_ = ~new_n2686_ | ~new_n2687_ | ~new_n2689_ | ~new_n2688_;
  assign new_n5620_ = ~new_n1221_ | ~pi112;
  assign new_n5621_ = ~new_n1220_ | ~pi120;
  assign new_n5622_ = ~new_n1219_ | ~pi128;
  assign new_n5623_ = ~new_n1218_ | ~pi136;
  assign new_n5624_ = ~new_n1216_ | ~pi144;
  assign new_n5625_ = ~new_n1215_ | ~pi152;
  assign new_n5626_ = ~new_n1214_ | ~pi160;
  assign new_n5627_ = ~new_n1213_ | ~pi168;
  assign new_n5628_ = ~new_n1211_ | ~pi176;
  assign new_n5629_ = ~new_n1210_ | ~pi184;
  assign new_n5630_ = ~new_n1209_ | ~pi192;
  assign new_n5631_ = ~new_n1208_ | ~pi200;
  assign new_n5632_ = ~new_n1206_ | ~pi208;
  assign new_n5633_ = ~new_n1205_ | ~pi216;
  assign new_n5634_ = ~new_n1204_ | ~pi224;
  assign new_n5635_ = ~new_n1203_ | ~pi232;
  assign new_n5636_ = ~new_n2690_ | ~new_n2691_ | ~new_n2693_ | ~new_n2692_;
  assign new_n5637_ = ~new_n1221_ | ~pi113;
  assign new_n5638_ = ~new_n1220_ | ~pi121;
  assign new_n5639_ = ~new_n1219_ | ~pi129;
  assign new_n5640_ = ~new_n1218_ | ~pi137;
  assign new_n5641_ = ~new_n1216_ | ~pi145;
  assign new_n5642_ = ~new_n1215_ | ~pi153;
  assign new_n5643_ = ~new_n1214_ | ~pi161;
  assign new_n5644_ = ~new_n1213_ | ~pi169;
  assign new_n5645_ = ~new_n1211_ | ~pi177;
  assign new_n5646_ = ~new_n1210_ | ~pi185;
  assign new_n5647_ = ~new_n1209_ | ~pi193;
  assign new_n5648_ = ~new_n1208_ | ~pi201;
  assign new_n5649_ = ~new_n1206_ | ~pi209;
  assign new_n5650_ = ~new_n1205_ | ~pi217;
  assign new_n5651_ = ~new_n1204_ | ~pi225;
  assign new_n5652_ = ~new_n1221_ | ~pi114;
  assign new_n5653_ = ~new_n1220_ | ~pi122;
  assign new_n5654_ = ~new_n1219_ | ~pi130;
  assign new_n5655_ = ~new_n1218_ | ~pi138;
  assign new_n5656_ = ~new_n1216_ | ~pi146;
  assign new_n5657_ = ~new_n1215_ | ~pi154;
  assign new_n5658_ = ~new_n1214_ | ~pi162;
  assign new_n5659_ = ~new_n1213_ | ~pi170;
  assign new_n5660_ = ~new_n1211_ | ~pi178;
  assign new_n5661_ = ~new_n1210_ | ~pi186;
  assign new_n5662_ = ~new_n1209_ | ~pi194;
  assign new_n5663_ = ~new_n1208_ | ~pi202;
  assign new_n5664_ = ~new_n1206_ | ~pi210;
  assign new_n5665_ = ~new_n1205_ | ~pi218;
  assign new_n5666_ = ~new_n1204_ | ~pi226;
  assign new_n5667_ = ~new_n1203_ | ~pi234;
  assign new_n5668_ = ~new_n2698_ | ~new_n2699_ | ~new_n2701_ | ~new_n2700_;
  assign new_n5669_ = ~new_n1221_ | ~pi115;
  assign new_n5670_ = ~new_n1220_ | ~pi123;
  assign new_n5671_ = ~new_n1219_ | ~pi131;
  assign new_n5672_ = ~new_n1218_ | ~pi139;
  assign new_n5673_ = ~new_n1216_ | ~pi147;
  assign new_n5674_ = ~new_n1215_ | ~pi155;
  assign new_n5675_ = ~new_n1214_ | ~pi163;
  assign new_n5676_ = ~new_n1213_ | ~pi171;
  assign new_n5677_ = ~new_n1211_ | ~pi179;
  assign new_n5678_ = ~new_n1210_ | ~pi187;
  assign new_n5679_ = ~new_n1209_ | ~pi195;
  assign new_n5680_ = ~new_n1208_ | ~pi203;
  assign new_n5681_ = ~new_n1206_ | ~pi211;
  assign new_n5682_ = ~new_n1205_ | ~pi219;
  assign new_n5683_ = ~new_n1204_ | ~pi227;
  assign new_n5684_ = ~new_n1203_ | ~pi235;
  assign new_n5685_ = ~new_n2702_ | ~new_n2703_ | ~new_n2705_ | ~new_n2704_;
  assign new_n5686_ = ~new_n2852_ | ~new_n1872_;
  assign new_n5687_ = ~new_n8659_ | ~new_n1012_;
  assign new_n5688_ = ~new_n7950_ | ~new_n1938_;
  assign new_n5689_ = ~new_n2852_ | ~new_n1871_;
  assign new_n5690_ = ~new_n8662_ | ~new_n1012_;
  assign new_n5691_ = ~new_n7951_ | ~new_n1938_;
  assign new_n5692_ = ~new_n2851_ | ~new_n1878_;
  assign new_n5693_ = ~new_n2837_ | ~pi230;
  assign new_n5694_ = ~new_n2851_ | ~new_n1877_;
  assign new_n5695_ = ~new_n2837_ | ~pi231;
  assign new_n5696_ = ~new_n2851_ | ~new_n1876_;
  assign new_n5697_ = ~new_n2837_ | ~pi232;
  assign new_n5698_ = ~new_n2851_ | ~new_n1875_;
  assign new_n5699_ = ~new_n2851_ | ~new_n1874_;
  assign new_n5700_ = ~new_n2837_ | ~pi234;
  assign new_n5701_ = ~new_n2851_ | ~new_n1873_;
  assign new_n5702_ = ~new_n2837_ | ~pi235;
  assign new_n5703_ = ~new_n2851_ | ~new_n1872_;
  assign new_n5704_ = ~new_n2837_ | ~pi236;
  assign new_n5705_ = ~new_n2851_ | ~new_n1871_;
  assign new_n5706_ = ~new_n1878_ | ~new_n3045_;
  assign new_n5707_ = ~new_n2837_ | ~pi237;
  assign new_n5708_ = ~new_n2072_ | ~new_n2071_;
  assign new_n5709_ = ~pi239 | ~new_n1908_;
  assign new_n5710_ = ~new_n2089_;
  assign new_n5711_ = ~new_n1239_ | ~pi166;
  assign new_n5712_ = ~new_n1238_ | ~pi158;
  assign new_n5713_ = ~new_n1237_ | ~pi150;
  assign new_n5714_ = ~new_n1236_ | ~pi142;
  assign new_n5715_ = ~new_n1234_ | ~pi134;
  assign new_n5716_ = ~new_n1233_ | ~pi126;
  assign new_n5717_ = ~new_n1232_ | ~pi118;
  assign new_n5718_ = ~new_n1231_ | ~pi110;
  assign new_n5719_ = ~new_n1230_ | ~pi230;
  assign new_n5720_ = ~new_n1229_ | ~pi222;
  assign new_n5721_ = ~new_n1228_ | ~pi214;
  assign new_n5722_ = ~new_n1227_ | ~pi206;
  assign new_n5723_ = ~new_n1225_ | ~pi198;
  assign new_n5724_ = ~new_n1224_ | ~pi190;
  assign new_n5725_ = ~new_n1223_ | ~pi182;
  assign new_n5726_ = ~new_n1222_ | ~pi174;
  assign new_n5727_ = ~new_n2708_ | ~new_n2709_ | ~new_n2711_ | ~new_n2710_;
  assign new_n5728_ = ~new_n2069_ | ~new_n2065_;
  assign new_n5729_ = ~new_n2718_ | ~new_n2836_;
  assign new_n5730_ = ~new_n5729_ | ~new_n2066_;
  assign new_n5731_ = ~new_n3148_ | ~new_n1922_;
  assign new_n5732_ = ~new_n1889_;
  assign new_n5733_ = ~new_n2038_ | ~new_n2799_ | ~new_n3045_ | ~new_n3148_;
  assign new_n5734_ = ~new_n2834_ | ~pi109;
  assign new_n5735_ = ~new_n2712_ | ~new_n1889_;
  assign new_n5736_ = ~new_n2095_;
  assign new_n5737_ = ~new_n6274_ | ~new_n2095_ | ~new_n4137_;
  assign new_n5738_ = ~new_n2839_ | ~new_n5737_;
  assign new_n5739_ = ~new_n2094_;
  assign new_n5740_ = ~pi244 | ~new_n1941_;
  assign new_n5741_ = ~pi239 | ~new_n2094_;
  assign new_n5742_ = ~new_n2848_ | ~new_n2004_;
  assign new_n5743_ = ~new_n1239_ | ~pi167;
  assign new_n5744_ = ~new_n1238_ | ~pi159;
  assign new_n5745_ = ~new_n1237_ | ~pi151;
  assign new_n5746_ = ~new_n1236_ | ~pi143;
  assign new_n5747_ = ~new_n1234_ | ~pi135;
  assign new_n5748_ = ~new_n1233_ | ~pi127;
  assign new_n5749_ = ~new_n1232_ | ~pi119;
  assign new_n5750_ = ~new_n1231_ | ~pi111;
  assign new_n5751_ = ~new_n1230_ | ~pi231;
  assign new_n5752_ = ~new_n1229_ | ~pi223;
  assign new_n5753_ = ~new_n1228_ | ~pi215;
  assign new_n5754_ = ~new_n1227_ | ~pi207;
  assign new_n5755_ = ~new_n1225_ | ~pi199;
  assign new_n5756_ = ~new_n1224_ | ~pi191;
  assign new_n5757_ = ~new_n1223_ | ~pi183;
  assign new_n5758_ = ~new_n1222_ | ~pi175;
  assign new_n5759_ = ~new_n2724_ | ~new_n2725_ | ~new_n2727_ | ~new_n2726_;
  assign new_n5760_ = ~new_n1239_ | ~pi168;
  assign new_n5761_ = ~new_n1238_ | ~pi160;
  assign new_n5762_ = ~new_n1237_ | ~pi152;
  assign new_n5763_ = ~new_n1236_ | ~pi144;
  assign new_n5764_ = ~new_n1234_ | ~pi136;
  assign new_n5765_ = ~new_n1233_ | ~pi128;
  assign new_n5766_ = ~new_n1232_ | ~pi120;
  assign new_n5767_ = ~new_n1231_ | ~pi112;
  assign new_n5768_ = ~new_n1230_ | ~pi232;
  assign new_n5769_ = ~new_n1229_ | ~pi224;
  assign new_n5770_ = ~new_n1228_ | ~pi216;
  assign new_n5771_ = ~new_n1227_ | ~pi208;
  assign new_n5772_ = ~new_n1225_ | ~pi200;
  assign new_n5773_ = ~new_n1224_ | ~pi192;
  assign new_n5774_ = ~new_n1223_ | ~pi184;
  assign new_n5775_ = ~new_n1222_ | ~pi176;
  assign new_n5776_ = ~new_n2728_ | ~new_n2729_ | ~new_n2731_ | ~new_n2730_;
  assign new_n5777_ = ~new_n1239_ | ~pi169;
  assign new_n5778_ = ~new_n1238_ | ~pi161;
  assign new_n5779_ = ~new_n1237_ | ~pi153;
  assign new_n5780_ = ~new_n1236_ | ~pi145;
  assign new_n5781_ = ~new_n1234_ | ~pi137;
  assign new_n5782_ = ~new_n1233_ | ~pi129;
  assign new_n5783_ = ~new_n1232_ | ~pi121;
  assign new_n5784_ = ~new_n1231_ | ~pi113;
  assign new_n5785_ = ~new_n1229_ | ~pi225;
  assign new_n5786_ = ~new_n1228_ | ~pi217;
  assign new_n5787_ = ~new_n1227_ | ~pi209;
  assign new_n5788_ = ~new_n1225_ | ~pi201;
  assign new_n5789_ = ~new_n1224_ | ~pi193;
  assign new_n5790_ = ~new_n1223_ | ~pi185;
  assign new_n5791_ = ~new_n1222_ | ~pi177;
  assign new_n5792_ = ~new_n1239_ | ~pi170;
  assign new_n5793_ = ~new_n1238_ | ~pi162;
  assign new_n5794_ = ~new_n1237_ | ~pi154;
  assign new_n5795_ = ~new_n1236_ | ~pi146;
  assign new_n5796_ = ~new_n1234_ | ~pi138;
  assign new_n5797_ = ~new_n1233_ | ~pi130;
  assign new_n5798_ = ~new_n1232_ | ~pi122;
  assign new_n5799_ = ~new_n1231_ | ~pi114;
  assign new_n5800_ = ~new_n1230_ | ~pi234;
  assign new_n5801_ = ~new_n1229_ | ~pi226;
  assign new_n5802_ = ~new_n1228_ | ~pi218;
  assign new_n5803_ = ~new_n1227_ | ~pi210;
  assign new_n5804_ = ~new_n1225_ | ~pi202;
  assign new_n5805_ = ~new_n1224_ | ~pi194;
  assign new_n5806_ = ~new_n1223_ | ~pi186;
  assign new_n5807_ = ~new_n1222_ | ~pi178;
  assign new_n5808_ = ~new_n2737_ | ~new_n2738_ | ~new_n2740_ | ~new_n2739_;
  assign new_n5809_ = ~new_n1239_ | ~pi171;
  assign new_n5810_ = ~new_n1238_ | ~pi163;
  assign new_n5811_ = ~new_n1237_ | ~pi155;
  assign new_n5812_ = ~new_n1236_ | ~pi147;
  assign new_n5813_ = ~new_n1234_ | ~pi139;
  assign new_n5814_ = ~new_n1233_ | ~pi131;
  assign new_n5815_ = ~new_n1232_ | ~pi123;
  assign new_n5816_ = ~new_n1231_ | ~pi115;
  assign new_n5817_ = ~new_n1230_ | ~pi235;
  assign new_n5818_ = ~new_n1229_ | ~pi227;
  assign new_n5819_ = ~new_n1228_ | ~pi219;
  assign new_n5820_ = ~new_n1227_ | ~pi211;
  assign new_n5821_ = ~new_n1225_ | ~pi203;
  assign new_n5822_ = ~new_n1224_ | ~pi195;
  assign new_n5823_ = ~new_n1223_ | ~pi187;
  assign new_n5824_ = ~new_n1222_ | ~pi179;
  assign new_n5825_ = ~new_n2741_ | ~new_n2742_ | ~new_n2744_ | ~new_n2743_;
  assign new_n5826_ = ~new_n1239_ | ~pi172;
  assign new_n5827_ = ~new_n1238_ | ~pi164;
  assign new_n5828_ = ~new_n1237_ | ~pi156;
  assign new_n5829_ = ~new_n1236_ | ~pi148;
  assign new_n5830_ = ~new_n1234_ | ~pi140;
  assign new_n5831_ = ~new_n1233_ | ~pi132;
  assign new_n5832_ = ~new_n1232_ | ~pi124;
  assign new_n5833_ = ~new_n1231_ | ~pi116;
  assign new_n5834_ = ~new_n1230_ | ~pi236;
  assign new_n5835_ = ~new_n1229_ | ~pi228;
  assign new_n5836_ = ~new_n1228_ | ~pi220;
  assign new_n5837_ = ~new_n1227_ | ~pi212;
  assign new_n5838_ = ~new_n1225_ | ~pi204;
  assign new_n5839_ = ~new_n1224_ | ~pi196;
  assign new_n5840_ = ~new_n1223_ | ~pi188;
  assign new_n5841_ = ~new_n1222_ | ~pi180;
  assign new_n5842_ = ~new_n2745_ | ~new_n2746_ | ~new_n2748_ | ~new_n2747_;
  assign new_n5843_ = ~new_n1239_ | ~pi173;
  assign new_n5844_ = ~new_n1238_ | ~pi165;
  assign new_n5845_ = ~new_n1237_ | ~pi157;
  assign new_n5846_ = ~new_n1236_ | ~pi149;
  assign new_n5847_ = ~new_n1234_ | ~pi141;
  assign new_n5848_ = ~new_n1233_ | ~pi133;
  assign new_n5849_ = ~new_n1232_ | ~pi125;
  assign new_n5850_ = ~new_n1231_ | ~pi117;
  assign new_n5851_ = ~new_n1230_ | ~pi237;
  assign new_n5852_ = ~new_n1229_ | ~pi229;
  assign new_n5853_ = ~new_n1228_ | ~pi221;
  assign new_n5854_ = ~new_n1227_ | ~pi213;
  assign new_n5855_ = ~new_n1225_ | ~pi205;
  assign new_n5856_ = ~new_n1224_ | ~pi197;
  assign new_n5857_ = ~new_n1223_ | ~pi189;
  assign new_n5858_ = ~new_n1222_ | ~pi181;
  assign new_n5859_ = ~new_n2749_ | ~new_n2750_ | ~new_n2752_ | ~new_n2751_;
  assign new_n5860_ = ~pi245 | ~new_n1941_;
  assign new_n5861_ = ~new_n2848_ | ~new_n2099_;
  assign new_n5862_ = ~pi246 | ~new_n1941_;
  assign new_n5863_ = ~new_n2848_ | ~new_n1879_;
  assign new_n5864_ = ~new_n2828_;
  assign new_n5865_ = ~new_n1259_ | ~pi166;
  assign new_n5866_ = ~new_n1258_ | ~pi158;
  assign new_n5867_ = ~new_n1257_ | ~pi150;
  assign new_n5868_ = ~new_n1256_ | ~pi142;
  assign new_n5869_ = ~new_n1254_ | ~pi134;
  assign new_n5870_ = ~new_n1253_ | ~pi126;
  assign new_n5871_ = ~new_n1252_ | ~pi118;
  assign new_n5872_ = ~new_n1251_ | ~pi110;
  assign new_n5873_ = ~new_n1249_ | ~pi230;
  assign new_n5874_ = ~new_n1248_ | ~pi222;
  assign new_n5875_ = ~new_n1247_ | ~pi214;
  assign new_n5876_ = ~new_n1246_ | ~pi206;
  assign new_n5877_ = ~new_n1244_ | ~pi198;
  assign new_n5878_ = ~new_n1243_ | ~pi190;
  assign new_n5879_ = ~new_n1242_ | ~pi182;
  assign new_n5880_ = ~new_n1241_ | ~pi174;
  assign new_n5881_ = ~new_n2766_ | ~new_n2767_ | ~new_n2769_ | ~new_n2768_;
  assign new_n5882_ = ~new_n1259_ | ~pi167;
  assign new_n5883_ = ~new_n1258_ | ~pi159;
  assign new_n5884_ = ~new_n1257_ | ~pi151;
  assign new_n5885_ = ~new_n1256_ | ~pi143;
  assign new_n5886_ = ~new_n1254_ | ~pi135;
  assign new_n5887_ = ~new_n1253_ | ~pi127;
  assign new_n5888_ = ~new_n1252_ | ~pi119;
  assign new_n5889_ = ~new_n1251_ | ~pi111;
  assign new_n5890_ = ~new_n1249_ | ~pi231;
  assign new_n5891_ = ~new_n1248_ | ~pi223;
  assign new_n5892_ = ~new_n1247_ | ~pi215;
  assign new_n5893_ = ~new_n1246_ | ~pi207;
  assign new_n5894_ = ~new_n1244_ | ~pi199;
  assign new_n5895_ = ~new_n1243_ | ~pi191;
  assign new_n5896_ = ~new_n1242_ | ~pi183;
  assign new_n5897_ = ~new_n1241_ | ~pi175;
  assign new_n5898_ = ~new_n2770_ | ~new_n2771_ | ~new_n2773_ | ~new_n2772_;
  assign new_n5899_ = ~new_n1259_ | ~pi168;
  assign new_n5900_ = ~new_n1258_ | ~pi160;
  assign new_n5901_ = ~new_n1257_ | ~pi152;
  assign new_n5902_ = ~new_n1256_ | ~pi144;
  assign new_n5903_ = ~new_n1254_ | ~pi136;
  assign new_n5904_ = ~new_n1253_ | ~pi128;
  assign new_n5905_ = ~new_n1252_ | ~pi120;
  assign new_n5906_ = ~new_n1251_ | ~pi112;
  assign new_n5907_ = ~new_n1249_ | ~pi232;
  assign new_n5908_ = ~new_n1248_ | ~pi224;
  assign new_n5909_ = ~new_n1247_ | ~pi216;
  assign new_n5910_ = ~new_n1246_ | ~pi208;
  assign new_n5911_ = ~new_n1244_ | ~pi200;
  assign new_n5912_ = ~new_n1243_ | ~pi192;
  assign new_n5913_ = ~new_n1242_ | ~pi184;
  assign new_n5914_ = ~new_n1241_ | ~pi176;
  assign new_n5915_ = ~new_n2774_ | ~new_n2775_ | ~new_n2777_ | ~new_n2776_;
  assign new_n5916_ = ~new_n1259_ | ~pi169;
  assign new_n5917_ = ~new_n1258_ | ~pi161;
  assign new_n5918_ = ~new_n1257_ | ~pi153;
  assign new_n5919_ = ~new_n1256_ | ~pi145;
  assign new_n5920_ = ~new_n1254_ | ~pi137;
  assign new_n5921_ = ~new_n1253_ | ~pi129;
  assign new_n5922_ = ~new_n1252_ | ~pi121;
  assign new_n5923_ = ~new_n1251_ | ~pi113;
  assign new_n5924_ = ~new_n1248_ | ~pi225;
  assign new_n5925_ = ~new_n1247_ | ~pi217;
  assign new_n5926_ = ~new_n1246_ | ~pi209;
  assign new_n5927_ = ~new_n1244_ | ~pi201;
  assign new_n5928_ = ~new_n1243_ | ~pi193;
  assign new_n5929_ = ~new_n1242_ | ~pi185;
  assign new_n5930_ = ~new_n1241_ | ~pi177;
  assign new_n5931_ = ~new_n1259_ | ~pi170;
  assign new_n5932_ = ~new_n1258_ | ~pi162;
  assign new_n5933_ = ~new_n1257_ | ~pi154;
  assign new_n5934_ = ~new_n1256_ | ~pi146;
  assign new_n5935_ = ~new_n1254_ | ~pi138;
  assign new_n5936_ = ~new_n1253_ | ~pi130;
  assign new_n5937_ = ~new_n1252_ | ~pi122;
  assign new_n5938_ = ~new_n1251_ | ~pi114;
  assign new_n5939_ = ~new_n1249_ | ~pi234;
  assign new_n5940_ = ~new_n1248_ | ~pi226;
  assign new_n5941_ = ~new_n1247_ | ~pi218;
  assign new_n5942_ = ~new_n1246_ | ~pi210;
  assign new_n5943_ = ~new_n1244_ | ~pi202;
  assign new_n5944_ = ~new_n1243_ | ~pi194;
  assign new_n5945_ = ~new_n1242_ | ~pi186;
  assign new_n5946_ = ~new_n1241_ | ~pi178;
  assign new_n5947_ = ~new_n2782_ | ~new_n2783_ | ~new_n2785_ | ~new_n2784_;
  assign new_n5948_ = ~new_n1259_ | ~pi171;
  assign new_n5949_ = ~new_n1258_ | ~pi163;
  assign new_n5950_ = ~new_n1257_ | ~pi155;
  assign new_n5951_ = ~new_n1256_ | ~pi147;
  assign new_n5952_ = ~new_n1254_ | ~pi139;
  assign new_n5953_ = ~new_n1253_ | ~pi131;
  assign new_n5954_ = ~new_n1252_ | ~pi123;
  assign new_n5955_ = ~new_n1251_ | ~pi115;
  assign new_n5956_ = ~new_n1249_ | ~pi235;
  assign new_n5957_ = ~new_n1248_ | ~pi227;
  assign new_n5958_ = ~new_n1247_ | ~pi219;
  assign new_n5959_ = ~new_n1246_ | ~pi211;
  assign new_n5960_ = ~new_n1244_ | ~pi203;
  assign new_n5961_ = ~new_n1243_ | ~pi195;
  assign new_n5962_ = ~new_n1242_ | ~pi187;
  assign new_n5963_ = ~new_n1241_ | ~pi179;
  assign new_n5964_ = ~new_n2786_ | ~new_n2787_ | ~new_n2789_ | ~new_n2788_;
  assign new_n5965_ = ~new_n1259_ | ~pi172;
  assign new_n5966_ = ~new_n1258_ | ~pi164;
  assign new_n5967_ = ~new_n1257_ | ~pi156;
  assign new_n5968_ = ~new_n1256_ | ~pi148;
  assign new_n5969_ = ~new_n1254_ | ~pi140;
  assign new_n5970_ = ~new_n1253_ | ~pi132;
  assign new_n5971_ = ~new_n1252_ | ~pi124;
  assign new_n5972_ = ~new_n1251_ | ~pi116;
  assign new_n5973_ = ~new_n1249_ | ~pi236;
  assign new_n5974_ = ~new_n1248_ | ~pi228;
  assign new_n5975_ = ~new_n1247_ | ~pi220;
  assign new_n5976_ = ~new_n1246_ | ~pi212;
  assign new_n5977_ = ~new_n1244_ | ~pi204;
  assign new_n5978_ = ~new_n1243_ | ~pi196;
  assign new_n5979_ = ~new_n1242_ | ~pi188;
  assign new_n5980_ = ~new_n1241_ | ~pi180;
  assign new_n5981_ = ~new_n2790_ | ~new_n2791_ | ~new_n2793_ | ~new_n2792_;
  assign new_n5982_ = ~new_n1259_ | ~pi173;
  assign new_n5983_ = ~new_n1258_ | ~pi165;
  assign new_n5984_ = ~new_n1257_ | ~pi157;
  assign new_n5985_ = ~new_n1256_ | ~pi149;
  assign new_n5986_ = ~new_n1254_ | ~pi141;
  assign new_n5987_ = ~new_n1253_ | ~pi133;
  assign new_n5988_ = ~new_n1252_ | ~pi125;
  assign new_n5989_ = ~new_n1251_ | ~pi117;
  assign new_n5990_ = ~new_n1249_ | ~pi237;
  assign new_n5991_ = ~new_n1248_ | ~pi229;
  assign new_n5992_ = ~new_n1247_ | ~pi221;
  assign new_n5993_ = ~new_n1246_ | ~pi213;
  assign new_n5994_ = ~new_n1244_ | ~pi205;
  assign new_n5995_ = ~new_n1243_ | ~pi197;
  assign new_n5996_ = ~new_n1242_ | ~pi189;
  assign new_n5997_ = ~new_n1241_ | ~pi181;
  assign new_n5998_ = ~new_n2794_ | ~new_n2795_ | ~new_n2797_ | ~new_n2796_;
  assign new_n5999_ = ~new_n2879_ | ~new_n2876_ | ~new_n1011_;
  assign new_n6000_ = ~new_n2798_ | ~new_n5732_;
  assign new_n6001_ = ~new_n2040_ | ~new_n2054_;
  assign new_n6002_ = ~new_n2879_ | ~new_n6001_;
  assign new_n6003_ = ~new_n2835_ | ~new_n1109_;
  assign new_n6004_ = ~new_n6000_ | ~new_n1915_;
  assign new_n6005_ = ~new_n2853_ | ~new_n5733_;
  assign new_n6006_ = ~new_n2805_ | ~new_n2853_;
  assign new_n6007_ = ~new_n1108_ | ~new_n2855_;
  assign new_n6008_ = ~new_n6006_ | ~new_n6007_ | ~new_n2840_ | ~new_n2064_ | ~new_n2078_;
  assign new_n6009_ = ~new_n8877_ | ~new_n6008_;
  assign new_n6010_ = ~new_n8938_ | ~new_n1011_;
  assign new_n6011_ = ~new_n8890_ | ~new_n6008_;
  assign new_n6012_ = ~new_n8951_ | ~new_n1011_;
  assign new_n6013_ = ~new_n8891_ | ~new_n6008_;
  assign new_n6014_ = ~new_n8952_ | ~new_n1011_;
  assign new_n6015_ = ~new_n8892_ | ~new_n6008_;
  assign new_n6016_ = ~new_n8953_ | ~new_n1011_;
  assign new_n6017_ = ~new_n8893_ | ~new_n6008_;
  assign new_n6018_ = ~new_n8954_ | ~new_n1011_;
  assign new_n6019_ = ~new_n8878_ | ~new_n6008_;
  assign new_n6020_ = ~new_n8939_ | ~new_n1011_;
  assign new_n6021_ = ~new_n8890_ | ~new_n2837_;
  assign new_n6022_ = ~pi238 | ~new_n1938_;
  assign new_n6023_ = ~new_n8891_ | ~new_n2837_;
  assign new_n6024_ = ~pi239 | ~new_n1938_;
  assign new_n6025_ = ~pi109 | ~new_n2818_;
  assign new_n6026_ = ~new_n2064_ | ~new_n6025_;
  assign new_n6027_ = ~new_n8892_ | ~new_n2837_;
  assign new_n6028_ = ~pi240 | ~new_n1938_;
  assign new_n6029_ = ~new_n1107_ | ~new_n1915_;
  assign new_n6030_ = ~new_n8893_ | ~new_n2837_;
  assign new_n6031_ = ~pi241 | ~new_n1938_;
  assign new_n6032_ = ~new_n1108_ | ~new_n1928_;
  assign new_n6033_ = ~new_n8878_ | ~new_n2837_;
  assign new_n6034_ = ~pi242 | ~new_n1938_;
  assign new_n6035_ = ~new_n2037_ | ~new_n1934_;
  assign new_n6036_ = ~new_n1928_ | ~new_n2093_;
  assign new_n6037_ = ~pi257 | ~new_n6036_;
  assign new_n6038_ = ~pi416 | ~new_n6035_;
  assign new_n6039_ = ~pi256 | ~new_n6036_;
  assign new_n6040_ = ~pi415 | ~new_n6035_;
  assign new_n6041_ = ~pi255 | ~new_n6036_;
  assign new_n6042_ = ~pi414 | ~new_n6035_;
  assign new_n6043_ = ~pi254 | ~new_n6036_;
  assign new_n6044_ = ~pi413 | ~new_n6035_;
  assign new_n6045_ = ~pi253 | ~new_n6036_;
  assign new_n6046_ = ~pi412 | ~new_n6035_;
  assign new_n6047_ = ~pi252 | ~new_n6036_;
  assign new_n6048_ = ~pi411 | ~new_n6035_;
  assign new_n6049_ = ~pi279 | ~new_n6036_;
  assign new_n6050_ = ~pi438 | ~new_n6035_;
  assign new_n6051_ = ~pi278 | ~new_n6036_;
  assign new_n6052_ = ~pi437 | ~new_n6035_;
  assign new_n6053_ = ~pi251 | ~new_n6036_;
  assign new_n6054_ = ~pi410 | ~new_n6035_;
  assign new_n6055_ = ~pi277 | ~new_n6036_;
  assign new_n6056_ = ~pi436 | ~new_n6035_;
  assign new_n6057_ = ~pi276 | ~new_n6036_;
  assign new_n6058_ = ~pi435 | ~new_n6035_;
  assign new_n6059_ = ~pi275 | ~new_n6036_;
  assign new_n6060_ = ~pi434 | ~new_n6035_;
  assign new_n6061_ = ~pi274 | ~new_n6036_;
  assign new_n6062_ = ~pi433 | ~new_n6035_;
  assign new_n6063_ = ~pi273 | ~new_n6036_;
  assign new_n6064_ = ~pi432 | ~new_n6035_;
  assign new_n6065_ = ~pi272 | ~new_n6036_;
  assign new_n6066_ = ~pi431 | ~new_n6035_;
  assign new_n6067_ = ~pi271 | ~new_n6036_;
  assign new_n6068_ = ~pi430 | ~new_n6035_;
  assign new_n6069_ = ~pi270 | ~new_n6036_;
  assign new_n6070_ = ~pi429 | ~new_n6035_;
  assign new_n6071_ = ~pi269 | ~new_n6036_;
  assign new_n6072_ = ~pi428 | ~new_n6035_;
  assign new_n6073_ = ~pi268 | ~new_n6036_;
  assign new_n6074_ = ~pi427 | ~new_n6035_;
  assign new_n6075_ = ~pi250 | ~new_n6036_;
  assign new_n6076_ = ~pi409 | ~new_n6035_;
  assign new_n6077_ = ~pi267 | ~new_n6036_;
  assign new_n6078_ = ~pi426 | ~new_n6035_;
  assign new_n6079_ = ~pi266 | ~new_n6036_;
  assign new_n6080_ = ~pi425 | ~new_n6035_;
  assign new_n6081_ = ~pi265 | ~new_n6036_;
  assign new_n6082_ = ~pi424 | ~new_n6035_;
  assign new_n6083_ = ~pi264 | ~new_n6036_;
  assign new_n6084_ = ~pi423 | ~new_n6035_;
  assign new_n6085_ = ~pi263 | ~new_n6036_;
  assign new_n6086_ = ~pi422 | ~new_n6035_;
  assign new_n6087_ = ~pi262 | ~new_n6036_;
  assign new_n6088_ = ~pi421 | ~new_n6035_;
  assign new_n6089_ = ~pi261 | ~new_n6036_;
  assign new_n6090_ = ~pi420 | ~new_n6035_;
  assign new_n6091_ = ~pi260 | ~new_n6036_;
  assign new_n6092_ = ~pi419 | ~new_n6035_;
  assign new_n6093_ = ~pi259 | ~new_n6036_;
  assign new_n6094_ = ~pi418 | ~new_n6035_;
  assign new_n6095_ = ~pi258 | ~new_n6036_;
  assign new_n6096_ = ~pi417 | ~new_n6035_;
  assign new_n6097_ = ~pi249 | ~new_n6036_;
  assign new_n6098_ = ~pi408 | ~new_n6035_;
  assign new_n6099_ = ~pi248 | ~new_n6036_;
  assign new_n6100_ = ~pi407 | ~new_n6035_;
  assign new_n6101_ = ~new_n3122_ | ~new_n3141_;
  assign new_n6102_ = ~new_n1087_ | ~pi238;
  assign new_n6103_ = ~new_n2133_ | ~new_n1906_;
  assign new_n6104_ = ~new_n1087_ | ~pi239;
  assign new_n6105_ = ~new_n2134_ | ~new_n1906_;
  assign new_n6106_ = ~new_n2114_ | ~pi476 | ~new_n1103_;
  assign new_n6107_ = ~new_n1087_ | ~pi240;
  assign new_n6108_ = ~new_n2135_ | ~new_n1906_;
  assign new_n6109_ = ~new_n6357_ | ~new_n1103_ | ~pi476;
  assign new_n6110_ = ~new_n1087_ | ~pi241;
  assign new_n6111_ = ~new_n2136_ | ~new_n1906_;
  assign new_n6112_ = ~new_n1087_ | ~pi242;
  assign new_n6113_ = ~pi073 | ~new_n2830_;
  assign new_n6114_ = pi035 | pi107;
  assign new_n6115_ = ~new_n2755_ | ~new_n5863_;
  assign new_n6116_ = ~new_n5729_ | ~new_n2066_;
  assign new_n6117_ = ~new_n2856_ | ~pi109;
  assign new_n6118_ = ~new_n2857_ | ~pi109;
  assign new_n6119_ = ~new_n2858_ | ~pi109;
  assign new_n6120_ = ~new_n2881_ | ~pi109;
  assign new_n6121_ = ~new_n2909_ | ~pi109;
  assign new_n6122_ = ~pi109 | ~new_n6277_;
  assign new_n6123_ = ~new_n1265_ | ~new_n1910_;
  assign new_n6124_ = ~new_n2765_ | ~new_n2763_ | ~new_n2762_ | ~new_n5738_;
  assign new_n6125_ = ~pi109 | ~new_n6277_;
  assign new_n6126_ = ~new_n1036_ | ~new_n2073_;
  assign new_n6127_ = ~new_n1026_ | ~new_n5012_;
  assign new_n6128_ = ~new_n2533_ | ~new_n1026_;
  assign new_n6129_ = ~new_n6127_ | ~new_n6126_ | ~new_n2874_;
  assign new_n6130_ = ~new_n6128_ | ~new_n2875_;
  assign new_n6131_ = ~new_n2839_ | ~new_n4136_ | ~new_n2816_;
  assign new_n6132_ = ~new_n5736_ | ~new_n2839_;
  assign new_n6133_ = ~new_n2839_ | ~new_n2036_;
  assign new_n6134_ = ~new_n2881_ | ~pi109;
  assign new_n6135_ = ~new_n2717_ | ~new_n6430_ | ~new_n6429_;
  assign new_n6136_ = ~new_n2753_ | ~new_n5861_;
  assign new_n6137_ = ~new_n2754_ | ~new_n5739_;
  assign new_n6138_ = ~new_n1923_;
  assign new_n6139_ = ~new_n1920_;
  assign new_n6140_ = ~new_n2713_ | ~new_n2714_ | ~new_n2715_ | ~new_n2716_ | ~new_n1264_;
  assign new_n6141_ = ~new_n2379_ | ~new_n6138_;
  assign new_n6142_ = ~new_n2380_ | ~new_n4114_;
  assign new_n6143_ = ~new_n1082_ | ~new_n6138_;
  assign new_n6144_ = ~new_n1082_ | ~new_n6138_;
  assign new_n6145_ = ~new_n6144_ | ~new_n5006_ | ~new_n5005_;
  assign new_n6146_ = ~new_n6138_ | ~new_n8624_;
  assign new_n6147_ = ~new_n8624_ | ~new_n6138_ | ~new_n2846_;
  assign new_n6148_ = ~new_n6147_ | ~new_n4794_;
  assign new_n6149_ = ~new_n6138_ | ~new_n5730_;
  assign new_n6150_ = ~new_n6138_ | ~new_n6116_;
  assign new_n6151_ = ~new_n2759_ | ~new_n2761_ | ~new_n2760_;
  assign new_n6152_ = ~new_n2404_ | ~new_n6138_;
  assign new_n6153_ = ~new_n2405_ | ~new_n2406_ | ~new_n4210_;
  assign new_n6154_ = ~new_n2391_ | ~new_n1176_;
  assign new_n6155_ = ~new_n6138_ | ~new_n4607_;
  assign new_n6156_ = ~new_n6138_ | ~new_n4610_;
  assign new_n6157_ = ~new_n6138_ | ~new_n4613_;
  assign new_n6158_ = ~new_n6138_ | ~new_n4616_;
  assign new_n6159_ = ~new_n6138_ | ~new_n4619_;
  assign new_n6160_ = ~new_n6138_ | ~new_n4622_;
  assign new_n6161_ = ~new_n6138_ | ~new_n4625_;
  assign new_n6162_ = ~new_n6138_ | ~new_n4628_;
  assign new_n6163_ = ~new_n6138_ | ~new_n4631_;
  assign new_n6164_ = ~new_n6138_ | ~new_n4634_;
  assign new_n6165_ = ~new_n6138_ | ~new_n4637_;
  assign new_n6166_ = ~new_n6138_ | ~new_n4640_;
  assign new_n6167_ = ~new_n6138_ | ~new_n4643_;
  assign new_n6168_ = ~new_n6138_ | ~new_n4646_;
  assign new_n6169_ = ~new_n6138_ | ~new_n4649_;
  assign new_n6170_ = ~new_n6138_ | ~new_n4652_;
  assign new_n6171_ = ~new_n6138_ | ~new_n4655_;
  assign new_n6172_ = ~new_n6138_ | ~new_n4658_;
  assign new_n6173_ = ~new_n6138_ | ~new_n4661_;
  assign new_n6174_ = ~new_n6138_ | ~new_n4664_;
  assign new_n6175_ = ~new_n6138_ | ~new_n4667_;
  assign new_n6176_ = ~new_n6138_ | ~new_n4670_;
  assign new_n6177_ = ~new_n6138_ | ~new_n4673_;
  assign new_n6178_ = ~new_n6138_ | ~new_n4676_;
  assign new_n6179_ = ~new_n6138_ | ~new_n4679_;
  assign new_n6180_ = ~new_n6138_ | ~new_n4682_;
  assign new_n6181_ = ~new_n6138_ | ~new_n4685_;
  assign new_n6182_ = ~new_n6138_ | ~new_n4688_;
  assign new_n6183_ = ~new_n6138_ | ~new_n4691_;
  assign new_n6184_ = ~new_n6138_ | ~new_n4694_;
  assign new_n6185_ = ~new_n6138_ | ~new_n4697_;
  assign new_n6186_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6187_ = ~pi342 | ~new_n6186_;
  assign new_n6188_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6189_ = ~pi341 | ~new_n6188_;
  assign new_n6190_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6191_ = ~pi340 | ~new_n6190_;
  assign new_n6192_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6193_ = ~pi339 | ~new_n6192_;
  assign new_n6194_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6195_ = ~pi338 | ~new_n6194_;
  assign new_n6196_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6197_ = ~pi337 | ~new_n6196_;
  assign new_n6198_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6199_ = ~pi336 | ~new_n6198_;
  assign new_n6200_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6201_ = ~pi335 | ~new_n6200_;
  assign new_n6202_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6203_ = ~pi334 | ~new_n6202_;
  assign new_n6204_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6205_ = ~pi333 | ~new_n6204_;
  assign new_n6206_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6207_ = ~pi332 | ~new_n6206_;
  assign new_n6208_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6209_ = ~pi331 | ~new_n6208_;
  assign new_n6210_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6211_ = ~pi330 | ~new_n6210_;
  assign new_n6212_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6213_ = ~pi329 | ~new_n6212_;
  assign new_n6214_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6215_ = ~pi328 | ~new_n6214_;
  assign new_n6216_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6217_ = ~pi327 | ~new_n6216_;
  assign new_n6218_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6219_ = ~pi326 | ~new_n6218_;
  assign new_n6220_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6221_ = ~pi325 | ~new_n6220_;
  assign new_n6222_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6223_ = ~pi324 | ~new_n6222_;
  assign new_n6224_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6225_ = ~pi323 | ~new_n6224_;
  assign new_n6226_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6227_ = ~pi322 | ~new_n6226_;
  assign new_n6228_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6229_ = ~pi321 | ~new_n6228_;
  assign new_n6230_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6231_ = ~pi320 | ~new_n6230_;
  assign new_n6232_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6233_ = ~pi319 | ~new_n6232_;
  assign new_n6234_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6235_ = ~pi318 | ~new_n6234_;
  assign new_n6236_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6237_ = ~pi317 | ~new_n6236_;
  assign new_n6238_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6239_ = ~pi316 | ~new_n6238_;
  assign new_n6240_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6241_ = ~pi315 | ~new_n6240_;
  assign new_n6242_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6243_ = ~pi314 | ~new_n6242_;
  assign new_n6244_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6245_ = ~pi313 | ~new_n6244_;
  assign new_n6246_ = ~new_n1014_ | ~new_n6138_;
  assign new_n6247_ = ~pi312 | ~new_n6246_;
  assign new_n6248_ = ~new_n2904_ | ~new_n6138_ | ~new_n2213_;
  assign new_n6249_ = ~new_n2226_ | ~new_n6329_ | ~new_n6328_;
  assign new_n6250_ = ~new_n2512_ | ~new_n6138_;
  assign new_n6251_ = ~new_n6250_ | ~new_n2072_;
  assign new_n6252_ = ~new_n2853_ | ~new_n6138_;
  assign new_n6253_ = ~new_n6252_ | ~new_n2091_;
  assign new_n6254_ = ~new_n1923_ | ~new_n2044_;
  assign new_n6255_ = ~new_n2399_ | ~new_n6138_;
  assign new_n6256_ = ~new_n2400_ | ~new_n6255_;
  assign new_n6257_ = ~pi233 | ~new_n4061_;
  assign new_n6258_ = ~new_n1180_ | ~pi233;
  assign new_n6259_ = ~new_n1203_ | ~pi233;
  assign new_n6260_ = ~new_n2694_ | ~new_n2695_ | ~new_n2697_ | ~new_n2696_;
  assign new_n6261_ = ~new_n2837_ | ~pi233;
  assign new_n6262_ = ~new_n1230_ | ~pi233;
  assign new_n6263_ = ~new_n2732_ | ~new_n2733_ | ~new_n2736_ | ~new_n2734_;
  assign new_n6264_ = ~new_n1249_ | ~pi233;
  assign new_n6265_ = ~new_n2778_ | ~new_n2779_ | ~new_n2781_ | ~new_n2780_;
  assign new_n6266_ = ~new_n1903_;
  assign new_n6267_ = ~new_n6266_ | ~new_n1905_;
  assign new_n6268_ = ~new_n3003_ | ~new_n3006_ | ~pi072;
  assign new_n6269_ = ~pi071 | ~new_n6113_;
  assign new_n6270_ = ~pi072 | ~new_n3003_;
  assign new_n6271_ = ~new_n3147_ | ~new_n3155_;
  assign new_n6272_ = ~new_n4132_ | ~new_n2816_;
  assign new_n6273_ = ~new_n1927_ | ~new_n1933_;
  assign new_n6274_ = ~new_n2036_;
  assign new_n6275_ = ~new_n2853_ | ~new_n6135_;
  assign new_n6276_ = ~new_n4132_ | ~new_n2816_;
  assign new_n6277_ = ~new_n6276_ | ~new_n6275_;
  assign new_n6278_ = ~pi037 | ~new_n1893_;
  assign new_n6279_ = ~pi471 | ~new_n2866_;
  assign new_n6280_ = ~pi038 | ~new_n1893_;
  assign new_n6281_ = ~pi472 | ~new_n2866_;
  assign new_n6282_ = ~pi039 | ~new_n1893_;
  assign new_n6283_ = ~pi473 | ~new_n2866_;
  assign new_n6284_ = ~pi040 | ~new_n1893_;
  assign new_n6285_ = ~pi474 | ~new_n2866_;
  assign new_n6286_ = ~new_n1895_ | ~pi073 | ~pi479;
  assign new_n6287_ = ~pi071 | ~new_n1903_;
  assign new_n6288_ = ~new_n6287_ | ~new_n6286_;
  assign new_n6289_ = ~pi072 | ~new_n6269_ | ~new_n3006_;
  assign new_n6290_ = ~new_n6288_ | ~new_n1892_;
  assign new_n6291_ = ~pi071 | ~pi073 | ~new_n1904_;
  assign new_n6292_ = ~new_n3016_ | ~new_n1895_;
  assign new_n6293_ = pi073 | pi072;
  assign new_n6294_ = ~pi073 | ~new_n2903_;
  assign new_n6295_ = ~new_n2106_;
  assign new_n6296_ = ~new_n6295_ | ~pi074;
  assign new_n6297_ = ~new_n2107_ | ~new_n2106_;
  assign new_n6298_ = ~new_n2106_ | ~new_n3021_;
  assign new_n6299_ = ~new_n6295_ | ~pi075;
  assign new_n6300_ = ~new_n1909_ | ~new_n2186_ | ~new_n2185_;
  assign new_n6301_ = ~pi241 | ~new_n1914_ | ~pi240 | ~pi177 | ~pi242;
  assign new_n6302_ = ~new_n1909_ | ~new_n1914_ | ~pi240 | ~pi193 | ~pi242;
  assign new_n6303_ = ~pi241 | ~new_n1910_ | ~new_n1908_ | ~pi217 | ~new_n1914_;
  assign new_n6304_ = ~new_n1914_ | ~new_n2188_ | ~new_n2187_;
  assign new_n6305_ = ~pi239 | ~new_n2190_ | ~new_n2189_;
  assign new_n6306_ = ~new_n1909_ | ~new_n2192_ | ~new_n2191_;
  assign new_n6307_ = ~pi241 | ~new_n2194_ | ~new_n2193_;
  assign new_n6308_ = ~new_n1910_ | ~new_n2196_ | ~new_n2195_;
  assign new_n6309_ = ~pi242 | ~pi240 | ~pi241 | ~pi113 | ~pi239;
  assign new_n6310_ = ~new_n1914_ | ~new_n1910_ | ~new_n1909_ | ~pi233 | ~new_n1908_;
  assign new_n6311_ = ~pi239 | ~new_n1910_ | ~new_n1909_ | ~pi169 | ~new_n1908_;
  assign new_n6312_ = ~new_n1910_ | ~new_n1908_ | ~pi241 | ~pi153 | ~pi239;
  assign new_n6313_ = ~pi242 | ~new_n2198_ | ~new_n2197_;
  assign new_n6314_ = ~new_n1914_ | ~new_n1908_ | ~pi241 | ~pi209 | ~pi242;
  assign new_n6315_ = ~pi239 | ~new_n1908_ | ~pi241 | ~pi145 | ~pi242;
  assign new_n6316_ = ~new_n1914_ | ~new_n1908_ | ~pi241 | ~pi208 | ~pi242;
  assign new_n6317_ = ~pi239 | ~new_n2174_ | ~new_n2173_;
  assign new_n6318_ = ~new_n1909_ | ~new_n1908_ | ~pi242 | ~pi159 | ~pi239;
  assign new_n6319_ = ~pi241 | ~new_n2180_ | ~new_n2179_;
  assign new_n6320_ = ~new_n1910_ | ~new_n1908_ | ~pi241 | ~pi151 | ~pi239;
  assign new_n6321_ = ~pi242 | ~new_n1908_ | ~pi241 | ~pi143 | ~pi239;
  assign new_n6322_ = ~new_n1914_ | ~new_n1910_ | ~new_n1909_ | ~pi231 | ~new_n1908_;
  assign new_n6323_ = ~pi239 | ~new_n1910_ | ~new_n1909_ | ~pi167 | ~new_n1908_;
  assign new_n6324_ = ~new_n3139_ | ~new_n2081_;
  assign new_n6325_ = ~new_n6146_ | ~new_n1928_;
  assign new_n6326_ = ~new_n2861_ | ~new_n8624_;
  assign new_n6327_ = ~new_n3151_ | ~new_n1917_;
  assign new_n6328_ = ~pi109 | ~new_n3157_;
  assign new_n6329_ = ~new_n3158_ | ~new_n1938_;
  assign new_n6330_ = ~pi106 | ~new_n1939_;
  assign new_n6331_ = ~new_n1085_ | ~new_n3159_;
  assign new_n6332_ = pi478 | pi109;
  assign new_n6333_ = ~pi109 | ~new_n6114_;
  assign new_n6334_ = ~pi109 | ~new_n3167_;
  assign new_n6335_ = ~new_n1938_ | ~new_n6249_ | ~new_n3166_;
  assign new_n6336_ = ~new_n8048_ | ~new_n1957_;
  assign new_n6337_ = ~new_n3173_ | ~new_n1955_;
  assign new_n6338_ = ~new_n2098_;
  assign new_n6339_ = ~pi245 | ~new_n1949_;
  assign new_n6340_ = ~new_n3178_ | ~new_n1948_;
  assign new_n6341_ = ~new_n2099_;
  assign new_n6342_ = ~new_n2861_ | ~new_n1917_;
  assign new_n6343_ = ~new_n8624_ | ~new_n6142_;
  assign new_n6344_ = ~new_n3077_ | ~new_n4111_;
  assign new_n6345_ = ~new_n4112_ | ~new_n2816_;
  assign new_n6346_ = ~new_n2111_ | ~new_n2817_;
  assign new_n6347_ = ~new_n4121_ | ~pi238;
  assign new_n6348_ = ~new_n3105_ | ~new_n1922_;
  assign new_n6349_ = ~new_n3060_ | ~new_n1921_;
  assign new_n6350_ = ~new_n1915_ | ~new_n2059_;
  assign new_n6351_ = ~new_n3122_ | ~new_n4138_;
  assign new_n6352_ = ~new_n6351_ | ~new_n6350_;
  assign new_n6353_ = ~new_n4121_ | ~pi239;
  assign new_n6354_ = ~new_n4154_ | ~new_n2817_;
  assign new_n6355_ = ~pi249 | ~new_n2819_;
  assign new_n6356_ = ~new_n8670_ | ~pi279;
  assign new_n6357_ = ~new_n2114_;
  assign new_n6358_ = ~pi248 | ~new_n2819_;
  assign new_n6359_ = ~pi248 | ~pi279;
  assign new_n6360_ = ~new_n2115_;
  assign new_n6361_ = ~new_n4156_ | ~new_n4146_;
  assign new_n6362_ = ~new_n2863_ | ~new_n2045_;
  assign new_n6363_ = ~pi241 | ~new_n1908_;
  assign new_n6364_ = ~pi240 | ~new_n1909_;
  assign new_n6365_ = ~new_n2100_;
  assign new_n6366_ = ~new_n4121_ | ~pi240;
  assign new_n6367_ = ~new_n4163_ | ~new_n2817_;
  assign new_n6368_ = ~new_n4121_ | ~pi241;
  assign new_n6369_ = ~new_n4174_ | ~new_n2817_;
  assign new_n6370_ = ~new_n2859_ | ~pi242;
  assign new_n6371_ = ~new_n4166_ | ~new_n1910_;
  assign new_n6372_ = ~new_n4121_ | ~pi242;
  assign new_n6373_ = ~new_n4180_ | ~new_n2817_;
  assign new_n6374_ = ~new_n4182_ | ~pi244;
  assign new_n6375_ = ~new_n4190_ | ~new_n2048_;
  assign new_n6376_ = ~new_n6338_ | ~new_n3172_;
  assign new_n6377_ = ~new_n2098_ | ~new_n1958_;
  assign new_n6378_ = ~new_n6377_ | ~new_n6376_;
  assign new_n6379_ = ~new_n4182_ | ~pi245;
  assign new_n6380_ = ~new_n4194_ | ~new_n2048_;
  assign new_n6381_ = ~new_n4182_ | ~pi246;
  assign new_n6382_ = ~new_n4199_ | ~new_n2048_;
  assign new_n6383_ = ~new_n4182_ | ~pi247;
  assign new_n6384_ = ~new_n4202_ | ~new_n2048_;
  assign new_n6385_ = ~new_n3122_ | ~new_n2032_;
  assign new_n6386_ = ~new_n1915_ | ~new_n1925_;
  assign new_n6387_ = ~new_n2816_ | ~new_n1901_ | ~new_n6386_ | ~new_n6385_;
  assign new_n6388_ = ~new_n3077_ | ~new_n8624_ | ~new_n6256_;
  assign new_n6389_ = ~pi406 | ~new_n2068_;
  assign new_n6390_ = ~new_n2123_ | ~new_n2868_;
  assign new_n6391_ = ~pi471 | ~new_n2077_;
  assign new_n6392_ = ~new_n2124_ | ~new_n2865_;
  assign new_n6393_ = pi074 | pi075;
  assign new_n6394_ = ~pi074 | ~new_n2057_;
  assign new_n6395_ = ~new_n6394_ | ~new_n6393_;
  assign new_n6396_ = ~new_n6395_ | ~new_n1897_;
  assign new_n6397_ = ~pi439 | ~pi440;
  assign new_n6398_ = ~new_n6397_ | ~new_n6396_;
  assign new_n6399_ = ~pi472 | ~new_n2077_;
  assign new_n6400_ = ~new_n6398_ | ~new_n2865_;
  assign new_n6401_ = ~pi473 | ~new_n2077_;
  assign new_n6402_ = ~new_n2865_ | ~pi440;
  assign new_n6403_ = ~pi474 | ~new_n2077_;
  assign new_n6404_ = ~new_n2865_ | ~new_n5244_;
  assign new_n6405_ = ~new_n2866_ | ~new_n2080_;
  assign new_n6406_ = ~pi475 | ~new_n1893_;
  assign new_n6407_ = ~pi477 | ~new_n2822_;
  assign new_n6408_ = ~new_n2882_ | ~new_n5245_;
  assign new_n6409_ = ~new_n6295_ | ~pi478;
  assign new_n6410_ = ~pi034 | ~new_n2106_;
  assign new_n6411_ = ~new_n5248_ | ~pi479;
  assign new_n6412_ = ~new_n5254_ | ~new_n2825_;
  assign new_n6413_ = ~new_n2866_ | ~new_n2079_;
  assign new_n6414_ = ~pi480 | ~new_n1893_;
  assign new_n6415_ = ~pi481 | ~new_n1893_;
  assign new_n6416_ = ~pi485 | ~new_n2866_;
  assign new_n6417_ = ~new_n5259_ | ~pi484;
  assign new_n6418_ = ~new_n5260_ | ~new_n2826_;
  assign new_n6419_ = ~new_n2132_ | ~new_n2827_;
  assign new_n6420_ = ~new_n4118_ | ~pi238;
  assign new_n6421_ = ~new_n4118_ | ~pi239;
  assign new_n6422_ = ~new_n4151_ | ~new_n2827_;
  assign new_n6423_ = ~new_n4118_ | ~pi240;
  assign new_n6424_ = ~new_n4159_ | ~new_n2827_;
  assign new_n6425_ = ~new_n4118_ | ~pi241;
  assign new_n6426_ = ~new_n4170_ | ~new_n2827_;
  assign new_n6427_ = ~new_n4118_ | ~pi242;
  assign new_n6428_ = ~new_n4176_ | ~new_n2827_;
  assign new_n6429_ = ~new_n1262_ | ~new_n1921_;
  assign new_n6430_ = ~new_n3105_ | ~new_n6140_;
  assign new_n6431_ = ~new_n2848_ | ~new_n1945_;
  assign new_n6432_ = ~pi247 | ~new_n1941_;
  assign new_n6433_ = ~pi239 | ~new_n2828_;
  assign new_n6434_ = ~new_n5864_ | ~new_n1914_;
  assign new_n6435_ = ~new_n2101_;
  assign new_n6436_ = ~new_n1920_ | ~new_n1928_;
  assign new_n6437_ = ~new_n6352_ | ~new_n3139_;
  assign new_n6438_ = ~new_n2137_ | ~new_n1906_;
  assign new_n6439_ = ~pi108 | ~pi476 | ~new_n6360_;
  assign new_n6440_ = ~new_n9324_ | ~new_n9246_;
  assign new_n6441_ = ~pi260 | ~new_n9245_;
  assign new_n6442_ = ~new_n9325_ | ~new_n9248_;
  assign new_n6443_ = ~pi261 | ~new_n9247_;
  assign new_n6444_ = ~new_n9326_ | ~new_n9250_;
  assign new_n6445_ = ~pi262 | ~new_n9249_;
  assign new_n6446_ = ~new_n9327_ | ~new_n9252_;
  assign new_n6447_ = ~pi263 | ~new_n9251_;
  assign new_n6448_ = ~new_n9328_ | ~new_n9254_;
  assign new_n6449_ = ~pi264 | ~new_n9253_;
  assign new_n6450_ = ~new_n9329_ | ~new_n9256_;
  assign new_n6451_ = ~pi265 | ~new_n9255_;
  assign new_n6452_ = ~new_n9330_ | ~new_n9258_;
  assign new_n6453_ = ~pi266 | ~new_n9257_;
  assign new_n6454_ = ~new_n9331_ | ~new_n9260_;
  assign new_n6455_ = ~pi267 | ~new_n9259_;
  assign new_n6456_ = ~new_n9332_ | ~new_n9262_;
  assign new_n6457_ = ~pi268 | ~new_n9261_;
  assign new_n6458_ = ~new_n9333_ | ~new_n9264_;
  assign new_n6459_ = ~pi269 | ~new_n9263_;
  assign new_n6460_ = ~new_n9334_ | ~new_n9266_;
  assign new_n6461_ = ~pi270 | ~new_n9265_;
  assign new_n6462_ = ~new_n9335_ | ~new_n9268_;
  assign new_n6463_ = ~pi271 | ~new_n9267_;
  assign new_n6464_ = ~new_n9336_ | ~new_n9270_;
  assign new_n6465_ = ~pi272 | ~new_n9269_;
  assign new_n6466_ = ~new_n9337_ | ~new_n9272_;
  assign new_n6467_ = ~pi248;
  assign new_n6468_ = ~pi250;
  assign new_n6469_ = ~pi249;
  assign new_n6470_ = ~pi252;
  assign new_n6471_ = ~pi251;
  assign new_n6472_ = ~pi249 | ~pi250 | ~pi248;
  assign new_n6473_ = ~pi254;
  assign new_n6474_ = ~pi253;
  assign new_n6475_ = ~new_n6544_ | ~new_n6573_;
  assign new_n6476_ = ~pi256;
  assign new_n6477_ = ~pi255;
  assign new_n6478_ = ~new_n6545_ | ~new_n6574_;
  assign new_n6479_ = ~new_n6546_ | ~new_n6580_;
  assign new_n6480_ = ~pi257;
  assign new_n6481_ = ~pi258;
  assign new_n6482_ = ~pi260;
  assign new_n6483_ = ~pi259;
  assign new_n6484_ = ~new_n6547_ | ~new_n6582_;
  assign new_n6485_ = ~pi262;
  assign new_n6486_ = ~pi261;
  assign new_n6487_ = ~new_n6548_ | ~new_n6575_;
  assign new_n6488_ = ~pi263;
  assign new_n6489_ = ~new_n6549_ | ~new_n6581_;
  assign new_n6490_ = ~pi264;
  assign new_n6491_ = ~pi266;
  assign new_n6492_ = ~pi265;
  assign new_n6493_ = ~new_n6550_ | ~new_n6586_;
  assign new_n6494_ = ~pi268;
  assign new_n6495_ = ~pi267;
  assign new_n6496_ = ~new_n6551_ | ~new_n6579_;
  assign new_n6497_ = ~pi269;
  assign new_n6498_ = ~new_n6552_ | ~new_n6576_;
  assign new_n6499_ = ~pi270;
  assign new_n6500_ = ~pi272;
  assign new_n6501_ = ~pi271;
  assign new_n6502_ = ~new_n6553_ | ~new_n6583_;
  assign new_n6503_ = ~pi274;
  assign new_n6504_ = ~pi273;
  assign new_n6505_ = ~new_n6554_ | ~new_n6577_;
  assign new_n6506_ = ~pi275;
  assign new_n6507_ = ~pi276;
  assign new_n6508_ = ~new_n6555_ | ~new_n6578_;
  assign new_n6509_ = ~pi277;
  assign new_n6510_ = ~new_n6556_ | ~new_n6584_;
  assign new_n6511_ = ~new_n6585_ | ~pi277;
  assign new_n6512_ = ~pi278;
  assign new_n6513_ = ~new_n6604_ | ~new_n6603_;
  assign new_n6514_ = ~new_n6606_ | ~new_n6605_;
  assign new_n6515_ = ~new_n6608_ | ~new_n6607_;
  assign new_n6516_ = ~new_n6610_ | ~new_n6609_;
  assign new_n6517_ = ~new_n6612_ | ~new_n6611_;
  assign new_n6518_ = ~new_n6614_ | ~new_n6613_;
  assign new_n6519_ = ~new_n6616_ | ~new_n6615_;
  assign new_n6520_ = ~new_n6618_ | ~new_n6617_;
  assign new_n6521_ = ~new_n6620_ | ~new_n6619_;
  assign new_n6522_ = ~new_n6622_ | ~new_n6621_;
  assign new_n6523_ = ~new_n6624_ | ~new_n6623_;
  assign new_n6524_ = ~new_n6626_ | ~new_n6625_;
  assign new_n6525_ = ~new_n6628_ | ~new_n6627_;
  assign new_n6526_ = ~new_n6630_ | ~new_n6629_;
  assign new_n6527_ = ~new_n6632_ | ~new_n6631_;
  assign new_n6528_ = ~new_n6634_ | ~new_n6633_;
  assign new_n6529_ = ~new_n6636_ | ~new_n6635_;
  assign new_n6530_ = ~new_n6638_ | ~new_n6637_;
  assign new_n6531_ = ~new_n6640_ | ~new_n6639_;
  assign new_n6532_ = ~new_n6642_ | ~new_n6641_;
  assign new_n6533_ = ~new_n6644_ | ~new_n6643_;
  assign new_n6534_ = ~new_n6646_ | ~new_n6645_;
  assign new_n6535_ = ~new_n6648_ | ~new_n6647_;
  assign new_n6536_ = ~new_n6650_ | ~new_n6649_;
  assign new_n6537_ = ~new_n6652_ | ~new_n6651_;
  assign new_n6538_ = ~new_n6654_ | ~new_n6653_;
  assign new_n6539_ = ~new_n6656_ | ~new_n6655_;
  assign new_n6540_ = ~new_n6658_ | ~new_n6657_;
  assign new_n6541_ = ~new_n6660_ | ~new_n6659_;
  assign new_n6542_ = ~new_n6662_ | ~new_n6661_;
  assign new_n6543_ = ~new_n6664_ | ~new_n6663_;
  assign new_n6544_ = pi251 & pi252;
  assign new_n6545_ = pi253 & pi254;
  assign new_n6546_ = pi255 & pi256;
  assign new_n6547_ = pi257 & pi258;
  assign new_n6548_ = pi259 & pi260;
  assign new_n6549_ = pi261 & pi262;
  assign new_n6550_ = pi264 & pi263;
  assign new_n6551_ = pi265 & pi266;
  assign new_n6552_ = pi267 & pi268;
  assign new_n6553_ = pi270 & pi269;
  assign new_n6554_ = pi271 & pi272;
  assign new_n6555_ = pi273 & pi274;
  assign new_n6556_ = pi276 & pi275;
  assign new_n6557_ = ~new_n6580_ | ~pi255;
  assign new_n6558_ = ~new_n6574_ | ~pi253;
  assign new_n6559_ = ~new_n6573_ | ~pi251;
  assign new_n6560_ = ~pi279;
  assign new_n6561_ = ~pi278 | ~new_n6590_;
  assign new_n6562_ = ~pi249 | ~pi248;
  assign new_n6563_ = ~new_n6584_ | ~pi275;
  assign new_n6564_ = ~new_n6578_ | ~pi273;
  assign new_n6565_ = ~new_n6577_ | ~pi271;
  assign new_n6566_ = ~new_n6583_ | ~pi269;
  assign new_n6567_ = ~new_n6576_ | ~pi267;
  assign new_n6568_ = ~new_n6579_ | ~pi265;
  assign new_n6569_ = ~new_n6586_ | ~pi263;
  assign new_n6570_ = ~new_n6581_ | ~pi261;
  assign new_n6571_ = ~new_n6575_ | ~pi259;
  assign new_n6572_ = ~pi257 | ~new_n6582_;
  assign new_n6573_ = ~new_n6472_;
  assign new_n6574_ = ~new_n6475_;
  assign new_n6575_ = ~new_n6484_;
  assign new_n6576_ = ~new_n6496_;
  assign new_n6577_ = ~new_n6502_;
  assign new_n6578_ = ~new_n6505_;
  assign new_n6579_ = ~new_n6493_;
  assign new_n6580_ = ~new_n6478_;
  assign new_n6581_ = ~new_n6487_;
  assign new_n6582_ = ~new_n6479_;
  assign new_n6583_ = ~new_n6498_;
  assign new_n6584_ = ~new_n6508_;
  assign new_n6585_ = ~new_n6510_;
  assign new_n6586_ = ~new_n6489_;
  assign new_n6587_ = ~new_n6557_;
  assign new_n6588_ = ~new_n6558_;
  assign new_n6589_ = ~new_n6559_;
  assign new_n6590_ = ~new_n6511_;
  assign new_n6591_ = ~new_n6561_;
  assign new_n6592_ = ~new_n6562_;
  assign new_n6593_ = ~new_n6563_;
  assign new_n6594_ = ~new_n6564_;
  assign new_n6595_ = ~new_n6565_;
  assign new_n6596_ = ~new_n6566_;
  assign new_n6597_ = ~new_n6567_;
  assign new_n6598_ = ~new_n6568_;
  assign new_n6599_ = ~new_n6569_;
  assign new_n6600_ = ~new_n6570_;
  assign new_n6601_ = ~new_n6571_;
  assign new_n6602_ = ~new_n6572_;
  assign new_n6603_ = ~new_n6582_ | ~new_n6480_;
  assign new_n6604_ = ~pi257 | ~new_n6479_;
  assign new_n6605_ = ~pi256 | ~new_n6557_;
  assign new_n6606_ = ~new_n6587_ | ~new_n6476_;
  assign new_n6607_ = ~new_n6580_ | ~new_n6477_;
  assign new_n6608_ = ~pi255 | ~new_n6478_;
  assign new_n6609_ = ~pi254 | ~new_n6558_;
  assign new_n6610_ = ~new_n6588_ | ~new_n6473_;
  assign new_n6611_ = ~new_n6574_ | ~new_n6474_;
  assign new_n6612_ = ~pi253 | ~new_n6475_;
  assign new_n6613_ = ~pi252 | ~new_n6559_;
  assign new_n6614_ = ~new_n6589_ | ~new_n6470_;
  assign new_n6615_ = ~new_n6573_ | ~new_n6471_;
  assign new_n6616_ = ~pi251 | ~new_n6472_;
  assign new_n6617_ = ~pi279 | ~new_n6561_;
  assign new_n6618_ = ~new_n6591_ | ~new_n6560_;
  assign new_n6619_ = ~pi278 | ~new_n6511_;
  assign new_n6620_ = ~new_n6590_ | ~new_n6512_;
  assign new_n6621_ = ~pi250 | ~new_n6562_;
  assign new_n6622_ = ~new_n6592_ | ~new_n6468_;
  assign new_n6623_ = ~new_n6585_ | ~new_n6509_;
  assign new_n6624_ = ~pi277 | ~new_n6510_;
  assign new_n6625_ = ~pi276 | ~new_n6563_;
  assign new_n6626_ = ~new_n6593_ | ~new_n6507_;
  assign new_n6627_ = ~new_n6584_ | ~new_n6506_;
  assign new_n6628_ = ~pi275 | ~new_n6508_;
  assign new_n6629_ = ~pi274 | ~new_n6564_;
  assign new_n6630_ = ~new_n6594_ | ~new_n6503_;
  assign new_n6631_ = ~new_n6578_ | ~new_n6504_;
  assign new_n6632_ = ~pi273 | ~new_n6505_;
  assign new_n6633_ = ~pi272 | ~new_n6565_;
  assign new_n6634_ = ~new_n6595_ | ~new_n6500_;
  assign new_n6635_ = ~new_n6577_ | ~new_n6501_;
  assign new_n6636_ = ~pi271 | ~new_n6502_;
  assign new_n6637_ = ~pi270 | ~new_n6566_;
  assign new_n6638_ = ~new_n6596_ | ~new_n6499_;
  assign new_n6639_ = ~new_n6583_ | ~new_n6497_;
  assign new_n6640_ = ~pi269 | ~new_n6498_;
  assign new_n6641_ = ~pi268 | ~new_n6567_;
  assign new_n6642_ = ~new_n6597_ | ~new_n6494_;
  assign new_n6643_ = ~pi248 | ~new_n6469_;
  assign new_n6644_ = ~pi249 | ~new_n6467_;
  assign new_n6645_ = ~new_n6576_ | ~new_n6495_;
  assign new_n6646_ = ~pi267 | ~new_n6496_;
  assign new_n6647_ = ~pi266 | ~new_n6568_;
  assign new_n6648_ = ~new_n6598_ | ~new_n6491_;
  assign new_n6649_ = ~new_n6579_ | ~new_n6492_;
  assign new_n6650_ = ~pi265 | ~new_n6493_;
  assign new_n6651_ = ~pi264 | ~new_n6569_;
  assign new_n6652_ = ~new_n6599_ | ~new_n6490_;
  assign new_n6653_ = ~new_n6586_ | ~new_n6488_;
  assign new_n6654_ = ~pi263 | ~new_n6489_;
  assign new_n6655_ = ~pi262 | ~new_n6570_;
  assign new_n6656_ = ~new_n6600_ | ~new_n6485_;
  assign new_n6657_ = ~new_n6581_ | ~new_n6486_;
  assign new_n6658_ = ~pi261 | ~new_n6487_;
  assign new_n6659_ = ~pi260 | ~new_n6571_;
  assign new_n6660_ = ~new_n6601_ | ~new_n6482_;
  assign new_n6661_ = ~new_n6575_ | ~new_n6483_;
  assign new_n6662_ = ~pi259 | ~new_n6484_;
  assign new_n6663_ = ~pi258 | ~new_n6572_;
  assign new_n6664_ = ~new_n6602_ | ~new_n6481_;
  assign new_n6665_ = new_n6877_ & new_n6875_;
  assign new_n6666_ = new_n6887_ & new_n6885_;
  assign new_n6667_ = new_n6666_ & new_n6868_;
  assign new_n6668_ = new_n6667_ & new_n6867_;
  assign new_n6669_ = new_n6895_ & new_n6891_;
  assign new_n6670_ = new_n6669_ & new_n6866_;
  assign new_n6671_ = new_n6670_ & new_n6865_;
  assign new_n6672_ = new_n6671_ & new_n6902_;
  assign new_n6673_ = new_n6672_ & new_n6864_;
  assign new_n6674_ = new_n6910_ & new_n6906_;
  assign new_n6675_ = new_n6674_ & new_n6913_;
  assign new_n6676_ = new_n6675_ & new_n6916_;
  assign new_n6677_ = new_n6952_ & new_n6679_;
  assign new_n6678_ = ~new_n1440_ | ~pi252;
  assign new_n6679_ = ~new_n1444_ | ~pi248;
  assign new_n6680_ = ~new_n1439_ | ~pi253;
  assign new_n6681_ = ~pi278;
  assign new_n6682_ = ~new_n1427_;
  assign new_n6683_ = ~new_n1427_ | ~pi267;
  assign new_n6684_ = ~new_n1428_ | ~pi264;
  assign new_n6685_ = ~new_n6700_ | ~new_n6867_;
  assign new_n6686_ = ~new_n1436_ | ~pi256;
  assign new_n6687_ = ~new_n1435_ | ~pi257;
  assign new_n6688_ = ~new_n1434_ | ~pi258;
  assign new_n6689_ = ~new_n1432_ | ~pi260;
  assign new_n6690_ = ~new_n1430_ | ~pi262;
  assign new_n6691_ = ~new_n1431_ | ~pi261;
  assign new_n6692_ = ~pi277;
  assign new_n6693_ = ~new_n1427_;
  assign new_n6694_ = ~pi276;
  assign new_n6695_ = ~new_n1427_;
  assign new_n6696_ = ~new_n1427_ | ~pi274;
  assign new_n6697_ = ~new_n6988_ | ~new_n6917_;
  assign new_n6698_ = ~new_n6985_ | ~new_n6914_;
  assign new_n6699_ = ~new_n6982_ | ~new_n6911_;
  assign new_n6700_ = ~new_n6966_ | ~new_n6889_;
  assign new_n6701_ = ~new_n6964_ | ~new_n6888_;
  assign new_n6702_ = ~new_n7062_ | ~new_n7061_;
  assign new_n6703_ = new_n6838_ & new_n6822_;
  assign new_n6704_ = new_n6963_ & new_n6839_;
  assign new_n6705_ = new_n6842_ & new_n6823_;
  assign new_n6706_ = new_n6962_ & new_n6961_;
  assign new_n6707_ = pi268 & new_n1427_;
  assign new_n6708_ = new_n6838_ & new_n6822_;
  assign new_n6709_ = new_n6997_ & new_n6839_;
  assign new_n6710_ = new_n6842_ & new_n6961_ & new_n6823_;
  assign new_n6711_ = new_n6849_ & new_n6845_;
  assign new_n6712_ = new_n6665_ & new_n6711_;
  assign new_n6713_ = new_n6846_ & new_n6849_;
  assign new_n6714_ = new_n6955_ & new_n6956_ & new_n6953_ & new_n6876_;
  assign new_n6715_ = new_n6869_ & new_n6881_ & new_n6871_ & new_n6873_;
  assign new_n6716_ = new_n6957_ & new_n6958_ & new_n6954_ & new_n6870_;
  assign new_n6717_ = new_n6673_ & new_n6668_;
  assign new_n6718_ = new_n6992_ & new_n6905_;
  assign new_n6719_ = new_n6718_ & new_n6993_ & new_n6980_;
  assign new_n6720_ = new_n6676_ & new_n6919_;
  assign new_n6721_ = new_n6991_ & new_n6920_;
  assign new_n6722_ = ~new_n7024_ | ~new_n7023_;
  assign new_n6723_ = ~new_n7029_ | ~new_n7028_;
  assign new_n6724_ = ~new_n7036_ | ~new_n7035_;
  assign new_n6725_ = ~new_n7041_ | ~new_n7040_;
  assign new_n6726_ = new_n6685_ & new_n6683_;
  assign new_n6727_ = new_n6978_ & new_n6903_;
  assign new_n6728_ = new_n6975_ & new_n6900_;
  assign new_n6729_ = new_n6972_ & new_n6898_;
  assign new_n6730_ = new_n6970_ & new_n6896_;
  assign new_n6731_ = new_n6955_ & new_n6956_ & new_n6953_ & new_n6876_;
  assign new_n6732_ = ~new_n6686_ | ~new_n6847_;
  assign new_n6733_ = ~new_n6849_ | ~new_n6687_;
  assign new_n6734_ = new_n7010_ & new_n7009_;
  assign new_n6735_ = ~new_n6705_ | ~new_n6706_ | ~new_n6843_;
  assign new_n6736_ = ~new_n6845_ | ~new_n6686_;
  assign new_n6737_ = new_n7012_ & new_n7011_;
  assign new_n6738_ = ~new_n6857_ | ~new_n6825_;
  assign new_n6739_ = ~new_n6822_ | ~new_n6823_;
  assign new_n6740_ = new_n7014_ & new_n7013_;
  assign new_n6741_ = ~new_n6680_ | ~new_n6855_;
  assign new_n6742_ = ~new_n6825_ | ~new_n6824_;
  assign new_n6743_ = new_n7016_ & new_n7015_;
  assign new_n6744_ = ~new_n6678_ | ~new_n6853_;
  assign new_n6745_ = ~new_n6839_ | ~new_n6680_;
  assign new_n6746_ = new_n7018_ & new_n7017_;
  assign new_n6747_ = ~new_n6835_ | ~new_n6836_;
  assign new_n6748_ = ~new_n6838_ | ~new_n6678_;
  assign new_n6749_ = new_n7020_ & new_n7019_;
  assign new_n6750_ = ~new_n6832_ | ~new_n6833_;
  assign new_n6751_ = ~new_n6826_ | ~new_n6835_;
  assign new_n6752_ = new_n7022_ & new_n7021_;
  assign new_n6753_ = ~new_n1426_;
  assign new_n6754_ = ~pi279;
  assign new_n6755_ = ~new_n6721_ | ~new_n6990_;
  assign new_n6756_ = new_n7027_ & new_n7026_;
  assign new_n6757_ = ~new_n6989_ | ~new_n6987_;
  assign new_n6758_ = new_n7032_ & new_n7031_;
  assign new_n6759_ = ~new_n6829_ | ~new_n6830_;
  assign new_n6760_ = ~new_n6827_ | ~new_n6832_;
  assign new_n6761_ = new_n7034_ & new_n7033_;
  assign new_n6762_ = ~new_n6986_ | ~new_n6984_;
  assign new_n6763_ = new_n7039_ & new_n7038_;
  assign new_n6764_ = ~new_n6983_ | ~new_n6981_;
  assign new_n6765_ = new_n7044_ & new_n7043_;
  assign new_n6766_ = ~new_n6696_ | ~new_n6908_;
  assign new_n6767_ = ~new_n6910_ | ~new_n6911_;
  assign new_n6768_ = new_n7046_ & new_n7045_;
  assign new_n6769_ = ~new_n6906_ | ~new_n6696_;
  assign new_n6770_ = ~new_n6719_ | ~new_n7007_;
  assign new_n6771_ = new_n7048_ & new_n7047_;
  assign new_n6772_ = ~new_n6727_ | ~new_n6976_;
  assign new_n6773_ = ~new_n6864_ | ~new_n6905_;
  assign new_n6774_ = new_n7050_ & new_n7049_;
  assign new_n6775_ = ~new_n6728_ | ~new_n6973_;
  assign new_n6776_ = ~new_n6903_ | ~new_n6902_;
  assign new_n6777_ = new_n7052_ & new_n7051_;
  assign new_n6778_ = ~new_n6729_ | ~new_n6971_;
  assign new_n6779_ = ~new_n6900_ | ~new_n6865_;
  assign new_n6780_ = new_n7054_ & new_n7053_;
  assign new_n6781_ = ~new_n6730_ | ~new_n6969_;
  assign new_n6782_ = ~new_n6898_ | ~new_n6866_;
  assign new_n6783_ = new_n7056_ & new_n7055_;
  assign new_n6784_ = ~new_n6892_ | ~new_n6893_;
  assign new_n6785_ = ~new_n6896_ | ~new_n6895_;
  assign new_n6786_ = new_n7058_ & new_n7057_;
  assign new_n6787_ = ~new_n6891_ | ~new_n6892_;
  assign new_n6788_ = ~new_n6726_ | ~new_n7005_;
  assign new_n6789_ = new_n7060_ & new_n7059_;
  assign new_n6790_ = ~new_n6828_ | ~new_n6829_;
  assign new_n6791_ = ~new_n6867_ | ~new_n6683_;
  assign new_n6792_ = ~new_n6967_ | ~new_n7003_;
  assign new_n6793_ = new_n7064_ & new_n7063_;
  assign new_n6794_ = ~new_n6868_ | ~new_n6889_;
  assign new_n6795_ = ~new_n6965_ | ~new_n7001_;
  assign new_n6796_ = new_n7066_ & new_n7065_;
  assign new_n6797_ = ~new_n6887_ | ~new_n6888_;
  assign new_n6798_ = ~new_n6999_ | ~new_n6684_;
  assign new_n6799_ = new_n7068_ & new_n7067_;
  assign new_n6800_ = ~new_n6883_ | ~new_n6716_;
  assign new_n6801_ = ~new_n6885_ | ~new_n6684_;
  assign new_n6802_ = new_n7070_ & new_n7069_;
  assign new_n6803_ = ~new_n6940_ | ~new_n6690_;
  assign new_n6804_ = ~new_n6869_ | ~new_n6870_;
  assign new_n6805_ = new_n7072_ & new_n7071_;
  assign new_n6806_ = ~new_n6691_ | ~new_n6938_;
  assign new_n6807_ = ~new_n6690_ | ~new_n6871_;
  assign new_n6808_ = new_n7074_ & new_n7073_;
  assign new_n6809_ = ~new_n6689_ | ~new_n6936_;
  assign new_n6810_ = ~new_n6873_ | ~new_n6691_;
  assign new_n6811_ = new_n7076_ & new_n7075_;
  assign new_n6812_ = ~new_n6879_ | ~new_n6731_;
  assign new_n6813_ = ~new_n6881_ | ~new_n6689_;
  assign new_n6814_ = new_n7078_ & new_n7077_;
  assign new_n6815_ = ~new_n6948_ | ~new_n6688_;
  assign new_n6816_ = ~new_n6875_ | ~new_n6876_;
  assign new_n6817_ = new_n7080_ & new_n7079_;
  assign new_n6818_ = ~new_n6687_ | ~new_n6946_;
  assign new_n6819_ = ~new_n6688_ | ~new_n6877_;
  assign new_n6820_ = new_n7082_ & new_n7081_;
  assign new_n6821_ = ~new_n6679_;
  assign new_n6822_ = pi255 | new_n1437_;
  assign new_n6823_ = ~new_n1437_ | ~pi255;
  assign new_n6824_ = pi254 | new_n1438_;
  assign new_n6825_ = ~new_n1438_ | ~pi254;
  assign new_n6826_ = pi251 | new_n1441_;
  assign new_n6827_ = pi250 | new_n1442_;
  assign new_n6828_ = pi249 | new_n1443_;
  assign new_n6829_ = ~new_n1443_ | ~pi249;
  assign new_n6830_ = ~new_n6821_ | ~new_n6828_;
  assign new_n6831_ = ~new_n6759_;
  assign new_n6832_ = ~new_n1442_ | ~pi250;
  assign new_n6833_ = ~new_n6759_ | ~new_n6959_;
  assign new_n6834_ = ~new_n6750_;
  assign new_n6835_ = ~new_n1441_ | ~pi251;
  assign new_n6836_ = ~new_n6960_ | ~new_n6826_;
  assign new_n6837_ = ~new_n6747_;
  assign new_n6838_ = pi252 | new_n1440_;
  assign new_n6839_ = pi253 | new_n1439_;
  assign new_n6840_ = ~new_n6680_;
  assign new_n6841_ = ~new_n6678_;
  assign new_n6842_ = ~new_n6822_ | ~new_n6824_ | ~new_n6841_ | ~new_n6839_;
  assign new_n6843_ = ~new_n6704_ | ~new_n6703_ | ~new_n6747_;
  assign new_n6844_ = ~new_n6735_;
  assign new_n6845_ = pi256 | new_n1436_;
  assign new_n6846_ = ~new_n6686_;
  assign new_n6847_ = ~new_n6845_ | ~new_n6735_;
  assign new_n6848_ = ~new_n6732_;
  assign new_n6849_ = pi257 | new_n1435_;
  assign new_n6850_ = ~new_n6687_;
  assign new_n6851_ = ~new_n6733_;
  assign new_n6852_ = ~new_n6736_;
  assign new_n6853_ = ~new_n6838_ | ~new_n6747_;
  assign new_n6854_ = ~new_n6744_;
  assign new_n6855_ = ~new_n6744_ | ~new_n6839_;
  assign new_n6856_ = ~new_n6741_;
  assign new_n6857_ = ~new_n6741_ | ~new_n6824_;
  assign new_n6858_ = ~new_n6738_;
  assign new_n6859_ = ~new_n6739_;
  assign new_n6860_ = ~new_n6742_;
  assign new_n6861_ = ~new_n6745_;
  assign new_n6862_ = ~new_n6748_;
  assign new_n6863_ = ~new_n6751_;
  assign new_n6864_ = pi273 | new_n1427_;
  assign new_n6865_ = pi271 | new_n1427_;
  assign new_n6866_ = pi270 | new_n1427_;
  assign new_n6867_ = pi267 | new_n1427_;
  assign new_n6868_ = pi266 | new_n1427_;
  assign new_n6869_ = pi263 | new_n1429_;
  assign new_n6870_ = ~new_n1429_ | ~pi263;
  assign new_n6871_ = pi262 | new_n1430_;
  assign new_n6872_ = ~new_n6690_;
  assign new_n6873_ = pi261 | new_n1431_;
  assign new_n6874_ = ~new_n6691_;
  assign new_n6875_ = pi259 | new_n1433_;
  assign new_n6876_ = ~new_n1433_ | ~pi259;
  assign new_n6877_ = pi258 | new_n1434_;
  assign new_n6878_ = ~new_n6688_;
  assign new_n6879_ = ~new_n6712_ | ~new_n6995_;
  assign new_n6880_ = ~new_n6812_;
  assign new_n6881_ = pi260 | new_n1432_;
  assign new_n6882_ = ~new_n6689_;
  assign new_n6883_ = ~new_n6715_ | ~new_n6998_;
  assign new_n6884_ = ~new_n6800_;
  assign new_n6885_ = pi264 | new_n1428_;
  assign new_n6886_ = ~new_n6684_;
  assign new_n6887_ = pi265 | new_n1427_;
  assign new_n6888_ = ~new_n1427_ | ~pi265;
  assign new_n6889_ = ~new_n1427_ | ~pi266;
  assign new_n6890_ = ~new_n6683_;
  assign new_n6891_ = pi268 | new_n1427_;
  assign new_n6892_ = ~new_n1427_ | ~pi268;
  assign new_n6893_ = ~new_n6891_ | ~new_n6788_;
  assign new_n6894_ = ~new_n6784_;
  assign new_n6895_ = pi269 | new_n1427_;
  assign new_n6896_ = ~new_n1427_ | ~pi269;
  assign new_n6897_ = ~new_n6781_;
  assign new_n6898_ = ~new_n1427_ | ~pi270;
  assign new_n6899_ = ~new_n6778_;
  assign new_n6900_ = ~new_n1427_ | ~pi271;
  assign new_n6901_ = ~new_n6775_;
  assign new_n6902_ = pi272 | new_n1427_;
  assign new_n6903_ = ~new_n1427_ | ~pi272;
  assign new_n6904_ = ~new_n6772_;
  assign new_n6905_ = ~new_n1427_ | ~pi273;
  assign new_n6906_ = pi274 | new_n1427_;
  assign new_n6907_ = ~new_n6696_;
  assign new_n6908_ = ~new_n6906_ | ~new_n6770_;
  assign new_n6909_ = ~new_n6766_;
  assign new_n6910_ = pi275 | new_n1427_;
  assign new_n6911_ = ~new_n1427_ | ~pi275;
  assign new_n6912_ = ~new_n6764_;
  assign new_n6913_ = pi276 | new_n1427_;
  assign new_n6914_ = ~new_n1427_ | ~pi276;
  assign new_n6915_ = ~new_n6762_;
  assign new_n6916_ = pi277 | new_n1427_;
  assign new_n6917_ = ~new_n1427_ | ~pi277;
  assign new_n6918_ = ~new_n6757_;
  assign new_n6919_ = pi278 | new_n1427_;
  assign new_n6920_ = ~new_n1427_ | ~pi278;
  assign new_n6921_ = ~new_n6755_;
  assign new_n6922_ = ~new_n6760_;
  assign new_n6923_ = ~new_n6767_;
  assign new_n6924_ = ~new_n6769_;
  assign new_n6925_ = ~new_n6773_;
  assign new_n6926_ = ~new_n6776_;
  assign new_n6927_ = ~new_n6779_;
  assign new_n6928_ = ~new_n6782_;
  assign new_n6929_ = ~new_n6785_;
  assign new_n6930_ = ~new_n6787_;
  assign new_n6931_ = ~new_n6790_;
  assign new_n6932_ = ~new_n6791_;
  assign new_n6933_ = ~new_n6794_;
  assign new_n6934_ = ~new_n6797_;
  assign new_n6935_ = ~new_n6801_;
  assign new_n6936_ = ~new_n6881_ | ~new_n6812_;
  assign new_n6937_ = ~new_n6809_;
  assign new_n6938_ = ~new_n6809_ | ~new_n6873_;
  assign new_n6939_ = ~new_n6806_;
  assign new_n6940_ = ~new_n6806_ | ~new_n6871_;
  assign new_n6941_ = ~new_n6803_;
  assign new_n6942_ = ~new_n6804_;
  assign new_n6943_ = ~new_n6807_;
  assign new_n6944_ = ~new_n6810_;
  assign new_n6945_ = ~new_n6813_;
  assign new_n6946_ = ~new_n6849_ | ~new_n6732_;
  assign new_n6947_ = ~new_n6818_;
  assign new_n6948_ = ~new_n6818_ | ~new_n6877_;
  assign new_n6949_ = ~new_n6815_;
  assign new_n6950_ = ~new_n6816_;
  assign new_n6951_ = ~new_n6819_;
  assign new_n6952_ = pi248 | new_n1444_;
  assign new_n6953_ = ~new_n6713_ | ~new_n6665_;
  assign new_n6954_ = ~new_n6869_ | ~new_n6871_ | ~new_n6882_ | ~new_n6873_;
  assign new_n6955_ = ~new_n6850_ | ~new_n6665_;
  assign new_n6956_ = ~new_n6878_ | ~new_n6665_;
  assign new_n6957_ = ~new_n6872_ | ~new_n6869_;
  assign new_n6958_ = ~new_n6869_ | ~new_n6871_ | ~new_n6874_;
  assign new_n6959_ = pi250 | new_n1442_;
  assign new_n6960_ = ~new_n6832_ | ~new_n6833_;
  assign new_n6961_ = ~new_n1438_ | ~pi254 | ~new_n6822_;
  assign new_n6962_ = ~new_n6824_ | ~new_n6840_ | ~new_n6822_;
  assign new_n6963_ = pi254 | new_n1438_;
  assign new_n6964_ = ~new_n6886_ | ~new_n6887_;
  assign new_n6965_ = ~new_n6701_;
  assign new_n6966_ = ~new_n6701_ | ~new_n6868_;
  assign new_n6967_ = ~new_n6700_;
  assign new_n6968_ = ~new_n6685_;
  assign new_n6969_ = ~new_n6669_ | ~new_n6788_;
  assign new_n6970_ = ~new_n6707_ | ~new_n6895_;
  assign new_n6971_ = ~new_n6670_ | ~new_n6788_;
  assign new_n6972_ = ~new_n6994_ | ~new_n6866_;
  assign new_n6973_ = ~new_n6671_ | ~new_n6788_;
  assign new_n6974_ = ~new_n6972_ | ~new_n6898_;
  assign new_n6975_ = ~new_n6974_ | ~new_n6865_;
  assign new_n6976_ = ~new_n6672_ | ~new_n6788_;
  assign new_n6977_ = ~new_n6975_ | ~new_n6900_;
  assign new_n6978_ = ~new_n6977_ | ~new_n6902_;
  assign new_n6979_ = ~new_n6978_ | ~new_n6903_;
  assign new_n6980_ = ~new_n6979_ | ~new_n6864_;
  assign new_n6981_ = ~new_n6674_ | ~new_n6770_;
  assign new_n6982_ = ~new_n6907_ | ~new_n6910_;
  assign new_n6983_ = ~new_n6699_;
  assign new_n6984_ = ~new_n6675_ | ~new_n6770_;
  assign new_n6985_ = ~new_n6699_ | ~new_n6913_;
  assign new_n6986_ = ~new_n6698_;
  assign new_n6987_ = ~new_n6676_ | ~new_n6770_;
  assign new_n6988_ = ~new_n6698_ | ~new_n6916_;
  assign new_n6989_ = ~new_n6697_;
  assign new_n6990_ = ~new_n6720_ | ~new_n6770_;
  assign new_n6991_ = ~new_n6697_ | ~new_n6919_;
  assign new_n6992_ = ~new_n6890_ | ~new_n6673_;
  assign new_n6993_ = ~new_n6968_ | ~new_n6673_;
  assign new_n6994_ = ~new_n6970_ | ~new_n6896_;
  assign new_n6995_ = ~new_n6710_ | ~new_n6996_ | ~new_n6962_;
  assign new_n6996_ = ~new_n6709_ | ~new_n6708_ | ~new_n6747_;
  assign new_n6997_ = pi254 | new_n1438_;
  assign new_n6998_ = ~new_n6879_ | ~new_n6714_;
  assign new_n6999_ = ~new_n6885_ | ~new_n6800_;
  assign new_n7000_ = ~new_n6798_;
  assign new_n7001_ = ~new_n6666_ | ~new_n6800_;
  assign new_n7002_ = ~new_n6795_;
  assign new_n7003_ = ~new_n6667_ | ~new_n6800_;
  assign new_n7004_ = ~new_n6792_;
  assign new_n7005_ = ~new_n6668_ | ~new_n6800_;
  assign new_n7006_ = ~new_n6788_;
  assign new_n7007_ = ~new_n6717_ | ~new_n6800_;
  assign new_n7008_ = ~new_n6770_;
  assign new_n7009_ = ~new_n6848_ | ~new_n6733_;
  assign new_n7010_ = ~new_n6851_ | ~new_n6732_;
  assign new_n7011_ = ~new_n6844_ | ~new_n6736_;
  assign new_n7012_ = ~new_n6852_ | ~new_n6735_;
  assign new_n7013_ = ~new_n6858_ | ~new_n6739_;
  assign new_n7014_ = ~new_n6859_ | ~new_n6738_;
  assign new_n7015_ = ~new_n6856_ | ~new_n6742_;
  assign new_n7016_ = ~new_n6860_ | ~new_n6741_;
  assign new_n7017_ = ~new_n6854_ | ~new_n6745_;
  assign new_n7018_ = ~new_n6861_ | ~new_n6744_;
  assign new_n7019_ = ~new_n6837_ | ~new_n6748_;
  assign new_n7020_ = ~new_n6862_ | ~new_n6747_;
  assign new_n7021_ = ~new_n6834_ | ~new_n6751_;
  assign new_n7022_ = ~new_n6863_ | ~new_n6750_;
  assign new_n7023_ = ~new_n1426_ | ~new_n6754_;
  assign new_n7024_ = ~pi279 | ~new_n6753_;
  assign new_n7025_ = ~new_n6722_;
  assign new_n7026_ = ~new_n6921_ | ~new_n7025_;
  assign new_n7027_ = ~new_n6722_ | ~new_n6755_;
  assign new_n7028_ = ~new_n1427_ | ~new_n6681_;
  assign new_n7029_ = ~pi278 | ~new_n6682_;
  assign new_n7030_ = ~new_n6723_;
  assign new_n7031_ = ~new_n6918_ | ~new_n7030_;
  assign new_n7032_ = ~new_n6723_ | ~new_n6757_;
  assign new_n7033_ = ~new_n6831_ | ~new_n6760_;
  assign new_n7034_ = ~new_n6922_ | ~new_n6759_;
  assign new_n7035_ = ~new_n1427_ | ~new_n6692_;
  assign new_n7036_ = ~pi277 | ~new_n6693_;
  assign new_n7037_ = ~new_n6724_;
  assign new_n7038_ = ~new_n6915_ | ~new_n7037_;
  assign new_n7039_ = ~new_n6724_ | ~new_n6762_;
  assign new_n7040_ = ~new_n1427_ | ~new_n6694_;
  assign new_n7041_ = ~pi276 | ~new_n6695_;
  assign new_n7042_ = ~new_n6725_;
  assign new_n7043_ = ~new_n6912_ | ~new_n7042_;
  assign new_n7044_ = ~new_n6725_ | ~new_n6764_;
  assign new_n7045_ = ~new_n6909_ | ~new_n6767_;
  assign new_n7046_ = ~new_n6923_ | ~new_n6766_;
  assign new_n7047_ = ~new_n6924_ | ~new_n6770_;
  assign new_n7048_ = ~new_n7008_ | ~new_n6769_;
  assign new_n7049_ = ~new_n6904_ | ~new_n6773_;
  assign new_n7050_ = ~new_n6925_ | ~new_n6772_;
  assign new_n7051_ = ~new_n6901_ | ~new_n6776_;
  assign new_n7052_ = ~new_n6926_ | ~new_n6775_;
  assign new_n7053_ = ~new_n6899_ | ~new_n6779_;
  assign new_n7054_ = ~new_n6927_ | ~new_n6778_;
  assign new_n7055_ = ~new_n6897_ | ~new_n6782_;
  assign new_n7056_ = ~new_n6928_ | ~new_n6781_;
  assign new_n7057_ = ~new_n6894_ | ~new_n6785_;
  assign new_n7058_ = ~new_n6929_ | ~new_n6784_;
  assign new_n7059_ = ~new_n6930_ | ~new_n6788_;
  assign new_n7060_ = ~new_n7006_ | ~new_n6787_;
  assign new_n7061_ = ~new_n6821_ | ~new_n6790_;
  assign new_n7062_ = ~new_n6931_ | ~new_n6679_;
  assign new_n7063_ = ~new_n6932_ | ~new_n6792_;
  assign new_n7064_ = ~new_n7004_ | ~new_n6791_;
  assign new_n7065_ = ~new_n6933_ | ~new_n6795_;
  assign new_n7066_ = ~new_n7002_ | ~new_n6794_;
  assign new_n7067_ = ~new_n6934_ | ~new_n6798_;
  assign new_n7068_ = ~new_n7000_ | ~new_n6797_;
  assign new_n7069_ = ~new_n6884_ | ~new_n6801_;
  assign new_n7070_ = ~new_n6935_ | ~new_n6800_;
  assign new_n7071_ = ~new_n6941_ | ~new_n6804_;
  assign new_n7072_ = ~new_n6942_ | ~new_n6803_;
  assign new_n7073_ = ~new_n6939_ | ~new_n6807_;
  assign new_n7074_ = ~new_n6943_ | ~new_n6806_;
  assign new_n7075_ = ~new_n6937_ | ~new_n6810_;
  assign new_n7076_ = ~new_n6944_ | ~new_n6809_;
  assign new_n7077_ = ~new_n6880_ | ~new_n6813_;
  assign new_n7078_ = ~new_n6945_ | ~new_n6812_;
  assign new_n7079_ = ~new_n6949_ | ~new_n6816_;
  assign new_n7080_ = ~new_n6950_ | ~new_n6815_;
  assign new_n7081_ = ~new_n6947_ | ~new_n6819_;
  assign new_n7082_ = ~new_n6951_ | ~new_n6818_;
  assign new_n7083_ = new_n7359_ & new_n7360_ & new_n7371_ & new_n7363_;
  assign new_n7084_ = new_n7407_ & new_n7403_;
  assign new_n7085_ = new_n7219_ & new_n7084_ & new_n7402_;
  assign new_n7086_ = new_n7213_ & new_n7083_;
  assign new_n7087_ = new_n7374_ & new_n7372_;
  assign new_n7088_ = new_n7382_ & new_n7331_;
  assign new_n7089_ = new_n7381_ & new_n7379_;
  assign new_n7090_ = new_n7086_ & new_n7085_;
  assign new_n7091_ = new_n7606_ & new_n7605_;
  assign new_n7092_ = new_n7457_ & new_n7456_;
  assign new_n7093_ = new_n7454_ & new_n7452_;
  assign new_n7094_ = new_n7448_ & new_n7445_;
  assign new_n7095_ = new_n7438_ & new_n7437_;
  assign new_n7096_ = new_n7432_ & new_n7430_;
  assign new_n7097_ = new_n7414_ & new_n7413_;
  assign new_n7098_ = new_n7354_ & new_n7352_;
  assign new_n7099_ = new_n7344_ & new_n7340_;
  assign new_n7100_ = ~new_n1009_;
  assign new_n7101_ = ~new_n1300_;
  assign new_n7102_ = ~new_n1301_;
  assign new_n7103_ = ~new_n1302_;
  assign new_n7104_ = ~new_n1303_;
  assign new_n7105_ = ~new_n1306_;
  assign new_n7106_ = ~new_n1305_;
  assign new_n7107_ = ~new_n1307_;
  assign new_n7108_ = ~new_n1304_;
  assign new_n7109_ = ~new_n1301_ | ~new_n7155_;
  assign new_n7110_ = ~new_n1299_;
  assign new_n7111_ = ~new_n1298_;
  assign new_n7112_ = ~new_n7324_ | ~new_n7337_;
  assign new_n7113_ = ~new_n1277_;
  assign new_n7114_ = ~new_n1282_;
  assign new_n7115_ = ~new_n1281_;
  assign new_n7116_ = ~new_n1279_;
  assign new_n7117_ = ~new_n1280_;
  assign new_n7118_ = ~new_n1278_;
  assign new_n7119_ = ~new_n1283_;
  assign new_n7120_ = ~new_n1284_;
  assign new_n7121_ = ~new_n1285_;
  assign new_n7122_ = ~new_n1286_;
  assign new_n7123_ = ~new_n1287_;
  assign new_n7124_ = ~new_n1287_ | ~new_n7156_;
  assign new_n7125_ = ~new_n1296_;
  assign new_n7126_ = ~new_n1297_;
  assign new_n7127_ = ~new_n1299_ | ~new_n7568_;
  assign new_n7128_ = ~new_n1294_;
  assign new_n7129_ = ~new_n1294_ | ~new_n7158_;
  assign new_n7130_ = ~new_n1295_;
  assign new_n7131_ = ~new_n1295_ | ~new_n7609_;
  assign new_n7132_ = ~new_n1293_;
  assign new_n7133_ = ~new_n7220_ | ~new_n7087_;
  assign new_n7134_ = ~new_n1288_;
  assign new_n7135_ = ~new_n1289_;
  assign new_n7136_ = ~new_n1290_;
  assign new_n7137_ = ~new_n1290_ | ~new_n7685_;
  assign new_n7138_ = ~new_n1291_;
  assign new_n7139_ = ~new_n1291_ | ~new_n7679_;
  assign new_n7140_ = ~new_n7516_ | ~new_n7398_;
  assign new_n7141_ = ~new_n7358_ | ~new_n7369_;
  assign new_n7142_ = ~new_n7311_ | ~new_n7348_;
  assign new_n7143_ = ~new_n7142_ | ~new_n7307_;
  assign new_n7144_ = ~new_n7495_ | ~new_n7394_;
  assign new_n7145_ = ~new_n7224_ | ~new_n7488_ | ~new_n7297_;
  assign new_n7146_ = ~new_n7496_ | ~new_n7494_;
  assign new_n7147_ = ~new_n7486_ | ~new_n7485_ | ~new_n7373_;
  assign new_n7148_ = ~new_n7391_ | ~new_n7145_;
  assign new_n7149_ = ~new_n1292_;
  assign new_n7150_ = ~new_n7129_ | ~new_n7442_;
  assign new_n7151_ = ~new_n7492_ | ~new_n7383_;
  assign new_n7152_ = ~new_n7501_ | ~new_n7491_;
  assign new_n7153_ = ~new_n7152_ | ~new_n7379_;
  assign new_n7154_ = ~new_n7519_ | ~new_n7518_;
  assign new_n7155_ = ~new_n7532_ | ~new_n7531_;
  assign new_n7156_ = ~new_n7630_ | ~new_n7629_;
  assign new_n7157_ = ~new_n7598_ | ~new_n7597_;
  assign new_n7158_ = ~new_n7603_ | ~new_n7602_;
  assign new_n7159_ = ~new_n7611_ | ~new_n7610_;
  assign new_n7160_ = ~new_n7732_ | ~new_n7731_;
  assign new_n7161_ = ~new_n7570_ | ~new_n7569_;
  assign new_n7162_ = new_n7127_ & new_n7331_;
  assign new_n7163_ = ~new_n7572_ | ~new_n7571_;
  assign new_n7164_ = ~new_n7577_ | ~new_n7576_;
  assign new_n7165_ = new_n7324_ & new_n7321_;
  assign new_n7166_ = ~new_n7579_ | ~new_n7578_;
  assign new_n7167_ = new_n7325_ & new_n7322_;
  assign new_n7168_ = ~new_n7581_ | ~new_n7580_;
  assign new_n7169_ = ~new_n7687_ | ~new_n7686_;
  assign new_n7170_ = new_n7356_ & new_n7355_;
  assign new_n7171_ = ~new_n7689_ | ~new_n7688_;
  assign new_n7172_ = new_n7358_ & new_n7357_;
  assign new_n7173_ = ~new_n7691_ | ~new_n7690_;
  assign new_n7174_ = new_n7366_ & new_n7359_;
  assign new_n7175_ = ~new_n7693_ | ~new_n7692_;
  assign new_n7176_ = new_n7367_ & new_n7360_;
  assign new_n7177_ = ~new_n7695_ | ~new_n7694_;
  assign new_n7178_ = new_n7363_ & new_n7362_;
  assign new_n7179_ = ~new_n7697_ | ~new_n7696_;
  assign new_n7180_ = new_n7371_ & new_n7361_;
  assign new_n7181_ = ~new_n7699_ | ~new_n7698_;
  assign new_n7182_ = new_n7398_ & new_n7397_;
  assign new_n7183_ = ~new_n7701_ | ~new_n7700_;
  assign new_n7184_ = new_n7400_ & new_n7399_;
  assign new_n7185_ = ~new_n7703_ | ~new_n7702_;
  assign new_n7186_ = new_n7402_ & new_n7401_;
  assign new_n7187_ = ~new_n7705_ | ~new_n7704_;
  assign new_n7188_ = ~new_n7710_ | ~new_n7709_;
  assign new_n7189_ = new_n7311_ & new_n7310_;
  assign new_n7190_ = ~new_n7712_ | ~new_n7711_;
  assign new_n7191_ = new_n7395_ & new_n7394_;
  assign new_n7192_ = ~new_n7714_ | ~new_n7713_;
  assign new_n7193_ = new_n7373_ & new_n7372_;
  assign new_n7194_ = ~new_n7716_ | ~new_n7715_;
  assign new_n7195_ = new_n7137_ & new_n7374_;
  assign new_n7196_ = ~new_n7718_ | ~new_n7717_;
  assign new_n7197_ = ~new_n7723_ | ~new_n7722_;
  assign new_n7198_ = ~new_n7728_ | ~new_n7727_;
  assign new_n7199_ = new_n7388_ & new_n7131_;
  assign new_n7200_ = ~new_n7730_ | ~new_n7729_;
  assign new_n7201_ = new_n7313_ & new_n7310_;
  assign new_n7202_ = new_n7309_ & new_n7307_;
  assign new_n7203_ = new_n7322_ & new_n7321_;
  assign new_n7204_ = new_n7327_ & new_n7323_;
  assign new_n7205_ = new_n7323_ & new_n7300_;
  assign new_n7206_ = new_n7343_ & new_n7109_;
  assign new_n7207_ = new_n7309_ & new_n7308_;
  assign new_n7208_ = new_n7363_ & new_n7360_;
  assign new_n7209_ = new_n7366_ & new_n7367_;
  assign new_n7210_ = new_n7359_ & new_n7357_;
  assign new_n7211_ = new_n7404_ & new_n7401_;
  assign new_n7212_ = new_n7400_ & new_n7397_;
  assign new_n7213_ = new_n7357_ & new_n7355_;
  assign new_n7214_ = new_n7089_ & new_n7088_;
  assign new_n7215_ = new_n7510_ & new_n7503_;
  assign new_n7216_ = new_n7388_ & new_n7302_;
  assign new_n7217_ = new_n7493_ & new_n7389_;
  assign new_n7218_ = new_n7498_ & new_n7489_;
  assign new_n7219_ = new_n7400_ & new_n7397_;
  assign new_n7220_ = new_n7395_ & new_n7391_;
  assign new_n7221_ = new_n7090_ & new_n7504_;
  assign new_n7222_ = new_n7480_ & new_n7356_;
  assign new_n7223_ = new_n7508_ & new_n7222_ & new_n7484_;
  assign new_n7224_ = new_n7498_ & new_n7489_;
  assign new_n7225_ = new_n7391_ & new_n7395_;
  assign new_n7226_ = new_n7085_ & new_n7227_;
  assign new_n7227_ = new_n7087_ & new_n7225_;
  assign new_n7228_ = new_n7500_ & new_n7517_;
  assign new_n7229_ = new_n7083_ & new_n7357_;
  assign new_n7230_ = new_n7371_ & new_n7363_ & new_n7360_;
  assign new_n7231_ = new_n7367_ & new_n7365_;
  assign new_n7232_ = new_n7362_ & new_n7361_;
  assign new_n7233_ = new_n7234_ & new_n7512_;
  assign new_n7234_ = new_n7084_ & new_n7402_;
  assign new_n7235_ = new_n7496_ & new_n7124_;
  assign new_n7236_ = new_n7084_ & new_n7404_;
  assign new_n7237_ = new_n7391_ & new_n7087_;
  assign new_n7238_ = new_n7378_ & new_n7377_ & new_n7302_;
  assign new_n7239_ = new_n7447_ & new_n7305_;
  assign new_n7240_ = new_n7381_ & new_n7380_;
  assign new_n7241_ = new_n7453_ & new_n7385_;
  assign new_n7242_ = ~new_n1269_;
  assign new_n7243_ = new_n7522_ & new_n7521_;
  assign new_n7244_ = ~new_n1267_;
  assign new_n7245_ = ~new_n1266_;
  assign new_n7246_ = ~new_n1324_;
  assign new_n7247_ = ~new_n1325_;
  assign new_n7248_ = ~new_n1327_;
  assign new_n7249_ = ~new_n1328_;
  assign new_n7250_ = ~new_n1329_;
  assign new_n7251_ = ~new_n1326_;
  assign new_n7252_ = ~new_n1268_;
  assign new_n7253_ = ~new_n7127_ | ~new_n7333_;
  assign new_n7254_ = ~new_n7204_ | ~new_n7329_ | ~new_n7328_;
  assign new_n7255_ = ~new_n7325_ | ~new_n7335_;
  assign new_n7256_ = ~new_n7308_ | ~new_n7318_;
  assign new_n7257_ = ~new_n1308_;
  assign new_n7258_ = new_n7583_ & new_n7582_;
  assign new_n7259_ = ~new_n1270_;
  assign new_n7260_ = ~new_n1271_;
  assign new_n7261_ = ~new_n1274_;
  assign new_n7262_ = ~new_n1272_;
  assign new_n7263_ = ~new_n1273_;
  assign new_n7264_ = ~new_n1275_;
  assign new_n7265_ = ~new_n1321_;
  assign new_n7266_ = ~new_n1322_;
  assign new_n7267_ = ~new_n1323_;
  assign new_n7268_ = ~new_n1320_;
  assign new_n7269_ = ~new_n1315_;
  assign new_n7270_ = ~new_n1316_;
  assign new_n7271_ = ~new_n1317_;
  assign new_n7272_ = ~new_n1318_;
  assign new_n7273_ = ~new_n1319_;
  assign new_n7274_ = ~new_n1311_;
  assign new_n7275_ = ~new_n1312_;
  assign new_n7276_ = ~new_n1313_;
  assign new_n7277_ = ~new_n1314_;
  assign new_n7278_ = ~new_n1309_;
  assign new_n7279_ = ~new_n1310_;
  assign new_n7280_ = ~new_n7223_ | ~new_n7507_;
  assign new_n7281_ = ~new_n7370_ | ~new_n7410_;
  assign new_n7282_ = ~new_n7416_ | ~new_n7415_;
  assign new_n7283_ = ~new_n7231_ | ~new_n7418_;
  assign new_n7284_ = ~new_n7422_ | ~new_n7363_;
  assign new_n7285_ = ~new_n7361_ | ~new_n7420_;
  assign new_n7286_ = ~new_n7228_ | ~new_n7499_;
  assign new_n7287_ = ~new_n7399_ | ~new_n7425_;
  assign new_n7288_ = ~new_n7423_ | ~new_n7515_;
  assign new_n7289_ = ~new_n7428_ | ~new_n7403_;
  assign new_n7290_ = ~new_n7314_ | ~new_n7346_;
  assign new_n7291_ = ~new_n7490_ | ~new_n7487_;
  assign new_n7292_ = ~new_n7434_ | ~new_n7137_;
  assign new_n7293_ = ~new_n7139_ | ~new_n7148_;
  assign new_n7294_ = ~new_n7131_ | ~new_n7439_;
  assign new_n7295_ = ~new_n7215_ | ~new_n7509_;
  assign new_n7296_ = ~new_n7314_ | ~new_n7313_;
  assign new_n7297_ = ~new_n7217_ | ~new_n7216_ | ~new_n7295_;
  assign new_n7298_ = ~new_n7289_;
  assign new_n7299_ = ~new_n7284_;
  assign new_n7300_ = ~new_n7482_ | ~new_n7481_;
  assign new_n7301_ = ~new_n7129_;
  assign new_n7302_ = ~new_n7599_ | ~new_n7132_;
  assign new_n7303_ = ~new_n7124_;
  assign new_n7304_ = ~new_n7427_ | ~new_n7407_;
  assign new_n7305_ = ~new_n1293_ | ~new_n7157_;
  assign new_n7306_ = ~new_n7109_;
  assign new_n7307_ = ~new_n7106_ | ~new_n7558_ | ~new_n7557_;
  assign new_n7308_ = ~new_n1304_ | ~new_n7563_;
  assign new_n7309_ = ~new_n7108_ | ~new_n7560_ | ~new_n7559_;
  assign new_n7310_ = ~new_n7105_ | ~new_n7554_ | ~new_n7553_;
  assign new_n7311_ = ~new_n1306_ | ~new_n7549_;
  assign new_n7312_ = ~new_n1305_ | ~new_n7546_;
  assign new_n7313_ = ~new_n7107_ | ~new_n7556_ | ~new_n7555_;
  assign new_n7314_ = ~new_n1307_ | ~new_n7552_;
  assign new_n7315_ = ~new_n7314_ | ~new_n7100_;
  assign new_n7316_ = ~new_n7201_ | ~new_n7315_;
  assign new_n7317_ = ~new_n7312_ | ~new_n7316_ | ~new_n7311_;
  assign new_n7318_ = ~new_n7202_ | ~new_n7317_;
  assign new_n7319_ = ~new_n7256_;
  assign new_n7320_ = ~new_n7101_ | ~new_n7530_ | ~new_n7529_;
  assign new_n7321_ = ~new_n7103_ | ~new_n7541_ | ~new_n7540_;
  assign new_n7322_ = ~new_n7104_ | ~new_n7543_ | ~new_n7542_;
  assign new_n7323_ = ~new_n1300_ | ~new_n7528_;
  assign new_n7324_ = ~new_n1302_ | ~new_n7536_;
  assign new_n7325_ = ~new_n1303_ | ~new_n7539_;
  assign new_n7326_ = ~new_n7325_ | ~new_n7324_;
  assign new_n7327_ = ~new_n7300_ | ~new_n7321_ | ~new_n7326_;
  assign new_n7328_ = ~new_n7300_ | ~new_n7256_ | ~new_n7203_;
  assign new_n7329_ = ~new_n7306_ | ~new_n7320_;
  assign new_n7330_ = ~new_n7254_;
  assign new_n7331_ = ~new_n7110_ | ~new_n7565_ | ~new_n7564_;
  assign new_n7332_ = ~new_n7127_;
  assign new_n7333_ = ~new_n7331_ | ~new_n7254_;
  assign new_n7334_ = ~new_n7253_;
  assign new_n7335_ = ~new_n7322_ | ~new_n7256_;
  assign new_n7336_ = ~new_n7255_;
  assign new_n7337_ = ~new_n7255_ | ~new_n7321_;
  assign new_n7338_ = ~new_n7112_;
  assign new_n7339_ = ~new_n7338_ | ~new_n7109_;
  assign new_n7340_ = ~new_n7205_ | ~new_n7339_;
  assign new_n7341_ = ~new_n7533_ | ~new_n7102_;
  assign new_n7342_ = ~new_n7341_ | ~new_n7112_;
  assign new_n7343_ = ~new_n7323_ | ~new_n7320_;
  assign new_n7344_ = ~new_n7206_ | ~new_n7342_;
  assign new_n7345_ = ~new_n7533_ | ~new_n7102_;
  assign new_n7346_ = ~new_n1009_ | ~new_n7313_;
  assign new_n7347_ = ~new_n7290_;
  assign new_n7348_ = ~new_n7290_ | ~new_n7310_;
  assign new_n7349_ = ~new_n7142_;
  assign new_n7350_ = ~new_n7143_;
  assign new_n7351_ = ~new_n7143_ | ~new_n7312_;
  assign new_n7352_ = ~new_n7207_ | ~new_n7351_;
  assign new_n7353_ = ~new_n7309_ | ~new_n7308_;
  assign new_n7354_ = ~new_n7353_ | ~new_n7143_ | ~new_n7312_;
  assign new_n7355_ = ~new_n7113_ | ~new_n7641_ | ~new_n7640_;
  assign new_n7356_ = ~new_n1277_ | ~new_n7658_;
  assign new_n7357_ = ~new_n7118_ | ~new_n7643_ | ~new_n7642_;
  assign new_n7358_ = ~new_n1278_ | ~new_n7673_;
  assign new_n7359_ = ~new_n7116_ | ~new_n7633_ | ~new_n7632_;
  assign new_n7360_ = ~new_n7117_ | ~new_n7635_ | ~new_n7634_;
  assign new_n7361_ = ~new_n1282_ | ~new_n7661_;
  assign new_n7362_ = ~new_n1281_ | ~new_n7664_;
  assign new_n7363_ = ~new_n7115_ | ~new_n7637_ | ~new_n7636_;
  assign new_n7364_ = ~new_n7362_ | ~new_n7361_;
  assign new_n7365_ = ~new_n7208_ | ~new_n7364_;
  assign new_n7366_ = ~new_n1279_ | ~new_n7670_;
  assign new_n7367_ = ~new_n1280_ | ~new_n7667_;
  assign new_n7368_ = ~new_n7209_ | ~new_n7365_;
  assign new_n7369_ = ~new_n7210_ | ~new_n7368_;
  assign new_n7370_ = ~new_n7141_;
  assign new_n7371_ = ~new_n7114_ | ~new_n7639_ | ~new_n7638_;
  assign new_n7372_ = ~new_n7135_ | ~new_n7614_ | ~new_n7613_;
  assign new_n7373_ = ~new_n1289_ | ~new_n7682_;
  assign new_n7374_ = ~new_n7136_ | ~new_n7616_ | ~new_n7615_;
  assign new_n7375_ = ~new_n7137_;
  assign new_n7376_ = ~new_n7139_;
  assign new_n7377_ = ~new_n7091_ | ~new_n7149_;
  assign new_n7378_ = ~new_n1292_ | ~new_n7159_;
  assign new_n7379_ = ~new_n7126_ | ~new_n7588_ | ~new_n7587_;
  assign new_n7380_ = ~new_n1296_ | ~new_n7593_;
  assign new_n7381_ = ~new_n7125_ | ~new_n7590_ | ~new_n7589_;
  assign new_n7382_ = ~new_n7520_ | ~new_n7111_;
  assign new_n7383_ = ~new_n1298_ | ~new_n7154_;
  assign new_n7384_ = ~new_n7152_;
  assign new_n7385_ = ~new_n1297_ | ~new_n7596_;
  assign new_n7386_ = ~new_n7295_;
  assign new_n7387_ = ~new_n7131_;
  assign new_n7388_ = ~new_n7130_ | ~new_n7601_ | ~new_n7600_;
  assign new_n7389_ = ~new_n7604_ | ~new_n7128_;
  assign new_n7390_ = ~new_n7145_;
  assign new_n7391_ = ~new_n7138_ | ~new_n7618_ | ~new_n7617_;
  assign new_n7392_ = ~new_n7148_;
  assign new_n7393_ = ~new_n7291_;
  assign new_n7394_ = ~new_n1288_ | ~new_n7676_;
  assign new_n7395_ = ~new_n7134_ | ~new_n7620_ | ~new_n7619_;
  assign new_n7396_ = ~new_n7146_;
  assign new_n7397_ = ~new_n7119_ | ~new_n7622_ | ~new_n7621_;
  assign new_n7398_ = ~new_n1283_ | ~new_n7646_;
  assign new_n7399_ = ~new_n1284_ | ~new_n7649_;
  assign new_n7400_ = ~new_n7120_ | ~new_n7624_ | ~new_n7623_;
  assign new_n7401_ = ~new_n1285_ | ~new_n7652_;
  assign new_n7402_ = ~new_n7121_ | ~new_n7626_ | ~new_n7625_;
  assign new_n7403_ = ~new_n7122_ | ~new_n7628_ | ~new_n7627_;
  assign new_n7404_ = ~new_n1286_ | ~new_n7655_;
  assign new_n7405_ = ~new_n7303_ | ~new_n7403_;
  assign new_n7406_ = ~new_n7515_ | ~new_n7399_;
  assign new_n7407_ = ~new_n7631_ | ~new_n7123_;
  assign new_n7408_ = ~new_n7280_;
  assign new_n7409_ = ~new_n7286_;
  assign new_n7410_ = ~new_n7229_ | ~new_n7286_;
  assign new_n7411_ = ~new_n7281_;
  assign new_n7412_ = ~new_n7312_ | ~new_n7307_;
  assign new_n7413_ = ~new_n7349_ | ~new_n7412_;
  assign new_n7414_ = ~new_n7350_ | ~new_n7312_;
  assign new_n7415_ = ~new_n7368_ | ~new_n7359_;
  assign new_n7416_ = ~new_n7083_ | ~new_n7286_;
  assign new_n7417_ = ~new_n7282_;
  assign new_n7418_ = ~new_n7230_ | ~new_n7286_;
  assign new_n7419_ = ~new_n7283_;
  assign new_n7420_ = ~new_n7286_ | ~new_n7371_;
  assign new_n7421_ = ~new_n7285_;
  assign new_n7422_ = ~new_n7232_ | ~new_n7420_;
  assign new_n7423_ = ~new_n7511_ | ~new_n7233_;
  assign new_n7424_ = ~new_n7288_;
  assign new_n7425_ = ~new_n7288_ | ~new_n7400_;
  assign new_n7426_ = ~new_n7287_;
  assign new_n7427_ = ~new_n7235_ | ~new_n7494_;
  assign new_n7428_ = ~new_n7404_ | ~new_n7304_;
  assign new_n7429_ = ~new_n7396_ | ~new_n7124_;
  assign new_n7430_ = ~new_n7236_ | ~new_n7429_;
  assign new_n7431_ = ~new_n7404_ | ~new_n7403_;
  assign new_n7432_ = ~new_n7304_ | ~new_n7431_;
  assign new_n7433_ = ~new_n7293_;
  assign new_n7434_ = ~new_n7293_ | ~new_n7374_;
  assign new_n7435_ = ~new_n7292_;
  assign new_n7436_ = ~new_n7391_ | ~new_n7139_;
  assign new_n7437_ = ~new_n7390_ | ~new_n7436_;
  assign new_n7438_ = ~new_n7392_ | ~new_n7139_;
  assign new_n7439_ = ~new_n7388_ | ~new_n7295_;
  assign new_n7440_ = ~new_n7294_;
  assign new_n7441_ = ~new_n7604_ | ~new_n7128_;
  assign new_n7442_ = ~new_n7441_ | ~new_n7294_;
  assign new_n7443_ = ~new_n7150_;
  assign new_n7444_ = ~new_n7443_ | ~new_n7305_;
  assign new_n7445_ = ~new_n7238_ | ~new_n7444_;
  assign new_n7446_ = ~new_n7150_ | ~new_n7302_;
  assign new_n7447_ = ~new_n7378_ | ~new_n7377_;
  assign new_n7448_ = ~new_n7239_ | ~new_n7446_;
  assign new_n7449_ = ~new_n7604_ | ~new_n7128_;
  assign new_n7450_ = ~new_n7153_;
  assign new_n7451_ = ~new_n7153_ | ~new_n7385_;
  assign new_n7452_ = ~new_n7240_ | ~new_n7451_;
  assign new_n7453_ = ~new_n7381_ | ~new_n7380_;
  assign new_n7454_ = ~new_n7241_ | ~new_n7153_;
  assign new_n7455_ = ~new_n7385_ | ~new_n7379_;
  assign new_n7456_ = ~new_n7384_ | ~new_n7455_;
  assign new_n7457_ = ~new_n7450_ | ~new_n7385_;
  assign new_n7458_ = ~new_n7296_;
  assign new_n7459_ = ~new_n7127_ | ~new_n7331_;
  assign new_n7460_ = ~new_n7345_ | ~new_n7109_;
  assign new_n7461_ = ~new_n7324_ | ~new_n7321_;
  assign new_n7462_ = ~new_n7325_ | ~new_n7322_;
  assign new_n7463_ = ~new_n7356_ | ~new_n7355_;
  assign new_n7464_ = ~new_n7358_ | ~new_n7357_;
  assign new_n7465_ = ~new_n7366_ | ~new_n7359_;
  assign new_n7466_ = ~new_n7367_ | ~new_n7360_;
  assign new_n7467_ = ~new_n7363_ | ~new_n7362_;
  assign new_n7468_ = ~new_n7371_ | ~new_n7361_;
  assign new_n7469_ = ~new_n7398_ | ~new_n7397_;
  assign new_n7470_ = ~new_n7400_ | ~new_n7399_;
  assign new_n7471_ = ~new_n7402_ | ~new_n7401_;
  assign new_n7472_ = ~new_n7407_ | ~new_n7124_;
  assign new_n7473_ = ~new_n7311_ | ~new_n7310_;
  assign new_n7474_ = ~new_n7395_ | ~new_n7394_;
  assign new_n7475_ = ~new_n7373_ | ~new_n7372_;
  assign new_n7476_ = ~new_n7137_ | ~new_n7374_;
  assign new_n7477_ = ~new_n7305_ | ~new_n7302_;
  assign new_n7478_ = ~new_n7449_ | ~new_n7129_;
  assign new_n7479_ = ~new_n7388_ | ~new_n7131_;
  assign new_n7480_ = ~new_n7141_ | ~new_n7355_;
  assign new_n7481_ = ~new_n7155_ | ~new_n7320_;
  assign new_n7482_ = ~new_n1301_ | ~new_n7320_;
  assign new_n7483_ = ~new_n1297_ | ~new_n7596_;
  assign new_n7484_ = ~new_n7086_ | ~new_n7140_;
  assign new_n7485_ = ~new_n7375_ | ~new_n7087_;
  assign new_n7486_ = ~new_n7376_ | ~new_n7087_;
  assign new_n7487_ = ~new_n7237_ | ~new_n7145_;
  assign new_n7488_ = ~new_n7377_ | ~new_n7301_ | ~new_n7302_;
  assign new_n7489_ = ~new_n7377_ | ~new_n7302_ | ~new_n7387_ | ~new_n7389_;
  assign new_n7490_ = ~new_n7147_;
  assign new_n7491_ = ~new_n7088_ | ~new_n7254_;
  assign new_n7492_ = ~new_n7332_ | ~new_n7382_;
  assign new_n7493_ = ~new_n7091_ | ~new_n7149_;
  assign new_n7494_ = ~new_n7504_ | ~new_n7145_;
  assign new_n7495_ = ~new_n7147_ | ~new_n7395_;
  assign new_n7496_ = ~new_n7144_;
  assign new_n7497_ = ~new_n7091_ | ~new_n7149_;
  assign new_n7498_ = ~new_n7506_ | ~new_n7505_ | ~new_n7497_;
  assign new_n7499_ = ~new_n7145_ | ~new_n7226_;
  assign new_n7500_ = ~new_n7144_ | ~new_n7085_;
  assign new_n7501_ = ~new_n7151_;
  assign new_n7502_ = ~new_n7483_ | ~new_n7380_;
  assign new_n7503_ = ~new_n7502_ | ~new_n7381_;
  assign new_n7504_ = ~new_n7133_;
  assign new_n7505_ = ~new_n7305_ | ~new_n7149_;
  assign new_n7506_ = ~new_n7612_ | ~new_n7305_;
  assign new_n7507_ = ~new_n7221_ | ~new_n7513_;
  assign new_n7508_ = ~new_n7090_ | ~new_n7144_;
  assign new_n7509_ = ~new_n7214_ | ~new_n7254_;
  assign new_n7510_ = ~new_n7089_ | ~new_n7151_;
  assign new_n7511_ = ~new_n7390_ | ~new_n7496_;
  assign new_n7512_ = ~new_n7496_ | ~new_n7133_;
  assign new_n7513_ = ~new_n7218_ | ~new_n7488_ | ~new_n7297_;
  assign new_n7514_ = ~new_n7211_ | ~new_n7405_;
  assign new_n7515_ = ~new_n7514_ | ~new_n7402_;
  assign new_n7516_ = ~new_n7212_ | ~new_n7406_;
  assign new_n7517_ = ~new_n7140_;
  assign new_n7518_ = ~new_n1009_ | ~new_n7242_;
  assign new_n7519_ = ~new_n1269_ | ~new_n7100_;
  assign new_n7520_ = ~new_n7154_;
  assign new_n7521_ = ~new_n7520_ | ~new_n1298_;
  assign new_n7522_ = ~new_n7154_ | ~new_n7111_;
  assign new_n7523_ = ~new_n7520_ | ~new_n1298_;
  assign new_n7524_ = ~new_n7154_ | ~new_n7111_;
  assign new_n7525_ = ~new_n7524_ | ~new_n7523_;
  assign new_n7526_ = ~new_n1009_ | ~new_n7244_;
  assign new_n7527_ = ~new_n1267_ | ~new_n7100_;
  assign new_n7528_ = ~new_n7527_ | ~new_n7526_;
  assign new_n7529_ = ~new_n1009_ | ~new_n7244_;
  assign new_n7530_ = ~new_n1267_ | ~new_n7100_;
  assign new_n7531_ = ~new_n1009_ | ~new_n7245_;
  assign new_n7532_ = ~new_n1266_ | ~new_n7100_;
  assign new_n7533_ = ~new_n7155_;
  assign new_n7534_ = ~new_n1009_ | ~new_n7246_;
  assign new_n7535_ = ~new_n1324_ | ~new_n7100_;
  assign new_n7536_ = ~new_n7535_ | ~new_n7534_;
  assign new_n7537_ = ~new_n1009_ | ~new_n7247_;
  assign new_n7538_ = ~new_n1325_ | ~new_n7100_;
  assign new_n7539_ = ~new_n7538_ | ~new_n7537_;
  assign new_n7540_ = ~new_n1009_ | ~new_n7246_;
  assign new_n7541_ = ~new_n1324_ | ~new_n7100_;
  assign new_n7542_ = ~new_n1009_ | ~new_n7247_;
  assign new_n7543_ = ~new_n1325_ | ~new_n7100_;
  assign new_n7544_ = ~new_n1009_ | ~new_n7248_;
  assign new_n7545_ = ~new_n1327_ | ~new_n7100_;
  assign new_n7546_ = ~new_n7545_ | ~new_n7544_;
  assign new_n7547_ = ~new_n1009_ | ~new_n7249_;
  assign new_n7548_ = ~new_n1328_ | ~new_n7100_;
  assign new_n7549_ = ~new_n7548_ | ~new_n7547_;
  assign new_n7550_ = ~new_n1009_ | ~new_n7250_;
  assign new_n7551_ = ~new_n1329_ | ~new_n7100_;
  assign new_n7552_ = ~new_n7551_ | ~new_n7550_;
  assign new_n7553_ = ~new_n1009_ | ~new_n7249_;
  assign new_n7554_ = ~new_n1328_ | ~new_n7100_;
  assign new_n7555_ = ~new_n1009_ | ~new_n7250_;
  assign new_n7556_ = ~new_n1329_ | ~new_n7100_;
  assign new_n7557_ = ~new_n1009_ | ~new_n7248_;
  assign new_n7558_ = ~new_n1327_ | ~new_n7100_;
  assign new_n7559_ = ~new_n1009_ | ~new_n7251_;
  assign new_n7560_ = ~new_n1326_ | ~new_n7100_;
  assign new_n7561_ = ~new_n1009_ | ~new_n7251_;
  assign new_n7562_ = ~new_n1326_ | ~new_n7100_;
  assign new_n7563_ = ~new_n7562_ | ~new_n7561_;
  assign new_n7564_ = ~new_n1009_ | ~new_n7252_;
  assign new_n7565_ = ~new_n1268_ | ~new_n7100_;
  assign new_n7566_ = ~new_n1009_ | ~new_n7252_;
  assign new_n7567_ = ~new_n1268_ | ~new_n7100_;
  assign new_n7568_ = ~new_n7567_ | ~new_n7566_;
  assign new_n7569_ = ~new_n7243_ | ~new_n7253_;
  assign new_n7570_ = ~new_n7334_ | ~new_n7525_;
  assign new_n7571_ = ~new_n7459_ | ~new_n7254_;
  assign new_n7572_ = ~new_n7162_ | ~new_n7330_;
  assign new_n7573_ = ~new_n7533_ | ~new_n1301_;
  assign new_n7574_ = ~new_n7155_ | ~new_n7102_;
  assign new_n7575_ = ~new_n7574_ | ~new_n7573_;
  assign new_n7576_ = ~new_n7460_ | ~new_n7112_;
  assign new_n7577_ = ~new_n7575_ | ~new_n7338_;
  assign new_n7578_ = ~new_n7461_ | ~new_n7255_;
  assign new_n7579_ = ~new_n7165_ | ~new_n7336_;
  assign new_n7580_ = ~new_n7462_ | ~new_n7256_;
  assign new_n7581_ = ~new_n7167_ | ~new_n7319_;
  assign new_n7582_ = ~new_n1009_ | ~new_n7257_;
  assign new_n7583_ = ~new_n1308_ | ~new_n7100_;
  assign new_n7584_ = ~new_n1009_ | ~new_n7257_;
  assign new_n7585_ = ~new_n1308_ | ~new_n7100_;
  assign new_n7586_ = ~new_n7585_ | ~new_n7584_;
  assign new_n7587_ = ~new_n1009_ | ~new_n7259_;
  assign new_n7588_ = ~new_n1270_ | ~new_n7100_;
  assign new_n7589_ = ~new_n1009_ | ~new_n7260_;
  assign new_n7590_ = ~new_n1271_ | ~new_n7100_;
  assign new_n7591_ = ~new_n1009_ | ~new_n7260_;
  assign new_n7592_ = ~new_n1271_ | ~new_n7100_;
  assign new_n7593_ = ~new_n7592_ | ~new_n7591_;
  assign new_n7594_ = ~new_n1009_ | ~new_n7259_;
  assign new_n7595_ = ~new_n1270_ | ~new_n7100_;
  assign new_n7596_ = ~new_n7595_ | ~new_n7594_;
  assign new_n7597_ = ~new_n1009_ | ~new_n7261_;
  assign new_n7598_ = ~new_n1274_ | ~new_n7100_;
  assign new_n7599_ = ~new_n7157_;
  assign new_n7600_ = ~new_n1009_ | ~new_n7262_;
  assign new_n7601_ = ~new_n1272_ | ~new_n7100_;
  assign new_n7602_ = ~new_n1009_ | ~new_n7263_;
  assign new_n7603_ = ~new_n1273_ | ~new_n7100_;
  assign new_n7604_ = ~new_n7158_;
  assign new_n7605_ = ~new_n1009_ | ~new_n7264_;
  assign new_n7606_ = ~new_n1275_ | ~new_n7100_;
  assign new_n7607_ = ~new_n1009_ | ~new_n7262_;
  assign new_n7608_ = ~new_n1272_ | ~new_n7100_;
  assign new_n7609_ = ~new_n7608_ | ~new_n7607_;
  assign new_n7610_ = ~new_n1009_ | ~new_n7264_;
  assign new_n7611_ = ~new_n1275_ | ~new_n7100_;
  assign new_n7612_ = ~new_n7159_;
  assign new_n7613_ = ~new_n1009_ | ~new_n7265_;
  assign new_n7614_ = ~new_n1321_ | ~new_n7100_;
  assign new_n7615_ = ~new_n1009_ | ~new_n7266_;
  assign new_n7616_ = ~new_n1322_ | ~new_n7100_;
  assign new_n7617_ = ~new_n1009_ | ~new_n7267_;
  assign new_n7618_ = ~new_n1323_ | ~new_n7100_;
  assign new_n7619_ = ~new_n1009_ | ~new_n7268_;
  assign new_n7620_ = ~new_n1320_ | ~new_n7100_;
  assign new_n7621_ = ~new_n1009_ | ~new_n7269_;
  assign new_n7622_ = ~new_n1315_ | ~new_n7100_;
  assign new_n7623_ = ~new_n1009_ | ~new_n7270_;
  assign new_n7624_ = ~new_n1316_ | ~new_n7100_;
  assign new_n7625_ = ~new_n1009_ | ~new_n7271_;
  assign new_n7626_ = ~new_n1317_ | ~new_n7100_;
  assign new_n7627_ = ~new_n1009_ | ~new_n7272_;
  assign new_n7628_ = ~new_n1318_ | ~new_n7100_;
  assign new_n7629_ = ~new_n1009_ | ~new_n7273_;
  assign new_n7630_ = ~new_n1319_ | ~new_n7100_;
  assign new_n7631_ = ~new_n7156_;
  assign new_n7632_ = ~new_n1009_ | ~new_n7274_;
  assign new_n7633_ = ~new_n1311_ | ~new_n7100_;
  assign new_n7634_ = ~new_n1009_ | ~new_n7275_;
  assign new_n7635_ = ~new_n1312_ | ~new_n7100_;
  assign new_n7636_ = ~new_n1009_ | ~new_n7276_;
  assign new_n7637_ = ~new_n1313_ | ~new_n7100_;
  assign new_n7638_ = ~new_n1009_ | ~new_n7277_;
  assign new_n7639_ = ~new_n1314_ | ~new_n7100_;
  assign new_n7640_ = ~new_n1009_ | ~new_n7278_;
  assign new_n7641_ = ~new_n1309_ | ~new_n7100_;
  assign new_n7642_ = ~new_n1009_ | ~new_n7279_;
  assign new_n7643_ = ~new_n1310_ | ~new_n7100_;
  assign new_n7644_ = ~new_n1009_ | ~new_n7269_;
  assign new_n7645_ = ~new_n1315_ | ~new_n7100_;
  assign new_n7646_ = ~new_n7645_ | ~new_n7644_;
  assign new_n7647_ = ~new_n1009_ | ~new_n7270_;
  assign new_n7648_ = ~new_n1316_ | ~new_n7100_;
  assign new_n7649_ = ~new_n7648_ | ~new_n7647_;
  assign new_n7650_ = ~new_n1009_ | ~new_n7271_;
  assign new_n7651_ = ~new_n1317_ | ~new_n7100_;
  assign new_n7652_ = ~new_n7651_ | ~new_n7650_;
  assign new_n7653_ = ~new_n1009_ | ~new_n7272_;
  assign new_n7654_ = ~new_n1318_ | ~new_n7100_;
  assign new_n7655_ = ~new_n7654_ | ~new_n7653_;
  assign new_n7656_ = ~new_n1009_ | ~new_n7278_;
  assign new_n7657_ = ~new_n1309_ | ~new_n7100_;
  assign new_n7658_ = ~new_n7657_ | ~new_n7656_;
  assign new_n7659_ = ~new_n1009_ | ~new_n7277_;
  assign new_n7660_ = ~new_n1314_ | ~new_n7100_;
  assign new_n7661_ = ~new_n7660_ | ~new_n7659_;
  assign new_n7662_ = ~new_n1009_ | ~new_n7276_;
  assign new_n7663_ = ~new_n1313_ | ~new_n7100_;
  assign new_n7664_ = ~new_n7663_ | ~new_n7662_;
  assign new_n7665_ = ~new_n1009_ | ~new_n7275_;
  assign new_n7666_ = ~new_n1312_ | ~new_n7100_;
  assign new_n7667_ = ~new_n7666_ | ~new_n7665_;
  assign new_n7668_ = ~new_n1009_ | ~new_n7274_;
  assign new_n7669_ = ~new_n1311_ | ~new_n7100_;
  assign new_n7670_ = ~new_n7669_ | ~new_n7668_;
  assign new_n7671_ = ~new_n1009_ | ~new_n7279_;
  assign new_n7672_ = ~new_n1310_ | ~new_n7100_;
  assign new_n7673_ = ~new_n7672_ | ~new_n7671_;
  assign new_n7674_ = ~new_n1009_ | ~new_n7268_;
  assign new_n7675_ = ~new_n1320_ | ~new_n7100_;
  assign new_n7676_ = ~new_n7675_ | ~new_n7674_;
  assign new_n7677_ = ~new_n1009_ | ~new_n7267_;
  assign new_n7678_ = ~new_n1323_ | ~new_n7100_;
  assign new_n7679_ = ~new_n7678_ | ~new_n7677_;
  assign new_n7680_ = ~new_n1009_ | ~new_n7265_;
  assign new_n7681_ = ~new_n1321_ | ~new_n7100_;
  assign new_n7682_ = ~new_n7681_ | ~new_n7680_;
  assign new_n7683_ = ~new_n1009_ | ~new_n7266_;
  assign new_n7684_ = ~new_n1322_ | ~new_n7100_;
  assign new_n7685_ = ~new_n7684_ | ~new_n7683_;
  assign new_n7686_ = ~new_n7258_ | ~new_n7280_;
  assign new_n7687_ = ~new_n7408_ | ~new_n7586_;
  assign new_n7688_ = ~new_n7463_ | ~new_n7281_;
  assign new_n7689_ = ~new_n7170_ | ~new_n7411_;
  assign new_n7690_ = ~new_n7464_ | ~new_n7282_;
  assign new_n7691_ = ~new_n7172_ | ~new_n7417_;
  assign new_n7692_ = ~new_n7465_ | ~new_n7283_;
  assign new_n7693_ = ~new_n7174_ | ~new_n7419_;
  assign new_n7694_ = ~new_n7299_ | ~new_n7466_;
  assign new_n7695_ = ~new_n7176_ | ~new_n7284_;
  assign new_n7696_ = ~new_n7467_ | ~new_n7285_;
  assign new_n7697_ = ~new_n7178_ | ~new_n7421_;
  assign new_n7698_ = ~new_n7468_ | ~new_n7286_;
  assign new_n7699_ = ~new_n7180_ | ~new_n7409_;
  assign new_n7700_ = ~new_n7469_ | ~new_n7287_;
  assign new_n7701_ = ~new_n7182_ | ~new_n7426_;
  assign new_n7702_ = ~new_n7470_ | ~new_n7288_;
  assign new_n7703_ = ~new_n7184_ | ~new_n7424_;
  assign new_n7704_ = ~new_n7298_ | ~new_n7471_;
  assign new_n7705_ = ~new_n7186_ | ~new_n7289_;
  assign new_n7706_ = ~new_n7631_ | ~new_n1287_;
  assign new_n7707_ = ~new_n7156_ | ~new_n7123_;
  assign new_n7708_ = ~new_n7707_ | ~new_n7706_;
  assign new_n7709_ = ~new_n7472_ | ~new_n7146_;
  assign new_n7710_ = ~new_n7708_ | ~new_n7396_;
  assign new_n7711_ = ~new_n7473_ | ~new_n7290_;
  assign new_n7712_ = ~new_n7189_ | ~new_n7347_;
  assign new_n7713_ = ~new_n7474_ | ~new_n7291_;
  assign new_n7714_ = ~new_n7191_ | ~new_n7393_;
  assign new_n7715_ = ~new_n7475_ | ~new_n7292_;
  assign new_n7716_ = ~new_n7193_ | ~new_n7435_;
  assign new_n7717_ = ~new_n7476_ | ~new_n7293_;
  assign new_n7718_ = ~new_n7195_ | ~new_n7433_;
  assign new_n7719_ = ~new_n7599_ | ~new_n1293_;
  assign new_n7720_ = ~new_n7157_ | ~new_n7132_;
  assign new_n7721_ = ~new_n7720_ | ~new_n7719_;
  assign new_n7722_ = ~new_n7477_ | ~new_n7150_;
  assign new_n7723_ = ~new_n7721_ | ~new_n7443_;
  assign new_n7724_ = ~new_n7604_ | ~new_n1294_;
  assign new_n7725_ = ~new_n7158_ | ~new_n7128_;
  assign new_n7726_ = ~new_n7725_ | ~new_n7724_;
  assign new_n7727_ = ~new_n7478_ | ~new_n7294_;
  assign new_n7728_ = ~new_n7440_ | ~new_n7726_;
  assign new_n7729_ = ~new_n7479_ | ~new_n7295_;
  assign new_n7730_ = ~new_n7199_ | ~new_n7386_;
  assign new_n7731_ = ~new_n1009_ | ~new_n7296_;
  assign new_n7732_ = ~new_n7458_ | ~new_n7100_;
  assign new_n7733_ = ~pi281;
  assign new_n7734_ = ~pi285;
  assign new_n7735_ = ~pi284;
  assign new_n7736_ = ~pi283;
  assign new_n7737_ = ~pi282;
  assign new_n7738_ = ~pi283 | ~pi282 | ~pi284 | ~pi285 | ~pi281;
  assign new_n7739_ = ~pi287;
  assign new_n7740_ = ~pi286;
  assign new_n7741_ = ~new_n7809_ | ~new_n7836_;
  assign new_n7742_ = ~pi288;
  assign new_n7743_ = ~pi289;
  assign new_n7744_ = ~pi282 | ~pi283 | ~pi281;
  assign new_n7745_ = ~new_n7810_ | ~new_n7838_;
  assign new_n7746_ = ~pi291;
  assign new_n7747_ = ~pi290;
  assign new_n7748_ = ~new_n7811_ | ~new_n7840_;
  assign new_n7749_ = ~pi293;
  assign new_n7750_ = ~pi292;
  assign new_n7751_ = ~new_n7812_ | ~new_n7842_;
  assign new_n7752_ = ~pi295;
  assign new_n7753_ = ~pi294;
  assign new_n7754_ = ~new_n7813_ | ~new_n7844_;
  assign new_n7755_ = ~pi297;
  assign new_n7756_ = ~pi296;
  assign new_n7757_ = ~new_n7814_ | ~new_n7846_;
  assign new_n7758_ = ~pi299;
  assign new_n7759_ = ~pi298;
  assign new_n7760_ = ~new_n7815_ | ~new_n7848_;
  assign new_n7761_ = ~pi301;
  assign new_n7762_ = ~pi300;
  assign new_n7763_ = ~new_n7816_ | ~new_n7850_;
  assign new_n7764_ = ~pi303;
  assign new_n7765_ = ~pi302;
  assign new_n7766_ = ~new_n7817_ | ~new_n7852_;
  assign new_n7767_ = ~pi305;
  assign new_n7768_ = ~pi304;
  assign new_n7769_ = ~new_n7818_ | ~new_n7854_;
  assign new_n7770_ = ~pi306;
  assign new_n7771_ = ~pi306 | ~new_n7856_;
  assign new_n7772_ = ~pi307;
  assign new_n7773_ = ~pi307 | ~new_n7857_;
  assign new_n7774_ = ~pi308;
  assign new_n7775_ = ~pi308 | ~new_n7858_;
  assign new_n7776_ = ~pi309;
  assign new_n7777_ = ~pi309 | ~new_n7859_;
  assign new_n7778_ = ~pi310;
  assign new_n7779_ = ~new_n7863_ | ~new_n7862_;
  assign new_n7780_ = ~new_n7865_ | ~new_n7864_;
  assign new_n7781_ = ~new_n7867_ | ~new_n7866_;
  assign new_n7782_ = ~new_n7869_ | ~new_n7868_;
  assign new_n7783_ = ~new_n7871_ | ~new_n7870_;
  assign new_n7784_ = ~new_n7873_ | ~new_n7872_;
  assign new_n7785_ = ~new_n7875_ | ~new_n7874_;
  assign new_n7786_ = ~new_n7877_ | ~new_n7876_;
  assign new_n7787_ = ~new_n7879_ | ~new_n7878_;
  assign new_n7788_ = ~new_n7881_ | ~new_n7880_;
  assign new_n7789_ = ~new_n7883_ | ~new_n7882_;
  assign new_n7790_ = ~new_n7885_ | ~new_n7884_;
  assign new_n7791_ = ~new_n7887_ | ~new_n7886_;
  assign new_n7792_ = ~new_n7889_ | ~new_n7888_;
  assign new_n7793_ = ~new_n7891_ | ~new_n7890_;
  assign new_n7794_ = ~new_n7893_ | ~new_n7892_;
  assign new_n7795_ = ~new_n7895_ | ~new_n7894_;
  assign new_n7796_ = ~new_n7897_ | ~new_n7896_;
  assign new_n7797_ = ~new_n7899_ | ~new_n7898_;
  assign new_n7798_ = ~new_n7901_ | ~new_n7900_;
  assign new_n7799_ = ~new_n7903_ | ~new_n7902_;
  assign new_n7800_ = ~new_n7905_ | ~new_n7904_;
  assign new_n7801_ = ~new_n7907_ | ~new_n7906_;
  assign new_n7802_ = ~new_n7909_ | ~new_n7908_;
  assign new_n7803_ = ~new_n7911_ | ~new_n7910_;
  assign new_n7804_ = ~new_n7913_ | ~new_n7912_;
  assign new_n7805_ = ~new_n7915_ | ~new_n7914_;
  assign new_n7806_ = ~new_n7917_ | ~new_n7916_;
  assign new_n7807_ = ~new_n7919_ | ~new_n7918_;
  assign new_n7808_ = ~new_n7921_ | ~new_n7920_;
  assign new_n7809_ = pi287 & pi286;
  assign new_n7810_ = pi288 & pi289;
  assign new_n7811_ = pi291 & pi290;
  assign new_n7812_ = pi293 & pi292;
  assign new_n7813_ = pi295 & pi294;
  assign new_n7814_ = pi297 & pi296;
  assign new_n7815_ = pi299 & pi298;
  assign new_n7816_ = pi301 & pi300;
  assign new_n7817_ = pi303 & pi302;
  assign new_n7818_ = pi305 & pi304;
  assign new_n7819_ = ~pi288 | ~new_n7838_;
  assign new_n7820_ = ~pi286 | ~new_n7836_;
  assign new_n7821_ = ~new_n7834_ | ~pi284;
  assign new_n7822_ = ~pi282 | ~pi281;
  assign new_n7823_ = ~pi311;
  assign new_n7824_ = ~pi310 | ~new_n7860_;
  assign new_n7825_ = ~pi304 | ~new_n7854_;
  assign new_n7826_ = ~pi302 | ~new_n7852_;
  assign new_n7827_ = ~pi300 | ~new_n7850_;
  assign new_n7828_ = ~pi298 | ~new_n7848_;
  assign new_n7829_ = ~pi296 | ~new_n7846_;
  assign new_n7830_ = ~pi294 | ~new_n7844_;
  assign new_n7831_ = ~pi292 | ~new_n7842_;
  assign new_n7832_ = ~pi290 | ~new_n7840_;
  assign new_n7833_ = ~new_n7822_;
  assign new_n7834_ = ~new_n7744_;
  assign new_n7835_ = ~new_n7821_;
  assign new_n7836_ = ~new_n7738_;
  assign new_n7837_ = ~new_n7820_;
  assign new_n7838_ = ~new_n7741_;
  assign new_n7839_ = ~new_n7819_;
  assign new_n7840_ = ~new_n7745_;
  assign new_n7841_ = ~new_n7832_;
  assign new_n7842_ = ~new_n7748_;
  assign new_n7843_ = ~new_n7831_;
  assign new_n7844_ = ~new_n7751_;
  assign new_n7845_ = ~new_n7830_;
  assign new_n7846_ = ~new_n7754_;
  assign new_n7847_ = ~new_n7829_;
  assign new_n7848_ = ~new_n7757_;
  assign new_n7849_ = ~new_n7828_;
  assign new_n7850_ = ~new_n7760_;
  assign new_n7851_ = ~new_n7827_;
  assign new_n7852_ = ~new_n7763_;
  assign new_n7853_ = ~new_n7826_;
  assign new_n7854_ = ~new_n7766_;
  assign new_n7855_ = ~new_n7825_;
  assign new_n7856_ = ~new_n7769_;
  assign new_n7857_ = ~new_n7771_;
  assign new_n7858_ = ~new_n7773_;
  assign new_n7859_ = ~new_n7775_;
  assign new_n7860_ = ~new_n7777_;
  assign new_n7861_ = ~new_n7824_;
  assign new_n7862_ = ~pi289 | ~new_n7819_;
  assign new_n7863_ = ~new_n7839_ | ~new_n7743_;
  assign new_n7864_ = ~pi288 | ~new_n7741_;
  assign new_n7865_ = ~new_n7838_ | ~new_n7742_;
  assign new_n7866_ = ~pi287 | ~new_n7820_;
  assign new_n7867_ = ~new_n7837_ | ~new_n7739_;
  assign new_n7868_ = ~pi286 | ~new_n7738_;
  assign new_n7869_ = ~new_n7836_ | ~new_n7740_;
  assign new_n7870_ = ~pi285 | ~new_n7821_;
  assign new_n7871_ = ~new_n7835_ | ~new_n7734_;
  assign new_n7872_ = ~pi284 | ~new_n7744_;
  assign new_n7873_ = ~new_n7834_ | ~new_n7735_;
  assign new_n7874_ = ~pi283 | ~new_n7822_;
  assign new_n7875_ = ~new_n7833_ | ~new_n7736_;
  assign new_n7876_ = ~pi311 | ~new_n7824_;
  assign new_n7877_ = ~new_n7861_ | ~new_n7823_;
  assign new_n7878_ = ~pi310 | ~new_n7777_;
  assign new_n7879_ = ~new_n7860_ | ~new_n7778_;
  assign new_n7880_ = ~pi281 | ~new_n7737_;
  assign new_n7881_ = ~pi282 | ~new_n7733_;
  assign new_n7882_ = ~pi309 | ~new_n7775_;
  assign new_n7883_ = ~new_n7859_ | ~new_n7776_;
  assign new_n7884_ = ~pi308 | ~new_n7773_;
  assign new_n7885_ = ~new_n7858_ | ~new_n7774_;
  assign new_n7886_ = ~pi307 | ~new_n7771_;
  assign new_n7887_ = ~new_n7857_ | ~new_n7772_;
  assign new_n7888_ = ~pi306 | ~new_n7769_;
  assign new_n7889_ = ~new_n7856_ | ~new_n7770_;
  assign new_n7890_ = ~pi305 | ~new_n7825_;
  assign new_n7891_ = ~new_n7855_ | ~new_n7767_;
  assign new_n7892_ = ~pi304 | ~new_n7766_;
  assign new_n7893_ = ~new_n7854_ | ~new_n7768_;
  assign new_n7894_ = ~pi303 | ~new_n7826_;
  assign new_n7895_ = ~new_n7853_ | ~new_n7764_;
  assign new_n7896_ = ~pi302 | ~new_n7763_;
  assign new_n7897_ = ~new_n7852_ | ~new_n7765_;
  assign new_n7898_ = ~pi301 | ~new_n7827_;
  assign new_n7899_ = ~new_n7851_ | ~new_n7761_;
  assign new_n7900_ = ~pi300 | ~new_n7760_;
  assign new_n7901_ = ~new_n7850_ | ~new_n7762_;
  assign new_n7902_ = ~pi299 | ~new_n7828_;
  assign new_n7903_ = ~new_n7849_ | ~new_n7758_;
  assign new_n7904_ = ~pi298 | ~new_n7757_;
  assign new_n7905_ = ~new_n7848_ | ~new_n7759_;
  assign new_n7906_ = ~pi297 | ~new_n7829_;
  assign new_n7907_ = ~new_n7847_ | ~new_n7755_;
  assign new_n7908_ = ~pi296 | ~new_n7754_;
  assign new_n7909_ = ~new_n7846_ | ~new_n7756_;
  assign new_n7910_ = ~pi295 | ~new_n7830_;
  assign new_n7911_ = ~new_n7845_ | ~new_n7752_;
  assign new_n7912_ = ~pi294 | ~new_n7751_;
  assign new_n7913_ = ~new_n7844_ | ~new_n7753_;
  assign new_n7914_ = ~pi293 | ~new_n7831_;
  assign new_n7915_ = ~new_n7843_ | ~new_n7749_;
  assign new_n7916_ = ~pi292 | ~new_n7748_;
  assign new_n7917_ = ~new_n7842_ | ~new_n7750_;
  assign new_n7918_ = ~pi291 | ~new_n7832_;
  assign new_n7919_ = ~new_n7841_ | ~new_n7746_;
  assign new_n7920_ = ~pi290 | ~new_n7745_;
  assign new_n7921_ = ~new_n7840_ | ~new_n7747_;
  assign new_n7922_ = new_n7964_ & new_n1397_;
  assign new_n7923_ = new_n7977_ & new_n7933_;
  assign new_n7924_ = ~new_n1401_;
  assign new_n7925_ = ~new_n1890_;
  assign new_n7926_ = ~new_n1890_ | ~new_n1401_;
  assign new_n7927_ = ~new_n1399_;
  assign new_n7928_ = ~new_n1398_;
  assign new_n7929_ = ~new_n1397_;
  assign new_n7930_ = ~new_n7952_ | ~new_n7958_;
  assign new_n7931_ = ~new_n1394_;
  assign new_n7932_ = ~new_n1395_;
  assign new_n7933_ = ~new_n1380_ | ~new_n1396_;
  assign new_n7934_ = ~new_n1393_;
  assign new_n7935_ = ~new_n1392_;
  assign new_n7936_ = ~new_n7953_ | ~new_n7966_;
  assign new_n7937_ = ~new_n1391_;
  assign new_n7938_ = ~new_n7954_ | ~new_n7963_;
  assign new_n7939_ = ~new_n7965_ | ~new_n1391_;
  assign new_n7940_ = ~new_n1390_;
  assign new_n7941_ = ~new_n7981_ | ~new_n7980_;
  assign new_n7942_ = ~new_n7983_ | ~new_n7982_;
  assign new_n7943_ = ~new_n7985_ | ~new_n7984_;
  assign new_n7944_ = ~new_n7989_ | ~new_n7988_;
  assign new_n7945_ = ~new_n7991_ | ~new_n7990_;
  assign new_n7946_ = ~new_n7993_ | ~new_n7992_;
  assign new_n7947_ = ~new_n7995_ | ~new_n7994_;
  assign new_n7948_ = ~new_n7997_ | ~new_n7996_;
  assign new_n7949_ = ~new_n7999_ | ~new_n7998_;
  assign new_n7950_ = ~new_n8001_ | ~new_n8000_;
  assign new_n7951_ = ~new_n8003_ | ~new_n8002_;
  assign new_n7952_ = new_n1399_ & new_n1398_;
  assign new_n7953_ = new_n1395_ & new_n1394_;
  assign new_n7954_ = new_n1392_ & new_n1393_;
  assign new_n7955_ = ~new_n1399_ | ~new_n7958_;
  assign new_n7956_ = ~new_n1389_;
  assign new_n7957_ = ~new_n1390_ | ~new_n7973_;
  assign new_n7958_ = ~new_n7969_ | ~new_n7970_;
  assign new_n7959_ = new_n7987_ & new_n7986_;
  assign new_n7960_ = ~new_n7963_ | ~new_n1393_;
  assign new_n7961_ = ~new_n7966_ | ~new_n1395_;
  assign new_n7962_ = ~new_n7968_ | ~new_n7979_;
  assign new_n7963_ = ~new_n7936_;
  assign new_n7964_ = ~new_n7930_;
  assign new_n7965_ = ~new_n7938_;
  assign new_n7966_ = ~new_n7933_;
  assign new_n7967_ = ~new_n7926_;
  assign new_n7968_ = new_n1400_ | new_n1388_;
  assign new_n7969_ = ~new_n1388_ | ~new_n1400_;
  assign new_n7970_ = ~new_n7967_ | ~new_n7968_;
  assign new_n7971_ = ~new_n7958_;
  assign new_n7972_ = ~new_n7955_;
  assign new_n7973_ = ~new_n7939_;
  assign new_n7974_ = ~new_n7957_;
  assign new_n7975_ = ~new_n7960_;
  assign new_n7976_ = ~new_n7961_;
  assign new_n7977_ = new_n1396_ | new_n1380_;
  assign new_n7978_ = ~new_n7962_;
  assign new_n7979_ = ~new_n1388_ | ~new_n1400_;
  assign new_n7980_ = ~new_n7964_ | ~new_n7929_;
  assign new_n7981_ = ~new_n1397_ | ~new_n7930_;
  assign new_n7982_ = ~new_n1398_ | ~new_n7955_;
  assign new_n7983_ = ~new_n7972_ | ~new_n7928_;
  assign new_n7984_ = ~new_n1389_ | ~new_n7957_;
  assign new_n7985_ = ~new_n7974_ | ~new_n7956_;
  assign new_n7986_ = ~new_n1399_ | ~new_n7958_;
  assign new_n7987_ = ~new_n7971_ | ~new_n7927_;
  assign new_n7988_ = ~new_n1390_ | ~new_n7939_;
  assign new_n7989_ = ~new_n7973_ | ~new_n7940_;
  assign new_n7990_ = ~new_n7965_ | ~new_n7937_;
  assign new_n7991_ = ~new_n1391_ | ~new_n7938_;
  assign new_n7992_ = ~new_n1392_ | ~new_n7960_;
  assign new_n7993_ = ~new_n7975_ | ~new_n7935_;
  assign new_n7994_ = ~new_n7963_ | ~new_n7934_;
  assign new_n7995_ = ~new_n1393_ | ~new_n7936_;
  assign new_n7996_ = ~new_n1394_ | ~new_n7961_;
  assign new_n7997_ = ~new_n7976_ | ~new_n7931_;
  assign new_n7998_ = ~new_n7966_ | ~new_n7932_;
  assign new_n7999_ = ~new_n1395_ | ~new_n7933_;
  assign new_n8000_ = ~new_n7967_ | ~new_n7962_;
  assign new_n8001_ = ~new_n7978_ | ~new_n7926_;
  assign new_n8002_ = ~new_n1890_ | ~new_n7924_;
  assign new_n8003_ = ~new_n1401_ | ~new_n7925_;
  assign new_n8004_ = new_n8103_ & new_n8102_;
  assign new_n8005_ = new_n8028_ & new_n8026_ & new_n8035_ & new_n8034_;
  assign new_n8006_ = new_n8103_ & new_n8080_;
  assign new_n8007_ = new_n8137_ & new_n8135_;
  assign new_n8008_ = new_n8127_ & new_n8126_;
  assign new_n8009_ = new_n8081_ & new_n8212_ & new_n8211_;
  assign new_n8010_ = ~new_n8143_ | ~new_n8145_;
  assign new_n8011_ = ~new_n1012_;
  assign new_n8012_ = ~new_n1407_;
  assign new_n8013_ = ~new_n1408_;
  assign new_n8014_ = ~new_n1409_;
  assign new_n8015_ = ~new_n1406_;
  assign new_n8016_ = ~new_n1402_;
  assign new_n8017_ = ~new_n1405_;
  assign new_n8018_ = ~new_n1405_ | ~new_n8177_;
  assign new_n8019_ = ~new_n1404_;
  assign new_n8020_ = ~new_n1404_ | ~new_n8169_;
  assign new_n8021_ = ~new_n1403_;
  assign new_n8022_ = ~new_n1403_ | ~new_n8172_;
  assign new_n8023_ = ~new_n8078_ | ~new_n8062_;
  assign new_n8024_ = ~new_n8005_ | ~new_n8078_;
  assign new_n8025_ = ~new_n8064_ | ~new_n8140_;
  assign new_n8026_ = ~new_n8205_ | ~new_n8204_;
  assign new_n8027_ = ~new_n8185_ | ~new_n8184_;
  assign new_n8028_ = ~new_n8202_ | ~new_n8201_;
  assign new_n8029_ = ~new_n8208_ | ~new_n8207_;
  assign new_n8030_ = ~new_n8223_ | ~new_n8222_;
  assign new_n8031_ = ~new_n8220_ | ~new_n8219_;
  assign new_n8032_ = ~new_n8226_ | ~new_n8225_;
  assign new_n8033_ = ~new_n8229_ | ~new_n8228_;
  assign new_n8034_ = ~new_n8232_ | ~new_n8231_;
  assign new_n8035_ = ~new_n8235_ | ~new_n8234_;
  assign new_n8036_ = ~new_n8247_ | ~new_n8246_;
  assign new_n8037_ = ~new_n8249_ | ~new_n8248_;
  assign new_n8038_ = ~new_n8251_ | ~new_n8250_;
  assign new_n8039_ = ~new_n8253_ | ~new_n8252_;
  assign new_n8040_ = ~new_n8255_ | ~new_n8254_;
  assign new_n8041_ = ~new_n8257_ | ~new_n8256_;
  assign new_n8042_ = ~new_n8259_ | ~new_n8258_;
  assign new_n8043_ = new_n8020_ & new_n8104_;
  assign new_n8044_ = ~new_n8216_ | ~new_n8215_;
  assign new_n8045_ = new_n8018_ & new_n8105_;
  assign new_n8046_ = ~new_n8218_ | ~new_n8217_;
  assign new_n8047_ = new_n8161_ & new_n8108_;
  assign new_n8048_ = ~new_n8238_ | ~new_n8237_;
  assign new_n8049_ = ~new_n8245_ | ~new_n8244_;
  assign new_n8050_ = new_n8109_ & new_n8108_;
  assign new_n8051_ = new_n8105_ & new_n8104_;
  assign new_n8052_ = new_n8006_ & new_n8051_;
  assign new_n8053_ = new_n8151_ & new_n8152_ & new_n8102_ & new_n8150_;
  assign new_n8054_ = new_n8108_ & new_n8105_;
  assign new_n8055_ = new_n8158_ & new_n8018_;
  assign new_n8056_ = new_n8155_ & new_n8020_;
  assign new_n8057_ = new_n8158_ & new_n8018_ & new_n8020_;
  assign new_n8058_ = new_n8004_ & new_n8104_;
  assign new_n8059_ = new_n8125_ & new_n8020_;
  assign new_n8060_ = new_n8022_ & new_n8080_;
  assign new_n8061_ = new_n8110_ & new_n8109_;
  assign new_n8062_ = new_n8005_ & new_n8063_;
  assign new_n8063_ = new_n8031_ & new_n8030_ & new_n8033_ & new_n8032_;
  assign new_n8064_ = new_n8033_ & new_n8032_;
  assign new_n8065_ = new_n8028_ & new_n8035_ & new_n8026_;
  assign new_n8066_ = new_n8028_ & new_n8026_;
  assign new_n8067_ = ~new_n1419_;
  assign new_n8068_ = ~new_n1418_;
  assign new_n8069_ = ~new_n1420_;
  assign new_n8070_ = ~new_n1421_;
  assign new_n8071_ = ~new_n1423_;
  assign new_n8072_ = ~new_n1424_;
  assign new_n8073_ = ~new_n1425_;
  assign new_n8074_ = ~new_n1422_;
  assign new_n8075_ = ~new_n1417_;
  assign new_n8076_ = ~new_n1416_;
  assign new_n8077_ = ~new_n8028_ | ~new_n8078_;
  assign new_n8078_ = ~new_n8098_ | ~new_n8053_;
  assign new_n8079_ = new_n8210_ & new_n8209_;
  assign new_n8080_ = ~new_n8021_ | ~new_n8164_ | ~new_n8163_;
  assign new_n8081_ = new_n8214_ & new_n8213_;
  assign new_n8082_ = ~new_n8055_ | ~new_n8157_;
  assign new_n8083_ = ~new_n8110_ | ~new_n8117_;
  assign new_n8084_ = ~new_n1411_;
  assign new_n8085_ = ~new_n1410_;
  assign new_n8086_ = ~new_n1412_;
  assign new_n8087_ = ~new_n1413_;
  assign new_n8088_ = ~new_n1414_;
  assign new_n8089_ = ~new_n1415_;
  assign new_n8090_ = ~new_n8099_ | ~new_n8131_;
  assign new_n8091_ = new_n8240_ & new_n8239_;
  assign new_n8092_ = ~new_n8128_ | ~new_n8112_;
  assign new_n8093_ = ~new_n8142_ | ~new_n8031_;
  assign new_n8094_ = ~new_n8140_ | ~new_n8033_;
  assign new_n8095_ = ~new_n8078_ | ~new_n8065_;
  assign new_n8096_ = ~new_n8066_ | ~new_n8078_;
  assign new_n8097_ = ~new_n8112_ | ~new_n8111_;
  assign new_n8098_ = ~new_n8052_ | ~new_n8083_;
  assign new_n8099_ = ~new_n1408_ | ~new_n8027_;
  assign new_n8100_ = ~new_n8023_;
  assign new_n8101_ = ~new_n8080_;
  assign new_n8102_ = ~new_n1402_ | ~new_n8180_;
  assign new_n8103_ = ~new_n8016_ | ~new_n8166_ | ~new_n8165_;
  assign new_n8104_ = ~new_n8019_ | ~new_n8174_ | ~new_n8173_;
  assign new_n8105_ = ~new_n8017_ | ~new_n8200_ | ~new_n8199_;
  assign new_n8106_ = ~new_n8020_;
  assign new_n8107_ = ~new_n8022_;
  assign new_n8108_ = ~new_n8012_ | ~new_n8193_ | ~new_n8192_;
  assign new_n8109_ = ~new_n8015_ | ~new_n8195_ | ~new_n8194_;
  assign new_n8110_ = ~new_n1406_ | ~new_n8198_;
  assign new_n8111_ = ~new_n8014_ | ~new_n8188_ | ~new_n8187_;
  assign new_n8112_ = ~new_n1409_ | ~new_n8191_;
  assign new_n8113_ = ~new_n8186_ | ~new_n8013_;
  assign new_n8114_ = ~new_n1012_ | ~new_n8111_;
  assign new_n8115_ = ~new_n1407_ | ~new_n8183_;
  assign new_n8116_ = ~new_n8154_ | ~new_n8156_;
  assign new_n8117_ = ~new_n8050_ | ~new_n8116_;
  assign new_n8118_ = ~new_n8083_;
  assign new_n8119_ = ~new_n8018_;
  assign new_n8120_ = ~new_n8078_;
  assign new_n8121_ = ~new_n8077_;
  assign new_n8122_ = ~new_n8082_;
  assign new_n8123_ = ~new_n8082_ | ~new_n8104_;
  assign new_n8124_ = ~new_n8020_ | ~new_n8123_;
  assign new_n8125_ = ~new_n8022_ | ~new_n8080_;
  assign new_n8126_ = ~new_n8059_ | ~new_n8123_;
  assign new_n8127_ = ~new_n8060_ | ~new_n8124_;
  assign new_n8128_ = ~new_n1012_ | ~new_n8111_;
  assign new_n8129_ = ~new_n8092_;
  assign new_n8130_ = ~new_n8186_ | ~new_n8013_;
  assign new_n8131_ = ~new_n8130_ | ~new_n8092_;
  assign new_n8132_ = ~new_n8090_;
  assign new_n8133_ = ~new_n8090_ | ~new_n8108_;
  assign new_n8134_ = ~new_n8133_ | ~new_n8115_;
  assign new_n8135_ = ~new_n8061_ | ~new_n8134_;
  assign new_n8136_ = ~new_n8160_ | ~new_n8109_;
  assign new_n8137_ = ~new_n8136_ | ~new_n8133_ | ~new_n8115_;
  assign new_n8138_ = ~new_n8096_;
  assign new_n8139_ = ~new_n8095_;
  assign new_n8140_ = ~new_n8024_;
  assign new_n8141_ = ~new_n8094_;
  assign new_n8142_ = ~new_n8025_;
  assign new_n8143_ = ~new_n1012_ | ~new_n8023_;
  assign new_n8144_ = ~new_n8143_;
  assign new_n8145_ = ~new_n8100_ | ~new_n8011_;
  assign new_n8146_ = ~new_n8093_;
  assign new_n8147_ = ~new_n8097_;
  assign new_n8148_ = ~new_n8020_ | ~new_n8104_;
  assign new_n8149_ = ~new_n8018_ | ~new_n8105_;
  assign new_n8150_ = ~new_n8006_ | ~new_n8119_ | ~new_n8104_;
  assign new_n8151_ = ~new_n8106_ | ~new_n8006_;
  assign new_n8152_ = ~new_n8107_ | ~new_n8006_;
  assign new_n8153_ = ~new_n8099_ | ~new_n8112_ | ~new_n8114_;
  assign new_n8154_ = ~new_n8153_ | ~new_n8113_;
  assign new_n8155_ = ~new_n8103_ | ~new_n8102_;
  assign new_n8156_ = ~new_n1407_ | ~new_n8183_;
  assign new_n8157_ = ~new_n8054_ | ~new_n8116_ | ~new_n8109_;
  assign new_n8158_ = ~new_n8198_ | ~new_n1406_ | ~new_n8105_;
  assign new_n8159_ = ~new_n8057_ | ~new_n8157_;
  assign new_n8160_ = ~new_n1406_ | ~new_n8198_;
  assign new_n8161_ = ~new_n1407_ | ~new_n8183_;
  assign new_n8162_ = ~new_n8115_ | ~new_n8108_;
  assign new_n8163_ = ~new_n1012_ | ~new_n8067_;
  assign new_n8164_ = ~new_n1419_ | ~new_n8011_;
  assign new_n8165_ = ~new_n1012_ | ~new_n8068_;
  assign new_n8166_ = ~new_n1418_ | ~new_n8011_;
  assign new_n8167_ = ~new_n1012_ | ~new_n8069_;
  assign new_n8168_ = ~new_n1420_ | ~new_n8011_;
  assign new_n8169_ = ~new_n8168_ | ~new_n8167_;
  assign new_n8170_ = ~new_n1012_ | ~new_n8067_;
  assign new_n8171_ = ~new_n1419_ | ~new_n8011_;
  assign new_n8172_ = ~new_n8171_ | ~new_n8170_;
  assign new_n8173_ = ~new_n1012_ | ~new_n8069_;
  assign new_n8174_ = ~new_n1420_ | ~new_n8011_;
  assign new_n8175_ = ~new_n1012_ | ~new_n8070_;
  assign new_n8176_ = ~new_n1421_ | ~new_n8011_;
  assign new_n8177_ = ~new_n8176_ | ~new_n8175_;
  assign new_n8178_ = ~new_n1012_ | ~new_n8068_;
  assign new_n8179_ = ~new_n1418_ | ~new_n8011_;
  assign new_n8180_ = ~new_n8179_ | ~new_n8178_;
  assign new_n8181_ = ~new_n1012_ | ~new_n8071_;
  assign new_n8182_ = ~new_n1423_ | ~new_n8011_;
  assign new_n8183_ = ~new_n8182_ | ~new_n8181_;
  assign new_n8184_ = ~new_n1012_ | ~new_n8072_;
  assign new_n8185_ = ~new_n1424_ | ~new_n8011_;
  assign new_n8186_ = ~new_n8027_;
  assign new_n8187_ = ~new_n1012_ | ~new_n8073_;
  assign new_n8188_ = ~new_n1425_ | ~new_n8011_;
  assign new_n8189_ = ~new_n1012_ | ~new_n8073_;
  assign new_n8190_ = ~new_n1425_ | ~new_n8011_;
  assign new_n8191_ = ~new_n8190_ | ~new_n8189_;
  assign new_n8192_ = ~new_n1012_ | ~new_n8071_;
  assign new_n8193_ = ~new_n1423_ | ~new_n8011_;
  assign new_n8194_ = ~new_n1012_ | ~new_n8074_;
  assign new_n8195_ = ~new_n1422_ | ~new_n8011_;
  assign new_n8196_ = ~new_n1012_ | ~new_n8074_;
  assign new_n8197_ = ~new_n1422_ | ~new_n8011_;
  assign new_n8198_ = ~new_n8197_ | ~new_n8196_;
  assign new_n8199_ = ~new_n1012_ | ~new_n8070_;
  assign new_n8200_ = ~new_n1421_ | ~new_n8011_;
  assign new_n8201_ = ~new_n1012_ | ~new_n8075_;
  assign new_n8202_ = ~new_n1417_ | ~new_n8011_;
  assign new_n8203_ = ~new_n8028_;
  assign new_n8204_ = ~new_n1012_ | ~new_n8076_;
  assign new_n8205_ = ~new_n1416_ | ~new_n8011_;
  assign new_n8206_ = ~new_n8026_;
  assign new_n8207_ = ~new_n8121_ | ~new_n8206_;
  assign new_n8208_ = ~new_n8026_ | ~new_n8077_;
  assign new_n8209_ = ~new_n8120_ | ~new_n8203_;
  assign new_n8210_ = ~new_n8028_ | ~new_n8078_;
  assign new_n8211_ = ~new_n8022_ | ~new_n8056_ | ~new_n8123_;
  assign new_n8212_ = ~new_n8004_ | ~new_n8107_;
  assign new_n8213_ = ~new_n8101_ | ~new_n8155_;
  assign new_n8214_ = ~new_n8080_ | ~new_n8058_ | ~new_n8159_;
  assign new_n8215_ = ~new_n8148_ | ~new_n8082_;
  assign new_n8216_ = ~new_n8043_ | ~new_n8122_;
  assign new_n8217_ = ~new_n8149_ | ~new_n8083_;
  assign new_n8218_ = ~new_n8045_ | ~new_n8118_;
  assign new_n8219_ = ~new_n1012_ | ~new_n8084_;
  assign new_n8220_ = ~new_n1411_ | ~new_n8011_;
  assign new_n8221_ = ~new_n8031_;
  assign new_n8222_ = ~new_n1012_ | ~new_n8085_;
  assign new_n8223_ = ~new_n1410_ | ~new_n8011_;
  assign new_n8224_ = ~new_n8030_;
  assign new_n8225_ = ~new_n1012_ | ~new_n8086_;
  assign new_n8226_ = ~new_n1412_ | ~new_n8011_;
  assign new_n8227_ = ~new_n8032_;
  assign new_n8228_ = ~new_n1012_ | ~new_n8087_;
  assign new_n8229_ = ~new_n1413_ | ~new_n8011_;
  assign new_n8230_ = ~new_n8033_;
  assign new_n8231_ = ~new_n1012_ | ~new_n8088_;
  assign new_n8232_ = ~new_n1414_ | ~new_n8011_;
  assign new_n8233_ = ~new_n8034_;
  assign new_n8234_ = ~new_n1012_ | ~new_n8089_;
  assign new_n8235_ = ~new_n1415_ | ~new_n8011_;
  assign new_n8236_ = ~new_n8035_;
  assign new_n8237_ = ~new_n8162_ | ~new_n8090_;
  assign new_n8238_ = ~new_n8047_ | ~new_n8132_;
  assign new_n8239_ = ~new_n8186_ | ~new_n1408_;
  assign new_n8240_ = ~new_n8027_ | ~new_n8013_;
  assign new_n8241_ = ~new_n8186_ | ~new_n1408_;
  assign new_n8242_ = ~new_n8027_ | ~new_n8013_;
  assign new_n8243_ = ~new_n8242_ | ~new_n8241_;
  assign new_n8244_ = ~new_n8091_ | ~new_n8092_;
  assign new_n8245_ = ~new_n8129_ | ~new_n8243_;
  assign new_n8246_ = ~new_n8146_ | ~new_n8224_;
  assign new_n8247_ = ~new_n8030_ | ~new_n8093_;
  assign new_n8248_ = ~new_n8221_ | ~new_n8142_;
  assign new_n8249_ = ~new_n8031_ | ~new_n8025_;
  assign new_n8250_ = ~new_n8141_ | ~new_n8227_;
  assign new_n8251_ = ~new_n8032_ | ~new_n8094_;
  assign new_n8252_ = ~new_n8230_ | ~new_n8140_;
  assign new_n8253_ = ~new_n8033_ | ~new_n8024_;
  assign new_n8254_ = ~new_n8139_ | ~new_n8233_;
  assign new_n8255_ = ~new_n8034_ | ~new_n8095_;
  assign new_n8256_ = ~new_n8138_ | ~new_n8236_;
  assign new_n8257_ = ~new_n8035_ | ~new_n8096_;
  assign new_n8258_ = ~new_n1012_ | ~new_n8097_;
  assign new_n8259_ = ~new_n8147_ | ~new_n8011_;
  assign new_n8260_ = new_n8262_ | new_n1330_;
  assign new_n8261_ = new_n8264_ & new_n8263_;
  assign new_n8262_ = ~new_n8265_ & ~new_n8261_ & ~new_n8266_;
  assign new_n8263_ = ~new_n1333_;
  assign new_n8264_ = ~new_n1334_;
  assign new_n8265_ = ~new_n1331_;
  assign new_n8266_ = ~new_n1332_;
  assign new_n8267_ = ~new_n2835_;
  assign new_n8268_ = ~new_n2834_;
  assign new_n8269_ = ~new_n1335_;
  assign new_n8270_ = ~new_n8351_ | ~new_n8400_;
  assign new_n8271_ = ~new_n8352_ | ~new_n8418_;
  assign new_n8272_ = ~new_n8353_ | ~new_n8420_;
  assign new_n8273_ = ~new_n8354_ | ~new_n8422_;
  assign new_n8274_ = ~new_n8355_ | ~new_n8424_;
  assign new_n8275_ = ~new_n8356_ | ~new_n8426_;
  assign new_n8276_ = ~new_n8357_ | ~new_n8428_;
  assign new_n8277_ = ~new_n8358_ | ~new_n8430_;
  assign new_n8278_ = ~new_n8432_ | ~new_n8318_;
  assign new_n8279_ = ~new_n8433_ | ~new_n8317_;
  assign new_n8280_ = ~new_n8434_ | ~new_n8316_;
  assign new_n8281_ = ~new_n8435_ | ~new_n8315_;
  assign new_n8282_ = ~new_n8436_ | ~new_n8314_;
  assign new_n8283_ = ~new_n8437_ | ~new_n8313_;
  assign new_n8284_ = ~new_n8438_ | ~new_n8312_;
  assign new_n8285_ = ~new_n8439_ | ~new_n8311_;
  assign new_n8286_ = ~new_n8440_ | ~new_n8310_;
  assign new_n8287_ = ~new_n8441_ | ~new_n8309_;
  assign new_n8288_ = ~new_n8442_ | ~new_n8308_;
  assign new_n8289_ = ~new_n8473_ | ~new_n8472_;
  assign new_n8290_ = ~new_n8446_ | ~new_n8445_;
  assign new_n8291_ = ~new_n8467_ | ~new_n8466_;
  assign new_n8292_ = ~new_n8470_ | ~new_n8469_;
  assign new_n8293_ = ~new_n8461_ | ~new_n8460_;
  assign new_n8294_ = ~new_n8464_ | ~new_n8463_;
  assign new_n8295_ = ~new_n8449_ | ~new_n8448_;
  assign new_n8296_ = ~new_n8452_ | ~new_n8451_;
  assign new_n8297_ = ~new_n8458_ | ~new_n8457_;
  assign new_n8298_ = ~new_n8455_ | ~new_n8454_;
  assign new_n8299_ = ~new_n8476_ | ~new_n8475_;
  assign new_n8300_ = ~new_n8478_ | ~new_n8477_;
  assign new_n8301_ = ~new_n8480_ | ~new_n8479_;
  assign new_n8302_ = ~new_n8482_ | ~new_n8481_;
  assign new_n8303_ = ~new_n8484_ | ~new_n8483_;
  assign new_n8304_ = ~new_n8486_ | ~new_n8485_;
  assign new_n8305_ = ~new_n8488_ | ~new_n8487_;
  assign new_n8306_ = ~new_n8547_ | ~new_n8546_;
  assign new_n8307_ = ~new_n8550_ | ~new_n8549_;
  assign new_n8308_ = ~new_n8490_ | ~new_n8489_;
  assign new_n8309_ = ~new_n8493_ | ~new_n8492_;
  assign new_n8310_ = ~new_n8496_ | ~new_n8495_;
  assign new_n8311_ = ~new_n8499_ | ~new_n8498_;
  assign new_n8312_ = ~new_n8502_ | ~new_n8501_;
  assign new_n8313_ = ~new_n8505_ | ~new_n8504_;
  assign new_n8314_ = ~new_n8508_ | ~new_n8507_;
  assign new_n8315_ = ~new_n8511_ | ~new_n8510_;
  assign new_n8316_ = ~new_n8514_ | ~new_n8513_;
  assign new_n8317_ = ~new_n8517_ | ~new_n8516_;
  assign new_n8318_ = ~new_n8520_ | ~new_n8519_;
  assign new_n8319_ = ~new_n8541_ | ~new_n8540_;
  assign new_n8320_ = ~new_n8544_ | ~new_n8543_;
  assign new_n8321_ = ~new_n8535_ | ~new_n8534_;
  assign new_n8322_ = ~new_n8538_ | ~new_n8537_;
  assign new_n8323_ = ~new_n8529_ | ~new_n8528_;
  assign new_n8324_ = ~new_n8532_ | ~new_n8531_;
  assign new_n8325_ = ~new_n8523_ | ~new_n8522_;
  assign new_n8326_ = ~new_n8526_ | ~new_n8525_;
  assign new_n8327_ = ~new_n8556_ | ~new_n8555_;
  assign new_n8328_ = ~new_n8558_ | ~new_n8557_;
  assign new_n8329_ = ~new_n8562_ | ~new_n8561_;
  assign new_n8330_ = ~new_n8564_ | ~new_n8563_;
  assign new_n8331_ = ~new_n8566_ | ~new_n8565_;
  assign new_n8332_ = ~new_n8568_ | ~new_n8567_;
  assign new_n8333_ = ~new_n8570_ | ~new_n8569_;
  assign new_n8334_ = ~new_n8572_ | ~new_n8571_;
  assign new_n8335_ = ~new_n8574_ | ~new_n8573_;
  assign new_n8336_ = ~new_n8576_ | ~new_n8575_;
  assign new_n8337_ = ~new_n8578_ | ~new_n8577_;
  assign new_n8338_ = ~new_n8580_ | ~new_n8579_;
  assign new_n8339_ = ~new_n8589_ | ~new_n8588_;
  assign new_n8340_ = ~new_n8591_ | ~new_n8590_;
  assign new_n8341_ = ~new_n8593_ | ~new_n8592_;
  assign new_n8342_ = ~new_n8595_ | ~new_n8594_;
  assign new_n8343_ = ~new_n8597_ | ~new_n8596_;
  assign new_n8344_ = ~new_n8599_ | ~new_n8598_;
  assign new_n8345_ = ~new_n8601_ | ~new_n8600_;
  assign new_n8346_ = ~new_n8603_ | ~new_n8602_;
  assign new_n8347_ = ~new_n8605_ | ~new_n8604_;
  assign new_n8348_ = ~new_n8607_ | ~new_n8606_;
  assign new_n8349_ = ~new_n8612_ | ~new_n8611_;
  assign new_n8350_ = ~new_n8587_ | ~new_n8586_;
  assign new_n8351_ = new_n8297_ & new_n8298_;
  assign new_n8352_ = new_n8294_ & new_n8293_;
  assign new_n8353_ = new_n8292_ & new_n8291_;
  assign new_n8354_ = new_n8289_ & new_n8290_;
  assign new_n8355_ = new_n8326_ & new_n8325_;
  assign new_n8356_ = new_n8324_ & new_n8323_;
  assign new_n8357_ = new_n8322_ & new_n8321_;
  assign new_n8358_ = new_n8320_ & new_n8319_;
  assign new_n8359_ = new_n8307_ & new_n8306_;
  assign new_n8360_ = ~new_n8553_ | ~new_n8552_;
  assign new_n8361_ = ~new_n8609_ | ~new_n8608_;
  assign new_n8362_ = ~new_n1359_;
  assign new_n8363_ = ~new_n1367_;
  assign new_n8364_ = ~new_n1366_;
  assign new_n8365_ = ~new_n1365_;
  assign new_n8366_ = ~new_n1364_;
  assign new_n8367_ = ~new_n1363_;
  assign new_n8368_ = ~new_n1362_;
  assign new_n8369_ = ~new_n1361_;
  assign new_n8370_ = ~new_n1360_;
  assign new_n8371_ = ~new_n1358_;
  assign new_n8372_ = ~new_n8422_ | ~new_n8290_;
  assign new_n8373_ = ~new_n8420_ | ~new_n8291_;
  assign new_n8374_ = ~new_n8418_ | ~new_n8293_;
  assign new_n8375_ = ~new_n8298_ | ~new_n8400_;
  assign new_n8376_ = ~new_n1339_;
  assign new_n8377_ = ~new_n1340_;
  assign new_n8378_ = ~new_n1341_;
  assign new_n8379_ = ~new_n1342_;
  assign new_n8380_ = ~new_n1343_;
  assign new_n8381_ = ~new_n1344_;
  assign new_n8382_ = ~new_n1345_;
  assign new_n8383_ = ~new_n1346_;
  assign new_n8384_ = ~new_n1347_;
  assign new_n8385_ = ~new_n1348_;
  assign new_n8386_ = ~new_n1349_;
  assign new_n8387_ = ~new_n1357_;
  assign new_n8388_ = ~new_n1356_;
  assign new_n8389_ = ~new_n1355_;
  assign new_n8390_ = ~new_n1354_;
  assign new_n8391_ = ~new_n1353_;
  assign new_n8392_ = ~new_n1352_;
  assign new_n8393_ = ~new_n1351_;
  assign new_n8394_ = ~new_n1350_;
  assign new_n8395_ = ~new_n1337_;
  assign new_n8396_ = ~new_n1338_;
  assign new_n8397_ = ~new_n1336_;
  assign new_n8398_ = ~new_n8359_ | ~new_n8443_;
  assign new_n8399_ = ~new_n8443_ | ~new_n8307_;
  assign new_n8400_ = ~new_n8415_ | ~new_n8414_;
  assign new_n8401_ = new_n8560_ & new_n8559_;
  assign new_n8402_ = new_n8582_ & new_n8581_;
  assign new_n8403_ = ~new_n8411_ | ~new_n8410_;
  assign new_n8404_ = ~new_n8430_ | ~new_n8319_;
  assign new_n8405_ = ~new_n8428_ | ~new_n8321_;
  assign new_n8406_ = ~new_n8426_ | ~new_n8323_;
  assign new_n8407_ = ~new_n8424_ | ~new_n8325_;
  assign new_n8408_ = ~new_n8398_;
  assign new_n8409_ = new_n2835_ | new_n2834_;
  assign new_n8410_ = ~new_n8295_ | ~new_n8409_;
  assign new_n8411_ = ~new_n2834_ | ~new_n2835_;
  assign new_n8412_ = ~new_n8403_;
  assign new_n8413_ = ~new_n8453_ | ~new_n8269_;
  assign new_n8414_ = ~new_n8413_ | ~new_n8403_;
  assign new_n8415_ = ~new_n1335_ | ~new_n8296_;
  assign new_n8416_ = ~new_n8400_;
  assign new_n8417_ = ~new_n8375_;
  assign new_n8418_ = ~new_n8270_;
  assign new_n8419_ = ~new_n8374_;
  assign new_n8420_ = ~new_n8271_;
  assign new_n8421_ = ~new_n8373_;
  assign new_n8422_ = ~new_n8272_;
  assign new_n8423_ = ~new_n8372_;
  assign new_n8424_ = ~new_n8273_;
  assign new_n8425_ = ~new_n8407_;
  assign new_n8426_ = ~new_n8274_;
  assign new_n8427_ = ~new_n8406_;
  assign new_n8428_ = ~new_n8275_;
  assign new_n8429_ = ~new_n8405_;
  assign new_n8430_ = ~new_n8276_;
  assign new_n8431_ = ~new_n8404_;
  assign new_n8432_ = ~new_n8277_;
  assign new_n8433_ = ~new_n8278_;
  assign new_n8434_ = ~new_n8279_;
  assign new_n8435_ = ~new_n8280_;
  assign new_n8436_ = ~new_n8281_;
  assign new_n8437_ = ~new_n8282_;
  assign new_n8438_ = ~new_n8283_;
  assign new_n8439_ = ~new_n8284_;
  assign new_n8440_ = ~new_n8285_;
  assign new_n8441_ = ~new_n8286_;
  assign new_n8442_ = ~new_n8287_;
  assign new_n8443_ = ~new_n8288_;
  assign new_n8444_ = ~new_n8399_;
  assign new_n8445_ = ~new_n2835_ | ~new_n8362_;
  assign new_n8446_ = ~new_n1359_ | ~new_n8267_;
  assign new_n8447_ = ~new_n8290_;
  assign new_n8448_ = ~new_n2835_ | ~new_n8363_;
  assign new_n8449_ = ~new_n1367_ | ~new_n8267_;
  assign new_n8450_ = ~new_n8295_;
  assign new_n8451_ = ~new_n2835_ | ~new_n8364_;
  assign new_n8452_ = ~new_n1366_ | ~new_n8267_;
  assign new_n8453_ = ~new_n8296_;
  assign new_n8454_ = ~new_n2835_ | ~new_n8365_;
  assign new_n8455_ = ~new_n1365_ | ~new_n8267_;
  assign new_n8456_ = ~new_n8298_;
  assign new_n8457_ = ~new_n2835_ | ~new_n8366_;
  assign new_n8458_ = ~new_n1364_ | ~new_n8267_;
  assign new_n8459_ = ~new_n8297_;
  assign new_n8460_ = ~new_n2835_ | ~new_n8367_;
  assign new_n8461_ = ~new_n1363_ | ~new_n8267_;
  assign new_n8462_ = ~new_n8293_;
  assign new_n8463_ = ~new_n2835_ | ~new_n8368_;
  assign new_n8464_ = ~new_n1362_ | ~new_n8267_;
  assign new_n8465_ = ~new_n8294_;
  assign new_n8466_ = ~new_n2835_ | ~new_n8369_;
  assign new_n8467_ = ~new_n1361_ | ~new_n8267_;
  assign new_n8468_ = ~new_n8291_;
  assign new_n8469_ = ~new_n2835_ | ~new_n8370_;
  assign new_n8470_ = ~new_n1360_ | ~new_n8267_;
  assign new_n8471_ = ~new_n8292_;
  assign new_n8472_ = ~new_n2835_ | ~new_n8371_;
  assign new_n8473_ = ~new_n1358_ | ~new_n8267_;
  assign new_n8474_ = ~new_n8289_;
  assign new_n8475_ = ~new_n8423_ | ~new_n8474_;
  assign new_n8476_ = ~new_n8289_ | ~new_n8372_;
  assign new_n8477_ = ~new_n8447_ | ~new_n8422_;
  assign new_n8478_ = ~new_n8290_ | ~new_n8272_;
  assign new_n8479_ = ~new_n8421_ | ~new_n8471_;
  assign new_n8480_ = ~new_n8292_ | ~new_n8373_;
  assign new_n8481_ = ~new_n8468_ | ~new_n8420_;
  assign new_n8482_ = ~new_n8291_ | ~new_n8271_;
  assign new_n8483_ = ~new_n8419_ | ~new_n8465_;
  assign new_n8484_ = ~new_n8294_ | ~new_n8374_;
  assign new_n8485_ = ~new_n8462_ | ~new_n8418_;
  assign new_n8486_ = ~new_n8293_ | ~new_n8270_;
  assign new_n8487_ = ~new_n8417_ | ~new_n8459_;
  assign new_n8488_ = ~new_n8297_ | ~new_n8375_;
  assign new_n8489_ = ~new_n2835_ | ~new_n8376_;
  assign new_n8490_ = ~new_n1339_ | ~new_n8267_;
  assign new_n8491_ = ~new_n8308_;
  assign new_n8492_ = ~new_n2835_ | ~new_n8377_;
  assign new_n8493_ = ~new_n1340_ | ~new_n8267_;
  assign new_n8494_ = ~new_n8309_;
  assign new_n8495_ = ~new_n2835_ | ~new_n8378_;
  assign new_n8496_ = ~new_n1341_ | ~new_n8267_;
  assign new_n8497_ = ~new_n8310_;
  assign new_n8498_ = ~new_n2835_ | ~new_n8379_;
  assign new_n8499_ = ~new_n1342_ | ~new_n8267_;
  assign new_n8500_ = ~new_n8311_;
  assign new_n8501_ = ~new_n2835_ | ~new_n8380_;
  assign new_n8502_ = ~new_n1343_ | ~new_n8267_;
  assign new_n8503_ = ~new_n8312_;
  assign new_n8504_ = ~new_n2835_ | ~new_n8381_;
  assign new_n8505_ = ~new_n1344_ | ~new_n8267_;
  assign new_n8506_ = ~new_n8313_;
  assign new_n8507_ = ~new_n2835_ | ~new_n8382_;
  assign new_n8508_ = ~new_n1345_ | ~new_n8267_;
  assign new_n8509_ = ~new_n8314_;
  assign new_n8510_ = ~new_n2835_ | ~new_n8383_;
  assign new_n8511_ = ~new_n1346_ | ~new_n8267_;
  assign new_n8512_ = ~new_n8315_;
  assign new_n8513_ = ~new_n2835_ | ~new_n8384_;
  assign new_n8514_ = ~new_n1347_ | ~new_n8267_;
  assign new_n8515_ = ~new_n8316_;
  assign new_n8516_ = ~new_n2835_ | ~new_n8385_;
  assign new_n8517_ = ~new_n1348_ | ~new_n8267_;
  assign new_n8518_ = ~new_n8317_;
  assign new_n8519_ = ~new_n2835_ | ~new_n8386_;
  assign new_n8520_ = ~new_n1349_ | ~new_n8267_;
  assign new_n8521_ = ~new_n8318_;
  assign new_n8522_ = ~new_n2835_ | ~new_n8387_;
  assign new_n8523_ = ~new_n1357_ | ~new_n8267_;
  assign new_n8524_ = ~new_n8325_;
  assign new_n8525_ = ~new_n2835_ | ~new_n8388_;
  assign new_n8526_ = ~new_n1356_ | ~new_n8267_;
  assign new_n8527_ = ~new_n8326_;
  assign new_n8528_ = ~new_n2835_ | ~new_n8389_;
  assign new_n8529_ = ~new_n1355_ | ~new_n8267_;
  assign new_n8530_ = ~new_n8323_;
  assign new_n8531_ = ~new_n2835_ | ~new_n8390_;
  assign new_n8532_ = ~new_n1354_ | ~new_n8267_;
  assign new_n8533_ = ~new_n8324_;
  assign new_n8534_ = ~new_n2835_ | ~new_n8391_;
  assign new_n8535_ = ~new_n1353_ | ~new_n8267_;
  assign new_n8536_ = ~new_n8321_;
  assign new_n8537_ = ~new_n2835_ | ~new_n8392_;
  assign new_n8538_ = ~new_n1352_ | ~new_n8267_;
  assign new_n8539_ = ~new_n8322_;
  assign new_n8540_ = ~new_n2835_ | ~new_n8393_;
  assign new_n8541_ = ~new_n1351_ | ~new_n8267_;
  assign new_n8542_ = ~new_n8319_;
  assign new_n8543_ = ~new_n2835_ | ~new_n8394_;
  assign new_n8544_ = ~new_n1350_ | ~new_n8267_;
  assign new_n8545_ = ~new_n8320_;
  assign new_n8546_ = ~new_n2835_ | ~new_n8395_;
  assign new_n8547_ = ~new_n1337_ | ~new_n8267_;
  assign new_n8548_ = ~new_n8306_;
  assign new_n8549_ = ~new_n2835_ | ~new_n8396_;
  assign new_n8550_ = ~new_n1338_ | ~new_n8267_;
  assign new_n8551_ = ~new_n8307_;
  assign new_n8552_ = ~new_n2835_ | ~new_n8397_;
  assign new_n8553_ = ~new_n1336_ | ~new_n8267_;
  assign new_n8554_ = ~new_n8360_;
  assign new_n8555_ = ~new_n8408_ | ~new_n8554_;
  assign new_n8556_ = ~new_n8360_ | ~new_n8398_;
  assign new_n8557_ = ~new_n8444_ | ~new_n8548_;
  assign new_n8558_ = ~new_n8306_ | ~new_n8399_;
  assign new_n8559_ = ~new_n8416_ | ~new_n8456_;
  assign new_n8560_ = ~new_n8298_ | ~new_n8400_;
  assign new_n8561_ = ~new_n8551_ | ~new_n8443_;
  assign new_n8562_ = ~new_n8307_ | ~new_n8288_;
  assign new_n8563_ = ~new_n8491_ | ~new_n8442_;
  assign new_n8564_ = ~new_n8308_ | ~new_n8287_;
  assign new_n8565_ = ~new_n8494_ | ~new_n8441_;
  assign new_n8566_ = ~new_n8309_ | ~new_n8286_;
  assign new_n8567_ = ~new_n8497_ | ~new_n8440_;
  assign new_n8568_ = ~new_n8310_ | ~new_n8285_;
  assign new_n8569_ = ~new_n8500_ | ~new_n8439_;
  assign new_n8570_ = ~new_n8311_ | ~new_n8284_;
  assign new_n8571_ = ~new_n8503_ | ~new_n8438_;
  assign new_n8572_ = ~new_n8312_ | ~new_n8283_;
  assign new_n8573_ = ~new_n8506_ | ~new_n8437_;
  assign new_n8574_ = ~new_n8313_ | ~new_n8282_;
  assign new_n8575_ = ~new_n8509_ | ~new_n8436_;
  assign new_n8576_ = ~new_n8314_ | ~new_n8281_;
  assign new_n8577_ = ~new_n8512_ | ~new_n8435_;
  assign new_n8578_ = ~new_n8315_ | ~new_n8280_;
  assign new_n8579_ = ~new_n8515_ | ~new_n8434_;
  assign new_n8580_ = ~new_n8316_ | ~new_n8279_;
  assign new_n8581_ = ~new_n8453_ | ~new_n1335_;
  assign new_n8582_ = ~new_n8296_ | ~new_n8269_;
  assign new_n8583_ = ~new_n8453_ | ~new_n1335_;
  assign new_n8584_ = ~new_n8296_ | ~new_n8269_;
  assign new_n8585_ = ~new_n8584_ | ~new_n8583_;
  assign new_n8586_ = ~new_n8402_ | ~new_n8403_;
  assign new_n8587_ = ~new_n8412_ | ~new_n8585_;
  assign new_n8588_ = ~new_n8518_ | ~new_n8433_;
  assign new_n8589_ = ~new_n8317_ | ~new_n8278_;
  assign new_n8590_ = ~new_n8521_ | ~new_n8432_;
  assign new_n8591_ = ~new_n8318_ | ~new_n8277_;
  assign new_n8592_ = ~new_n8431_ | ~new_n8545_;
  assign new_n8593_ = ~new_n8320_ | ~new_n8404_;
  assign new_n8594_ = ~new_n8542_ | ~new_n8430_;
  assign new_n8595_ = ~new_n8319_ | ~new_n8276_;
  assign new_n8596_ = ~new_n8429_ | ~new_n8539_;
  assign new_n8597_ = ~new_n8322_ | ~new_n8405_;
  assign new_n8598_ = ~new_n8536_ | ~new_n8428_;
  assign new_n8599_ = ~new_n8321_ | ~new_n8275_;
  assign new_n8600_ = ~new_n8427_ | ~new_n8533_;
  assign new_n8601_ = ~new_n8324_ | ~new_n8406_;
  assign new_n8602_ = ~new_n8530_ | ~new_n8426_;
  assign new_n8603_ = ~new_n8323_ | ~new_n8274_;
  assign new_n8604_ = ~new_n8425_ | ~new_n8527_;
  assign new_n8605_ = ~new_n8326_ | ~new_n8407_;
  assign new_n8606_ = ~new_n8524_ | ~new_n8424_;
  assign new_n8607_ = ~new_n8325_ | ~new_n8273_;
  assign new_n8608_ = ~new_n2834_ | ~new_n8267_;
  assign new_n8609_ = ~new_n2835_ | ~new_n8268_;
  assign new_n8610_ = ~new_n8361_;
  assign new_n8611_ = ~new_n8295_ | ~new_n8610_;
  assign new_n8612_ = ~new_n8361_ | ~new_n8450_;
  assign new_n8613_ = ~new_n1373_;
  assign new_n8614_ = ~new_n1371_;
  assign new_n8615_ = ~new_n1377_;
  assign new_n8616_ = ~new_n1376_;
  assign new_n8617_ = ~new_n1370_;
  assign new_n8618_ = ~new_n1369_;
  assign new_n8619_ = ~new_n1375_;
  assign new_n8620_ = ~new_n1374_;
  assign new_n8621_ = ~new_n1368_;
  assign new_n8622_ = ~new_n1013_;
  assign new_n8623_ = ~pi109;
  assign new_n8624_ = ~new_n8657_ | ~new_n8656_;
  assign new_n8625_ = new_n8636_ & new_n8637_;
  assign new_n8626_ = new_n8639_ & new_n8640_;
  assign new_n8627_ = new_n8642_ & new_n8643_;
  assign new_n8628_ = new_n8645_ & new_n8646_;
  assign new_n8629_ = ~new_n1378_;
  assign new_n8630_ = ~new_n1379_;
  assign new_n8631_ = ~new_n1372_ | ~new_n8630_;
  assign new_n8632_ = ~new_n1372_ | ~new_n8629_;
  assign new_n8633_ = new_n1378_ | new_n1379_;
  assign new_n8634_ = ~new_n1371_ | ~new_n8615_;
  assign new_n8635_ = ~new_n8631_ | ~new_n8632_ | ~new_n8634_ | ~new_n8633_;
  assign new_n8636_ = ~new_n1377_ | ~new_n8614_;
  assign new_n8637_ = ~new_n1376_ | ~new_n8617_;
  assign new_n8638_ = ~new_n8625_ | ~new_n8635_;
  assign new_n8639_ = ~new_n1370_ | ~new_n8616_;
  assign new_n8640_ = ~new_n1369_ | ~new_n8619_;
  assign new_n8641_ = ~new_n8626_ | ~new_n8638_;
  assign new_n8642_ = ~new_n1375_ | ~new_n8618_;
  assign new_n8643_ = ~new_n1374_ | ~new_n8621_;
  assign new_n8644_ = ~new_n8627_ | ~new_n8641_;
  assign new_n8645_ = ~new_n1368_ | ~new_n8620_;
  assign new_n8646_ = ~new_n1013_ | ~new_n8613_;
  assign new_n8647_ = ~new_n8628_ | ~new_n8644_;
  assign new_n8648_ = ~new_n1373_ | ~new_n8622_;
  assign new_n8649_ = ~new_n8647_ | ~new_n8648_;
  assign new_n8650_ = ~new_n1373_ | ~new_n8623_;
  assign new_n8651_ = ~new_n8649_ | ~new_n8613_;
  assign new_n8652_ = ~new_n8651_ | ~new_n8650_;
  assign new_n8653_ = ~pi109 | ~new_n8613_;
  assign new_n8654_ = ~new_n1373_ | ~new_n8649_;
  assign new_n8655_ = ~new_n8654_ | ~new_n8653_;
  assign new_n8656_ = ~new_n8652_ | ~new_n8622_;
  assign new_n8657_ = ~new_n1013_ | ~new_n8655_;
  assign new_n8658_ = ~new_n1877_;
  assign new_n8659_ = ~new_n1872_;
  assign new_n8660_ = ~new_n1878_;
  assign new_n8661_ = ~new_n1876_;
  assign new_n8662_ = ~new_n1871_;
  assign new_n8663_ = ~new_n1874_;
  assign new_n8664_ = ~new_n1873_;
  assign new_n8665_ = ~new_n1875_;
  assign new_n8666_ = new_n8669_ & new_n8668_;
  assign new_n8667_ = ~new_n1330_;
  assign new_n8668_ = ~new_n8265_ | ~new_n8667_;
  assign new_n8669_ = ~new_n8266_ | ~new_n8667_;
  assign new_n8670_ = ~new_n8674_ | ~new_n8673_;
  assign new_n8671_ = ~pi249;
  assign new_n8672_ = ~pi248;
  assign new_n8673_ = ~pi249 | ~new_n8672_;
  assign new_n8674_ = ~pi248 | ~new_n8671_;
  assign new_n8675_ = ~pi440;
  assign new_n8676_ = ~pi441;
  assign new_n8677_ = ~pi441 | ~pi440;
  assign new_n8678_ = ~pi442;
  assign new_n8679_ = ~pi442 | ~new_n8765_;
  assign new_n8680_ = ~pi443;
  assign new_n8681_ = ~pi443 | ~new_n8766_;
  assign new_n8682_ = ~pi444;
  assign new_n8683_ = ~pi444 | ~new_n8767_;
  assign new_n8684_ = ~pi445;
  assign new_n8685_ = ~pi445 | ~new_n8768_;
  assign new_n8686_ = ~pi446;
  assign new_n8687_ = ~pi446 | ~new_n8769_;
  assign new_n8688_ = ~pi447;
  assign new_n8689_ = ~pi448;
  assign new_n8690_ = ~pi447 | ~new_n8770_;
  assign new_n8691_ = ~new_n8771_ | ~pi448;
  assign new_n8692_ = ~pi449;
  assign new_n8693_ = ~pi449 | ~new_n8772_;
  assign new_n8694_ = ~pi450;
  assign new_n8695_ = ~pi450 | ~new_n8773_;
  assign new_n8696_ = ~pi451;
  assign new_n8697_ = ~pi451 | ~new_n8774_;
  assign new_n8698_ = ~pi452;
  assign new_n8699_ = ~pi452 | ~new_n8775_;
  assign new_n8700_ = ~pi453;
  assign new_n8701_ = ~pi453 | ~new_n8776_;
  assign new_n8702_ = ~pi454;
  assign new_n8703_ = ~pi454 | ~new_n8777_;
  assign new_n8704_ = ~pi455;
  assign new_n8705_ = ~pi455 | ~new_n8778_;
  assign new_n8706_ = ~pi456;
  assign new_n8707_ = ~pi456 | ~new_n8779_;
  assign new_n8708_ = ~pi457;
  assign new_n8709_ = ~pi457 | ~new_n8780_;
  assign new_n8710_ = ~pi458;
  assign new_n8711_ = ~pi458 | ~new_n8781_;
  assign new_n8712_ = ~pi459;
  assign new_n8713_ = ~pi459 | ~new_n8782_;
  assign new_n8714_ = ~pi460;
  assign new_n8715_ = ~pi460 | ~new_n8783_;
  assign new_n8716_ = ~pi461;
  assign new_n8717_ = ~pi461 | ~new_n8784_;
  assign new_n8718_ = ~pi462;
  assign new_n8719_ = ~pi462 | ~new_n8785_;
  assign new_n8720_ = ~pi463;
  assign new_n8721_ = ~pi463 | ~new_n8786_;
  assign new_n8722_ = ~pi464;
  assign new_n8723_ = ~pi464 | ~new_n8787_;
  assign new_n8724_ = ~pi465;
  assign new_n8725_ = ~pi465 | ~new_n8788_;
  assign new_n8726_ = ~pi466;
  assign new_n8727_ = ~pi466 | ~new_n8789_;
  assign new_n8728_ = ~pi467;
  assign new_n8729_ = ~pi467 | ~new_n8790_;
  assign new_n8730_ = ~pi468;
  assign new_n8731_ = ~pi468 | ~new_n8791_;
  assign new_n8732_ = ~pi469;
  assign new_n8733_ = ~new_n8795_ | ~new_n8794_;
  assign new_n8734_ = ~new_n8797_ | ~new_n8796_;
  assign new_n8735_ = ~new_n8799_ | ~new_n8798_;
  assign new_n8736_ = ~new_n8801_ | ~new_n8800_;
  assign new_n8737_ = ~new_n8803_ | ~new_n8802_;
  assign new_n8738_ = ~new_n8805_ | ~new_n8804_;
  assign new_n8739_ = ~new_n8807_ | ~new_n8806_;
  assign new_n8740_ = ~new_n8809_ | ~new_n8808_;
  assign new_n8741_ = ~new_n8811_ | ~new_n8810_;
  assign new_n8742_ = ~new_n8813_ | ~new_n8812_;
  assign new_n8743_ = ~new_n8815_ | ~new_n8814_;
  assign new_n8744_ = ~new_n8817_ | ~new_n8816_;
  assign new_n8745_ = ~new_n8819_ | ~new_n8818_;
  assign new_n8746_ = ~new_n8821_ | ~new_n8820_;
  assign new_n8747_ = ~new_n8823_ | ~new_n8822_;
  assign new_n8748_ = ~new_n8825_ | ~new_n8824_;
  assign new_n8749_ = ~new_n8827_ | ~new_n8826_;
  assign new_n8750_ = ~new_n8829_ | ~new_n8828_;
  assign new_n8751_ = ~new_n8831_ | ~new_n8830_;
  assign new_n8752_ = ~new_n8833_ | ~new_n8832_;
  assign new_n8753_ = ~new_n8835_ | ~new_n8834_;
  assign new_n8754_ = ~new_n8837_ | ~new_n8836_;
  assign new_n8755_ = ~new_n8839_ | ~new_n8838_;
  assign new_n8756_ = ~new_n8841_ | ~new_n8840_;
  assign new_n8757_ = ~new_n8843_ | ~new_n8842_;
  assign new_n8758_ = ~new_n8845_ | ~new_n8844_;
  assign new_n8759_ = ~new_n8847_ | ~new_n8846_;
  assign new_n8760_ = ~new_n8849_ | ~new_n8848_;
  assign new_n8761_ = ~new_n8851_ | ~new_n8850_;
  assign new_n8762_ = ~new_n8853_ | ~new_n8852_;
  assign new_n8763_ = ~pi470;
  assign new_n8764_ = ~pi469 | ~new_n8792_;
  assign new_n8765_ = ~new_n8677_;
  assign new_n8766_ = ~new_n8679_;
  assign new_n8767_ = ~new_n8681_;
  assign new_n8768_ = ~new_n8683_;
  assign new_n8769_ = ~new_n8685_;
  assign new_n8770_ = ~new_n8687_;
  assign new_n8771_ = ~new_n8690_;
  assign new_n8772_ = ~new_n8691_;
  assign new_n8773_ = ~new_n8693_;
  assign new_n8774_ = ~new_n8695_;
  assign new_n8775_ = ~new_n8697_;
  assign new_n8776_ = ~new_n8699_;
  assign new_n8777_ = ~new_n8701_;
  assign new_n8778_ = ~new_n8703_;
  assign new_n8779_ = ~new_n8705_;
  assign new_n8780_ = ~new_n8707_;
  assign new_n8781_ = ~new_n8709_;
  assign new_n8782_ = ~new_n8711_;
  assign new_n8783_ = ~new_n8713_;
  assign new_n8784_ = ~new_n8715_;
  assign new_n8785_ = ~new_n8717_;
  assign new_n8786_ = ~new_n8719_;
  assign new_n8787_ = ~new_n8721_;
  assign new_n8788_ = ~new_n8723_;
  assign new_n8789_ = ~new_n8725_;
  assign new_n8790_ = ~new_n8727_;
  assign new_n8791_ = ~new_n8729_;
  assign new_n8792_ = ~new_n8731_;
  assign new_n8793_ = ~new_n8764_;
  assign new_n8794_ = ~pi448 | ~new_n8690_;
  assign new_n8795_ = ~new_n8771_ | ~new_n8689_;
  assign new_n8796_ = ~pi447 | ~new_n8687_;
  assign new_n8797_ = ~new_n8770_ | ~new_n8688_;
  assign new_n8798_ = ~pi446 | ~new_n8685_;
  assign new_n8799_ = ~new_n8769_ | ~new_n8686_;
  assign new_n8800_ = ~pi445 | ~new_n8683_;
  assign new_n8801_ = ~new_n8768_ | ~new_n8684_;
  assign new_n8802_ = ~pi444 | ~new_n8681_;
  assign new_n8803_ = ~new_n8767_ | ~new_n8682_;
  assign new_n8804_ = ~pi443 | ~new_n8679_;
  assign new_n8805_ = ~new_n8766_ | ~new_n8680_;
  assign new_n8806_ = ~pi442 | ~new_n8677_;
  assign new_n8807_ = ~new_n8765_ | ~new_n8678_;
  assign new_n8808_ = ~pi470 | ~new_n8764_;
  assign new_n8809_ = ~new_n8793_ | ~new_n8763_;
  assign new_n8810_ = ~pi469 | ~new_n8731_;
  assign new_n8811_ = ~new_n8792_ | ~new_n8732_;
  assign new_n8812_ = ~pi441 | ~new_n8675_;
  assign new_n8813_ = ~pi440 | ~new_n8676_;
  assign new_n8814_ = ~pi468 | ~new_n8729_;
  assign new_n8815_ = ~new_n8791_ | ~new_n8730_;
  assign new_n8816_ = ~pi467 | ~new_n8727_;
  assign new_n8817_ = ~new_n8790_ | ~new_n8728_;
  assign new_n8818_ = ~pi466 | ~new_n8725_;
  assign new_n8819_ = ~new_n8789_ | ~new_n8726_;
  assign new_n8820_ = ~pi465 | ~new_n8723_;
  assign new_n8821_ = ~new_n8788_ | ~new_n8724_;
  assign new_n8822_ = ~pi464 | ~new_n8721_;
  assign new_n8823_ = ~new_n8787_ | ~new_n8722_;
  assign new_n8824_ = ~pi463 | ~new_n8719_;
  assign new_n8825_ = ~new_n8786_ | ~new_n8720_;
  assign new_n8826_ = ~pi462 | ~new_n8717_;
  assign new_n8827_ = ~new_n8785_ | ~new_n8718_;
  assign new_n8828_ = ~pi461 | ~new_n8715_;
  assign new_n8829_ = ~new_n8784_ | ~new_n8716_;
  assign new_n8830_ = ~pi460 | ~new_n8713_;
  assign new_n8831_ = ~new_n8783_ | ~new_n8714_;
  assign new_n8832_ = ~pi459 | ~new_n8711_;
  assign new_n8833_ = ~new_n8782_ | ~new_n8712_;
  assign new_n8834_ = ~pi458 | ~new_n8709_;
  assign new_n8835_ = ~new_n8781_ | ~new_n8710_;
  assign new_n8836_ = ~pi457 | ~new_n8707_;
  assign new_n8837_ = ~new_n8780_ | ~new_n8708_;
  assign new_n8838_ = ~pi456 | ~new_n8705_;
  assign new_n8839_ = ~new_n8779_ | ~new_n8706_;
  assign new_n8840_ = ~pi455 | ~new_n8703_;
  assign new_n8841_ = ~new_n8778_ | ~new_n8704_;
  assign new_n8842_ = ~pi454 | ~new_n8701_;
  assign new_n8843_ = ~new_n8777_ | ~new_n8702_;
  assign new_n8844_ = ~pi453 | ~new_n8699_;
  assign new_n8845_ = ~new_n8776_ | ~new_n8700_;
  assign new_n8846_ = ~pi452 | ~new_n8697_;
  assign new_n8847_ = ~new_n8775_ | ~new_n8698_;
  assign new_n8848_ = ~pi451 | ~new_n8695_;
  assign new_n8849_ = ~new_n8774_ | ~new_n8696_;
  assign new_n8850_ = ~pi450 | ~new_n8693_;
  assign new_n8851_ = ~new_n8773_ | ~new_n8694_;
  assign new_n8852_ = ~pi449 | ~new_n8691_;
  assign new_n8853_ = ~new_n8772_ | ~new_n8692_;
  assign new_n8854_ = new_n8875_ & new_n8874_;
  assign new_n8855_ = ~pi245;
  assign new_n8856_ = ~new_n2135_;
  assign new_n8857_ = ~new_n2134_;
  assign new_n8858_ = ~pi244;
  assign new_n8859_ = ~pi243;
  assign new_n8860_ = ~new_n2133_;
  assign new_n8861_ = new_n8869_ & new_n8870_;
  assign new_n8862_ = new_n8872_ & new_n8873_;
  assign new_n8863_ = ~new_n2136_;
  assign new_n8864_ = ~new_n2137_;
  assign new_n8865_ = ~pi247 | ~new_n8864_ | ~new_n8863_;
  assign new_n8866_ = ~pi246 | ~new_n8863_;
  assign new_n8867_ = ~pi245 | ~new_n8856_;
  assign new_n8868_ = ~new_n8865_ | ~new_n8866_ | ~new_n8876_ | ~new_n8867_;
  assign new_n8869_ = ~new_n2135_ | ~new_n8855_;
  assign new_n8870_ = ~new_n2134_ | ~new_n8858_;
  assign new_n8871_ = ~new_n8861_ | ~new_n8868_;
  assign new_n8872_ = ~pi244 | ~new_n8857_;
  assign new_n8873_ = ~pi243 | ~new_n8860_;
  assign new_n8874_ = ~new_n8862_ | ~new_n8871_;
  assign new_n8875_ = ~new_n2133_ | ~new_n8859_;
  assign new_n8876_ = ~new_n8864_ | ~pi247 | ~pi246;
  assign new_n8877_ = ~new_n8916_ | ~new_n8915_;
  assign new_n8878_ = ~new_n8880_ | ~new_n8917_;
  assign new_n8879_ = ~pi242;
  assign new_n8880_ = ~pi242 | ~new_n8889_;
  assign new_n8881_ = ~pi246;
  assign new_n8882_ = ~pi240;
  assign new_n8883_ = ~pi245;
  assign new_n8884_ = ~pi239;
  assign new_n8885_ = ~pi244;
  assign new_n8886_ = ~pi243;
  assign new_n8887_ = ~new_n8912_ | ~new_n8911_;
  assign new_n8888_ = ~pi238;
  assign new_n8889_ = ~pi247;
  assign new_n8890_ = ~new_n8922_ | ~new_n8921_;
  assign new_n8891_ = ~new_n8927_ | ~new_n8926_;
  assign new_n8892_ = ~new_n8932_ | ~new_n8931_;
  assign new_n8893_ = ~new_n8937_ | ~new_n8936_;
  assign new_n8894_ = ~new_n8919_ | ~new_n8918_;
  assign new_n8895_ = ~new_n8924_ | ~new_n8923_;
  assign new_n8896_ = ~new_n8929_ | ~new_n8928_;
  assign new_n8897_ = ~new_n8934_ | ~new_n8933_;
  assign new_n8898_ = ~new_n8908_ | ~new_n8907_;
  assign new_n8899_ = ~new_n8904_ | ~new_n8903_;
  assign new_n8900_ = ~pi241;
  assign new_n8901_ = ~new_n8880_;
  assign new_n8902_ = ~new_n8901_ | ~new_n8881_;
  assign new_n8903_ = ~new_n8902_ | ~new_n8900_;
  assign new_n8904_ = ~pi246 | ~new_n8880_;
  assign new_n8905_ = ~new_n8899_;
  assign new_n8906_ = ~pi240 | ~new_n8883_;
  assign new_n8907_ = ~new_n8906_ | ~new_n8899_;
  assign new_n8908_ = ~pi245 | ~new_n8882_;
  assign new_n8909_ = ~new_n8898_;
  assign new_n8910_ = ~pi239 | ~new_n8885_;
  assign new_n8911_ = ~new_n8910_ | ~new_n8898_;
  assign new_n8912_ = ~pi244 | ~new_n8884_;
  assign new_n8913_ = ~new_n8887_;
  assign new_n8914_ = ~pi243 | ~new_n8888_;
  assign new_n8915_ = ~new_n8913_ | ~new_n8914_;
  assign new_n8916_ = ~pi238 | ~new_n8886_;
  assign new_n8917_ = ~pi247 | ~new_n8879_;
  assign new_n8918_ = ~pi238 | ~new_n8886_;
  assign new_n8919_ = ~pi243 | ~new_n8888_;
  assign new_n8920_ = ~new_n8894_;
  assign new_n8921_ = ~new_n8920_ | ~new_n8913_;
  assign new_n8922_ = ~new_n8894_ | ~new_n8887_;
  assign new_n8923_ = ~pi239 | ~new_n8885_;
  assign new_n8924_ = ~pi244 | ~new_n8884_;
  assign new_n8925_ = ~new_n8895_;
  assign new_n8926_ = ~new_n8909_ | ~new_n8925_;
  assign new_n8927_ = ~new_n8895_ | ~new_n8898_;
  assign new_n8928_ = ~pi240 | ~new_n8883_;
  assign new_n8929_ = ~pi245 | ~new_n8882_;
  assign new_n8930_ = ~new_n8896_;
  assign new_n8931_ = ~new_n8905_ | ~new_n8930_;
  assign new_n8932_ = ~new_n8896_ | ~new_n8899_;
  assign new_n8933_ = ~pi241 | ~new_n8881_;
  assign new_n8934_ = ~pi246 | ~new_n8900_;
  assign new_n8935_ = ~new_n8897_;
  assign new_n8936_ = ~new_n8935_ | ~new_n8901_;
  assign new_n8937_ = ~new_n8897_ | ~new_n8880_;
  assign new_n8938_ = ~new_n8977_ | ~new_n8976_;
  assign new_n8939_ = ~new_n8941_ | ~new_n8978_;
  assign new_n8940_ = ~pi242;
  assign new_n8941_ = ~pi242 | ~new_n8950_;
  assign new_n8942_ = ~pi246;
  assign new_n8943_ = ~pi240;
  assign new_n8944_ = ~pi245;
  assign new_n8945_ = ~pi239;
  assign new_n8946_ = ~pi244;
  assign new_n8947_ = ~pi243;
  assign new_n8948_ = ~new_n8973_ | ~new_n8972_;
  assign new_n8949_ = ~pi238;
  assign new_n8950_ = ~pi247;
  assign new_n8951_ = ~new_n8983_ | ~new_n8982_;
  assign new_n8952_ = ~new_n8988_ | ~new_n8987_;
  assign new_n8953_ = ~new_n8993_ | ~new_n8992_;
  assign new_n8954_ = ~new_n8998_ | ~new_n8997_;
  assign new_n8955_ = ~new_n8980_ | ~new_n8979_;
  assign new_n8956_ = ~new_n8985_ | ~new_n8984_;
  assign new_n8957_ = ~new_n8990_ | ~new_n8989_;
  assign new_n8958_ = ~new_n8995_ | ~new_n8994_;
  assign new_n8959_ = ~new_n8969_ | ~new_n8968_;
  assign new_n8960_ = ~new_n8965_ | ~new_n8964_;
  assign new_n8961_ = ~pi241;
  assign new_n8962_ = ~new_n8941_;
  assign new_n8963_ = ~new_n8962_ | ~new_n8942_;
  assign new_n8964_ = ~new_n8963_ | ~new_n8961_;
  assign new_n8965_ = ~pi246 | ~new_n8941_;
  assign new_n8966_ = ~new_n8960_;
  assign new_n8967_ = ~pi240 | ~new_n8944_;
  assign new_n8968_ = ~new_n8967_ | ~new_n8960_;
  assign new_n8969_ = ~pi245 | ~new_n8943_;
  assign new_n8970_ = ~new_n8959_;
  assign new_n8971_ = ~pi239 | ~new_n8946_;
  assign new_n8972_ = ~new_n8971_ | ~new_n8959_;
  assign new_n8973_ = ~pi244 | ~new_n8945_;
  assign new_n8974_ = ~new_n8948_;
  assign new_n8975_ = ~pi243 | ~new_n8949_;
  assign new_n8976_ = ~new_n8974_ | ~new_n8975_;
  assign new_n8977_ = ~pi238 | ~new_n8947_;
  assign new_n8978_ = ~pi247 | ~new_n8940_;
  assign new_n8979_ = ~pi238 | ~new_n8947_;
  assign new_n8980_ = ~pi243 | ~new_n8949_;
  assign new_n8981_ = ~new_n8955_;
  assign new_n8982_ = ~new_n8981_ | ~new_n8974_;
  assign new_n8983_ = ~new_n8955_ | ~new_n8948_;
  assign new_n8984_ = ~pi239 | ~new_n8946_;
  assign new_n8985_ = ~pi244 | ~new_n8945_;
  assign new_n8986_ = ~new_n8956_;
  assign new_n8987_ = ~new_n8970_ | ~new_n8986_;
  assign new_n8988_ = ~new_n8956_ | ~new_n8959_;
  assign new_n8989_ = ~pi240 | ~new_n8944_;
  assign new_n8990_ = ~pi245 | ~new_n8943_;
  assign new_n8991_ = ~new_n8957_;
  assign new_n8992_ = ~new_n8966_ | ~new_n8991_;
  assign new_n8993_ = ~new_n8957_ | ~new_n8960_;
  assign new_n8994_ = ~pi241 | ~new_n8942_;
  assign new_n8995_ = ~pi246 | ~new_n8961_;
  assign new_n8996_ = ~new_n8958_;
  assign new_n8997_ = ~new_n8996_ | ~new_n8962_;
  assign new_n8998_ = ~new_n8958_ | ~new_n8941_;
  assign new_n8999_ = ~new_n1871_;
  assign new_n9000_ = ~new_n9019_ | ~new_n9027_;
  assign new_n9001_ = new_n9017_ & new_n9025_;
  assign new_n9002_ = ~new_n1872_;
  assign new_n9003_ = ~new_n1874_;
  assign new_n9004_ = ~new_n1874_ | ~new_n9019_;
  assign new_n9005_ = ~new_n1875_;
  assign new_n9006_ = ~new_n1875_ | ~new_n9023_;
  assign new_n9007_ = ~new_n1876_;
  assign new_n9008_ = ~new_n1876_ | ~new_n9024_;
  assign new_n9009_ = ~new_n1878_;
  assign new_n9010_ = ~new_n1877_;
  assign new_n9011_ = ~new_n1873_;
  assign new_n9012_ = ~new_n9029_ | ~new_n9028_;
  assign new_n9013_ = ~new_n9031_ | ~new_n9030_;
  assign new_n9014_ = ~new_n9033_ | ~new_n9032_;
  assign new_n9015_ = ~new_n9035_ | ~new_n9034_;
  assign new_n9016_ = ~new_n9039_ | ~new_n9038_;
  assign new_n9017_ = new_n1878_ & new_n1877_;
  assign new_n9018_ = ~new_n1877_ | ~new_n9025_;
  assign new_n9019_ = ~new_n9011_ | ~new_n9021_;
  assign new_n9020_ = new_n9037_ & new_n9036_;
  assign new_n9021_ = ~new_n1872_ | ~new_n1871_;
  assign new_n9022_ = ~new_n9019_;
  assign new_n9023_ = ~new_n9004_;
  assign new_n9024_ = ~new_n9006_;
  assign new_n9025_ = ~new_n9008_;
  assign new_n9026_ = ~new_n9018_;
  assign new_n9027_ = ~new_n1873_ | ~new_n1872_ | ~new_n1871_;
  assign new_n9028_ = ~new_n1878_ | ~new_n9018_;
  assign new_n9029_ = ~new_n9026_ | ~new_n9009_;
  assign new_n9030_ = ~new_n1877_ | ~new_n9008_;
  assign new_n9031_ = ~new_n9025_ | ~new_n9010_;
  assign new_n9032_ = ~new_n1876_ | ~new_n9006_;
  assign new_n9033_ = ~new_n9024_ | ~new_n9007_;
  assign new_n9034_ = ~new_n1875_ | ~new_n9004_;
  assign new_n9035_ = ~new_n9023_ | ~new_n9005_;
  assign new_n9036_ = ~new_n1874_ | ~new_n9019_;
  assign new_n9037_ = ~new_n9022_ | ~new_n9003_;
  assign new_n9038_ = ~new_n1872_ | ~new_n8999_;
  assign new_n9039_ = ~new_n1871_ | ~new_n9002_;
  assign new_n9040_ = ~pi248;
  assign new_n9041_ = ~new_n9128_ | ~new_n9162_;
  assign new_n9042_ = ~pi249;
  assign new_n9043_ = ~pi251;
  assign new_n9044_ = ~pi251 | ~new_n9128_;
  assign new_n9045_ = ~pi252;
  assign new_n9046_ = ~pi252 | ~new_n9134_;
  assign new_n9047_ = ~pi253;
  assign new_n9048_ = ~pi253 | ~new_n9135_;
  assign new_n9049_ = ~pi254;
  assign new_n9050_ = ~pi254 | ~new_n9136_;
  assign new_n9051_ = ~pi255;
  assign new_n9052_ = ~pi255 | ~new_n9137_;
  assign new_n9053_ = ~pi256;
  assign new_n9054_ = ~pi257;
  assign new_n9055_ = ~pi256 | ~new_n9138_;
  assign new_n9056_ = ~new_n9139_ | ~pi257;
  assign new_n9057_ = ~pi258;
  assign new_n9058_ = ~pi258 | ~new_n9140_;
  assign new_n9059_ = ~pi259;
  assign new_n9060_ = ~pi259 | ~new_n9141_;
  assign new_n9061_ = ~pi260;
  assign new_n9062_ = ~pi260 | ~new_n9142_;
  assign new_n9063_ = ~pi261;
  assign new_n9064_ = ~pi261 | ~new_n9143_;
  assign new_n9065_ = ~pi262;
  assign new_n9066_ = ~pi262 | ~new_n9144_;
  assign new_n9067_ = ~pi263;
  assign new_n9068_ = ~pi263 | ~new_n9145_;
  assign new_n9069_ = ~pi264;
  assign new_n9070_ = ~pi264 | ~new_n9146_;
  assign new_n9071_ = ~pi265;
  assign new_n9072_ = ~pi265 | ~new_n9147_;
  assign new_n9073_ = ~pi266;
  assign new_n9074_ = ~pi266 | ~new_n9148_;
  assign new_n9075_ = ~pi267;
  assign new_n9076_ = ~pi267 | ~new_n9149_;
  assign new_n9077_ = ~pi268;
  assign new_n9078_ = ~pi268 | ~new_n9150_;
  assign new_n9079_ = ~pi269;
  assign new_n9080_ = ~pi269 | ~new_n9151_;
  assign new_n9081_ = ~pi270;
  assign new_n9082_ = ~pi270 | ~new_n9152_;
  assign new_n9083_ = ~pi271;
  assign new_n9084_ = ~pi271 | ~new_n9153_;
  assign new_n9085_ = ~pi272;
  assign new_n9086_ = ~pi272 | ~new_n9154_;
  assign new_n9087_ = ~pi273;
  assign new_n9088_ = ~pi273 | ~new_n9155_;
  assign new_n9089_ = ~pi274;
  assign new_n9090_ = ~pi274 | ~new_n9156_;
  assign new_n9091_ = ~pi275;
  assign new_n9092_ = ~pi275 | ~new_n9157_;
  assign new_n9093_ = ~pi276;
  assign new_n9094_ = ~pi276 | ~new_n9158_;
  assign new_n9095_ = ~pi277;
  assign new_n9096_ = ~pi277 | ~new_n9159_;
  assign new_n9097_ = ~pi278;
  assign new_n9098_ = ~pi250;
  assign new_n9099_ = ~new_n9164_ | ~new_n9163_;
  assign new_n9100_ = ~new_n9166_ | ~new_n9165_;
  assign new_n9101_ = ~new_n9168_ | ~new_n9167_;
  assign new_n9102_ = ~new_n9170_ | ~new_n9169_;
  assign new_n9103_ = ~new_n9172_ | ~new_n9171_;
  assign new_n9104_ = ~new_n9174_ | ~new_n9173_;
  assign new_n9105_ = ~new_n9178_ | ~new_n9177_;
  assign new_n9106_ = ~new_n9180_ | ~new_n9179_;
  assign new_n9107_ = ~new_n9182_ | ~new_n9181_;
  assign new_n9108_ = ~new_n9184_ | ~new_n9183_;
  assign new_n9109_ = ~new_n9186_ | ~new_n9185_;
  assign new_n9110_ = ~new_n9188_ | ~new_n9187_;
  assign new_n9111_ = ~new_n9190_ | ~new_n9189_;
  assign new_n9112_ = ~new_n9192_ | ~new_n9191_;
  assign new_n9113_ = ~new_n9194_ | ~new_n9193_;
  assign new_n9114_ = ~new_n9196_ | ~new_n9195_;
  assign new_n9115_ = ~new_n9198_ | ~new_n9197_;
  assign new_n9116_ = ~new_n9200_ | ~new_n9199_;
  assign new_n9117_ = ~new_n9202_ | ~new_n9201_;
  assign new_n9118_ = ~new_n9204_ | ~new_n9203_;
  assign new_n9119_ = ~new_n9206_ | ~new_n9205_;
  assign new_n9120_ = ~new_n9208_ | ~new_n9207_;
  assign new_n9121_ = ~new_n9210_ | ~new_n9209_;
  assign new_n9122_ = ~new_n9212_ | ~new_n9211_;
  assign new_n9123_ = ~new_n9214_ | ~new_n9213_;
  assign new_n9124_ = ~new_n9216_ | ~new_n9215_;
  assign new_n9125_ = ~new_n9218_ | ~new_n9217_;
  assign new_n9126_ = ~new_n9220_ | ~new_n9219_;
  assign new_n9127_ = ~new_n9222_ | ~new_n9221_;
  assign new_n9128_ = ~new_n9098_ | ~new_n9132_;
  assign new_n9129_ = new_n9176_ & new_n9175_;
  assign new_n9130_ = ~pi279;
  assign new_n9131_ = ~pi278 | ~new_n9160_;
  assign new_n9132_ = ~pi249 | ~pi248;
  assign new_n9133_ = ~new_n9128_;
  assign new_n9134_ = ~new_n9044_;
  assign new_n9135_ = ~new_n9046_;
  assign new_n9136_ = ~new_n9048_;
  assign new_n9137_ = ~new_n9050_;
  assign new_n9138_ = ~new_n9052_;
  assign new_n9139_ = ~new_n9055_;
  assign new_n9140_ = ~new_n9056_;
  assign new_n9141_ = ~new_n9058_;
  assign new_n9142_ = ~new_n9060_;
  assign new_n9143_ = ~new_n9062_;
  assign new_n9144_ = ~new_n9064_;
  assign new_n9145_ = ~new_n9066_;
  assign new_n9146_ = ~new_n9068_;
  assign new_n9147_ = ~new_n9070_;
  assign new_n9148_ = ~new_n9072_;
  assign new_n9149_ = ~new_n9074_;
  assign new_n9150_ = ~new_n9076_;
  assign new_n9151_ = ~new_n9078_;
  assign new_n9152_ = ~new_n9080_;
  assign new_n9153_ = ~new_n9082_;
  assign new_n9154_ = ~new_n9084_;
  assign new_n9155_ = ~new_n9086_;
  assign new_n9156_ = ~new_n9088_;
  assign new_n9157_ = ~new_n9090_;
  assign new_n9158_ = ~new_n9092_;
  assign new_n9159_ = ~new_n9094_;
  assign new_n9160_ = ~new_n9096_;
  assign new_n9161_ = ~new_n9131_;
  assign new_n9162_ = ~pi250 | ~pi249 | ~pi248;
  assign new_n9163_ = ~pi257 | ~new_n9055_;
  assign new_n9164_ = ~new_n9139_ | ~new_n9054_;
  assign new_n9165_ = ~pi256 | ~new_n9052_;
  assign new_n9166_ = ~new_n9138_ | ~new_n9053_;
  assign new_n9167_ = ~pi255 | ~new_n9050_;
  assign new_n9168_ = ~new_n9137_ | ~new_n9051_;
  assign new_n9169_ = ~pi254 | ~new_n9048_;
  assign new_n9170_ = ~new_n9136_ | ~new_n9049_;
  assign new_n9171_ = ~pi253 | ~new_n9046_;
  assign new_n9172_ = ~new_n9135_ | ~new_n9047_;
  assign new_n9173_ = ~pi252 | ~new_n9044_;
  assign new_n9174_ = ~new_n9134_ | ~new_n9045_;
  assign new_n9175_ = ~pi251 | ~new_n9128_;
  assign new_n9176_ = ~new_n9133_ | ~new_n9043_;
  assign new_n9177_ = ~pi279 | ~new_n9131_;
  assign new_n9178_ = ~new_n9161_ | ~new_n9130_;
  assign new_n9179_ = ~pi278 | ~new_n9096_;
  assign new_n9180_ = ~new_n9160_ | ~new_n9097_;
  assign new_n9181_ = ~pi277 | ~new_n9094_;
  assign new_n9182_ = ~new_n9159_ | ~new_n9095_;
  assign new_n9183_ = ~pi276 | ~new_n9092_;
  assign new_n9184_ = ~new_n9158_ | ~new_n9093_;
  assign new_n9185_ = ~pi275 | ~new_n9090_;
  assign new_n9186_ = ~new_n9157_ | ~new_n9091_;
  assign new_n9187_ = ~pi274 | ~new_n9088_;
  assign new_n9188_ = ~new_n9156_ | ~new_n9089_;
  assign new_n9189_ = ~pi273 | ~new_n9086_;
  assign new_n9190_ = ~new_n9155_ | ~new_n9087_;
  assign new_n9191_ = ~pi272 | ~new_n9084_;
  assign new_n9192_ = ~new_n9154_ | ~new_n9085_;
  assign new_n9193_ = ~pi271 | ~new_n9082_;
  assign new_n9194_ = ~new_n9153_ | ~new_n9083_;
  assign new_n9195_ = ~pi270 | ~new_n9080_;
  assign new_n9196_ = ~new_n9152_ | ~new_n9081_;
  assign new_n9197_ = ~pi269 | ~new_n9078_;
  assign new_n9198_ = ~new_n9151_ | ~new_n9079_;
  assign new_n9199_ = ~pi268 | ~new_n9076_;
  assign new_n9200_ = ~new_n9150_ | ~new_n9077_;
  assign new_n9201_ = ~pi249 | ~new_n9040_;
  assign new_n9202_ = ~pi248 | ~new_n9042_;
  assign new_n9203_ = ~pi267 | ~new_n9074_;
  assign new_n9204_ = ~new_n9149_ | ~new_n9075_;
  assign new_n9205_ = ~pi266 | ~new_n9072_;
  assign new_n9206_ = ~new_n9148_ | ~new_n9073_;
  assign new_n9207_ = ~pi265 | ~new_n9070_;
  assign new_n9208_ = ~new_n9147_ | ~new_n9071_;
  assign new_n9209_ = ~pi264 | ~new_n9068_;
  assign new_n9210_ = ~new_n9146_ | ~new_n9069_;
  assign new_n9211_ = ~pi263 | ~new_n9066_;
  assign new_n9212_ = ~new_n9145_ | ~new_n9067_;
  assign new_n9213_ = ~pi262 | ~new_n9064_;
  assign new_n9214_ = ~new_n9144_ | ~new_n9065_;
  assign new_n9215_ = ~pi261 | ~new_n9062_;
  assign new_n9216_ = ~new_n9143_ | ~new_n9063_;
  assign new_n9217_ = ~pi260 | ~new_n9060_;
  assign new_n9218_ = ~new_n9142_ | ~new_n9061_;
  assign new_n9219_ = ~pi259 | ~new_n9058_;
  assign new_n9220_ = ~new_n9141_ | ~new_n9059_;
  assign new_n9221_ = ~pi258 | ~new_n9056_;
  assign new_n9222_ = ~new_n9140_ | ~new_n9057_;
  assign new_n9223_ = ~new_n8877_ & ~new_n9224_;
  assign new_n9224_ = ~new_n8891_ & ~new_n8892_ & ~new_n8893_ & ~new_n8890_;
  assign new_n9225_ = ~pi249;
  assign new_n9226_ = ~pi250;
  assign new_n9227_ = ~pi250 | ~pi249;
  assign new_n9228_ = ~pi251;
  assign new_n9229_ = ~pi251 | ~new_n9315_;
  assign new_n9230_ = ~pi252;
  assign new_n9231_ = ~pi252 | ~new_n9316_;
  assign new_n9232_ = ~pi253;
  assign new_n9233_ = ~pi253 | ~new_n9317_;
  assign new_n9234_ = ~pi254;
  assign new_n9235_ = ~pi254 | ~new_n9318_;
  assign new_n9236_ = ~pi255;
  assign new_n9237_ = ~pi255 | ~new_n9319_;
  assign new_n9238_ = ~pi256;
  assign new_n9239_ = ~pi257;
  assign new_n9240_ = ~pi256 | ~new_n9320_;
  assign new_n9241_ = ~new_n9321_ | ~pi257;
  assign new_n9242_ = ~pi258;
  assign new_n9243_ = ~pi258 | ~new_n9322_;
  assign new_n9244_ = ~pi259;
  assign new_n9245_ = ~pi259 | ~new_n9323_;
  assign new_n9246_ = ~pi260;
  assign new_n9247_ = ~pi260 | ~new_n9324_;
  assign new_n9248_ = ~pi261;
  assign new_n9249_ = ~pi261 | ~new_n9325_;
  assign new_n9250_ = ~pi262;
  assign new_n9251_ = ~pi262 | ~new_n9326_;
  assign new_n9252_ = ~pi263;
  assign new_n9253_ = ~pi263 | ~new_n9327_;
  assign new_n9254_ = ~pi264;
  assign new_n9255_ = ~pi264 | ~new_n9328_;
  assign new_n9256_ = ~pi265;
  assign new_n9257_ = ~pi265 | ~new_n9329_;
  assign new_n9258_ = ~pi266;
  assign new_n9259_ = ~pi266 | ~new_n9330_;
  assign new_n9260_ = ~pi267;
  assign new_n9261_ = ~pi267 | ~new_n9331_;
  assign new_n9262_ = ~pi268;
  assign new_n9263_ = ~pi268 | ~new_n9332_;
  assign new_n9264_ = ~pi269;
  assign new_n9265_ = ~pi269 | ~new_n9333_;
  assign new_n9266_ = ~pi270;
  assign new_n9267_ = ~pi270 | ~new_n9334_;
  assign new_n9268_ = ~pi271;
  assign new_n9269_ = ~pi271 | ~new_n9335_;
  assign new_n9270_ = ~pi272;
  assign new_n9271_ = ~pi272 | ~new_n9336_;
  assign new_n9272_ = ~pi273;
  assign new_n9273_ = ~pi273 | ~new_n9337_;
  assign new_n9274_ = ~pi274;
  assign new_n9275_ = ~pi274 | ~new_n9338_;
  assign new_n9276_ = ~pi275;
  assign new_n9277_ = ~pi275 | ~new_n9339_;
  assign new_n9278_ = ~pi276;
  assign new_n9279_ = ~pi276 | ~new_n9340_;
  assign new_n9280_ = ~pi277;
  assign new_n9281_ = ~pi277 | ~new_n9341_;
  assign new_n9282_ = ~pi278;
  assign new_n9283_ = ~new_n9345_ | ~new_n9344_;
  assign new_n9284_ = ~new_n9347_ | ~new_n9346_;
  assign new_n9285_ = ~new_n9349_ | ~new_n9348_;
  assign new_n9286_ = ~new_n9351_ | ~new_n9350_;
  assign new_n9287_ = ~new_n9353_ | ~new_n9352_;
  assign new_n9288_ = ~new_n9355_ | ~new_n9354_;
  assign new_n9289_ = ~new_n9357_ | ~new_n9356_;
  assign new_n9290_ = ~new_n9359_ | ~new_n9358_;
  assign new_n9291_ = ~new_n9361_ | ~new_n9360_;
  assign new_n9292_ = ~new_n9363_ | ~new_n9362_;
  assign new_n9293_ = ~new_n9365_ | ~new_n9364_;
  assign new_n9294_ = ~new_n9367_ | ~new_n9366_;
  assign new_n9295_ = ~new_n9369_ | ~new_n9368_;
  assign new_n9296_ = ~new_n9371_ | ~new_n9370_;
  assign new_n9297_ = ~new_n6466_ | ~new_n9372_;
  assign new_n9298_ = ~new_n6464_ | ~new_n6465_;
  assign new_n9299_ = ~new_n6462_ | ~new_n6463_;
  assign new_n9300_ = ~new_n6460_ | ~new_n6461_;
  assign new_n9301_ = ~new_n6458_ | ~new_n6459_;
  assign new_n9302_ = ~new_n6456_ | ~new_n6457_;
  assign new_n9303_ = ~new_n6454_ | ~new_n6455_;
  assign new_n9304_ = ~new_n6452_ | ~new_n6453_;
  assign new_n9305_ = ~new_n6450_ | ~new_n6451_;
  assign new_n9306_ = ~new_n6448_ | ~new_n6449_;
  assign new_n9307_ = ~new_n6446_ | ~new_n6447_;
  assign new_n9308_ = ~new_n6444_ | ~new_n6445_;
  assign new_n9309_ = ~new_n6442_ | ~new_n6443_;
  assign new_n9310_ = ~new_n6440_ | ~new_n6441_;
  assign new_n9311_ = ~new_n1008_ | ~new_n1276_;
  assign new_n9312_ = ~new_n1006_ | ~new_n1007_;
  assign new_n9313_ = ~pi279;
  assign new_n9314_ = ~pi278 | ~new_n9342_;
  assign new_n9315_ = ~new_n9227_;
  assign new_n9316_ = ~new_n9229_;
  assign new_n9317_ = ~new_n9231_;
  assign new_n9318_ = ~new_n9233_;
  assign new_n9319_ = ~new_n9235_;
  assign new_n9320_ = ~new_n9237_;
  assign new_n9321_ = ~new_n9240_;
  assign new_n9322_ = ~new_n9241_;
  assign new_n9323_ = ~new_n9243_;
  assign new_n9324_ = ~new_n9245_;
  assign new_n9325_ = ~new_n9247_;
  assign new_n9326_ = ~new_n9249_;
  assign new_n9327_ = ~new_n9251_;
  assign new_n9328_ = ~new_n9253_;
  assign new_n9329_ = ~new_n9255_;
  assign new_n9330_ = ~new_n9257_;
  assign new_n9331_ = ~new_n9259_;
  assign new_n9332_ = ~new_n9261_;
  assign new_n9333_ = ~new_n9263_;
  assign new_n9334_ = ~new_n9265_;
  assign new_n9335_ = ~new_n9267_;
  assign new_n9336_ = ~new_n9269_;
  assign new_n9337_ = ~new_n9271_;
  assign new_n9338_ = ~new_n9273_;
  assign new_n9339_ = ~new_n9275_;
  assign new_n9340_ = ~new_n9277_;
  assign new_n9341_ = ~new_n9279_;
  assign new_n9342_ = ~new_n9281_;
  assign new_n9343_ = ~new_n9314_;
  assign new_n9344_ = ~pi257 | ~new_n9240_;
  assign new_n9345_ = ~new_n9321_ | ~new_n9239_;
  assign new_n9346_ = ~pi256 | ~new_n9237_;
  assign new_n9347_ = ~new_n9320_ | ~new_n9238_;
  assign new_n9348_ = ~pi255 | ~new_n9235_;
  assign new_n9349_ = ~new_n9319_ | ~new_n9236_;
  assign new_n9350_ = ~pi254 | ~new_n9233_;
  assign new_n9351_ = ~new_n9318_ | ~new_n9234_;
  assign new_n9352_ = ~pi253 | ~new_n9231_;
  assign new_n9353_ = ~new_n9317_ | ~new_n9232_;
  assign new_n9354_ = ~pi252 | ~new_n9229_;
  assign new_n9355_ = ~new_n9316_ | ~new_n9230_;
  assign new_n9356_ = ~pi251 | ~new_n9227_;
  assign new_n9357_ = ~new_n9315_ | ~new_n9228_;
  assign new_n9358_ = ~pi279 | ~new_n9314_;
  assign new_n9359_ = ~new_n9343_ | ~new_n9313_;
  assign new_n9360_ = ~pi278 | ~new_n9281_;
  assign new_n9361_ = ~new_n9342_ | ~new_n9282_;
  assign new_n9362_ = ~pi250 | ~new_n9225_;
  assign new_n9363_ = ~pi249 | ~new_n9226_;
  assign new_n9364_ = ~pi277 | ~new_n9279_;
  assign new_n9365_ = ~new_n9341_ | ~new_n9280_;
  assign new_n9366_ = ~pi276 | ~new_n9277_;
  assign new_n9367_ = ~new_n9340_ | ~new_n9278_;
  assign new_n9368_ = ~pi275 | ~new_n9275_;
  assign new_n9369_ = ~new_n9339_ | ~new_n9276_;
  assign new_n9370_ = ~pi274 | ~new_n9273_;
  assign new_n9371_ = ~new_n9338_ | ~new_n9274_;
  assign new_n9372_ = ~pi273 | ~new_n9271_;
  assign po000 = pi037;
  assign po001 = pi038;
  assign po002 = pi039;
  assign po003 = pi040;
  assign po004 = pi041;
  assign po005 = pi042;
  assign po006 = pi043;
  assign po007 = pi044;
  assign po008 = pi045;
  assign po009 = pi046;
  assign po010 = pi047;
  assign po011 = pi048;
  assign po012 = pi049;
  assign po013 = pi050;
  assign po014 = pi051;
  assign po015 = pi052;
  assign po016 = pi053;
  assign po017 = pi054;
  assign po018 = pi055;
  assign po019 = pi056;
  assign po020 = pi057;
  assign po021 = pi058;
  assign po022 = pi059;
  assign po023 = pi060;
  assign po024 = pi061;
  assign po025 = pi062;
  assign po026 = pi063;
  assign po027 = pi064;
  assign po028 = pi065;
  assign po029 = pi066;
  assign po030 = pi067;
  assign po031 = pi068;
  assign po032 = pi069;
  assign po033 = pi070;
  assign po034 = pi475;
  assign po035 = pi480;
  assign po036 = pi481;
  assign po037 = pi483;
  assign po038 = pi374;
  assign po039 = pi373;
  assign po040 = pi372;
  assign po041 = pi371;
  assign po042 = pi370;
  assign po043 = pi369;
  assign po044 = pi368;
  assign po045 = pi367;
  assign po046 = pi366;
  assign po047 = pi365;
  assign po048 = pi364;
  assign po049 = pi363;
  assign po050 = pi362;
  assign po051 = pi361;
  assign po052 = pi360;
  assign po053 = pi359;
  assign po054 = pi358;
  assign po055 = pi357;
  assign po056 = pi356;
  assign po057 = pi355;
  assign po058 = pi354;
  assign po059 = pi353;
  assign po060 = pi352;
  assign po061 = pi351;
  assign po062 = pi350;
  assign po063 = pi349;
  assign po064 = pi348;
  assign po065 = pi347;
  assign po066 = pi346;
  assign po067 = pi345;
  assign po068 = pi344;
  assign po069 = pi343;
endmodule


